
module ALU_VARIABLE ( a, b, op, c_in, result, c_out, z, n, v );
  input [31:0] a;
  input [31:0] b;
  input [3:0] op;
  output [31:0] result;
  input c_in;
  output c_out, z, n, v;
  wire   mult_x_18_n726, mult_x_18_n725, mult_x_18_n724, mult_x_18_n723,
         mult_x_18_n722, mult_x_18_n721, mult_x_18_n720, mult_x_18_n719,
         mult_x_18_n718, mult_x_18_n717, mult_x_18_n716, mult_x_18_n715,
         mult_x_18_n714, mult_x_18_n713, mult_x_18_n712, mult_x_18_n711,
         mult_x_18_n710, mult_x_18_n709, mult_x_18_n708, mult_x_18_n707,
         mult_x_18_n706, mult_x_18_n705, mult_x_18_n704, mult_x_18_n699,
         mult_x_18_n698, mult_x_18_n697, mult_x_18_n696, mult_x_18_n695,
         mult_x_18_n694, mult_x_18_n693, mult_x_18_n692, mult_x_18_n691,
         mult_x_18_n690, mult_x_18_n689, mult_x_18_n688, mult_x_18_n687,
         mult_x_18_n686, mult_x_18_n685, mult_x_18_n684, mult_x_18_n683,
         mult_x_18_n682, mult_x_18_n681, mult_x_18_n680, mult_x_18_n679,
         mult_x_18_n678, mult_x_18_n677, mult_x_18_n669, mult_x_18_n668,
         mult_x_18_n667, mult_x_18_n666, mult_x_18_n665, mult_x_18_n664,
         mult_x_18_n663, mult_x_18_n662, mult_x_18_n661, mult_x_18_n660,
         mult_x_18_n659, mult_x_18_n658, mult_x_18_n657, mult_x_18_n656,
         mult_x_18_n655, mult_x_18_n654, mult_x_18_n653, mult_x_18_n648,
         mult_x_18_n647, mult_x_18_n646, mult_x_18_n645, mult_x_18_n644,
         mult_x_18_n643, mult_x_18_n642, mult_x_18_n641, mult_x_18_n640,
         mult_x_18_n639, mult_x_18_n638, mult_x_18_n637, mult_x_18_n636,
         mult_x_18_n635, mult_x_18_n634, mult_x_18_n633, mult_x_18_n632,
         mult_x_18_n624, mult_x_18_n623, mult_x_18_n622, mult_x_18_n621,
         mult_x_18_n620, mult_x_18_n619, mult_x_18_n618, mult_x_18_n617,
         mult_x_18_n616, mult_x_18_n615, mult_x_18_n614, mult_x_18_n609,
         mult_x_18_n608, mult_x_18_n607, mult_x_18_n606, mult_x_18_n605,
         mult_x_18_n604, mult_x_18_n603, mult_x_18_n602, mult_x_18_n601,
         mult_x_18_n600, mult_x_18_n599, mult_x_18_n591, mult_x_18_n590,
         mult_x_18_n589, mult_x_18_n588, mult_x_18_n587, mult_x_18_n582,
         mult_x_18_n581, mult_x_18_n580, mult_x_18_n579, mult_x_18_n578,
         mult_x_18_n467, mult_x_18_n465, mult_x_18_n464, mult_x_18_n462,
         mult_x_18_n461, mult_x_18_n460, mult_x_18_n459, mult_x_18_n457,
         mult_x_18_n456, mult_x_18_n455, mult_x_18_n454, mult_x_18_n452,
         mult_x_18_n451, mult_x_18_n450, mult_x_18_n447, mult_x_18_n445,
         mult_x_18_n444, mult_x_18_n443, mult_x_18_n440, mult_x_18_n438,
         mult_x_18_n437, mult_x_18_n436, mult_x_18_n434, mult_x_18_n433,
         mult_x_18_n432, mult_x_18_n431, mult_x_18_n430, mult_x_18_n429,
         mult_x_18_n428, mult_x_18_n426, mult_x_18_n425, mult_x_18_n424,
         mult_x_18_n423, mult_x_18_n422, mult_x_18_n421, mult_x_18_n420,
         mult_x_18_n418, mult_x_18_n417, mult_x_18_n416, mult_x_18_n415,
         mult_x_18_n414, mult_x_18_n413, mult_x_18_n412, mult_x_18_n410,
         mult_x_18_n409, mult_x_18_n408, mult_x_18_n407, mult_x_18_n406,
         mult_x_18_n405, mult_x_18_n402, mult_x_18_n400, mult_x_18_n399,
         mult_x_18_n398, mult_x_18_n397, mult_x_18_n396, mult_x_18_n395,
         mult_x_18_n392, mult_x_18_n390, mult_x_18_n389, mult_x_18_n388,
         mult_x_18_n387, mult_x_18_n386, mult_x_18_n385, mult_x_18_n383,
         mult_x_18_n382, mult_x_18_n381, mult_x_18_n380, mult_x_18_n379,
         mult_x_18_n378, mult_x_18_n377, mult_x_18_n376, mult_x_18_n375,
         mult_x_18_n374, mult_x_18_n372, mult_x_18_n371, mult_x_18_n370,
         mult_x_18_n369, mult_x_18_n368, mult_x_18_n367, mult_x_18_n366,
         mult_x_18_n365, mult_x_18_n364, mult_x_18_n363, mult_x_18_n361,
         mult_x_18_n360, mult_x_18_n359, mult_x_18_n358, mult_x_18_n357,
         mult_x_18_n356, mult_x_18_n355, mult_x_18_n354, mult_x_18_n353,
         mult_x_18_n352, mult_x_18_n350, mult_x_18_n349, mult_x_18_n348,
         mult_x_18_n347, mult_x_18_n346, mult_x_18_n345, mult_x_18_n344,
         mult_x_18_n343, mult_x_18_n342, mult_x_18_n339, mult_x_18_n337,
         mult_x_18_n336, mult_x_18_n335, mult_x_18_n334, mult_x_18_n333,
         mult_x_18_n332, mult_x_18_n331, mult_x_18_n330, mult_x_18_n329,
         mult_x_18_n326, mult_x_18_n324, mult_x_18_n323, mult_x_18_n322,
         mult_x_18_n321, mult_x_18_n320, mult_x_18_n319, mult_x_18_n318,
         mult_x_18_n317, mult_x_18_n316, mult_x_18_n314, mult_x_18_n313,
         mult_x_18_n312, mult_x_18_n311, mult_x_18_n310, mult_x_18_n309,
         mult_x_18_n308, mult_x_18_n307, mult_x_18_n306, mult_x_18_n305,
         mult_x_18_n304, mult_x_18_n303, mult_x_18_n302, mult_x_18_n300,
         mult_x_18_n299, mult_x_18_n298, mult_x_18_n297, mult_x_18_n296,
         mult_x_18_n295, mult_x_18_n294, mult_x_18_n293, mult_x_18_n292,
         mult_x_18_n291, mult_x_18_n290, mult_x_18_n289, mult_x_18_n288,
         mult_x_18_n286, mult_x_18_n285, mult_x_18_n284, mult_x_18_n283,
         mult_x_18_n282, mult_x_18_n281, mult_x_18_n280, mult_x_18_n279,
         mult_x_18_n278, mult_x_18_n277, mult_x_18_n276, mult_x_18_n275,
         mult_x_18_n274, mult_x_18_n272, mult_x_18_n271, mult_x_18_n270,
         mult_x_18_n269, mult_x_18_n268, mult_x_18_n267, mult_x_18_n266,
         mult_x_18_n265, mult_x_18_n264, mult_x_18_n263, mult_x_18_n262,
         mult_x_18_n261, mult_x_18_n258, mult_x_18_n256, mult_x_18_n255,
         mult_x_18_n254, mult_x_18_n253, mult_x_18_n252, mult_x_18_n251,
         mult_x_18_n250, mult_x_18_n249, mult_x_18_n248, mult_x_18_n247,
         mult_x_18_n246, mult_x_18_n245, mult_x_18_n242, mult_x_18_n240,
         mult_x_18_n239, mult_x_18_n238, mult_x_18_n237, mult_x_18_n236,
         mult_x_18_n235, mult_x_18_n234, mult_x_18_n233, mult_x_18_n232,
         mult_x_18_n231, mult_x_18_n230, mult_x_18_n229, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008;

  CMPE42D1BWP12T mult_x_18_U294 ( .A(mult_x_18_n699), .B(mult_x_18_n464), .C(
        mult_x_18_n467), .CIX(mult_x_18_n465), .D(mult_x_18_n726), .CO(
        mult_x_18_n461), .COX(mult_x_18_n460), .S(mult_x_18_n462) );
  CMPE42D1BWP12T mult_x_18_U292 ( .A(mult_x_18_n459), .B(mult_x_18_n698), .C(
        mult_x_18_n460), .CIX(mult_x_18_n461), .D(mult_x_18_n725), .CO(
        mult_x_18_n456), .COX(mult_x_18_n455), .S(mult_x_18_n457) );
  CMPE42D1BWP12T mult_x_18_U290 ( .A(mult_x_18_n697), .B(mult_x_18_n454), .C(
        mult_x_18_n455), .CIX(mult_x_18_n456), .D(mult_x_18_n724), .CO(
        mult_x_18_n451), .COX(mult_x_18_n450), .S(mult_x_18_n452) );
  CMPE42D1BWP12T mult_x_18_U287 ( .A(mult_x_18_n696), .B(mult_x_18_n447), .C(
        mult_x_18_n450), .CIX(mult_x_18_n451), .D(mult_x_18_n723), .CO(
        mult_x_18_n444), .COX(mult_x_18_n443), .S(mult_x_18_n445) );
  CMPE42D1BWP12T mult_x_18_U284 ( .A(mult_x_18_n695), .B(mult_x_18_n440), .C(
        mult_x_18_n443), .CIX(mult_x_18_n444), .D(mult_x_18_n722), .CO(
        mult_x_18_n437), .COX(mult_x_18_n436), .S(mult_x_18_n438) );
  CMPE42D1BWP12T mult_x_18_U281 ( .A(mult_x_18_n694), .B(mult_x_18_n433), .C(
        mult_x_18_n436), .CIX(mult_x_18_n437), .D(mult_x_18_n721), .CO(
        mult_x_18_n430), .COX(mult_x_18_n429), .S(mult_x_18_n431) );
  CMPE42D1BWP12T mult_x_18_U279 ( .A(mult_x_18_n648), .B(mult_x_18_n428), .C(
        mult_x_18_n434), .CIX(mult_x_18_n432), .D(mult_x_18_n669), .CO(
        mult_x_18_n425), .COX(mult_x_18_n424), .S(mult_x_18_n426) );
  CMPE42D1BWP12T mult_x_18_U278 ( .A(mult_x_18_n693), .B(mult_x_18_n426), .C(
        mult_x_18_n429), .CIX(mult_x_18_n430), .D(mult_x_18_n720), .CO(
        mult_x_18_n422), .COX(mult_x_18_n421), .S(mult_x_18_n423) );
  CMPE42D1BWP12T mult_x_18_U276 ( .A(mult_x_18_n420), .B(mult_x_18_n647), .C(
        mult_x_18_n424), .CIX(mult_x_18_n425), .D(mult_x_18_n668), .CO(
        mult_x_18_n417), .COX(mult_x_18_n416), .S(mult_x_18_n418) );
  CMPE42D1BWP12T mult_x_18_U275 ( .A(mult_x_18_n692), .B(mult_x_18_n418), .C(
        mult_x_18_n421), .CIX(mult_x_18_n422), .D(mult_x_18_n719), .CO(
        mult_x_18_n414), .COX(mult_x_18_n413), .S(mult_x_18_n415) );
  CMPE42D1BWP12T mult_x_18_U273 ( .A(mult_x_18_n646), .B(mult_x_18_n412), .C(
        mult_x_18_n416), .CIX(mult_x_18_n417), .D(mult_x_18_n667), .CO(
        mult_x_18_n409), .COX(mult_x_18_n408), .S(mult_x_18_n410) );
  CMPE42D1BWP12T mult_x_18_U272 ( .A(mult_x_18_n691), .B(mult_x_18_n410), .C(
        mult_x_18_n413), .CIX(mult_x_18_n414), .D(mult_x_18_n718), .CO(
        mult_x_18_n406), .COX(mult_x_18_n405), .S(mult_x_18_n407) );
  CMPE42D1BWP12T mult_x_18_U269 ( .A(mult_x_18_n645), .B(mult_x_18_n402), .C(
        mult_x_18_n408), .CIX(mult_x_18_n409), .D(mult_x_18_n666), .CO(
        mult_x_18_n399), .COX(mult_x_18_n398), .S(mult_x_18_n400) );
  CMPE42D1BWP12T mult_x_18_U268 ( .A(mult_x_18_n690), .B(mult_x_18_n400), .C(
        mult_x_18_n405), .CIX(mult_x_18_n406), .D(mult_x_18_n717), .CO(
        mult_x_18_n396), .COX(mult_x_18_n395), .S(mult_x_18_n397) );
  CMPE42D1BWP12T mult_x_18_U265 ( .A(mult_x_18_n644), .B(mult_x_18_n392), .C(
        mult_x_18_n398), .CIX(mult_x_18_n399), .D(mult_x_18_n665), .CO(
        mult_x_18_n389), .COX(mult_x_18_n388), .S(mult_x_18_n390) );
  CMPE42D1BWP12T mult_x_18_U264 ( .A(mult_x_18_n689), .B(mult_x_18_n390), .C(
        mult_x_18_n395), .CIX(mult_x_18_n396), .D(mult_x_18_n716), .CO(
        mult_x_18_n386), .COX(mult_x_18_n385), .S(mult_x_18_n387) );
  CMPE42D1BWP12T mult_x_18_U261 ( .A(mult_x_18_n643), .B(mult_x_18_n382), .C(
        mult_x_18_n388), .CIX(mult_x_18_n389), .D(mult_x_18_n664), .CO(
        mult_x_18_n379), .COX(mult_x_18_n378), .S(mult_x_18_n380) );
  CMPE42D1BWP12T mult_x_18_U260 ( .A(mult_x_18_n688), .B(mult_x_18_n380), .C(
        mult_x_18_n385), .CIX(mult_x_18_n386), .D(mult_x_18_n715), .CO(
        mult_x_18_n376), .COX(mult_x_18_n375), .S(mult_x_18_n377) );
  CMPE42D1BWP12T mult_x_18_U258 ( .A(mult_x_18_n609), .B(mult_x_18_n374), .C(
        mult_x_18_n383), .CIX(mult_x_18_n381), .D(mult_x_18_n624), .CO(
        mult_x_18_n371), .COX(mult_x_18_n370), .S(mult_x_18_n372) );
  CMPE42D1BWP12T mult_x_18_U257 ( .A(mult_x_18_n642), .B(mult_x_18_n372), .C(
        mult_x_18_n378), .CIX(mult_x_18_n379), .D(mult_x_18_n663), .CO(
        mult_x_18_n368), .COX(mult_x_18_n367), .S(mult_x_18_n369) );
  CMPE42D1BWP12T mult_x_18_U256 ( .A(mult_x_18_n687), .B(mult_x_18_n369), .C(
        mult_x_18_n375), .CIX(mult_x_18_n376), .D(mult_x_18_n714), .CO(
        mult_x_18_n365), .COX(mult_x_18_n364), .S(mult_x_18_n366) );
  CMPE42D1BWP12T mult_x_18_U254 ( .A(mult_x_18_n363), .B(mult_x_18_n608), .C(
        mult_x_18_n370), .CIX(mult_x_18_n371), .D(mult_x_18_n623), .CO(
        mult_x_18_n360), .COX(mult_x_18_n359), .S(mult_x_18_n361) );
  CMPE42D1BWP12T mult_x_18_U253 ( .A(mult_x_18_n641), .B(mult_x_18_n361), .C(
        mult_x_18_n367), .CIX(mult_x_18_n368), .D(mult_x_18_n662), .CO(
        mult_x_18_n357), .COX(mult_x_18_n356), .S(mult_x_18_n358) );
  CMPE42D1BWP12T mult_x_18_U252 ( .A(mult_x_18_n686), .B(mult_x_18_n358), .C(
        mult_x_18_n364), .CIX(mult_x_18_n365), .D(mult_x_18_n713), .CO(
        mult_x_18_n354), .COX(mult_x_18_n353), .S(mult_x_18_n355) );
  CMPE42D1BWP12T mult_x_18_U250 ( .A(mult_x_18_n607), .B(mult_x_18_n352), .C(
        mult_x_18_n359), .CIX(mult_x_18_n360), .D(mult_x_18_n622), .CO(
        mult_x_18_n349), .COX(mult_x_18_n348), .S(mult_x_18_n350) );
  CMPE42D1BWP12T mult_x_18_U249 ( .A(mult_x_18_n640), .B(mult_x_18_n350), .C(
        mult_x_18_n356), .CIX(mult_x_18_n357), .D(mult_x_18_n661), .CO(
        mult_x_18_n346), .COX(mult_x_18_n345), .S(mult_x_18_n347) );
  CMPE42D1BWP12T mult_x_18_U248 ( .A(mult_x_18_n685), .B(mult_x_18_n347), .C(
        mult_x_18_n353), .CIX(mult_x_18_n354), .D(mult_x_18_n712), .CO(
        mult_x_18_n343), .COX(mult_x_18_n342), .S(mult_x_18_n344) );
  CMPE42D1BWP12T mult_x_18_U245 ( .A(mult_x_18_n606), .B(mult_x_18_n339), .C(
        mult_x_18_n348), .CIX(mult_x_18_n349), .D(mult_x_18_n621), .CO(
        mult_x_18_n336), .COX(mult_x_18_n335), .S(mult_x_18_n337) );
  CMPE42D1BWP12T mult_x_18_U244 ( .A(mult_x_18_n639), .B(mult_x_18_n337), .C(
        mult_x_18_n345), .CIX(mult_x_18_n346), .D(mult_x_18_n660), .CO(
        mult_x_18_n333), .COX(mult_x_18_n332), .S(mult_x_18_n334) );
  CMPE42D1BWP12T mult_x_18_U243 ( .A(mult_x_18_n684), .B(mult_x_18_n334), .C(
        mult_x_18_n342), .CIX(mult_x_18_n343), .D(mult_x_18_n711), .CO(
        mult_x_18_n330), .COX(mult_x_18_n329), .S(mult_x_18_n331) );
  CMPE42D1BWP12T mult_x_18_U240 ( .A(mult_x_18_n605), .B(mult_x_18_n326), .C(
        mult_x_18_n335), .CIX(mult_x_18_n336), .D(mult_x_18_n620), .CO(
        mult_x_18_n323), .COX(mult_x_18_n322), .S(mult_x_18_n324) );
  CMPE42D1BWP12T mult_x_18_U239 ( .A(mult_x_18_n638), .B(mult_x_18_n324), .C(
        mult_x_18_n332), .CIX(mult_x_18_n333), .D(mult_x_18_n659), .CO(
        mult_x_18_n320), .COX(mult_x_18_n319), .S(mult_x_18_n321) );
  CMPE42D1BWP12T mult_x_18_U238 ( .A(mult_x_18_n683), .B(mult_x_18_n321), .C(
        mult_x_18_n329), .CIX(mult_x_18_n330), .D(mult_x_18_n710), .CO(
        mult_x_18_n317), .COX(mult_x_18_n316), .S(mult_x_18_n318) );
  CMPE42D1BWP12T mult_x_18_U235 ( .A(mult_x_18_n604), .B(mult_x_18_n313), .C(
        mult_x_18_n322), .CIX(mult_x_18_n323), .D(mult_x_18_n619), .CO(
        mult_x_18_n310), .COX(mult_x_18_n309), .S(mult_x_18_n311) );
  CMPE42D1BWP12T mult_x_18_U234 ( .A(mult_x_18_n637), .B(mult_x_18_n311), .C(
        mult_x_18_n319), .CIX(mult_x_18_n320), .D(mult_x_18_n658), .CO(
        mult_x_18_n307), .COX(mult_x_18_n306), .S(mult_x_18_n308) );
  CMPE42D1BWP12T mult_x_18_U233 ( .A(mult_x_18_n682), .B(mult_x_18_n308), .C(
        mult_x_18_n316), .CIX(mult_x_18_n317), .D(mult_x_18_n709), .CO(
        mult_x_18_n304), .COX(mult_x_18_n303), .S(mult_x_18_n305) );
  CMPE42D1BWP12T mult_x_18_U231 ( .A(mult_x_18_n582), .B(mult_x_18_n302), .C(
        mult_x_18_n314), .CIX(mult_x_18_n312), .D(mult_x_18_n591), .CO(
        mult_x_18_n299), .COX(mult_x_18_n298), .S(mult_x_18_n300) );
  CMPE42D1BWP12T mult_x_18_U230 ( .A(mult_x_18_n603), .B(mult_x_18_n300), .C(
        mult_x_18_n309), .CIX(mult_x_18_n310), .D(mult_x_18_n618), .CO(
        mult_x_18_n296), .COX(mult_x_18_n295), .S(mult_x_18_n297) );
  CMPE42D1BWP12T mult_x_18_U229 ( .A(mult_x_18_n636), .B(mult_x_18_n297), .C(
        mult_x_18_n306), .CIX(mult_x_18_n307), .D(mult_x_18_n657), .CO(
        mult_x_18_n293), .COX(mult_x_18_n292), .S(mult_x_18_n294) );
  CMPE42D1BWP12T mult_x_18_U228 ( .A(mult_x_18_n294), .B(mult_x_18_n681), .C(
        mult_x_18_n303), .CIX(mult_x_18_n304), .D(mult_x_18_n708), .CO(
        mult_x_18_n290), .COX(mult_x_18_n289), .S(mult_x_18_n291) );
  CMPE42D1BWP12T mult_x_18_U226 ( .A(mult_x_18_n288), .B(mult_x_18_n581), .C(
        mult_x_18_n298), .CIX(mult_x_18_n299), .D(mult_x_18_n590), .CO(
        mult_x_18_n285), .COX(mult_x_18_n284), .S(mult_x_18_n286) );
  CMPE42D1BWP12T mult_x_18_U225 ( .A(mult_x_18_n602), .B(mult_x_18_n286), .C(
        mult_x_18_n295), .CIX(mult_x_18_n296), .D(mult_x_18_n617), .CO(
        mult_x_18_n282), .COX(mult_x_18_n281), .S(mult_x_18_n283) );
  CMPE42D1BWP12T mult_x_18_U224 ( .A(mult_x_18_n635), .B(mult_x_18_n283), .C(
        mult_x_18_n292), .CIX(mult_x_18_n293), .D(mult_x_18_n656), .CO(
        mult_x_18_n279), .COX(mult_x_18_n278), .S(mult_x_18_n280) );
  CMPE42D1BWP12T mult_x_18_U223 ( .A(mult_x_18_n280), .B(mult_x_18_n680), .C(
        mult_x_18_n289), .CIX(mult_x_18_n290), .D(mult_x_18_n707), .CO(
        mult_x_18_n276), .COX(mult_x_18_n275), .S(mult_x_18_n277) );
  CMPE42D1BWP12T mult_x_18_U221 ( .A(mult_x_18_n580), .B(mult_x_18_n274), .C(
        mult_x_18_n284), .CIX(mult_x_18_n285), .D(mult_x_18_n589), .CO(
        mult_x_18_n271), .COX(mult_x_18_n270), .S(mult_x_18_n272) );
  CMPE42D1BWP12T mult_x_18_U220 ( .A(mult_x_18_n601), .B(mult_x_18_n272), .C(
        mult_x_18_n281), .CIX(mult_x_18_n282), .D(mult_x_18_n616), .CO(
        mult_x_18_n268), .COX(mult_x_18_n267), .S(mult_x_18_n269) );
  CMPE42D1BWP12T mult_x_18_U219 ( .A(mult_x_18_n634), .B(mult_x_18_n269), .C(
        mult_x_18_n278), .CIX(mult_x_18_n279), .D(mult_x_18_n655), .CO(
        mult_x_18_n265), .COX(mult_x_18_n264), .S(mult_x_18_n266) );
  CMPE42D1BWP12T mult_x_18_U218 ( .A(mult_x_18_n266), .B(mult_x_18_n679), .C(
        mult_x_18_n275), .CIX(mult_x_18_n276), .D(mult_x_18_n706), .CO(
        mult_x_18_n262), .COX(mult_x_18_n261), .S(mult_x_18_n263) );
  CMPE42D1BWP12T mult_x_18_U215 ( .A(mult_x_18_n579), .B(mult_x_18_n258), .C(
        mult_x_18_n270), .CIX(mult_x_18_n271), .D(mult_x_18_n588), .CO(
        mult_x_18_n255), .COX(mult_x_18_n254), .S(mult_x_18_n256) );
  CMPE42D1BWP12T mult_x_18_U214 ( .A(mult_x_18_n600), .B(mult_x_18_n256), .C(
        mult_x_18_n267), .CIX(mult_x_18_n268), .D(mult_x_18_n615), .CO(
        mult_x_18_n252), .COX(mult_x_18_n251), .S(mult_x_18_n253) );
  CMPE42D1BWP12T mult_x_18_U213 ( .A(mult_x_18_n633), .B(mult_x_18_n253), .C(
        mult_x_18_n264), .CIX(mult_x_18_n265), .D(mult_x_18_n654), .CO(
        mult_x_18_n249), .COX(mult_x_18_n248), .S(mult_x_18_n250) );
  CMPE42D1BWP12T mult_x_18_U212 ( .A(mult_x_18_n250), .B(mult_x_18_n678), .C(
        mult_x_18_n261), .CIX(mult_x_18_n262), .D(mult_x_18_n705), .CO(
        mult_x_18_n246), .COX(mult_x_18_n245), .S(mult_x_18_n247) );
  CMPE42D1BWP12T mult_x_18_U209 ( .A(mult_x_18_n578), .B(mult_x_18_n242), .C(
        mult_x_18_n254), .CIX(mult_x_18_n255), .D(mult_x_18_n587), .CO(
        mult_x_18_n239), .COX(mult_x_18_n238), .S(mult_x_18_n240) );
  CMPE42D1BWP12T mult_x_18_U208 ( .A(mult_x_18_n599), .B(mult_x_18_n240), .C(
        mult_x_18_n251), .CIX(mult_x_18_n252), .D(mult_x_18_n614), .CO(
        mult_x_18_n236), .COX(mult_x_18_n235), .S(mult_x_18_n237) );
  CMPE42D1BWP12T mult_x_18_U207 ( .A(mult_x_18_n632), .B(mult_x_18_n237), .C(
        mult_x_18_n248), .CIX(mult_x_18_n249), .D(mult_x_18_n653), .CO(
        mult_x_18_n233), .COX(mult_x_18_n232), .S(mult_x_18_n234) );
  CMPE42D1BWP12T mult_x_18_U206 ( .A(mult_x_18_n234), .B(mult_x_18_n677), .C(
        mult_x_18_n245), .CIX(mult_x_18_n246), .D(mult_x_18_n704), .CO(
        mult_x_18_n230), .COX(mult_x_18_n229), .S(mult_x_18_n231) );
  CKND0BWP12T U1364 ( .I(n3219), .ZN(n1326) );
  AOI22D0BWP12T U1365 ( .A1(n2692), .A2(n3784), .B1(n2708), .B2(n1326), .ZN(
        n1327) );
  OAI211D0BWP12T U1366 ( .A1(n2886), .A2(n2691), .B(n3144), .C(n1327), .ZN(
        n3609) );
  MAOI22D0BWP12T U1367 ( .A1(n3165), .A2(n2594), .B1(n2593), .B2(n3155), .ZN(
        n2622) );
  AOI22D0BWP12T U1368 ( .A1(n2774), .A2(a[21]), .B1(a[24]), .B2(n3725), .ZN(
        n1328) );
  NR3D0BWP12T U1369 ( .A1(n2752), .A2(n3522), .A3(n3494), .ZN(n1329) );
  OAI22D0BWP12T U1370 ( .A1(a[19]), .A2(n3598), .B1(a[25]), .B2(n3757), .ZN(
        n1330) );
  NR2D0BWP12T U1371 ( .A1(a[30]), .A2(n3912), .ZN(n1331) );
  INR4D0BWP12T U1372 ( .A1(n2769), .B1(n2768), .B2(n3271), .B3(n2767), .ZN(
        n1332) );
  NR4D0BWP12T U1373 ( .A1(n2764), .A2(n2766), .A3(n2765), .A4(n2763), .ZN(
        n1333) );
  NR4D0BWP12T U1374 ( .A1(n3444), .A2(n2762), .A3(n2761), .A4(n2760), .ZN(
        n1334) );
  NR4D0BWP12T U1375 ( .A1(n3296), .A2(n3328), .A3(n2757), .A4(n2758), .ZN(
        n1335) );
  ND4D0BWP12T U1376 ( .A1(n1332), .A2(n1333), .A3(n1334), .A4(n1335), .ZN(
        n1336) );
  ND4D0BWP12T U1377 ( .A1(n3027), .A2(n3823), .A3(n2756), .A4(n2755), .ZN(
        n1337) );
  OR4D0BWP12T U1378 ( .A1(n2770), .A2(n1331), .A3(n1336), .A4(n1337), .Z(n1338) );
  NR4D0BWP12T U1379 ( .A1(n3678), .A2(n2753), .A3(n1330), .A4(n1338), .ZN(
        n1339) );
  OAI211D0BWP12T U1380 ( .A1(a[18]), .A2(n2751), .B(n1329), .C(n1339), .ZN(
        n1340) );
  OAI32D0BWP12T U1381 ( .A1(n3758), .A2(n2773), .A3(n3650), .B1(n1340), .B2(
        n3758), .ZN(n1341) );
  ND4D0BWP12T U1382 ( .A1(n2775), .A2(n2776), .A3(n1328), .A4(n1341), .ZN(
        n1342) );
  IAO21D0BWP12T U1383 ( .A1(b[30]), .A2(n3932), .B(n1342), .ZN(n2924) );
  ND4D0BWP12T U1384 ( .A1(a[23]), .A2(a[9]), .A3(a[30]), .A4(a[0]), .ZN(n1343)
         );
  ND4D0BWP12T U1385 ( .A1(a[25]), .A2(a[24]), .A3(a[27]), .A4(a[28]), .ZN(
        n1344) );
  NR3D0BWP12T U1386 ( .A1(n3995), .A2(n1343), .A3(n1344), .ZN(n2928) );
  NR2D0BWP12T U1387 ( .A1(n3814), .A2(n2531), .ZN(n1345) );
  OAI22D0BWP12T U1388 ( .A1(b[4]), .A2(n3702), .B1(n3603), .B2(n2532), .ZN(
        n1346) );
  AOI211D0BWP12T U1389 ( .A1(n2575), .A2(n2533), .B(n1345), .C(n1346), .ZN(
        n3703) );
  INR2D0BWP12T U1390 ( .A1(n3268), .B1(n3269), .ZN(n3996) );
  ND4D0BWP12T U1391 ( .A1(n3653), .A2(n3732), .A3(n3825), .A4(n2443), .ZN(
        n1347) );
  CKND2D0BWP12T U1392 ( .A1(n3581), .A2(n3791), .ZN(n1348) );
  NR3D0BWP12T U1393 ( .A1(n1348), .A2(n1347), .A3(n2567), .ZN(n1349) );
  ND4D0BWP12T U1394 ( .A1(n3702), .A2(n3558), .A3(n2577), .A4(n1349), .ZN(
        n1350) );
  AOI211D0BWP12T U1395 ( .A1(n3199), .A2(n1350), .B(n3308), .C(n3189), .ZN(
        n2462) );
  NR4D0BWP12T U1396 ( .A1(a[20]), .A2(a[26]), .A3(a[31]), .A4(a[29]), .ZN(
        n1351) );
  ND3D0BWP12T U1397 ( .A1(n2719), .A2(n2720), .A3(n1351), .ZN(n1352) );
  ND4D0BWP12T U1398 ( .A1(n3479), .A2(n3701), .A3(n3428), .A4(n3193), .ZN(
        n1353) );
  NR4D0BWP12T U1399 ( .A1(n2721), .A2(n2722), .A3(n1352), .A4(n1353), .ZN(
        n1354) );
  NR4D0BWP12T U1400 ( .A1(n2717), .A2(n2718), .A3(n2716), .A4(n2715), .ZN(
        n1355) );
  ND4D0BWP12T U1401 ( .A1(n3940), .A2(n2723), .A3(n1354), .A4(n1355), .ZN(
        n1356) );
  NR4D0BWP12T U1402 ( .A1(n3297), .A2(n3737), .A3(n2724), .A4(n1356), .ZN(
        n2734) );
  OAI22D0BWP12T U1403 ( .A1(n3976), .A2(n3977), .B1(n3975), .B2(n3974), .ZN(
        n1357) );
  AOI21D0BWP12T U1404 ( .A1(n3982), .A2(n3983), .B(n1357), .ZN(n1358) );
  AOI22D0BWP12T U1405 ( .A1(n3987), .A2(n3986), .B1(n3984), .B2(n3985), .ZN(
        n1359) );
  OAI21D0BWP12T U1406 ( .A1(b[3]), .A2(n3989), .B(n3988), .ZN(n1360) );
  AOI211D0BWP12T U1407 ( .A1(n3992), .A2(a[3]), .B(n3990), .C(n3991), .ZN(
        n1361) );
  OAI22D0BWP12T U1408 ( .A1(a[3]), .A2(n3995), .B1(n3994), .B2(n3993), .ZN(
        n1362) );
  AOI211D0BWP12T U1409 ( .A1(a[3]), .A2(n1360), .B(n1361), .C(n1362), .ZN(
        n1363) );
  AOI22D0BWP12T U1410 ( .A1(n3997), .A2(n3996), .B1(n3999), .B2(n3998), .ZN(
        n1364) );
  OAI211D0BWP12T U1411 ( .A1(n4001), .A2(n4000), .B(n1363), .C(n1364), .ZN(
        n1365) );
  AOI211D0BWP12T U1412 ( .A1(n4003), .A2(n4004), .B(n4002), .C(n1365), .ZN(
        n1366) );
  AOI32D0BWP12T U1413 ( .A1(n3980), .A2(n3981), .A3(n3979), .B1(n3978), .B2(
        n3981), .ZN(n1367) );
  ND4D0BWP12T U1414 ( .A1(n1358), .A2(n1359), .A3(n1366), .A4(n1367), .ZN(
        result[3]) );
  OAI31D0BWP12T U1415 ( .A1(n3165), .A2(n2847), .A3(n2429), .B(n3219), .ZN(
        n1368) );
  OAI22D0BWP12T U1416 ( .A1(n2886), .A2(n2568), .B1(n2399), .B2(n2455), .ZN(
        n1369) );
  AO211D0BWP12T U1417 ( .A1(n2906), .A2(n2448), .B(n1368), .C(n1369), .Z(n1370) );
  OAI21D0BWP12T U1418 ( .A1(n3219), .A2(n2440), .B(n1370), .ZN(n2500) );
  AOI22D0BWP12T U1419 ( .A1(b[6]), .A2(n2074), .B1(b[5]), .B2(n2112), .ZN(
        n1371) );
  AOI22D0BWP12T U1420 ( .A1(b[7]), .A2(n2086), .B1(n2085), .B2(n2021), .ZN(
        n1372) );
  CKND2D0BWP12T U1421 ( .A1(n1371), .A2(n1372), .ZN(n1373) );
  MOAI22D0BWP12T U1422 ( .A1(a[2]), .A2(n1373), .B1(a[2]), .B2(n1373), .ZN(
        n1374) );
  MAOI22D0BWP12T U1423 ( .A1(n1374), .A2(n2830), .B1(n1374), .B2(n2830), .ZN(
        n1375) );
  MAOI22D0BWP12T U1424 ( .A1(n2052), .A2(n1375), .B1(n2052), .B2(n1375), .ZN(
        n3289) );
  CKND0BWP12T U1425 ( .I(n2830), .ZN(n1376) );
  MAOI222D0BWP12T U1426 ( .A(n1374), .B(n2052), .C(n1376), .ZN(n2829) );
  OAI22D0BWP12T U1427 ( .A1(n3836), .A2(n3816), .B1(n3818), .B2(n3817), .ZN(
        n1377) );
  MOAI22D0BWP12T U1428 ( .A1(n3814), .A2(n3815), .B1(n3980), .B2(n3813), .ZN(
        n1378) );
  NR4D0BWP12T U1429 ( .A1(n3891), .A2(n3812), .A3(n1377), .A4(n1378), .ZN(
        n1379) );
  NR2D0BWP12T U1430 ( .A1(n3920), .A2(n3819), .ZN(n1380) );
  AOI211D0BWP12T U1431 ( .A1(n3828), .A2(n3999), .B(n1379), .C(n1380), .ZN(
        n1381) );
  AOI211D0BWP12T U1432 ( .A1(n3811), .A2(a[27]), .B(n3990), .C(n3852), .ZN(
        n1382) );
  OAI21D0BWP12T U1433 ( .A1(n3899), .A2(n3820), .B(n3996), .ZN(n1383) );
  OAI211D0BWP12T U1434 ( .A1(a[27]), .A2(op[2]), .B(b[27]), .C(n3833), .ZN(
        n1384) );
  OAI211D0BWP12T U1435 ( .A1(n3989), .A2(n3821), .B(n1383), .C(n1384), .ZN(
        n1385) );
  AOI22D0BWP12T U1436 ( .A1(a[27]), .A2(n3940), .B1(n4003), .B2(n3822), .ZN(
        n1386) );
  AOI32D0BWP12T U1437 ( .A1(b[27]), .A2(n3824), .A3(n3823), .B1(n3959), .B2(
        n3824), .ZN(n1387) );
  OAI211D0BWP12T U1438 ( .A1(n3922), .A2(n3825), .B(n1386), .C(n1387), .ZN(
        n1388) );
  OAI22D0BWP12T U1439 ( .A1(n3956), .A2(n3826), .B1(n3975), .B2(n3827), .ZN(
        n1389) );
  NR4D0BWP12T U1440 ( .A1(n1382), .A2(n1385), .A3(n1388), .A4(n1389), .ZN(
        n1390) );
  OAI211D0BWP12T U1441 ( .A1(n3976), .A2(n3829), .B(n1381), .C(n1390), .ZN(
        result[27]) );
  MOAI22D0BWP12T U1442 ( .A1(n1832), .A2(n1831), .B1(n1832), .B2(n1831), .ZN(
        n1912) );
  IOA21D0BWP12T U1443 ( .A1(n2123), .A2(n2124), .B(a[31]), .ZN(n2125) );
  ND4D0BWP12T U1444 ( .A1(a[12]), .A2(a[13]), .A3(a[1]), .A4(a[2]), .ZN(n1391)
         );
  ND4D0BWP12T U1445 ( .A1(a[15]), .A2(a[16]), .A3(a[11]), .A4(a[10]), .ZN(
        n1392) );
  NR2D0BWP12T U1446 ( .A1(n1391), .A2(n1392), .ZN(n2929) );
  ND4D0BWP12T U1447 ( .A1(a[26]), .A2(a[29]), .A3(a[14]), .A4(a[17]), .ZN(
        n1393) );
  ND4D0BWP12T U1448 ( .A1(a[3]), .A2(a[4]), .A3(a[19]), .A4(a[18]), .ZN(n1394)
         );
  NR2D0BWP12T U1449 ( .A1(n1393), .A2(n1394), .ZN(n2930) );
  ND4D0BWP12T U1450 ( .A1(a[5]), .A2(a[8]), .A3(a[20]), .A4(a[31]), .ZN(n1395)
         );
  ND4D0BWP12T U1451 ( .A1(a[6]), .A2(a[7]), .A3(a[22]), .A4(a[21]), .ZN(n1396)
         );
  NR2D0BWP12T U1452 ( .A1(n1395), .A2(n1396), .ZN(n2931) );
  ND4D0BWP12T U1453 ( .A1(n3651), .A2(n3672), .A3(n3698), .A4(n3727), .ZN(
        n1397) );
  AOI22D0BWP12T U1454 ( .A1(b[27]), .A2(a[27]), .B1(b[28]), .B2(a[28]), .ZN(
        n1398) );
  ND3D0BWP12T U1455 ( .A1(n3574), .A2(n3608), .A3(n3556), .ZN(n1399) );
  ND4D0BWP12T U1456 ( .A1(n3531), .A2(n2725), .A3(n3918), .A4(n3866), .ZN(
        n1400) );
  AOI211D0BWP12T U1457 ( .A1(a[20]), .A2(b[20]), .B(n1399), .C(n1400), .ZN(
        n1401) );
  ND4D0BWP12T U1458 ( .A1(n3788), .A2(n3759), .A3(n1398), .A4(n1401), .ZN(
        n1402) );
  NR2D0BWP12T U1459 ( .A1(n1397), .A2(n1402), .ZN(n2733) );
  AOI22D0BWP12T U1460 ( .A1(b[7]), .A2(n2074), .B1(b[6]), .B2(n2112), .ZN(
        n1403) );
  AOI22D0BWP12T U1461 ( .A1(b[8]), .A2(n2086), .B1(n2085), .B2(n2163), .ZN(
        n1404) );
  CKND2D0BWP12T U1462 ( .A1(n1403), .A2(n1404), .ZN(n1405) );
  MOAI22D0BWP12T U1463 ( .A1(a[2]), .A2(n1405), .B1(a[2]), .B2(n1405), .ZN(
        n1406) );
  CKND0BWP12T U1464 ( .I(n2829), .ZN(n1407) );
  MAOI222D0BWP12T U1465 ( .A(n1406), .B(n2056), .C(n1407), .ZN(n2827) );
  MAOI22D0BWP12T U1466 ( .A1(n1406), .A2(n2829), .B1(n1406), .B2(n2829), .ZN(
        n1408) );
  MAOI22D0BWP12T U1467 ( .A1(n2056), .A2(n1408), .B1(n2056), .B2(n1408), .ZN(
        n3317) );
  IAO21D0BWP12T U1468 ( .A1(n3194), .A2(n2906), .B(n2907), .ZN(n3909) );
  INVD1BWP12T U1469 ( .I(a[4]), .ZN(n3218) );
  OAI22D1BWP12T U1470 ( .A1(n3247), .A2(n3218), .B1(a[4]), .B2(a[5]), .ZN(
        n1411) );
  INVD1BWP12T U1471 ( .I(a[3]), .ZN(n2471) );
  OAI22D1BWP12T U1472 ( .A1(n2471), .A2(a[2]), .B1(n3961), .B2(a[3]), .ZN(
        n1410) );
  ND2D1BWP12T U1473 ( .A1(n1411), .A2(n1410), .ZN(n1881) );
  INVD1BWP12T U1474 ( .I(n1881), .ZN(n2197) );
  INVD1BWP12T U1475 ( .I(n1410), .ZN(n2025) );
  OAI22D1BWP12T U1476 ( .A1(n3218), .A2(a[3]), .B1(n2471), .B2(a[4]), .ZN(
        n1409) );
  ND2D1BWP12T U1477 ( .A1(n2025), .A2(n1409), .ZN(n1882) );
  INVD1BWP12T U1478 ( .I(n1882), .ZN(n2196) );
  AOI22D1BWP12T U1479 ( .A1(b[28]), .A2(n2197), .B1(b[27]), .B2(n2196), .ZN(
        n1414) );
  NR3D1BWP12T U1480 ( .A1(n1410), .A2(n1409), .A3(n1411), .ZN(n2200) );
  NR2D1BWP12T U1481 ( .A1(n2025), .A2(n1411), .ZN(n2198) );
  INVD1BWP12T U1482 ( .I(n2198), .ZN(n1883) );
  INVD1BWP12T U1483 ( .I(b[4]), .ZN(n3219) );
  ND2D1BWP12T U1484 ( .A1(n3219), .A2(n2886), .ZN(n2914) );
  INVD1BWP12T U1485 ( .I(n2914), .ZN(n3784) );
  INVD1BWP12T U1486 ( .I(b[1]), .ZN(n3165) );
  INVD1BWP12T U1487 ( .I(b[0]), .ZN(n3170) );
  NR2D1BWP12T U1488 ( .A1(n3165), .A2(n3170), .ZN(n1622) );
  NR2D1BWP12T U1489 ( .A1(b[2]), .A2(n1622), .ZN(n1666) );
  INVD1BWP12T U1490 ( .I(n1666), .ZN(n2382) );
  INVD1BWP12T U1491 ( .I(b[2]), .ZN(n2652) );
  NR2D1BWP12T U1492 ( .A1(n2652), .A2(n3165), .ZN(n1665) );
  AOI21D1BWP12T U1493 ( .A1(b[3]), .A2(n2382), .B(n1665), .ZN(n1614) );
  INVD1BWP12T U1494 ( .I(b[3]), .ZN(n2886) );
  NR2D1BWP12T U1495 ( .A1(n3219), .A2(n2886), .ZN(n2625) );
  INVD1BWP12T U1496 ( .I(n2625), .ZN(n1412) );
  OAI21D1BWP12T U1497 ( .A1(n3784), .A2(n1614), .B(n1412), .ZN(n1686) );
  AOI22D1BWP12T U1498 ( .A1(b[26]), .A2(n2200), .B1(n2198), .B2(n2081), .ZN(
        n1413) );
  ND2D1BWP12T U1499 ( .A1(n1414), .A2(n1413), .ZN(n1415) );
  MAOI22D0BWP12T U1500 ( .A1(a[5]), .A2(n1415), .B1(a[5]), .B2(n1415), .ZN(
        mult_x_18_n704) );
  AOI22D1BWP12T U1501 ( .A1(b[24]), .A2(n2197), .B1(b[23]), .B2(n2196), .ZN(
        n1418) );
  FA1D0BWP12T U1502 ( .A(b[23]), .B(b[24]), .CI(n1416), .CO(n1521), .S(n2073)
         );
  AOI22D1BWP12T U1503 ( .A1(b[22]), .A2(n2200), .B1(n2198), .B2(n2073), .ZN(
        n1417) );
  ND2D1BWP12T U1504 ( .A1(n1418), .A2(n1417), .ZN(n1419) );
  MAOI22D0BWP12T U1505 ( .A1(a[5]), .A2(n1419), .B1(a[5]), .B2(n1419), .ZN(
        mult_x_18_n708) );
  INVD1BWP12T U1506 ( .I(a[11]), .ZN(n4005) );
  INVD1BWP12T U1507 ( .I(a[10]), .ZN(n3380) );
  OAI22D1BWP12T U1508 ( .A1(n4005), .A2(n3380), .B1(a[10]), .B2(a[11]), .ZN(
        n1421) );
  INVD1BWP12T U1509 ( .I(a[9]), .ZN(n3346) );
  INVD1BWP12T U1510 ( .I(a[8]), .ZN(n3321) );
  OAI22D1BWP12T U1511 ( .A1(n3346), .A2(n3321), .B1(a[8]), .B2(a[9]), .ZN(
        n1921) );
  INR2D1BWP12T U1512 ( .A1(n1421), .B1(n1921), .ZN(n2185) );
  AOI22D1BWP12T U1513 ( .A1(a[10]), .A2(n3346), .B1(a[9]), .B2(n3380), .ZN(
        n1420) );
  INR2D1BWP12T U1514 ( .A1(n1921), .B1(n1420), .ZN(n2186) );
  AOI22D1BWP12T U1515 ( .A1(b[22]), .A2(n2185), .B1(b[21]), .B2(n2186), .ZN(
        n1424) );
  ND2D1BWP12T U1516 ( .A1(n1921), .A2(n1420), .ZN(n2724) );
  NR2D1BWP12T U1517 ( .A1(n1421), .A2(n2724), .ZN(n2189) );
  NR2D1BWP12T U1518 ( .A1(n1921), .A2(n1421), .ZN(n2187) );
  FA1D0BWP12T U1519 ( .A(b[21]), .B(b[22]), .CI(n1422), .CO(n1538), .S(n1995)
         );
  AOI22D1BWP12T U1520 ( .A1(b[20]), .A2(n2189), .B1(n2187), .B2(n1995), .ZN(
        n1423) );
  ND2D1BWP12T U1521 ( .A1(n1424), .A2(n1423), .ZN(n1425) );
  MAOI22D0BWP12T U1522 ( .A1(a[11]), .A2(n1425), .B1(a[11]), .B2(n1425), .ZN(
        mult_x_18_n653) );
  AOI22D1BWP12T U1523 ( .A1(b[18]), .A2(n2185), .B1(b[17]), .B2(n2186), .ZN(
        n1428) );
  FA1D0BWP12T U1524 ( .A(b[17]), .B(b[18]), .CI(n1426), .CO(n1459), .S(n2008)
         );
  AOI22D1BWP12T U1525 ( .A1(b[16]), .A2(n2189), .B1(n2187), .B2(n2008), .ZN(
        n1427) );
  ND2D1BWP12T U1526 ( .A1(n1428), .A2(n1427), .ZN(n1429) );
  MAOI22D0BWP12T U1527 ( .A1(a[11]), .A2(n1429), .B1(a[11]), .B2(n1429), .ZN(
        mult_x_18_n657) );
  INVD1BWP12T U1528 ( .I(a[17]), .ZN(n3565) );
  INVD1BWP12T U1529 ( .I(a[16]), .ZN(n3529) );
  OAI22D1BWP12T U1530 ( .A1(n3565), .A2(n3529), .B1(a[16]), .B2(a[17]), .ZN(
        n1432) );
  INVD1BWP12T U1531 ( .I(a[15]), .ZN(n2485) );
  OAI22D1BWP12T U1532 ( .A1(n2485), .A2(a[14]), .B1(n3479), .B2(a[15]), .ZN(
        n1431) );
  ND2D1BWP12T U1533 ( .A1(n1432), .A2(n1431), .ZN(n1621) );
  INVD1BWP12T U1534 ( .I(n1621), .ZN(n2179) );
  INVD1BWP12T U1535 ( .I(n1431), .ZN(n1718) );
  OAI22D1BWP12T U1536 ( .A1(n3529), .A2(a[15]), .B1(n2485), .B2(a[16]), .ZN(
        n1430) );
  ND2D1BWP12T U1537 ( .A1(n1718), .A2(n1430), .ZN(n1620) );
  INVD1BWP12T U1538 ( .I(n1620), .ZN(n2178) );
  AOI22D1BWP12T U1539 ( .A1(b[16]), .A2(n2179), .B1(b[15]), .B2(n2178), .ZN(
        n1435) );
  NR3D1BWP12T U1540 ( .A1(n1431), .A2(n1430), .A3(n1432), .ZN(n2182) );
  NR2D1BWP12T U1541 ( .A1(n1718), .A2(n1432), .ZN(n2180) );
  FA1D0BWP12T U1542 ( .A(b[15]), .B(b[16]), .CI(n1433), .CO(n1475), .S(n2070)
         );
  AOI22D1BWP12T U1543 ( .A1(b[14]), .A2(n2182), .B1(n2180), .B2(n2070), .ZN(
        n1434) );
  ND2D1BWP12T U1544 ( .A1(n1435), .A2(n1434), .ZN(n1436) );
  MAOI22D0BWP12T U1545 ( .A1(a[17]), .A2(n1436), .B1(a[17]), .B2(n1436), .ZN(
        mult_x_18_n614) );
  AOI22D1BWP12T U1546 ( .A1(b[12]), .A2(n2179), .B1(b[11]), .B2(n2178), .ZN(
        n1439) );
  FA1D0BWP12T U1547 ( .A(b[11]), .B(b[12]), .CI(n1437), .CO(n1534), .S(n2059)
         );
  AOI22D1BWP12T U1548 ( .A1(b[10]), .A2(n2182), .B1(n2180), .B2(n2059), .ZN(
        n1438) );
  ND2D1BWP12T U1549 ( .A1(n1439), .A2(n1438), .ZN(n1440) );
  MAOI22D0BWP12T U1550 ( .A1(a[17]), .A2(n1440), .B1(a[17]), .B2(n1440), .ZN(
        mult_x_18_n618) );
  INVD1BWP12T U1551 ( .I(a[22]), .ZN(n3684) );
  INVD1BWP12T U1552 ( .I(a[23]), .ZN(n3701) );
  OAI22D1BWP12T U1553 ( .A1(n3684), .A2(n3701), .B1(a[23]), .B2(a[22]), .ZN(
        n1443) );
  INVD1BWP12T U1554 ( .I(a[21]), .ZN(n3685) );
  OAI22D1BWP12T U1555 ( .A1(n3685), .A2(a[20]), .B1(n3632), .B2(a[21]), .ZN(
        n1442) );
  ND2D1BWP12T U1556 ( .A1(n1443), .A2(n1442), .ZN(n1862) );
  INVD1BWP12T U1557 ( .I(n1862), .ZN(n2152) );
  INVD1BWP12T U1558 ( .I(n1442), .ZN(n1853) );
  OAI22D1BWP12T U1559 ( .A1(n3684), .A2(a[21]), .B1(n3685), .B2(a[22]), .ZN(
        n1441) );
  ND2D1BWP12T U1560 ( .A1(n1853), .A2(n1441), .ZN(n1863) );
  INVD1BWP12T U1561 ( .I(n1863), .ZN(n2151) );
  AOI22D1BWP12T U1562 ( .A1(b[10]), .A2(n2152), .B1(b[9]), .B2(n2151), .ZN(
        n1446) );
  NR3D1BWP12T U1563 ( .A1(n1442), .A2(n1441), .A3(n1443), .ZN(n2155) );
  NR2D1BWP12T U1564 ( .A1(n1443), .A2(n1853), .ZN(n2153) );
  FA1D0BWP12T U1565 ( .A(b[9]), .B(b[10]), .CI(n1444), .CO(n1517), .S(n2013)
         );
  AOI22D1BWP12T U1566 ( .A1(b[8]), .A2(n2155), .B1(n2153), .B2(n2013), .ZN(
        n1445) );
  ND2D1BWP12T U1567 ( .A1(n1446), .A2(n1445), .ZN(n1447) );
  MAOI22D0BWP12T U1568 ( .A1(a[23]), .A2(n1447), .B1(a[23]), .B2(n1447), .ZN(
        mult_x_18_n587) );
  AOI22D1BWP12T U1569 ( .A1(b[6]), .A2(n2152), .B1(b[5]), .B2(n2151), .ZN(
        n1450) );
  FA1D0BWP12T U1570 ( .A(b[5]), .B(b[6]), .CI(n1448), .CO(n1467), .S(n2043) );
  AOI22D1BWP12T U1571 ( .A1(b[4]), .A2(n2155), .B1(n2153), .B2(n2043), .ZN(
        n1449) );
  ND2D1BWP12T U1572 ( .A1(n1450), .A2(n1449), .ZN(n1451) );
  MAOI22D0BWP12T U1573 ( .A1(a[23]), .A2(n1451), .B1(a[23]), .B2(n1451), .ZN(
        mult_x_18_n591) );
  AOI22D1BWP12T U1574 ( .A1(b[6]), .A2(n2197), .B1(b[5]), .B2(n2196), .ZN(
        n1453) );
  CKBD1BWP12T U1575 ( .I(n2200), .Z(n1602) );
  AOI22D1BWP12T U1576 ( .A1(b[4]), .A2(n1602), .B1(n2198), .B2(n2043), .ZN(
        n1452) );
  ND2D1BWP12T U1577 ( .A1(n1453), .A2(n1452), .ZN(n1454) );
  MAOI22D0BWP12T U1578 ( .A1(a[5]), .A2(n1454), .B1(a[5]), .B2(n1454), .ZN(
        mult_x_18_n726) );
  AOI22D1BWP12T U1579 ( .A1(b[27]), .A2(n2197), .B1(b[26]), .B2(n2196), .ZN(
        n1457) );
  FA1D0BWP12T U1580 ( .A(b[26]), .B(b[27]), .CI(n1455), .CO(n1974), .S(n1985)
         );
  AOI22D1BWP12T U1581 ( .A1(b[25]), .A2(n2200), .B1(n2198), .B2(n1985), .ZN(
        n1456) );
  ND2D1BWP12T U1582 ( .A1(n1457), .A2(n1456), .ZN(n1458) );
  MAOI22D0BWP12T U1583 ( .A1(a[5]), .A2(n1458), .B1(a[5]), .B2(n1458), .ZN(
        mult_x_18_n705) );
  AOI22D1BWP12T U1584 ( .A1(b[19]), .A2(n2197), .B1(b[18]), .B2(n2196), .ZN(
        n1461) );
  FA1D0BWP12T U1585 ( .A(b[18]), .B(b[19]), .CI(n1459), .CO(n1497), .S(n2004)
         );
  AOI22D1BWP12T U1586 ( .A1(b[17]), .A2(n2200), .B1(n2198), .B2(n2004), .ZN(
        n1460) );
  ND2D1BWP12T U1587 ( .A1(n1461), .A2(n1460), .ZN(n1462) );
  MAOI22D0BWP12T U1588 ( .A1(a[5]), .A2(n1462), .B1(a[5]), .B2(n1462), .ZN(
        mult_x_18_n713) );
  AOI22D1BWP12T U1589 ( .A1(b[21]), .A2(n2185), .B1(b[20]), .B2(n2186), .ZN(
        n1465) );
  FA1D0BWP12T U1590 ( .A(b[20]), .B(b[21]), .CI(n1463), .CO(n1422), .S(n1998)
         );
  AOI22D1BWP12T U1591 ( .A1(b[19]), .A2(n2189), .B1(n2187), .B2(n1998), .ZN(
        n1464) );
  ND2D1BWP12T U1592 ( .A1(n1465), .A2(n1464), .ZN(n1466) );
  MAOI22D0BWP12T U1593 ( .A1(a[11]), .A2(n1466), .B1(a[11]), .B2(n1466), .ZN(
        mult_x_18_n654) );
  AOI22D1BWP12T U1594 ( .A1(b[7]), .A2(n2197), .B1(b[6]), .B2(n2196), .ZN(
        n1469) );
  FA1D0BWP12T U1595 ( .A(b[6]), .B(b[7]), .CI(n1467), .CO(n1483), .S(n2021) );
  AOI22D1BWP12T U1596 ( .A1(b[5]), .A2(n1602), .B1(n2198), .B2(n2021), .ZN(
        n1468) );
  ND2D1BWP12T U1597 ( .A1(n1469), .A2(n1468), .ZN(n1470) );
  MAOI22D0BWP12T U1598 ( .A1(a[5]), .A2(n1470), .B1(a[5]), .B2(n1470), .ZN(
        mult_x_18_n725) );
  AOI22D1BWP12T U1599 ( .A1(b[15]), .A2(n2179), .B1(b[14]), .B2(n2178), .ZN(
        n1473) );
  FA1D0BWP12T U1600 ( .A(b[14]), .B(b[15]), .CI(n1471), .CO(n1433), .S(n2067)
         );
  AOI22D1BWP12T U1601 ( .A1(b[13]), .A2(n2182), .B1(n2180), .B2(n2067), .ZN(
        n1472) );
  ND2D1BWP12T U1602 ( .A1(n1473), .A2(n1472), .ZN(n1474) );
  MAOI22D0BWP12T U1603 ( .A1(a[17]), .A2(n1474), .B1(a[17]), .B2(n1474), .ZN(
        mult_x_18_n615) );
  AOI22D1BWP12T U1604 ( .A1(b[17]), .A2(n2185), .B1(b[16]), .B2(n2186), .ZN(
        n1477) );
  FA1D0BWP12T U1605 ( .A(b[16]), .B(b[17]), .CI(n1475), .CO(n1426), .S(n2181)
         );
  AOI22D1BWP12T U1606 ( .A1(b[15]), .A2(n2189), .B1(n2181), .B2(n2187), .ZN(
        n1476) );
  ND2D1BWP12T U1607 ( .A1(n1477), .A2(n1476), .ZN(n1478) );
  MAOI22D0BWP12T U1608 ( .A1(a[11]), .A2(n1478), .B1(a[11]), .B2(n1478), .ZN(
        mult_x_18_n658) );
  AOI22D1BWP12T U1609 ( .A1(b[9]), .A2(n2152), .B1(b[8]), .B2(n2151), .ZN(
        n1481) );
  FA1D0BWP12T U1610 ( .A(b[8]), .B(b[9]), .CI(n1479), .CO(n1444), .S(n2017) );
  AOI22D1BWP12T U1611 ( .A1(b[7]), .A2(n2155), .B1(n2153), .B2(n2017), .ZN(
        n1480) );
  ND2D1BWP12T U1612 ( .A1(n1481), .A2(n1480), .ZN(n1482) );
  MAOI22D0BWP12T U1613 ( .A1(a[23]), .A2(n1482), .B1(a[23]), .B2(n1482), .ZN(
        mult_x_18_n588) );
  AOI22D1BWP12T U1614 ( .A1(b[8]), .A2(n2197), .B1(b[7]), .B2(n2196), .ZN(
        n1485) );
  FA1D0BWP12T U1615 ( .A(b[7]), .B(b[8]), .CI(n1483), .CO(n1479), .S(n2163) );
  AOI22D1BWP12T U1616 ( .A1(b[6]), .A2(n1602), .B1(n2163), .B2(n2198), .ZN(
        n1484) );
  ND2D1BWP12T U1617 ( .A1(n1485), .A2(n1484), .ZN(n1486) );
  MAOI22D0BWP12T U1618 ( .A1(a[5]), .A2(n1486), .B1(a[5]), .B2(n1486), .ZN(
        mult_x_18_n724) );
  AOI22D1BWP12T U1619 ( .A1(b[9]), .A2(n2185), .B1(b[8]), .B2(n2186), .ZN(
        n1488) );
  AOI22D1BWP12T U1620 ( .A1(b[7]), .A2(n2189), .B1(n2187), .B2(n2017), .ZN(
        n1487) );
  ND2D1BWP12T U1621 ( .A1(n1488), .A2(n1487), .ZN(n1489) );
  MAOI22D0BWP12T U1622 ( .A1(a[11]), .A2(n1489), .B1(a[11]), .B2(n1489), .ZN(
        mult_x_18_n666) );
  AOI22D1BWP12T U1623 ( .A1(b[26]), .A2(n2197), .B1(b[25]), .B2(n2196), .ZN(
        n1492) );
  FA1D0BWP12T U1624 ( .A(b[25]), .B(b[26]), .CI(n1490), .CO(n1455), .S(n2147)
         );
  AOI22D1BWP12T U1625 ( .A1(b[24]), .A2(n2200), .B1(n2147), .B2(n2198), .ZN(
        n1491) );
  ND2D1BWP12T U1626 ( .A1(n1492), .A2(n1491), .ZN(n1493) );
  MAOI22D0BWP12T U1627 ( .A1(a[5]), .A2(n1493), .B1(a[5]), .B2(n1493), .ZN(
        mult_x_18_n706) );
  AOI22D1BWP12T U1628 ( .A1(b[9]), .A2(n2197), .B1(b[8]), .B2(n2196), .ZN(
        n1495) );
  AOI22D1BWP12T U1629 ( .A1(b[7]), .A2(n1602), .B1(n2198), .B2(n2017), .ZN(
        n1494) );
  ND2D1BWP12T U1630 ( .A1(n1495), .A2(n1494), .ZN(n1496) );
  MAOI22D0BWP12T U1631 ( .A1(a[5]), .A2(n1496), .B1(a[5]), .B2(n1496), .ZN(
        mult_x_18_n723) );
  AOI22D1BWP12T U1632 ( .A1(b[20]), .A2(n2185), .B1(b[19]), .B2(n2186), .ZN(
        n1499) );
  FA1D0BWP12T U1633 ( .A(b[19]), .B(b[20]), .CI(n1497), .CO(n1463), .S(n2095)
         );
  AOI22D1BWP12T U1634 ( .A1(b[18]), .A2(n2189), .B1(n2095), .B2(n2187), .ZN(
        n1498) );
  ND2D1BWP12T U1635 ( .A1(n1499), .A2(n1498), .ZN(n1500) );
  MAOI22D0BWP12T U1636 ( .A1(a[11]), .A2(n1500), .B1(a[11]), .B2(n1500), .ZN(
        mult_x_18_n655) );
  AOI22D1BWP12T U1637 ( .A1(b[16]), .A2(n2185), .B1(b[15]), .B2(n2186), .ZN(
        n1502) );
  AOI22D1BWP12T U1638 ( .A1(b[14]), .A2(n2189), .B1(n2187), .B2(n2070), .ZN(
        n1501) );
  ND2D1BWP12T U1639 ( .A1(n1502), .A2(n1501), .ZN(n1503) );
  MAOI22D0BWP12T U1640 ( .A1(a[11]), .A2(n1503), .B1(a[11]), .B2(n1503), .ZN(
        mult_x_18_n659) );
  AOI22D1BWP12T U1641 ( .A1(b[14]), .A2(n2179), .B1(b[13]), .B2(n2178), .ZN(
        n1506) );
  FA1D0BWP12T U1642 ( .A(b[13]), .B(b[14]), .CI(n1504), .CO(n1471), .S(n2174)
         );
  AOI22D1BWP12T U1643 ( .A1(b[12]), .A2(n2182), .B1(n2174), .B2(n2180), .ZN(
        n1505) );
  ND2D1BWP12T U1644 ( .A1(n1506), .A2(n1505), .ZN(n1507) );
  MAOI22D0BWP12T U1645 ( .A1(a[17]), .A2(n1507), .B1(a[17]), .B2(n1507), .ZN(
        mult_x_18_n616) );
  AOI22D1BWP12T U1646 ( .A1(b[10]), .A2(n2197), .B1(b[9]), .B2(n2196), .ZN(
        n1509) );
  AOI22D1BWP12T U1647 ( .A1(b[8]), .A2(n1602), .B1(n2198), .B2(n2013), .ZN(
        n1508) );
  ND2D1BWP12T U1648 ( .A1(n1509), .A2(n1508), .ZN(n1510) );
  MAOI22D0BWP12T U1649 ( .A1(a[5]), .A2(n1510), .B1(a[5]), .B2(n1510), .ZN(
        mult_x_18_n722) );
  AOI22D1BWP12T U1650 ( .A1(b[8]), .A2(n2152), .B1(b[7]), .B2(n2151), .ZN(
        n1512) );
  AOI22D1BWP12T U1651 ( .A1(b[6]), .A2(n2155), .B1(n2163), .B2(n2153), .ZN(
        n1511) );
  ND2D1BWP12T U1652 ( .A1(n1512), .A2(n1511), .ZN(n1513) );
  MAOI22D0BWP12T U1653 ( .A1(a[23]), .A2(n1513), .B1(a[23]), .B2(n1513), .ZN(
        mult_x_18_n589) );
  AOI22D1BWP12T U1654 ( .A1(b[14]), .A2(n2185), .B1(b[13]), .B2(n2186), .ZN(
        n1515) );
  AOI22D1BWP12T U1655 ( .A1(b[12]), .A2(n2189), .B1(n2174), .B2(n2187), .ZN(
        n1514) );
  ND2D1BWP12T U1656 ( .A1(n1515), .A2(n1514), .ZN(n1516) );
  MAOI22D0BWP12T U1657 ( .A1(a[11]), .A2(n1516), .B1(a[11]), .B2(n1516), .ZN(
        mult_x_18_n661) );
  AOI22D1BWP12T U1658 ( .A1(b[11]), .A2(n2197), .B1(b[10]), .B2(n2196), .ZN(
        n1519) );
  FA1D0BWP12T U1659 ( .A(b[10]), .B(b[11]), .CI(n1517), .CO(n1437), .S(n2154)
         );
  AOI22D1BWP12T U1660 ( .A1(b[9]), .A2(n1602), .B1(n2154), .B2(n2198), .ZN(
        n1518) );
  ND2D1BWP12T U1661 ( .A1(n1519), .A2(n1518), .ZN(n1520) );
  MAOI22D0BWP12T U1662 ( .A1(a[5]), .A2(n1520), .B1(a[5]), .B2(n1520), .ZN(
        mult_x_18_n721) );
  AOI22D1BWP12T U1663 ( .A1(b[25]), .A2(n2197), .B1(b[24]), .B2(n2196), .ZN(
        n1523) );
  FA1D0BWP12T U1664 ( .A(b[24]), .B(b[25]), .CI(n1521), .CO(n1490), .S(n1988)
         );
  AOI22D1BWP12T U1665 ( .A1(b[23]), .A2(n2200), .B1(n2198), .B2(n1988), .ZN(
        n1522) );
  ND2D1BWP12T U1666 ( .A1(n1523), .A2(n1522), .ZN(n1524) );
  MAOI22D0BWP12T U1667 ( .A1(a[5]), .A2(n1524), .B1(a[5]), .B2(n1524), .ZN(
        mult_x_18_n707) );
  AOI22D1BWP12T U1668 ( .A1(b[15]), .A2(n2185), .B1(b[14]), .B2(n2186), .ZN(
        n1526) );
  AOI22D1BWP12T U1669 ( .A1(b[13]), .A2(n2189), .B1(n2187), .B2(n2067), .ZN(
        n1525) );
  ND2D1BWP12T U1670 ( .A1(n1526), .A2(n1525), .ZN(n1527) );
  MAOI22D0BWP12T U1671 ( .A1(a[11]), .A2(n1527), .B1(a[11]), .B2(n1527), .ZN(
        mult_x_18_n660) );
  AOI22D1BWP12T U1672 ( .A1(b[19]), .A2(n2185), .B1(b[18]), .B2(n2186), .ZN(
        n1529) );
  AOI22D1BWP12T U1673 ( .A1(b[17]), .A2(n2189), .B1(n2187), .B2(n2004), .ZN(
        n1528) );
  ND2D1BWP12T U1674 ( .A1(n1529), .A2(n1528), .ZN(n1530) );
  MAOI22D0BWP12T U1675 ( .A1(a[11]), .A2(n1530), .B1(a[11]), .B2(n1530), .ZN(
        mult_x_18_n656) );
  AOI22D1BWP12T U1676 ( .A1(b[9]), .A2(n2179), .B1(b[8]), .B2(n2178), .ZN(
        n1532) );
  AOI22D1BWP12T U1677 ( .A1(b[7]), .A2(n2182), .B1(n2180), .B2(n2017), .ZN(
        n1531) );
  ND2D1BWP12T U1678 ( .A1(n1532), .A2(n1531), .ZN(n1533) );
  MAOI22D0BWP12T U1679 ( .A1(a[17]), .A2(n1533), .B1(a[17]), .B2(n1533), .ZN(
        mult_x_18_n621) );
  AOI22D1BWP12T U1680 ( .A1(b[13]), .A2(n2179), .B1(b[12]), .B2(n2178), .ZN(
        n1536) );
  FA1D0BWP12T U1681 ( .A(b[12]), .B(b[13]), .CI(n1534), .CO(n1504), .S(n2062)
         );
  AOI22D1BWP12T U1682 ( .A1(b[11]), .A2(n2182), .B1(n2180), .B2(n2062), .ZN(
        n1535) );
  ND2D1BWP12T U1683 ( .A1(n1536), .A2(n1535), .ZN(n1537) );
  MAOI22D0BWP12T U1684 ( .A1(a[17]), .A2(n1537), .B1(a[17]), .B2(n1537), .ZN(
        mult_x_18_n617) );
  AOI22D1BWP12T U1685 ( .A1(b[22]), .A2(n2196), .B1(b[23]), .B2(n2197), .ZN(
        n1540) );
  FA1D0BWP12T U1686 ( .A(b[22]), .B(b[23]), .CI(n1538), .CO(n1416), .S(n2188)
         );
  AOI22D1BWP12T U1687 ( .A1(b[21]), .A2(n2200), .B1(n2198), .B2(n2188), .ZN(
        n1539) );
  ND2D1BWP12T U1688 ( .A1(n1540), .A2(n1539), .ZN(n1541) );
  MAOI22D0BWP12T U1689 ( .A1(a[5]), .A2(n1541), .B1(a[5]), .B2(n1541), .ZN(
        mult_x_18_n709) );
  AOI22D1BWP12T U1690 ( .A1(b[7]), .A2(n2152), .B1(b[6]), .B2(n2151), .ZN(
        n1543) );
  AOI22D1BWP12T U1691 ( .A1(b[5]), .A2(n2155), .B1(n2153), .B2(n2021), .ZN(
        n1542) );
  ND2D1BWP12T U1692 ( .A1(n1543), .A2(n1542), .ZN(n1544) );
  MAOI22D0BWP12T U1693 ( .A1(a[23]), .A2(n1544), .B1(a[23]), .B2(n1544), .ZN(
        mult_x_18_n590) );
  AOI22D1BWP12T U1694 ( .A1(b[6]), .A2(n2185), .B1(b[5]), .B2(n2186), .ZN(
        n1546) );
  AOI22D1BWP12T U1695 ( .A1(b[4]), .A2(n2189), .B1(n2187), .B2(n2043), .ZN(
        n1545) );
  ND2D1BWP12T U1696 ( .A1(n1546), .A2(n1545), .ZN(n1547) );
  MAOI22D0BWP12T U1697 ( .A1(a[11]), .A2(n1547), .B1(a[11]), .B2(n1547), .ZN(
        mult_x_18_n669) );
  AOI22D1BWP12T U1698 ( .A1(b[12]), .A2(n2197), .B1(b[11]), .B2(n2196), .ZN(
        n1549) );
  AOI22D1BWP12T U1699 ( .A1(b[10]), .A2(n1602), .B1(n2198), .B2(n2059), .ZN(
        n1548) );
  ND2D1BWP12T U1700 ( .A1(n1549), .A2(n1548), .ZN(n1550) );
  MAOI22D0BWP12T U1701 ( .A1(a[5]), .A2(n1550), .B1(a[5]), .B2(n1550), .ZN(
        mult_x_18_n720) );
  AOI22D1BWP12T U1702 ( .A1(b[12]), .A2(n2185), .B1(b[11]), .B2(n2186), .ZN(
        n1552) );
  AOI22D1BWP12T U1703 ( .A1(b[10]), .A2(n2189), .B1(n2187), .B2(n2059), .ZN(
        n1551) );
  ND2D1BWP12T U1704 ( .A1(n1552), .A2(n1551), .ZN(n1553) );
  MAOI22D0BWP12T U1705 ( .A1(a[11]), .A2(n1553), .B1(a[11]), .B2(n1553), .ZN(
        mult_x_18_n663) );
  AOI22D1BWP12T U1706 ( .A1(b[8]), .A2(n2179), .B1(b[7]), .B2(n2178), .ZN(
        n1555) );
  AOI22D1BWP12T U1707 ( .A1(b[6]), .A2(n2182), .B1(n2163), .B2(n2180), .ZN(
        n1554) );
  ND2D1BWP12T U1708 ( .A1(n1555), .A2(n1554), .ZN(n1556) );
  MAOI22D0BWP12T U1709 ( .A1(a[17]), .A2(n1556), .B1(a[17]), .B2(n1556), .ZN(
        mult_x_18_n622) );
  AOI22D1BWP12T U1710 ( .A1(b[18]), .A2(n2197), .B1(b[17]), .B2(n2196), .ZN(
        n1558) );
  AOI22D1BWP12T U1711 ( .A1(b[16]), .A2(n2200), .B1(n2198), .B2(n2008), .ZN(
        n1557) );
  ND2D1BWP12T U1712 ( .A1(n1558), .A2(n1557), .ZN(n1559) );
  MAOI22D0BWP12T U1713 ( .A1(a[5]), .A2(n1559), .B1(a[5]), .B2(n1559), .ZN(
        mult_x_18_n714) );
  AOI22D1BWP12T U1714 ( .A1(b[7]), .A2(n2185), .B1(b[6]), .B2(n2186), .ZN(
        n1561) );
  AOI22D1BWP12T U1715 ( .A1(b[5]), .A2(n2189), .B1(n2187), .B2(n2021), .ZN(
        n1560) );
  ND2D1BWP12T U1716 ( .A1(n1561), .A2(n1560), .ZN(n1562) );
  MAOI22D0BWP12T U1717 ( .A1(a[11]), .A2(n1562), .B1(a[11]), .B2(n1562), .ZN(
        mult_x_18_n668) );
  AOI22D1BWP12T U1718 ( .A1(b[8]), .A2(n2185), .B1(b[7]), .B2(n2186), .ZN(
        n1564) );
  AOI22D1BWP12T U1719 ( .A1(b[6]), .A2(n2189), .B1(n2163), .B2(n2187), .ZN(
        n1563) );
  ND2D1BWP12T U1720 ( .A1(n1564), .A2(n1563), .ZN(n1565) );
  MAOI22D0BWP12T U1721 ( .A1(a[11]), .A2(n1565), .B1(a[11]), .B2(n1565), .ZN(
        mult_x_18_n667) );
  AOI22D1BWP12T U1722 ( .A1(b[13]), .A2(n2197), .B1(b[12]), .B2(n2196), .ZN(
        n1567) );
  AOI22D1BWP12T U1723 ( .A1(b[11]), .A2(n1602), .B1(n2198), .B2(n2062), .ZN(
        n1566) );
  ND2D1BWP12T U1724 ( .A1(n1567), .A2(n1566), .ZN(n1568) );
  MAOI22D0BWP12T U1725 ( .A1(a[5]), .A2(n1568), .B1(a[5]), .B2(n1568), .ZN(
        mult_x_18_n719) );
  AOI22D1BWP12T U1726 ( .A1(b[13]), .A2(n2185), .B1(b[12]), .B2(n2186), .ZN(
        n1570) );
  AOI22D1BWP12T U1727 ( .A1(b[11]), .A2(n2189), .B1(n2187), .B2(n2062), .ZN(
        n1569) );
  ND2D1BWP12T U1728 ( .A1(n1570), .A2(n1569), .ZN(n1571) );
  MAOI22D0BWP12T U1729 ( .A1(a[11]), .A2(n1571), .B1(a[11]), .B2(n1571), .ZN(
        mult_x_18_n662) );
  AOI22D1BWP12T U1730 ( .A1(b[10]), .A2(n2179), .B1(b[9]), .B2(n2178), .ZN(
        n1573) );
  AOI22D1BWP12T U1731 ( .A1(b[8]), .A2(n2182), .B1(n2180), .B2(n2013), .ZN(
        n1572) );
  ND2D1BWP12T U1732 ( .A1(n1573), .A2(n1572), .ZN(n1574) );
  MAOI22D0BWP12T U1733 ( .A1(a[17]), .A2(n1574), .B1(a[17]), .B2(n1574), .ZN(
        mult_x_18_n620) );
  AOI22D1BWP12T U1734 ( .A1(b[16]), .A2(n2197), .B1(b[15]), .B2(n2196), .ZN(
        n1576) );
  AOI22D1BWP12T U1735 ( .A1(b[14]), .A2(n1602), .B1(n2198), .B2(n2070), .ZN(
        n1575) );
  ND2D1BWP12T U1736 ( .A1(n1576), .A2(n1575), .ZN(n1577) );
  MAOI22D0BWP12T U1737 ( .A1(a[5]), .A2(n1577), .B1(a[5]), .B2(n1577), .ZN(
        mult_x_18_n716) );
  AOI22D1BWP12T U1738 ( .A1(b[11]), .A2(n2179), .B1(b[10]), .B2(n2178), .ZN(
        n1579) );
  AOI22D1BWP12T U1739 ( .A1(b[9]), .A2(n2182), .B1(n2154), .B2(n2180), .ZN(
        n1578) );
  ND2D1BWP12T U1740 ( .A1(n1579), .A2(n1578), .ZN(n1580) );
  MAOI22D0BWP12T U1741 ( .A1(a[17]), .A2(n1580), .B1(a[17]), .B2(n1580), .ZN(
        mult_x_18_n619) );
  AOI22D1BWP12T U1742 ( .A1(b[7]), .A2(n2179), .B1(b[6]), .B2(n2178), .ZN(
        n1582) );
  AOI22D1BWP12T U1743 ( .A1(b[5]), .A2(n2182), .B1(n2180), .B2(n2021), .ZN(
        n1581) );
  ND2D1BWP12T U1744 ( .A1(n1582), .A2(n1581), .ZN(n1583) );
  MAOI22D0BWP12T U1745 ( .A1(a[17]), .A2(n1583), .B1(a[17]), .B2(n1583), .ZN(
        mult_x_18_n623) );
  AOI22D1BWP12T U1746 ( .A1(b[11]), .A2(n2185), .B1(b[10]), .B2(n2186), .ZN(
        n1585) );
  AOI22D1BWP12T U1747 ( .A1(b[9]), .A2(n2189), .B1(n2154), .B2(n2187), .ZN(
        n1584) );
  ND2D1BWP12T U1748 ( .A1(n1585), .A2(n1584), .ZN(n1586) );
  MAOI22D0BWP12T U1749 ( .A1(a[11]), .A2(n1586), .B1(a[11]), .B2(n1586), .ZN(
        mult_x_18_n664) );
  AOI22D1BWP12T U1750 ( .A1(b[14]), .A2(n2197), .B1(b[13]), .B2(n2196), .ZN(
        n1588) );
  AOI22D1BWP12T U1751 ( .A1(b[12]), .A2(n1602), .B1(n2198), .B2(n2174), .ZN(
        n1587) );
  ND2D1BWP12T U1752 ( .A1(n1588), .A2(n1587), .ZN(n1589) );
  MAOI22D0BWP12T U1753 ( .A1(a[5]), .A2(n1589), .B1(a[5]), .B2(n1589), .ZN(
        mult_x_18_n718) );
  AOI22D1BWP12T U1754 ( .A1(b[17]), .A2(n2197), .B1(b[16]), .B2(n2196), .ZN(
        n1591) );
  AOI22D1BWP12T U1755 ( .A1(b[15]), .A2(n1602), .B1(n2198), .B2(n2181), .ZN(
        n1590) );
  ND2D1BWP12T U1756 ( .A1(n1591), .A2(n1590), .ZN(n1592) );
  MAOI22D0BWP12T U1757 ( .A1(a[5]), .A2(n1592), .B1(a[5]), .B2(n1592), .ZN(
        mult_x_18_n715) );
  AOI22D1BWP12T U1758 ( .A1(b[20]), .A2(n2197), .B1(b[19]), .B2(n2196), .ZN(
        n1594) );
  AOI22D1BWP12T U1759 ( .A1(b[18]), .A2(n2200), .B1(n2095), .B2(n2198), .ZN(
        n1593) );
  ND2D1BWP12T U1760 ( .A1(n1594), .A2(n1593), .ZN(n1595) );
  MAOI22D0BWP12T U1761 ( .A1(a[5]), .A2(n1595), .B1(a[5]), .B2(n1595), .ZN(
        mult_x_18_n712) );
  AOI22D1BWP12T U1762 ( .A1(b[10]), .A2(n2185), .B1(b[9]), .B2(n2186), .ZN(
        n1597) );
  AOI22D1BWP12T U1763 ( .A1(b[8]), .A2(n2189), .B1(n2187), .B2(n2013), .ZN(
        n1596) );
  ND2D1BWP12T U1764 ( .A1(n1597), .A2(n1596), .ZN(n1598) );
  MAOI22D0BWP12T U1765 ( .A1(a[11]), .A2(n1598), .B1(a[11]), .B2(n1598), .ZN(
        mult_x_18_n665) );
  AOI22D1BWP12T U1766 ( .A1(b[22]), .A2(n2197), .B1(b[21]), .B2(n2196), .ZN(
        n1600) );
  AOI22D1BWP12T U1767 ( .A1(b[20]), .A2(n2200), .B1(n2198), .B2(n1995), .ZN(
        n1599) );
  ND2D1BWP12T U1768 ( .A1(n1600), .A2(n1599), .ZN(n1601) );
  MAOI22D0BWP12T U1769 ( .A1(a[5]), .A2(n1601), .B1(a[5]), .B2(n1601), .ZN(
        mult_x_18_n710) );
  AOI22D1BWP12T U1770 ( .A1(b[15]), .A2(n2197), .B1(b[14]), .B2(n2196), .ZN(
        n1604) );
  AOI22D1BWP12T U1771 ( .A1(b[13]), .A2(n1602), .B1(n2198), .B2(n2067), .ZN(
        n1603) );
  ND2D1BWP12T U1772 ( .A1(n1604), .A2(n1603), .ZN(n1605) );
  MAOI22D0BWP12T U1773 ( .A1(a[5]), .A2(n1605), .B1(a[5]), .B2(n1605), .ZN(
        mult_x_18_n717) );
  AOI22D1BWP12T U1774 ( .A1(b[21]), .A2(n2197), .B1(b[20]), .B2(n2196), .ZN(
        n1607) );
  AOI22D1BWP12T U1775 ( .A1(b[19]), .A2(n2200), .B1(n2198), .B2(n1998), .ZN(
        n1606) );
  ND2D1BWP12T U1776 ( .A1(n1607), .A2(n1606), .ZN(n1608) );
  MAOI22D0BWP12T U1777 ( .A1(a[5]), .A2(n1608), .B1(a[5]), .B2(n1608), .ZN(
        mult_x_18_n711) );
  AOI22D1BWP12T U1778 ( .A1(b[6]), .A2(n2179), .B1(b[5]), .B2(n2178), .ZN(
        n1610) );
  AOI22D1BWP12T U1779 ( .A1(b[4]), .A2(n2182), .B1(n2180), .B2(n2043), .ZN(
        n1609) );
  ND2D1BWP12T U1780 ( .A1(n1610), .A2(n1609), .ZN(n1611) );
  MAOI22D0BWP12T U1781 ( .A1(a[17]), .A2(n1611), .B1(a[17]), .B2(n1611), .ZN(
        mult_x_18_n624) );
  INVD1BWP12T U1782 ( .I(a[7]), .ZN(n3292) );
  INVD1BWP12T U1783 ( .I(a[6]), .ZN(n3276) );
  OAI22D1BWP12T U1784 ( .A1(n3292), .A2(a[6]), .B1(n3276), .B2(a[7]), .ZN(
        n1616) );
  INVD1BWP12T U1785 ( .I(a[5]), .ZN(n3247) );
  OAI22D1BWP12T U1786 ( .A1(n3276), .A2(a[5]), .B1(n3247), .B2(a[6]), .ZN(
        n1888) );
  INVD1BWP12T U1787 ( .I(n1888), .ZN(n2047) );
  AN2D1BWP12T U1788 ( .A1(n1616), .A2(n2047), .Z(n2144) );
  OAI22D1BWP12T U1789 ( .A1(n3321), .A2(n3292), .B1(a[7]), .B2(a[8]), .ZN(
        n1615) );
  NR2D1BWP12T U1790 ( .A1(n2047), .A2(n1615), .ZN(n2146) );
  ND2D1BWP12T U1791 ( .A1(n3219), .A2(b[3]), .ZN(n2662) );
  INVD1BWP12T U1792 ( .I(n2662), .ZN(n2912) );
  AOI221D1BWP12T U1793 ( .A1(b[3]), .A2(n1666), .B1(n2886), .B2(n1665), .C(
        n3219), .ZN(n1613) );
  NR2D1BWP12T U1794 ( .A1(n2914), .A2(n1614), .ZN(n1612) );
  AOI211D1BWP12T U1795 ( .A1(n1614), .A2(n2912), .B(n1613), .C(n1612), .ZN(
        n2033) );
  INVD1BWP12T U1796 ( .I(n2033), .ZN(n1933) );
  AOI22D1BWP12T U1797 ( .A1(b[3]), .A2(n2144), .B1(n2146), .B2(n1933), .ZN(
        n1618) );
  AN2D1BWP12T U1798 ( .A1(n1615), .A2(n1888), .Z(n2145) );
  NR3D1BWP12T U1799 ( .A1(n1888), .A2(n1616), .A3(n1615), .ZN(n2148) );
  AOI22D1BWP12T U1800 ( .A1(b[4]), .A2(n2145), .B1(b[2]), .B2(n2148), .ZN(
        n1617) );
  ND2D1BWP12T U1801 ( .A1(n1618), .A2(n1617), .ZN(n1619) );
  MAOI22D0BWP12T U1802 ( .A1(a[8]), .A2(n1619), .B1(a[8]), .B2(n1619), .ZN(
        mult_x_18_n698) );
  NR2D1BWP12T U1803 ( .A1(n3170), .A2(n1718), .ZN(mult_x_18_n428) );
  NR2D1BWP12T U1804 ( .A1(b[1]), .A2(b[0]), .ZN(n2512) );
  NR2D1BWP12T U1805 ( .A1(n2512), .A2(n1622), .ZN(n2570) );
  CKBD1BWP12T U1806 ( .I(n2570), .Z(n3881) );
  INVD1BWP12T U1807 ( .I(n3881), .ZN(n3878) );
  INVD1BWP12T U1808 ( .I(n2180), .ZN(n1819) );
  OAI222D1BWP12T U1809 ( .A1(n3878), .A2(n1819), .B1(n1621), .B2(n3165), .C1(
        n3170), .C2(n1620), .ZN(n1719) );
  NR3D1BWP12T U1810 ( .A1(mult_x_18_n428), .A2(n3565), .A3(n1719), .ZN(n1815)
         );
  NR2D1BWP12T U1811 ( .A1(n1815), .A2(n3565), .ZN(n1625) );
  ND2D1BWP12T U1812 ( .A1(b[2]), .A2(n1622), .ZN(n2445) );
  NR2D1BWP12T U1813 ( .A1(b[2]), .A2(b[1]), .ZN(n2849) );
  AOI31D1BWP12T U1814 ( .A1(n2445), .A2(n2382), .A3(b[1]), .B(n2849), .ZN(
        n1941) );
  AOI22D1BWP12T U1815 ( .A1(b[1]), .A2(n2178), .B1(n2180), .B2(n1941), .ZN(
        n1624) );
  AOI22D1BWP12T U1816 ( .A1(b[2]), .A2(n2179), .B1(b[0]), .B2(n2182), .ZN(
        n1623) );
  ND2D1BWP12T U1817 ( .A1(n1624), .A2(n1623), .ZN(n1816) );
  MAOI22D0BWP12T U1818 ( .A1(n1625), .A2(n1816), .B1(n1625), .B2(n1816), .ZN(
        mult_x_18_n412) );
  INVD1BWP12T U1819 ( .I(a[13]), .ZN(n3446) );
  INVD1BWP12T U1820 ( .I(a[12]), .ZN(n3428) );
  OAI22D1BWP12T U1821 ( .A1(n3446), .A2(a[12]), .B1(n3428), .B2(a[13]), .ZN(
        n1628) );
  OAI22D1BWP12T U1822 ( .A1(n3428), .A2(a[11]), .B1(n4005), .B2(a[12]), .ZN(
        n1833) );
  INVD1BWP12T U1823 ( .I(n1833), .ZN(n1626) );
  AN2D1BWP12T U1824 ( .A1(n1628), .A2(n1626), .Z(n2092) );
  OAI22D1BWP12T U1825 ( .A1(n3479), .A2(n3446), .B1(a[13]), .B2(a[14]), .ZN(
        n1627) );
  NR2D1BWP12T U1826 ( .A1(n1626), .A2(n1627), .ZN(n2094) );
  AOI22D1BWP12T U1827 ( .A1(b[3]), .A2(n2092), .B1(n2094), .B2(n1933), .ZN(
        n1630) );
  AN2D1BWP12T U1828 ( .A1(n1627), .A2(n1833), .Z(n2093) );
  NR3D1BWP12T U1829 ( .A1(n1833), .A2(n1628), .A3(n1627), .ZN(n2096) );
  AOI22D1BWP12T U1830 ( .A1(b[4]), .A2(n2093), .B1(b[2]), .B2(n2096), .ZN(
        n1629) );
  ND2D1BWP12T U1831 ( .A1(n1630), .A2(n1629), .ZN(n1631) );
  MAOI22D0BWP12T U1832 ( .A1(a[14]), .A2(n1631), .B1(a[14]), .B2(n1631), .ZN(
        mult_x_18_n647) );
  INVD1BWP12T U1833 ( .I(a[19]), .ZN(n3618) );
  INVD1BWP12T U1834 ( .I(a[18]), .ZN(n3578) );
  OAI22D1BWP12T U1835 ( .A1(n3618), .A2(a[18]), .B1(n3578), .B2(a[19]), .ZN(
        n1634) );
  OAI22D1BWP12T U1836 ( .A1(n3578), .A2(a[17]), .B1(n3565), .B2(a[18]), .ZN(
        n1811) );
  INVD1BWP12T U1837 ( .I(n1811), .ZN(n1632) );
  AN2D1BWP12T U1838 ( .A1(n1634), .A2(n1632), .Z(n2171) );
  OAI22D1BWP12T U1839 ( .A1(n3632), .A2(n3618), .B1(a[19]), .B2(a[20]), .ZN(
        n1633) );
  NR2D1BWP12T U1840 ( .A1(n1632), .A2(n1633), .ZN(n2173) );
  AOI22D1BWP12T U1841 ( .A1(b[3]), .A2(n2171), .B1(n2173), .B2(n1933), .ZN(
        n1636) );
  AN2D1BWP12T U1842 ( .A1(n1633), .A2(n1811), .Z(n2172) );
  NR3D1BWP12T U1843 ( .A1(n1811), .A2(n1634), .A3(n1633), .ZN(n2175) );
  AOI22D1BWP12T U1844 ( .A1(b[4]), .A2(n2172), .B1(b[2]), .B2(n2175), .ZN(
        n1635) );
  ND2D1BWP12T U1845 ( .A1(n1636), .A2(n1635), .ZN(n1637) );
  MAOI22D0BWP12T U1846 ( .A1(a[20]), .A2(n1637), .B1(a[20]), .B2(n1637), .ZN(
        mult_x_18_n608) );
  AOI22D1BWP12T U1847 ( .A1(b[25]), .A2(n2145), .B1(b[24]), .B2(n2144), .ZN(
        n1639) );
  AOI22D1BWP12T U1848 ( .A1(b[23]), .A2(n2148), .B1(n2146), .B2(n1988), .ZN(
        n1638) );
  ND2D1BWP12T U1849 ( .A1(n1639), .A2(n1638), .ZN(n1640) );
  MAOI22D0BWP12T U1850 ( .A1(a[8]), .A2(n1640), .B1(a[8]), .B2(n1640), .ZN(
        mult_x_18_n677) );
  AOI22D1BWP12T U1851 ( .A1(b[21]), .A2(n2145), .B1(b[20]), .B2(n2144), .ZN(
        n1642) );
  AOI22D1BWP12T U1852 ( .A1(b[19]), .A2(n2148), .B1(n2146), .B2(n1998), .ZN(
        n1641) );
  ND2D1BWP12T U1853 ( .A1(n1642), .A2(n1641), .ZN(n1643) );
  MAOI22D0BWP12T U1854 ( .A1(a[8]), .A2(n1643), .B1(a[8]), .B2(n1643), .ZN(
        mult_x_18_n681) );
  AOI22D1BWP12T U1855 ( .A1(b[24]), .A2(n2145), .B1(b[23]), .B2(n2144), .ZN(
        n1645) );
  AOI22D1BWP12T U1856 ( .A1(b[22]), .A2(n2148), .B1(n2146), .B2(n2073), .ZN(
        n1644) );
  ND2D1BWP12T U1857 ( .A1(n1645), .A2(n1644), .ZN(n1646) );
  MAOI22D0BWP12T U1858 ( .A1(a[8]), .A2(n1646), .B1(a[8]), .B2(n1646), .ZN(
        mult_x_18_n678) );
  INVD1BWP12T U1859 ( .I(a[25]), .ZN(n3768) );
  INVD1BWP12T U1860 ( .I(a[24]), .ZN(n2518) );
  OAI22D1BWP12T U1861 ( .A1(n3768), .A2(a[24]), .B1(n2518), .B2(a[25]), .ZN(
        n1649) );
  OAI22D1BWP12T U1862 ( .A1(n2518), .A2(a[23]), .B1(n3701), .B2(a[24]), .ZN(
        n1860) );
  INVD1BWP12T U1863 ( .I(n1860), .ZN(n1647) );
  AN2D1BWP12T U1864 ( .A1(n1649), .A2(n1647), .Z(n2160) );
  INVD1BWP12T U1865 ( .I(a[26]), .ZN(n3790) );
  OAI22D1BWP12T U1866 ( .A1(n3790), .A2(n3768), .B1(a[25]), .B2(a[26]), .ZN(
        n1648) );
  NR2D1BWP12T U1867 ( .A1(n1647), .A2(n1648), .ZN(n2162) );
  AOI22D1BWP12T U1868 ( .A1(b[3]), .A2(n2160), .B1(n2162), .B2(n1933), .ZN(
        n1651) );
  AN2D1BWP12T U1869 ( .A1(n1648), .A2(n1860), .Z(n2161) );
  NR3D1BWP12T U1870 ( .A1(n1860), .A2(n1649), .A3(n1648), .ZN(n2164) );
  AOI22D1BWP12T U1871 ( .A1(b[4]), .A2(n2161), .B1(b[2]), .B2(n2164), .ZN(
        n1650) );
  ND2D1BWP12T U1872 ( .A1(n1651), .A2(n1650), .ZN(n1652) );
  MAOI22D0BWP12T U1873 ( .A1(a[26]), .A2(n1652), .B1(a[26]), .B2(n1652), .ZN(
        mult_x_18_n581) );
  AOI22D1BWP12T U1874 ( .A1(b[22]), .A2(n2145), .B1(b[21]), .B2(n2144), .ZN(
        n1654) );
  AOI22D1BWP12T U1875 ( .A1(b[20]), .A2(n2148), .B1(n2146), .B2(n1995), .ZN(
        n1653) );
  ND2D1BWP12T U1876 ( .A1(n1654), .A2(n1653), .ZN(n1655) );
  MAOI22D0BWP12T U1877 ( .A1(a[8]), .A2(n1655), .B1(a[8]), .B2(n1655), .ZN(
        mult_x_18_n680) );
  AOI22D1BWP12T U1878 ( .A1(b[22]), .A2(n2144), .B1(b[23]), .B2(n2145), .ZN(
        n1657) );
  AOI22D1BWP12T U1879 ( .A1(b[21]), .A2(n2148), .B1(n2146), .B2(n2188), .ZN(
        n1656) );
  ND2D1BWP12T U1880 ( .A1(n1657), .A2(n1656), .ZN(n1658) );
  MAOI22D0BWP12T U1881 ( .A1(a[8]), .A2(n1658), .B1(a[8]), .B2(n1658), .ZN(
        mult_x_18_n679) );
  AOI22D1BWP12T U1882 ( .A1(b[19]), .A2(n2093), .B1(b[18]), .B2(n2092), .ZN(
        n1660) );
  AOI22D1BWP12T U1883 ( .A1(b[17]), .A2(n2096), .B1(n2094), .B2(n2004), .ZN(
        n1659) );
  ND2D1BWP12T U1884 ( .A1(n1660), .A2(n1659), .ZN(n1661) );
  MAOI22D0BWP12T U1885 ( .A1(a[14]), .A2(n1661), .B1(a[14]), .B2(n1661), .ZN(
        mult_x_18_n632) );
  AOI22D1BWP12T U1886 ( .A1(b[12]), .A2(n2172), .B1(b[11]), .B2(n2171), .ZN(
        n1663) );
  AOI22D1BWP12T U1887 ( .A1(b[10]), .A2(n2175), .B1(n2173), .B2(n2059), .ZN(
        n1662) );
  ND2D1BWP12T U1888 ( .A1(n1663), .A2(n1662), .ZN(n1664) );
  MAOI22D0BWP12T U1889 ( .A1(a[20]), .A2(n1664), .B1(a[20]), .B2(n1664), .ZN(
        mult_x_18_n600) );
  NR2D1BWP12T U1890 ( .A1(n1666), .A2(n1665), .ZN(n1667) );
  MAOI22D0BWP12T U1891 ( .A1(b[3]), .A2(n1667), .B1(b[3]), .B2(n1667), .ZN(
        n2026) );
  AOI22D1BWP12T U1892 ( .A1(b[2]), .A2(n2144), .B1(n2146), .B2(n2026), .ZN(
        n1669) );
  AOI22D1BWP12T U1893 ( .A1(b[3]), .A2(n2145), .B1(b[1]), .B2(n2148), .ZN(
        n1668) );
  ND2D1BWP12T U1894 ( .A1(n1669), .A2(n1668), .ZN(n1670) );
  MAOI22D0BWP12T U1895 ( .A1(a[8]), .A2(n1670), .B1(a[8]), .B2(n1670), .ZN(
        mult_x_18_n699) );
  AOI22D1BWP12T U1896 ( .A1(b[13]), .A2(n2172), .B1(b[12]), .B2(n2171), .ZN(
        n1672) );
  AOI22D1BWP12T U1897 ( .A1(b[11]), .A2(n2175), .B1(n2173), .B2(n2062), .ZN(
        n1671) );
  ND2D1BWP12T U1898 ( .A1(n1672), .A2(n1671), .ZN(n1673) );
  MAOI22D0BWP12T U1899 ( .A1(a[20]), .A2(n1673), .B1(a[20]), .B2(n1673), .ZN(
        mult_x_18_n599) );
  AOI22D1BWP12T U1900 ( .A1(b[11]), .A2(n2172), .B1(b[10]), .B2(n2171), .ZN(
        n1675) );
  AOI22D1BWP12T U1901 ( .A1(b[9]), .A2(n2175), .B1(n2154), .B2(n2173), .ZN(
        n1674) );
  ND2D1BWP12T U1902 ( .A1(n1675), .A2(n1674), .ZN(n1676) );
  MAOI22D0BWP12T U1903 ( .A1(a[20]), .A2(n1676), .B1(a[20]), .B2(n1676), .ZN(
        mult_x_18_n601) );
  AOI22D1BWP12T U1904 ( .A1(b[7]), .A2(n2161), .B1(b[6]), .B2(n2160), .ZN(
        n1678) );
  AOI22D1BWP12T U1905 ( .A1(b[5]), .A2(n2164), .B1(n2162), .B2(n2021), .ZN(
        n1677) );
  ND2D1BWP12T U1906 ( .A1(n1678), .A2(n1677), .ZN(n1679) );
  MAOI22D0BWP12T U1907 ( .A1(a[26]), .A2(n1679), .B1(a[26]), .B2(n1679), .ZN(
        mult_x_18_n578) );
  AOI22D1BWP12T U1908 ( .A1(b[6]), .A2(n2145), .B1(b[5]), .B2(n2144), .ZN(
        n1681) );
  AOI22D1BWP12T U1909 ( .A1(b[4]), .A2(n2148), .B1(n2146), .B2(n2043), .ZN(
        n1680) );
  ND2D1BWP12T U1910 ( .A1(n1681), .A2(n1680), .ZN(n1682) );
  MAOI22D0BWP12T U1911 ( .A1(a[8]), .A2(n1682), .B1(a[8]), .B2(n1682), .ZN(
        mult_x_18_n696) );
  AOI22D1BWP12T U1912 ( .A1(b[8]), .A2(n2145), .B1(b[7]), .B2(n2144), .ZN(
        n1684) );
  AOI22D1BWP12T U1913 ( .A1(b[6]), .A2(n2148), .B1(n2163), .B2(n2146), .ZN(
        n1683) );
  ND2D1BWP12T U1914 ( .A1(n1684), .A2(n1683), .ZN(n1685) );
  MAOI22D0BWP12T U1915 ( .A1(a[8]), .A2(n1685), .B1(a[8]), .B2(n1685), .ZN(
        mult_x_18_n694) );
  AOI22D1BWP12T U1916 ( .A1(b[5]), .A2(n2161), .B1(b[4]), .B2(n2160), .ZN(
        n1688) );
  FA1D0BWP12T U1917 ( .A(b[4]), .B(b[5]), .CI(n1686), .CO(n1448), .S(n2140) );
  AOI22D1BWP12T U1918 ( .A1(b[3]), .A2(n2164), .B1(n2140), .B2(n2162), .ZN(
        n1687) );
  ND2D1BWP12T U1919 ( .A1(n1688), .A2(n1687), .ZN(n1689) );
  MAOI22D0BWP12T U1920 ( .A1(a[26]), .A2(n1689), .B1(a[26]), .B2(n1689), .ZN(
        mult_x_18_n580) );
  AOI22D1BWP12T U1921 ( .A1(b[18]), .A2(n2093), .B1(b[17]), .B2(n2092), .ZN(
        n1691) );
  AOI22D1BWP12T U1922 ( .A1(b[16]), .A2(n2096), .B1(n2094), .B2(n2008), .ZN(
        n1690) );
  ND2D1BWP12T U1923 ( .A1(n1691), .A2(n1690), .ZN(n1692) );
  MAOI22D0BWP12T U1924 ( .A1(a[14]), .A2(n1692), .B1(a[14]), .B2(n1692), .ZN(
        mult_x_18_n633) );
  AOI22D1BWP12T U1925 ( .A1(b[2]), .A2(n2092), .B1(n2094), .B2(n2026), .ZN(
        n1694) );
  AOI22D1BWP12T U1926 ( .A1(b[3]), .A2(n2093), .B1(b[1]), .B2(n2096), .ZN(
        n1693) );
  ND2D1BWP12T U1927 ( .A1(n1694), .A2(n1693), .ZN(n1695) );
  MAOI22D0BWP12T U1928 ( .A1(a[14]), .A2(n1695), .B1(a[14]), .B2(n1695), .ZN(
        mult_x_18_n648) );
  AOI22D1BWP12T U1929 ( .A1(b[5]), .A2(n2145), .B1(b[4]), .B2(n2144), .ZN(
        n1697) );
  AOI22D1BWP12T U1930 ( .A1(b[3]), .A2(n2148), .B1(n2140), .B2(n2146), .ZN(
        n1696) );
  ND2D1BWP12T U1931 ( .A1(n1697), .A2(n1696), .ZN(n1698) );
  MAOI22D0BWP12T U1932 ( .A1(a[8]), .A2(n1698), .B1(a[8]), .B2(n1698), .ZN(
        mult_x_18_n697) );
  AOI22D1BWP12T U1933 ( .A1(b[16]), .A2(n2093), .B1(b[15]), .B2(n2092), .ZN(
        n1700) );
  AOI22D1BWP12T U1934 ( .A1(b[14]), .A2(n2096), .B1(n2094), .B2(n2070), .ZN(
        n1699) );
  ND2D1BWP12T U1935 ( .A1(n1700), .A2(n1699), .ZN(n1701) );
  MAOI22D0BWP12T U1936 ( .A1(a[14]), .A2(n1701), .B1(a[14]), .B2(n1701), .ZN(
        mult_x_18_n635) );
  AOI22D1BWP12T U1937 ( .A1(b[10]), .A2(n2172), .B1(b[9]), .B2(n2171), .ZN(
        n1703) );
  AOI22D1BWP12T U1938 ( .A1(b[8]), .A2(n2175), .B1(n2173), .B2(n2013), .ZN(
        n1702) );
  ND2D1BWP12T U1939 ( .A1(n1703), .A2(n1702), .ZN(n1704) );
  MAOI22D0BWP12T U1940 ( .A1(a[20]), .A2(n1704), .B1(a[20]), .B2(n1704), .ZN(
        mult_x_18_n602) );
  AOI22D1BWP12T U1941 ( .A1(b[6]), .A2(n2161), .B1(b[5]), .B2(n2160), .ZN(
        n1706) );
  AOI22D1BWP12T U1942 ( .A1(b[4]), .A2(n2164), .B1(n2162), .B2(n2043), .ZN(
        n1705) );
  ND2D1BWP12T U1943 ( .A1(n1706), .A2(n1705), .ZN(n1707) );
  MAOI22D0BWP12T U1944 ( .A1(a[26]), .A2(n1707), .B1(a[26]), .B2(n1707), .ZN(
        mult_x_18_n579) );
  AOI22D1BWP12T U1945 ( .A1(b[9]), .A2(n2145), .B1(b[8]), .B2(n2144), .ZN(
        n1709) );
  AOI22D1BWP12T U1946 ( .A1(b[7]), .A2(n2148), .B1(n2146), .B2(n2017), .ZN(
        n1708) );
  ND2D1BWP12T U1947 ( .A1(n1709), .A2(n1708), .ZN(n1710) );
  MAOI22D0BWP12T U1948 ( .A1(a[8]), .A2(n1710), .B1(a[8]), .B2(n1710), .ZN(
        mult_x_18_n693) );
  AOI22D1BWP12T U1949 ( .A1(b[17]), .A2(n2093), .B1(b[16]), .B2(n2092), .ZN(
        n1712) );
  AOI22D1BWP12T U1950 ( .A1(b[15]), .A2(n2096), .B1(n2094), .B2(n2181), .ZN(
        n1711) );
  ND2D1BWP12T U1951 ( .A1(n1712), .A2(n1711), .ZN(n1713) );
  MAOI22D0BWP12T U1952 ( .A1(a[14]), .A2(n1713), .B1(a[14]), .B2(n1713), .ZN(
        mult_x_18_n634) );
  AOI22D1BWP12T U1953 ( .A1(b[7]), .A2(n2145), .B1(b[6]), .B2(n2144), .ZN(
        n1715) );
  AOI22D1BWP12T U1954 ( .A1(b[5]), .A2(n2148), .B1(n2146), .B2(n2021), .ZN(
        n1714) );
  ND2D1BWP12T U1955 ( .A1(n1715), .A2(n1714), .ZN(n1716) );
  MAOI22D0BWP12T U1956 ( .A1(a[8]), .A2(n1716), .B1(a[8]), .B2(n1716), .ZN(
        mult_x_18_n695) );
  ND2D1BWP12T U1957 ( .A1(a[17]), .A2(b[0]), .ZN(n1717) );
  NR2D1BWP12T U1958 ( .A1(n1718), .A2(n1717), .ZN(n1720) );
  MAOI22D0BWP12T U1959 ( .A1(n1720), .A2(n1719), .B1(n1720), .B2(n1719), .ZN(
        mult_x_18_n420) );
  AOI22D1BWP12T U1960 ( .A1(b[15]), .A2(n2093), .B1(b[14]), .B2(n2092), .ZN(
        n1722) );
  AOI22D1BWP12T U1961 ( .A1(b[13]), .A2(n2096), .B1(n2094), .B2(n2067), .ZN(
        n1721) );
  ND2D1BWP12T U1962 ( .A1(n1722), .A2(n1721), .ZN(n1723) );
  MAOI22D0BWP12T U1963 ( .A1(a[14]), .A2(n1723), .B1(a[14]), .B2(n1723), .ZN(
        mult_x_18_n636) );
  AOI22D1BWP12T U1964 ( .A1(b[10]), .A2(n2093), .B1(b[9]), .B2(n2092), .ZN(
        n1725) );
  AOI22D1BWP12T U1965 ( .A1(b[8]), .A2(n2096), .B1(n2094), .B2(n2013), .ZN(
        n1724) );
  ND2D1BWP12T U1966 ( .A1(n1725), .A2(n1724), .ZN(n1726) );
  MAOI22D0BWP12T U1967 ( .A1(a[14]), .A2(n1726), .B1(a[14]), .B2(n1726), .ZN(
        mult_x_18_n641) );
  AOI22D1BWP12T U1968 ( .A1(b[9]), .A2(n2172), .B1(b[8]), .B2(n2171), .ZN(
        n1728) );
  AOI22D1BWP12T U1969 ( .A1(b[7]), .A2(n2175), .B1(n2173), .B2(n2017), .ZN(
        n1727) );
  ND2D1BWP12T U1970 ( .A1(n1728), .A2(n1727), .ZN(n1729) );
  MAOI22D0BWP12T U1971 ( .A1(a[20]), .A2(n1729), .B1(a[20]), .B2(n1729), .ZN(
        mult_x_18_n603) );
  AOI22D1BWP12T U1972 ( .A1(b[10]), .A2(n2145), .B1(b[9]), .B2(n2144), .ZN(
        n1731) );
  AOI22D1BWP12T U1973 ( .A1(b[8]), .A2(n2148), .B1(n2146), .B2(n2013), .ZN(
        n1730) );
  ND2D1BWP12T U1974 ( .A1(n1731), .A2(n1730), .ZN(n1732) );
  MAOI22D0BWP12T U1975 ( .A1(a[8]), .A2(n1732), .B1(a[8]), .B2(n1732), .ZN(
        mult_x_18_n692) );
  AOI22D1BWP12T U1976 ( .A1(b[5]), .A2(n2093), .B1(b[4]), .B2(n2092), .ZN(
        n1734) );
  AOI22D1BWP12T U1977 ( .A1(b[3]), .A2(n2096), .B1(n2094), .B2(n2140), .ZN(
        n1733) );
  ND2D1BWP12T U1978 ( .A1(n1734), .A2(n1733), .ZN(n1735) );
  MAOI22D0BWP12T U1979 ( .A1(a[14]), .A2(n1735), .B1(a[14]), .B2(n1735), .ZN(
        mult_x_18_n646) );
  AOI22D1BWP12T U1980 ( .A1(b[2]), .A2(n2160), .B1(n2162), .B2(n2026), .ZN(
        n1737) );
  AOI22D1BWP12T U1981 ( .A1(b[3]), .A2(n2161), .B1(b[1]), .B2(n2164), .ZN(
        n1736) );
  ND2D1BWP12T U1982 ( .A1(n1737), .A2(n1736), .ZN(n1738) );
  MAOI22D0BWP12T U1983 ( .A1(a[26]), .A2(n1738), .B1(a[26]), .B2(n1738), .ZN(
        mult_x_18_n582) );
  AOI22D1BWP12T U1984 ( .A1(b[20]), .A2(n2145), .B1(b[19]), .B2(n2144), .ZN(
        n1740) );
  AOI22D1BWP12T U1985 ( .A1(b[18]), .A2(n2148), .B1(n2095), .B2(n2146), .ZN(
        n1739) );
  ND2D1BWP12T U1986 ( .A1(n1740), .A2(n1739), .ZN(n1741) );
  MAOI22D0BWP12T U1987 ( .A1(a[8]), .A2(n1741), .B1(a[8]), .B2(n1741), .ZN(
        mult_x_18_n682) );
  AOI22D1BWP12T U1988 ( .A1(b[11]), .A2(n2145), .B1(b[10]), .B2(n2144), .ZN(
        n1743) );
  AOI22D1BWP12T U1989 ( .A1(b[9]), .A2(n2148), .B1(n2146), .B2(n2154), .ZN(
        n1742) );
  ND2D1BWP12T U1990 ( .A1(n1743), .A2(n1742), .ZN(n1744) );
  MAOI22D0BWP12T U1991 ( .A1(a[8]), .A2(n1744), .B1(a[8]), .B2(n1744), .ZN(
        mult_x_18_n691) );
  AOI22D1BWP12T U1992 ( .A1(b[14]), .A2(n2093), .B1(b[13]), .B2(n2092), .ZN(
        n1746) );
  AOI22D1BWP12T U1993 ( .A1(b[12]), .A2(n2096), .B1(n2094), .B2(n2174), .ZN(
        n1745) );
  ND2D1BWP12T U1994 ( .A1(n1746), .A2(n1745), .ZN(n1747) );
  MAOI22D0BWP12T U1995 ( .A1(a[14]), .A2(n1747), .B1(a[14]), .B2(n1747), .ZN(
        mult_x_18_n637) );
  AOI22D1BWP12T U1996 ( .A1(b[6]), .A2(n2093), .B1(b[5]), .B2(n2092), .ZN(
        n1749) );
  AOI22D1BWP12T U1997 ( .A1(b[4]), .A2(n2096), .B1(n2094), .B2(n2043), .ZN(
        n1748) );
  ND2D1BWP12T U1998 ( .A1(n1749), .A2(n1748), .ZN(n1750) );
  MAOI22D0BWP12T U1999 ( .A1(a[14]), .A2(n1750), .B1(a[14]), .B2(n1750), .ZN(
        mult_x_18_n645) );
  AOI22D1BWP12T U2000 ( .A1(b[8]), .A2(n2172), .B1(b[7]), .B2(n2171), .ZN(
        n1752) );
  AOI22D1BWP12T U2001 ( .A1(b[6]), .A2(n2175), .B1(n2163), .B2(n2173), .ZN(
        n1751) );
  ND2D1BWP12T U2002 ( .A1(n1752), .A2(n1751), .ZN(n1753) );
  MAOI22D0BWP12T U2003 ( .A1(a[20]), .A2(n1753), .B1(a[20]), .B2(n1753), .ZN(
        mult_x_18_n604) );
  AOI22D1BWP12T U2004 ( .A1(b[12]), .A2(n2145), .B1(b[11]), .B2(n2144), .ZN(
        n1755) );
  AOI22D1BWP12T U2005 ( .A1(b[10]), .A2(n2148), .B1(n2146), .B2(n2059), .ZN(
        n1754) );
  ND2D1BWP12T U2006 ( .A1(n1755), .A2(n1754), .ZN(n1756) );
  MAOI22D0BWP12T U2007 ( .A1(a[8]), .A2(n1756), .B1(a[8]), .B2(n1756), .ZN(
        mult_x_18_n690) );
  AOI22D1BWP12T U2008 ( .A1(b[19]), .A2(n2145), .B1(b[18]), .B2(n2144), .ZN(
        n1758) );
  AOI22D1BWP12T U2009 ( .A1(b[17]), .A2(n2148), .B1(n2146), .B2(n2004), .ZN(
        n1757) );
  ND2D1BWP12T U2010 ( .A1(n1758), .A2(n1757), .ZN(n1759) );
  MAOI22D0BWP12T U2011 ( .A1(a[8]), .A2(n1759), .B1(a[8]), .B2(n1759), .ZN(
        mult_x_18_n683) );
  AOI22D1BWP12T U2012 ( .A1(b[7]), .A2(n2093), .B1(b[6]), .B2(n2092), .ZN(
        n1761) );
  AOI22D1BWP12T U2013 ( .A1(b[5]), .A2(n2096), .B1(n2094), .B2(n2021), .ZN(
        n1760) );
  ND2D1BWP12T U2014 ( .A1(n1761), .A2(n1760), .ZN(n1762) );
  MAOI22D0BWP12T U2015 ( .A1(a[14]), .A2(n1762), .B1(a[14]), .B2(n1762), .ZN(
        mult_x_18_n644) );
  AOI22D1BWP12T U2016 ( .A1(b[13]), .A2(n2093), .B1(b[12]), .B2(n2092), .ZN(
        n1764) );
  AOI22D1BWP12T U2017 ( .A1(b[11]), .A2(n2096), .B1(n2094), .B2(n2062), .ZN(
        n1763) );
  ND2D1BWP12T U2018 ( .A1(n1764), .A2(n1763), .ZN(n1765) );
  MAOI22D0BWP12T U2019 ( .A1(a[14]), .A2(n1765), .B1(a[14]), .B2(n1765), .ZN(
        mult_x_18_n638) );
  AOI22D1BWP12T U2020 ( .A1(b[13]), .A2(n2145), .B1(b[12]), .B2(n2144), .ZN(
        n1767) );
  AOI22D1BWP12T U2021 ( .A1(b[11]), .A2(n2148), .B1(n2146), .B2(n2062), .ZN(
        n1766) );
  ND2D1BWP12T U2022 ( .A1(n1767), .A2(n1766), .ZN(n1768) );
  MAOI22D0BWP12T U2023 ( .A1(a[8]), .A2(n1768), .B1(a[8]), .B2(n1768), .ZN(
        mult_x_18_n689) );
  AOI22D1BWP12T U2024 ( .A1(b[7]), .A2(n2172), .B1(b[6]), .B2(n2171), .ZN(
        n1770) );
  AOI22D1BWP12T U2025 ( .A1(b[5]), .A2(n2175), .B1(n2173), .B2(n2021), .ZN(
        n1769) );
  ND2D1BWP12T U2026 ( .A1(n1770), .A2(n1769), .ZN(n1771) );
  MAOI22D0BWP12T U2027 ( .A1(a[20]), .A2(n1771), .B1(a[20]), .B2(n1771), .ZN(
        mult_x_18_n605) );
  AOI22D1BWP12T U2028 ( .A1(b[8]), .A2(n2093), .B1(b[7]), .B2(n2092), .ZN(
        n1773) );
  AOI22D1BWP12T U2029 ( .A1(b[6]), .A2(n2096), .B1(n2094), .B2(n2163), .ZN(
        n1772) );
  ND2D1BWP12T U2030 ( .A1(n1773), .A2(n1772), .ZN(n1774) );
  MAOI22D0BWP12T U2031 ( .A1(a[14]), .A2(n1774), .B1(a[14]), .B2(n1774), .ZN(
        mult_x_18_n643) );
  AOI22D1BWP12T U2032 ( .A1(b[18]), .A2(n2145), .B1(b[17]), .B2(n2144), .ZN(
        n1776) );
  AOI22D1BWP12T U2033 ( .A1(b[16]), .A2(n2148), .B1(n2146), .B2(n2008), .ZN(
        n1775) );
  ND2D1BWP12T U2034 ( .A1(n1776), .A2(n1775), .ZN(n1777) );
  MAOI22D0BWP12T U2035 ( .A1(a[8]), .A2(n1777), .B1(a[8]), .B2(n1777), .ZN(
        mult_x_18_n684) );
  AOI22D1BWP12T U2036 ( .A1(b[12]), .A2(n2093), .B1(b[11]), .B2(n2092), .ZN(
        n1779) );
  AOI22D1BWP12T U2037 ( .A1(b[10]), .A2(n2096), .B1(n2094), .B2(n2059), .ZN(
        n1778) );
  ND2D1BWP12T U2038 ( .A1(n1779), .A2(n1778), .ZN(n1780) );
  MAOI22D0BWP12T U2039 ( .A1(a[14]), .A2(n1780), .B1(a[14]), .B2(n1780), .ZN(
        mult_x_18_n639) );
  AOI22D1BWP12T U2040 ( .A1(b[14]), .A2(n2145), .B1(b[13]), .B2(n2144), .ZN(
        n1782) );
  AOI22D1BWP12T U2041 ( .A1(b[12]), .A2(n2148), .B1(n2146), .B2(n2174), .ZN(
        n1781) );
  ND2D1BWP12T U2042 ( .A1(n1782), .A2(n1781), .ZN(n1783) );
  MAOI22D0BWP12T U2043 ( .A1(a[8]), .A2(n1783), .B1(a[8]), .B2(n1783), .ZN(
        mult_x_18_n688) );
  AOI22D1BWP12T U2044 ( .A1(b[2]), .A2(n2171), .B1(n2173), .B2(n2026), .ZN(
        n1785) );
  AOI22D1BWP12T U2045 ( .A1(b[3]), .A2(n2172), .B1(b[1]), .B2(n2175), .ZN(
        n1784) );
  ND2D1BWP12T U2046 ( .A1(n1785), .A2(n1784), .ZN(n1786) );
  MAOI22D0BWP12T U2047 ( .A1(a[20]), .A2(n1786), .B1(a[20]), .B2(n1786), .ZN(
        mult_x_18_n609) );
  AOI22D1BWP12T U2048 ( .A1(b[15]), .A2(n2145), .B1(b[14]), .B2(n2144), .ZN(
        n1788) );
  AOI22D1BWP12T U2049 ( .A1(b[13]), .A2(n2148), .B1(n2146), .B2(n2067), .ZN(
        n1787) );
  ND2D1BWP12T U2050 ( .A1(n1788), .A2(n1787), .ZN(n1789) );
  MAOI22D0BWP12T U2051 ( .A1(a[8]), .A2(n1789), .B1(a[8]), .B2(n1789), .ZN(
        mult_x_18_n687) );
  AOI22D1BWP12T U2052 ( .A1(b[6]), .A2(n2172), .B1(b[5]), .B2(n2171), .ZN(
        n1791) );
  AOI22D1BWP12T U2053 ( .A1(b[4]), .A2(n2175), .B1(n2173), .B2(n2043), .ZN(
        n1790) );
  ND2D1BWP12T U2054 ( .A1(n1791), .A2(n1790), .ZN(n1792) );
  MAOI22D0BWP12T U2055 ( .A1(a[20]), .A2(n1792), .B1(a[20]), .B2(n1792), .ZN(
        mult_x_18_n606) );
  AOI22D1BWP12T U2056 ( .A1(b[17]), .A2(n2145), .B1(b[16]), .B2(n2144), .ZN(
        n1794) );
  AOI22D1BWP12T U2057 ( .A1(b[15]), .A2(n2148), .B1(n2146), .B2(n2181), .ZN(
        n1793) );
  ND2D1BWP12T U2058 ( .A1(n1794), .A2(n1793), .ZN(n1795) );
  MAOI22D0BWP12T U2059 ( .A1(a[8]), .A2(n1795), .B1(a[8]), .B2(n1795), .ZN(
        mult_x_18_n685) );
  AOI22D1BWP12T U2060 ( .A1(b[11]), .A2(n2093), .B1(b[10]), .B2(n2092), .ZN(
        n1797) );
  AOI22D1BWP12T U2061 ( .A1(b[9]), .A2(n2096), .B1(n2094), .B2(n2154), .ZN(
        n1796) );
  ND2D1BWP12T U2062 ( .A1(n1797), .A2(n1796), .ZN(n1798) );
  MAOI22D0BWP12T U2063 ( .A1(a[14]), .A2(n1798), .B1(a[14]), .B2(n1798), .ZN(
        mult_x_18_n640) );
  AOI22D1BWP12T U2064 ( .A1(b[9]), .A2(n2093), .B1(b[8]), .B2(n2092), .ZN(
        n1800) );
  AOI22D1BWP12T U2065 ( .A1(b[7]), .A2(n2096), .B1(n2094), .B2(n2017), .ZN(
        n1799) );
  ND2D1BWP12T U2066 ( .A1(n1800), .A2(n1799), .ZN(n1801) );
  MAOI22D0BWP12T U2067 ( .A1(a[14]), .A2(n1801), .B1(a[14]), .B2(n1801), .ZN(
        mult_x_18_n642) );
  AOI22D1BWP12T U2068 ( .A1(b[5]), .A2(n2172), .B1(b[4]), .B2(n2171), .ZN(
        n1803) );
  AOI22D1BWP12T U2069 ( .A1(b[3]), .A2(n2175), .B1(n2140), .B2(n2173), .ZN(
        n1802) );
  ND2D1BWP12T U2070 ( .A1(n1803), .A2(n1802), .ZN(n1804) );
  MAOI22D0BWP12T U2071 ( .A1(a[20]), .A2(n1804), .B1(a[20]), .B2(n1804), .ZN(
        mult_x_18_n607) );
  AOI22D1BWP12T U2072 ( .A1(b[16]), .A2(n2145), .B1(b[15]), .B2(n2144), .ZN(
        n1806) );
  AOI22D1BWP12T U2073 ( .A1(b[14]), .A2(n2148), .B1(n2146), .B2(n2070), .ZN(
        n1805) );
  ND2D1BWP12T U2074 ( .A1(n1806), .A2(n1805), .ZN(n1807) );
  MAOI22D0BWP12T U2075 ( .A1(a[8]), .A2(n1807), .B1(a[8]), .B2(n1807), .ZN(
        mult_x_18_n686) );
  AOI22D1BWP12T U2076 ( .A1(b[5]), .A2(n2179), .B1(b[4]), .B2(n2178), .ZN(
        n1809) );
  AOI22D1BWP12T U2077 ( .A1(b[3]), .A2(n2182), .B1(n2140), .B2(n2180), .ZN(
        n1808) );
  ND2D1BWP12T U2078 ( .A1(n1809), .A2(n1808), .ZN(n1810) );
  MAOI22D0BWP12T U2079 ( .A1(n3565), .A2(n1810), .B1(n3565), .B2(n1810), .ZN(
        n1924) );
  ND2D1BWP12T U2080 ( .A1(b[0]), .A2(n1811), .ZN(n1919) );
  AOI22D1BWP12T U2081 ( .A1(b[2]), .A2(n2178), .B1(n2180), .B2(n2026), .ZN(
        n1813) );
  AOI22D1BWP12T U2082 ( .A1(b[3]), .A2(n2179), .B1(b[1]), .B2(n2182), .ZN(
        n1812) );
  ND2D1BWP12T U2083 ( .A1(n1813), .A2(n1812), .ZN(n1814) );
  MAOI22D0BWP12T U2084 ( .A1(n3565), .A2(n1814), .B1(n3565), .B2(n1814), .ZN(
        n1918) );
  IND2D1BWP12T U2085 ( .A1(n1816), .B1(n1815), .ZN(n1917) );
  AOI22D1BWP12T U2086 ( .A1(b[3]), .A2(n2178), .B1(b[2]), .B2(n2182), .ZN(
        n1818) );
  ND2D1BWP12T U2087 ( .A1(b[4]), .A2(n2179), .ZN(n1817) );
  OAI211D1BWP12T U2088 ( .A1(n2033), .A2(n1819), .B(n1818), .C(n1817), .ZN(
        n1820) );
  MAOI22D0BWP12T U2089 ( .A1(n3565), .A2(n1820), .B1(n3565), .B2(n1820), .ZN(
        n1927) );
  AOI222D1BWP12T U2090 ( .A1(b[1]), .A2(n2172), .B1(b[0]), .B2(n2171), .C1(
        n2173), .C2(n3881), .ZN(n1821) );
  INVD1BWP12T U2091 ( .I(a[20]), .ZN(n3632) );
  OAI21D1BWP12T U2092 ( .A1(n3632), .A2(n1919), .B(n1821), .ZN(n1899) );
  OAI31D1BWP12T U2093 ( .A1(n1821), .A2(n1919), .A3(n3632), .B(n1899), .ZN(
        n1926) );
  ND2D1BWP12T U2094 ( .A1(a[20]), .A2(n1899), .ZN(n1824) );
  AOI22D1BWP12T U2095 ( .A1(b[1]), .A2(n2171), .B1(n2173), .B2(n1941), .ZN(
        n1823) );
  AOI22D1BWP12T U2096 ( .A1(b[2]), .A2(n2172), .B1(b[0]), .B2(n2175), .ZN(
        n1822) );
  ND2D1BWP12T U2097 ( .A1(n1823), .A2(n1822), .ZN(n1898) );
  MAOI22D0BWP12T U2098 ( .A1(n1824), .A2(n1898), .B1(n1824), .B2(n1898), .ZN(
        n1922) );
  INVD1BWP12T U2099 ( .I(n1825), .ZN(mult_x_18_n381) );
  ND2D1BWP12T U2100 ( .A1(a[11]), .A2(b[0]), .ZN(n1826) );
  NR2D1BWP12T U2101 ( .A1(n1921), .A2(n1826), .ZN(n1969) );
  INVD1BWP12T U2102 ( .I(n2187), .ZN(n1836) );
  INVD1BWP12T U2103 ( .I(n2185), .ZN(n1838) );
  INVD1BWP12T U2104 ( .I(n2186), .ZN(n1837) );
  OAI222D1BWP12T U2105 ( .A1(n3878), .A2(n1836), .B1(n1838), .B2(n3165), .C1(
        n1837), .C2(n3170), .ZN(n1968) );
  NR2D1BWP12T U2106 ( .A1(n1969), .A2(n1968), .ZN(n4006) );
  NR2D1BWP12T U2107 ( .A1(n3165), .A2(n1837), .ZN(n1828) );
  INVD1BWP12T U2108 ( .I(n2189), .ZN(n1835) );
  INVD1BWP12T U2109 ( .I(n1941), .ZN(n2027) );
  OAI22D1BWP12T U2110 ( .A1(n2534), .A2(n1835), .B1(n1836), .B2(n2027), .ZN(
        n1827) );
  AOI211D1BWP12T U2111 ( .A1(n2185), .A2(b[2]), .B(n1828), .C(n1827), .ZN(
        n4008) );
  AOI21D1BWP12T U2112 ( .A1(n4006), .A2(n4008), .B(n4005), .ZN(n1832) );
  AOI22D1BWP12T U2113 ( .A1(b[1]), .A2(n2189), .B1(n2187), .B2(n2026), .ZN(
        n1830) );
  AOI22D1BWP12T U2114 ( .A1(b[3]), .A2(n2185), .B1(b[2]), .B2(n2186), .ZN(
        n1829) );
  ND2D1BWP12T U2115 ( .A1(n1830), .A2(n1829), .ZN(n1831) );
  NR2D1BWP12T U2116 ( .A1(n1832), .A2(n1831), .ZN(n1834) );
  ND2D1BWP12T U2117 ( .A1(b[0]), .A2(n1833), .ZN(n1911) );
  NR2D1BWP12T U2118 ( .A1(n1912), .A2(n1911), .ZN(n1910) );
  AOI21D1BWP12T U2119 ( .A1(n1834), .A2(a[11]), .B(n1910), .ZN(n1915) );
  OAI22D1BWP12T U2120 ( .A1(n2033), .A2(n1836), .B1(n2652), .B2(n1835), .ZN(
        n1840) );
  OAI22D1BWP12T U2121 ( .A1(n3219), .A2(n1838), .B1(n2886), .B2(n1837), .ZN(
        n1839) );
  NR2D1BWP12T U2122 ( .A1(n1840), .A2(n1839), .ZN(n1841) );
  MAOI22D0BWP12T U2123 ( .A1(a[11]), .A2(n1841), .B1(a[11]), .B2(n1841), .ZN(
        n1914) );
  AOI222D1BWP12T U2124 ( .A1(b[1]), .A2(n2093), .B1(b[0]), .B2(n2092), .C1(
        n2094), .C2(n3881), .ZN(n1842) );
  INVD1BWP12T U2125 ( .I(a[14]), .ZN(n3479) );
  OAI21D1BWP12T U2126 ( .A1(n3479), .A2(n1911), .B(n1842), .ZN(n1903) );
  OAI31D1BWP12T U2127 ( .A1(n1842), .A2(n1911), .A3(n3479), .B(n1903), .ZN(
        n1913) );
  ND2D1BWP12T U2128 ( .A1(a[14]), .A2(n1903), .ZN(n1845) );
  AOI22D1BWP12T U2129 ( .A1(b[1]), .A2(n2092), .B1(n2094), .B2(n1941), .ZN(
        n1844) );
  AOI22D1BWP12T U2130 ( .A1(b[2]), .A2(n2093), .B1(b[0]), .B2(n2096), .ZN(
        n1843) );
  ND2D1BWP12T U2131 ( .A1(n1844), .A2(n1843), .ZN(n1902) );
  MAOI22D0BWP12T U2132 ( .A1(n1845), .A2(n1902), .B1(n1845), .B2(n1902), .ZN(
        n1907) );
  AOI22D1BWP12T U2133 ( .A1(b[5]), .A2(n2185), .B1(b[4]), .B2(n2186), .ZN(
        n1847) );
  AOI22D1BWP12T U2134 ( .A1(b[3]), .A2(n2189), .B1(n2140), .B2(n2187), .ZN(
        n1846) );
  ND2D1BWP12T U2135 ( .A1(n1847), .A2(n1846), .ZN(n1848) );
  MAOI22D0BWP12T U2136 ( .A1(n4005), .A2(n1848), .B1(n4005), .B2(n1848), .ZN(
        n1906) );
  INVD1BWP12T U2137 ( .I(n1849), .ZN(mult_x_18_n432) );
  AOI22D1BWP12T U2138 ( .A1(b[5]), .A2(n2152), .B1(b[4]), .B2(n2151), .ZN(
        n1851) );
  AOI22D1BWP12T U2139 ( .A1(b[3]), .A2(n2155), .B1(n2140), .B2(n2153), .ZN(
        n1850) );
  ND2D1BWP12T U2140 ( .A1(n1851), .A2(n1850), .ZN(n1852) );
  MAOI22D0BWP12T U2141 ( .A1(n3701), .A2(n1852), .B1(n3701), .B2(n1852), .ZN(
        n1960) );
  NR2D1BWP12T U2142 ( .A1(n3170), .A2(n1853), .ZN(mult_x_18_n374) );
  INVD1BWP12T U2143 ( .I(n2153), .ZN(n1864) );
  OAI222D1BWP12T U2144 ( .A1(n3878), .A2(n1864), .B1(n1862), .B2(n3165), .C1(
        n1863), .C2(n3170), .ZN(n1973) );
  AOI21D1BWP12T U2145 ( .A1(a[23]), .A2(mult_x_18_n374), .B(n1973), .ZN(n1972)
         );
  NR2D1BWP12T U2146 ( .A1(n1972), .A2(n3701), .ZN(n1932) );
  AOI22D1BWP12T U2147 ( .A1(b[2]), .A2(n2152), .B1(b[1]), .B2(n2151), .ZN(
        n1855) );
  ND2D1BWP12T U2148 ( .A1(b[0]), .A2(n2155), .ZN(n1854) );
  OAI211D1BWP12T U2149 ( .A1(n2027), .A2(n1864), .B(n1855), .C(n1854), .ZN(
        n1931) );
  NR2D1BWP12T U2150 ( .A1(n1932), .A2(n1931), .ZN(n1930) );
  NR2D1BWP12T U2151 ( .A1(n1930), .A2(n3701), .ZN(n1859) );
  AOI22D1BWP12T U2152 ( .A1(b[2]), .A2(n2151), .B1(n2153), .B2(n2026), .ZN(
        n1857) );
  AOI22D1BWP12T U2153 ( .A1(b[3]), .A2(n2152), .B1(b[1]), .B2(n2155), .ZN(
        n1856) );
  ND2D1BWP12T U2154 ( .A1(n1857), .A2(n1856), .ZN(n1858) );
  NR2D1BWP12T U2155 ( .A1(n1859), .A2(n1858), .ZN(n1861) );
  MOAI22D0BWP12T U2156 ( .A1(n1859), .A2(n1858), .B1(n1859), .B2(n1858), .ZN(
        n1964) );
  ND2D1BWP12T U2157 ( .A1(b[0]), .A2(n1860), .ZN(n1963) );
  NR2D1BWP12T U2158 ( .A1(n1964), .A2(n1963), .ZN(n1962) );
  AOI21D1BWP12T U2159 ( .A1(n1861), .A2(a[23]), .B(n1962), .ZN(n1954) );
  NR2D1BWP12T U2160 ( .A1(n3219), .A2(n1862), .ZN(n1866) );
  OAI22D1BWP12T U2161 ( .A1(n2033), .A2(n1864), .B1(n2886), .B2(n1863), .ZN(
        n1865) );
  AOI211D1BWP12T U2162 ( .A1(n2155), .A2(b[2]), .B(n1866), .C(n1865), .ZN(
        n1867) );
  MAOI22D0BWP12T U2163 ( .A1(a[23]), .A2(n1867), .B1(a[23]), .B2(n1867), .ZN(
        n1953) );
  AOI222D1BWP12T U2164 ( .A1(b[1]), .A2(n2161), .B1(b[0]), .B2(n2160), .C1(
        n2162), .C2(n3881), .ZN(n1868) );
  OAI21D1BWP12T U2165 ( .A1(n3790), .A2(n1963), .B(n1868), .ZN(n1905) );
  OAI31D1BWP12T U2166 ( .A1(n1868), .A2(n1963), .A3(n3790), .B(n1905), .ZN(
        n1952) );
  ND2D1BWP12T U2167 ( .A1(a[26]), .A2(n1905), .ZN(n1871) );
  AOI22D1BWP12T U2168 ( .A1(b[1]), .A2(n2160), .B1(n2162), .B2(n1941), .ZN(
        n1870) );
  AOI22D1BWP12T U2169 ( .A1(b[2]), .A2(n2161), .B1(b[0]), .B2(n2164), .ZN(
        n1869) );
  ND2D1BWP12T U2170 ( .A1(n1870), .A2(n1869), .ZN(n1904) );
  MAOI22D0BWP12T U2171 ( .A1(n1871), .A2(n1904), .B1(n1871), .B2(n1904), .ZN(
        n1958) );
  INVD1BWP12T U2172 ( .I(n1872), .ZN(mult_x_18_n312) );
  ND2D1BWP12T U2173 ( .A1(a[5]), .A2(b[0]), .ZN(n1873) );
  NR2D1BWP12T U2174 ( .A1(n2025), .A2(n1873), .ZN(n2039) );
  OAI222D1BWP12T U2175 ( .A1(n3878), .A2(n1883), .B1(n1881), .B2(n3165), .C1(
        n1882), .C2(n3170), .ZN(n2038) );
  NR2D1BWP12T U2176 ( .A1(n2039), .A2(n2038), .ZN(n2037) );
  NR2D1BWP12T U2177 ( .A1(n2037), .A2(n3247), .ZN(n2042) );
  AOI22D1BWP12T U2178 ( .A1(b[1]), .A2(n2196), .B1(n2198), .B2(n1941), .ZN(
        n1875) );
  AOI22D1BWP12T U2179 ( .A1(b[2]), .A2(n2197), .B1(b[0]), .B2(n2200), .ZN(
        n1874) );
  ND2D1BWP12T U2180 ( .A1(n1875), .A2(n1874), .ZN(n2041) );
  NR2D1BWP12T U2181 ( .A1(n2042), .A2(n2041), .ZN(n2040) );
  NR2D1BWP12T U2182 ( .A1(n2040), .A2(n3247), .ZN(n1879) );
  AOI22D1BWP12T U2183 ( .A1(b[2]), .A2(n2196), .B1(n2198), .B2(n2026), .ZN(
        n1877) );
  AOI22D1BWP12T U2184 ( .A1(b[3]), .A2(n2197), .B1(b[1]), .B2(n2200), .ZN(
        n1876) );
  ND2D1BWP12T U2185 ( .A1(n1877), .A2(n1876), .ZN(n1878) );
  NR2D1BWP12T U2186 ( .A1(n1879), .A2(n1878), .ZN(n1880) );
  MOAI22D0BWP12T U2187 ( .A1(n1879), .A2(n1878), .B1(n1879), .B2(n1878), .ZN(
        n2046) );
  NR3D1BWP12T U2188 ( .A1(n3170), .A2(n2047), .A3(n2046), .ZN(n2048) );
  AOI21D1BWP12T U2189 ( .A1(n1880), .A2(a[5]), .B(n2048), .ZN(n2051) );
  NR2D1BWP12T U2190 ( .A1(n3219), .A2(n1881), .ZN(n1885) );
  OAI22D1BWP12T U2191 ( .A1(n2033), .A2(n1883), .B1(n2886), .B2(n1882), .ZN(
        n1884) );
  AOI211D1BWP12T U2192 ( .A1(n2200), .A2(b[2]), .B(n1885), .C(n1884), .ZN(
        n1886) );
  MAOI22D0BWP12T U2193 ( .A1(a[5]), .A2(n1886), .B1(a[5]), .B2(n1886), .ZN(
        n2050) );
  AOI222D1BWP12T U2194 ( .A1(b[1]), .A2(n2145), .B1(b[0]), .B2(n2144), .C1(
        n2146), .C2(n3881), .ZN(n1890) );
  NR2D1BWP12T U2195 ( .A1(n3321), .A2(n3170), .ZN(n1887) );
  ND2D1BWP12T U2196 ( .A1(n1888), .A2(n1887), .ZN(n1889) );
  ND2D1BWP12T U2197 ( .A1(n1890), .A2(n1889), .ZN(n1901) );
  OAI21D1BWP12T U2198 ( .A1(n1890), .A2(n1889), .B(n1901), .ZN(n2049) );
  ND2D1BWP12T U2199 ( .A1(a[8]), .A2(n1901), .ZN(n1893) );
  AOI22D1BWP12T U2200 ( .A1(b[1]), .A2(n2144), .B1(n2146), .B2(n1941), .ZN(
        n1892) );
  AOI22D1BWP12T U2201 ( .A1(b[2]), .A2(n2145), .B1(b[0]), .B2(n2148), .ZN(
        n1891) );
  ND2D1BWP12T U2202 ( .A1(n1892), .A2(n1891), .ZN(n1900) );
  MAOI22D0BWP12T U2203 ( .A1(n1893), .A2(n1900), .B1(n1893), .B2(n1900), .ZN(
        n2054) );
  AOI22D1BWP12T U2204 ( .A1(b[5]), .A2(n2197), .B1(b[4]), .B2(n2196), .ZN(
        n1895) );
  AOI22D1BWP12T U2205 ( .A1(b[3]), .A2(n2200), .B1(n2140), .B2(n2198), .ZN(
        n1894) );
  ND2D1BWP12T U2206 ( .A1(n1895), .A2(n1894), .ZN(n1896) );
  MAOI22D0BWP12T U2207 ( .A1(n3247), .A2(n1896), .B1(n3247), .B2(n1896), .ZN(
        n2053) );
  INVD1BWP12T U2208 ( .I(n1897), .ZN(mult_x_18_n465) );
  NR3D1BWP12T U2209 ( .A1(n3632), .A2(n1899), .A3(n1898), .ZN(mult_x_18_n383)
         );
  NR3D1BWP12T U2210 ( .A1(n3321), .A2(n1901), .A3(n1900), .ZN(mult_x_18_n467)
         );
  NR3D1BWP12T U2211 ( .A1(n3479), .A2(n1903), .A3(n1902), .ZN(mult_x_18_n434)
         );
  NR3D1BWP12T U2212 ( .A1(n3790), .A2(n1905), .A3(n1904), .ZN(mult_x_18_n314)
         );
  FA1D0BWP12T U2213 ( .A(n1908), .B(n1907), .CI(n1906), .CO(n1849), .S(n1909)
         );
  INVD1BWP12T U2214 ( .I(n1909), .ZN(mult_x_18_n433) );
  AOI21D1BWP12T U2215 ( .A1(n1912), .A2(n1911), .B(n1910), .ZN(mult_x_18_n447)
         );
  FA1D0BWP12T U2216 ( .A(n1915), .B(n1914), .CI(n1913), .CO(n1908), .S(n1916)
         );
  INVD1BWP12T U2217 ( .I(n1916), .ZN(mult_x_18_n440) );
  FA1D0BWP12T U2218 ( .A(n1919), .B(n1918), .CI(n1917), .CO(n1928), .S(n1920)
         );
  INVD1BWP12T U2219 ( .I(n1920), .ZN(mult_x_18_n402) );
  NR2D1BWP12T U2220 ( .A1(n3170), .A2(n1921), .ZN(mult_x_18_n464) );
  FA1D0BWP12T U2221 ( .A(n1924), .B(n1923), .CI(n1922), .CO(n1825), .S(n1925)
         );
  INVD1BWP12T U2222 ( .I(n1925), .ZN(mult_x_18_n382) );
  FA1D0BWP12T U2223 ( .A(n1928), .B(n1927), .CI(n1926), .CO(n1923), .S(n1929)
         );
  INVD1BWP12T U2224 ( .I(n1929), .ZN(mult_x_18_n392) );
  AOI21D1BWP12T U2225 ( .A1(n1932), .A2(n1931), .B(n1930), .ZN(mult_x_18_n352)
         );
  INVD1BWP12T U2226 ( .I(a[29]), .ZN(n3869) );
  INVD1BWP12T U2227 ( .I(a[28]), .ZN(n3851) );
  INVD1BWP12T U2228 ( .I(a[27]), .ZN(n3824) );
  OAI22D1BWP12T U2229 ( .A1(n3851), .A2(a[27]), .B1(n3824), .B2(a[28]), .ZN(
        n1935) );
  OAI22D1BWP12T U2230 ( .A1(n3824), .A2(a[26]), .B1(n3790), .B2(a[27]), .ZN(
        n1936) );
  INVD1BWP12T U2231 ( .I(n1936), .ZN(n1940) );
  AN2D1BWP12T U2232 ( .A1(n1935), .A2(n1940), .Z(n2137) );
  OAI22D1BWP12T U2233 ( .A1(n3869), .A2(n3851), .B1(a[28]), .B2(a[29]), .ZN(
        n1934) );
  NR2D1BWP12T U2234 ( .A1(n1934), .A2(n1940), .ZN(n2139) );
  AOI22D1BWP12T U2235 ( .A1(b[3]), .A2(n2137), .B1(n2139), .B2(n1933), .ZN(
        n1938) );
  AN2D1BWP12T U2236 ( .A1(n1934), .A2(n1936), .Z(n2138) );
  NR3D1BWP12T U2237 ( .A1(n1936), .A2(n1935), .A3(n1934), .ZN(n2141) );
  AOI22D1BWP12T U2238 ( .A1(b[4]), .A2(n2138), .B1(b[2]), .B2(n2141), .ZN(
        n1937) );
  ND2D1BWP12T U2239 ( .A1(n1938), .A2(n1937), .ZN(n1939) );
  MAOI22D0BWP12T U2240 ( .A1(n3869), .A2(n1939), .B1(n3869), .B2(n1939), .ZN(
        n2101) );
  NR2D1BWP12T U2241 ( .A1(n3170), .A2(n1940), .ZN(mult_x_18_n302) );
  AO222D1BWP12T U2242 ( .A1(b[1]), .A2(n2138), .B1(n2139), .B2(n2570), .C1(
        n2137), .C2(b[0]), .Z(n1971) );
  AOI21D1BWP12T U2243 ( .A1(a[29]), .A2(mult_x_18_n302), .B(n1971), .ZN(n1970)
         );
  NR2D1BWP12T U2244 ( .A1(n1970), .A2(n3869), .ZN(n1967) );
  AOI22D1BWP12T U2245 ( .A1(b[1]), .A2(n2137), .B1(n2139), .B2(n1941), .ZN(
        n1943) );
  AOI22D1BWP12T U2246 ( .A1(b[2]), .A2(n2138), .B1(b[0]), .B2(n2141), .ZN(
        n1942) );
  ND2D1BWP12T U2247 ( .A1(n1943), .A2(n1942), .ZN(n1966) );
  NR2D1BWP12T U2248 ( .A1(n1967), .A2(n1966), .ZN(n1965) );
  NR2D1BWP12T U2249 ( .A1(n1965), .A2(n3869), .ZN(n1947) );
  AOI22D1BWP12T U2250 ( .A1(b[2]), .A2(n2137), .B1(n2139), .B2(n2026), .ZN(
        n1945) );
  AOI22D1BWP12T U2251 ( .A1(b[3]), .A2(n2138), .B1(b[1]), .B2(n2141), .ZN(
        n1944) );
  ND2D1BWP12T U2252 ( .A1(n1945), .A2(n1944), .ZN(n1946) );
  NR2D1BWP12T U2253 ( .A1(n1947), .A2(n1946), .ZN(n1948) );
  INVD1BWP12T U2254 ( .I(a[30]), .ZN(n3932) );
  AOI22D1BWP12T U2255 ( .A1(a[30]), .A2(a[29]), .B1(n3869), .B2(n3932), .ZN(
        n2091) );
  ND2D1BWP12T U2256 ( .A1(b[0]), .A2(n2091), .ZN(n2123) );
  MOAI22D0BWP12T U2257 ( .A1(n1947), .A2(n1946), .B1(n1947), .B2(n1946), .ZN(
        n1957) );
  NR2D1BWP12T U2258 ( .A1(n2123), .A2(n1957), .ZN(n1956) );
  AOI21D1BWP12T U2259 ( .A1(n1948), .A2(a[29]), .B(n1956), .ZN(n2100) );
  INVD1BWP12T U2260 ( .I(a[31]), .ZN(n3194) );
  ND2D1BWP12T U2261 ( .A1(a[30]), .A2(a[29]), .ZN(n1949) );
  OAI32D1BWP12T U2262 ( .A1(n3194), .A2(a[30]), .A3(a[29]), .B1(a[31]), .B2(
        n1949), .ZN(n2090) );
  AOI22D1BWP12T U2263 ( .A1(b[1]), .A2(n2091), .B1(b[0]), .B2(n2090), .ZN(
        n2124) );
  NR2D1BWP12T U2264 ( .A1(n3194), .A2(n2123), .ZN(n1950) );
  MAOI22D0BWP12T U2265 ( .A1(n2124), .A2(n1950), .B1(n2124), .B2(n1950), .ZN(
        n2099) );
  INVD1BWP12T U2266 ( .I(n1951), .ZN(mult_x_18_n242) );
  FA1D0BWP12T U2267 ( .A(n1954), .B(n1953), .CI(n1952), .CO(n1959), .S(n1955)
         );
  INVD1BWP12T U2268 ( .I(n1955), .ZN(mult_x_18_n326) );
  AOI21D1BWP12T U2269 ( .A1(n2123), .A2(n1957), .B(n1956), .ZN(mult_x_18_n258)
         );
  FA1D0BWP12T U2270 ( .A(n1960), .B(n1959), .CI(n1958), .CO(n1872), .S(n1961)
         );
  INVD1BWP12T U2271 ( .I(n1961), .ZN(mult_x_18_n313) );
  AOI21D1BWP12T U2272 ( .A1(n1964), .A2(n1963), .B(n1962), .ZN(mult_x_18_n339)
         );
  AOI21D1BWP12T U2273 ( .A1(n1967), .A2(n1966), .B(n1965), .ZN(mult_x_18_n274)
         );
  AOI21D1BWP12T U2274 ( .A1(n1969), .A2(n1968), .B(n4006), .ZN(mult_x_18_n459)
         );
  AOI31D1BWP12T U2275 ( .A1(mult_x_18_n302), .A2(a[29]), .A3(n1971), .B(n1970), 
        .ZN(mult_x_18_n288) );
  AOI31D1BWP12T U2276 ( .A1(mult_x_18_n374), .A2(a[23]), .A3(n1973), .B(n1972), 
        .ZN(mult_x_18_n363) );
  INVD1BWP12T U2277 ( .I(b[31]), .ZN(n3193) );
  NR2D1BWP12T U2278 ( .A1(a[31]), .A2(n3193), .ZN(n3143) );
  INVD1BWP12T U2279 ( .I(op[2]), .ZN(n3627) );
  NR2D1BWP12T U2280 ( .A1(op[3]), .A2(n3627), .ZN(n3268) );
  INR2D1BWP12T U2281 ( .A1(op[1]), .B1(op[0]), .ZN(n2772) );
  ND2D1BWP12T U2282 ( .A1(n3268), .A2(n2772), .ZN(n3949) );
  INVD1BWP12T U2283 ( .I(op[0]), .ZN(n2288) );
  INR2D1BWP12T U2284 ( .A1(op[3]), .B1(op[2]), .ZN(n2228) );
  ND2D1BWP12T U2285 ( .A1(op[1]), .A2(n2228), .ZN(n2287) );
  INVD1BWP12T U2286 ( .I(n2287), .ZN(n3152) );
  ND2D1BWP12T U2287 ( .A1(n2288), .A2(n3152), .ZN(n3976) );
  ND2D1BWP12T U2288 ( .A1(n3949), .A2(n3976), .ZN(n2211) );
  NR2D1BWP12T U2289 ( .A1(op[1]), .A2(n2288), .ZN(n3102) );
  ND2D1BWP12T U2290 ( .A1(op[3]), .A2(op[2]), .ZN(n2927) );
  INVD1BWP12T U2291 ( .I(n2927), .ZN(n2771) );
  ND2D1BWP12T U2292 ( .A1(n3102), .A2(n2771), .ZN(n3958) );
  INVD1BWP12T U2293 ( .I(b[30]), .ZN(n3912) );
  INVD1BWP12T U2294 ( .I(a[1]), .ZN(n2470) );
  NR2D1BWP12T U2295 ( .A1(n2470), .A2(a[0]), .ZN(n2074) );
  INVD1BWP12T U2296 ( .I(n2074), .ZN(n2113) );
  INVD1BWP12T U2297 ( .I(a[2]), .ZN(n3961) );
  NR2D1BWP12T U2298 ( .A1(a[1]), .A2(a[0]), .ZN(n3174) );
  INVD1BWP12T U2299 ( .I(n3174), .ZN(n2087) );
  NR2D1BWP12T U2300 ( .A1(n3961), .A2(n2087), .ZN(n2112) );
  INVD1BWP12T U2301 ( .I(a[0]), .ZN(n3169) );
  AOI22D1BWP12T U2302 ( .A1(a[2]), .A2(n2470), .B1(a[1]), .B2(n3961), .ZN(
        n1976) );
  NR2D1BWP12T U2303 ( .A1(n3169), .A2(n1976), .ZN(n2085) );
  FA1D0BWP12T U2304 ( .A(b[27]), .B(b[28]), .CI(n1974), .CO(n2084), .S(n2081)
         );
  AOI22D1BWP12T U2305 ( .A1(b[29]), .A2(n2112), .B1(n2085), .B2(n1975), .ZN(
        n1978) );
  ND2D1BWP12T U2306 ( .A1(a[0]), .A2(n1976), .ZN(n2115) );
  INVD1BWP12T U2307 ( .I(n2115), .ZN(n2086) );
  ND2D1BWP12T U2308 ( .A1(b[31]), .A2(n2086), .ZN(n1977) );
  OAI211D1BWP12T U2309 ( .A1(n3912), .A2(n2113), .B(n1978), .C(n1977), .ZN(
        n1979) );
  MAOI22D0BWP12T U2310 ( .A1(a[2]), .A2(n1979), .B1(a[2]), .B2(n1979), .ZN(
        n2117) );
  FA1D0BWP12T U2311 ( .A(b[29]), .B(b[30]), .CI(n1980), .CO(n2110), .S(n1981)
         );
  AOI22D1BWP12T U2312 ( .A1(b[30]), .A2(n2086), .B1(n2085), .B2(n1981), .ZN(
        n1983) );
  AOI22D1BWP12T U2313 ( .A1(b[29]), .A2(n2074), .B1(b[28]), .B2(n2112), .ZN(
        n1982) );
  ND2D1BWP12T U2314 ( .A1(n1983), .A2(n1982), .ZN(n1984) );
  MAOI22D0BWP12T U2315 ( .A1(a[2]), .A2(n1984), .B1(a[2]), .B2(n1984), .ZN(
        n2782) );
  AOI222D1BWP12T U2316 ( .A1(b[27]), .A2(n2086), .B1(b[26]), .B2(n2074), .C1(
        n2085), .C2(n1985), .ZN(n1987) );
  INVD1BWP12T U2317 ( .I(b[25]), .ZN(n3757) );
  OAI211D1BWP12T U2318 ( .A1(n2087), .A2(n3757), .B(a[2]), .C(n1987), .ZN(
        n1986) );
  OAI21D1BWP12T U2319 ( .A1(n1987), .A2(a[2]), .B(n1986), .ZN(n2789) );
  AOI22D1BWP12T U2320 ( .A1(b[25]), .A2(n2086), .B1(n2085), .B2(n1988), .ZN(
        n1990) );
  AOI22D1BWP12T U2321 ( .A1(b[24]), .A2(n2074), .B1(b[23]), .B2(n2112), .ZN(
        n1989) );
  ND2D1BWP12T U2322 ( .A1(n1990), .A2(n1989), .ZN(n1991) );
  MAOI22D0BWP12T U2323 ( .A1(a[2]), .A2(n1991), .B1(a[2]), .B2(n1991), .ZN(
        n2793) );
  AOI22D1BWP12T U2324 ( .A1(b[23]), .A2(n2086), .B1(n2085), .B2(n2188), .ZN(
        n1993) );
  AOI22D1BWP12T U2325 ( .A1(b[22]), .A2(n2074), .B1(b[21]), .B2(n2112), .ZN(
        n1992) );
  ND2D1BWP12T U2326 ( .A1(n1993), .A2(n1992), .ZN(n1994) );
  MAOI22D0BWP12T U2327 ( .A1(a[2]), .A2(n1994), .B1(a[2]), .B2(n1994), .ZN(
        n2797) );
  INVD1BWP12T U2328 ( .I(n2085), .ZN(n2034) );
  AOI222D1BWP12T U2329 ( .A1(b[22]), .A2(n2086), .B1(b[21]), .B2(n2074), .C1(
        n2085), .C2(n1995), .ZN(n1997) );
  INVD1BWP12T U2330 ( .I(b[20]), .ZN(n3628) );
  OAI211D1BWP12T U2331 ( .A1(n2087), .A2(n3628), .B(a[2]), .C(n1997), .ZN(
        n1996) );
  OAI21D1BWP12T U2332 ( .A1(n1997), .A2(a[2]), .B(n1996), .ZN(n2799) );
  AOI22D1BWP12T U2333 ( .A1(b[21]), .A2(n2086), .B1(n2085), .B2(n1998), .ZN(
        n2000) );
  AOI22D1BWP12T U2334 ( .A1(b[20]), .A2(n2074), .B1(b[19]), .B2(n2112), .ZN(
        n1999) );
  ND2D1BWP12T U2335 ( .A1(n2000), .A2(n1999), .ZN(n2001) );
  MAOI22D0BWP12T U2336 ( .A1(a[2]), .A2(n2001), .B1(a[2]), .B2(n2001), .ZN(
        n2801) );
  AOI222D1BWP12T U2337 ( .A1(b[20]), .A2(n2086), .B1(b[19]), .B2(n2074), .C1(
        n2095), .C2(n2085), .ZN(n2003) );
  INVD1BWP12T U2338 ( .I(b[18]), .ZN(n2751) );
  OAI211D1BWP12T U2339 ( .A1(n2087), .A2(n2751), .B(a[2]), .C(n2003), .ZN(
        n2002) );
  OAI21D1BWP12T U2340 ( .A1(n2003), .A2(a[2]), .B(n2002), .ZN(n2803) );
  AOI22D1BWP12T U2341 ( .A1(b[19]), .A2(n2086), .B1(n2085), .B2(n2004), .ZN(
        n2006) );
  AOI22D1BWP12T U2342 ( .A1(b[18]), .A2(n2074), .B1(b[17]), .B2(n2112), .ZN(
        n2005) );
  ND2D1BWP12T U2343 ( .A1(n2006), .A2(n2005), .ZN(n2007) );
  MAOI22D0BWP12T U2344 ( .A1(a[2]), .A2(n2007), .B1(a[2]), .B2(n2007), .ZN(
        n2808) );
  AOI222D1BWP12T U2345 ( .A1(b[18]), .A2(n2086), .B1(b[17]), .B2(n2074), .C1(
        n2085), .C2(n2008), .ZN(n2010) );
  INVD1BWP12T U2346 ( .I(b[16]), .ZN(n2232) );
  OAI211D1BWP12T U2347 ( .A1(n2087), .A2(n2232), .B(a[2]), .C(n2010), .ZN(
        n2009) );
  OAI21D1BWP12T U2348 ( .A1(n2010), .A2(a[2]), .B(n2009), .ZN(n2810) );
  AOI222D1BWP12T U2349 ( .A1(b[17]), .A2(n2086), .B1(b[16]), .B2(n2074), .C1(
        n2085), .C2(n2181), .ZN(n2012) );
  INVD1BWP12T U2350 ( .I(b[15]), .ZN(n2231) );
  OAI211D1BWP12T U2351 ( .A1(n2087), .A2(n2231), .B(a[2]), .C(n2012), .ZN(
        n2011) );
  OAI21D1BWP12T U2352 ( .A1(n2012), .A2(a[2]), .B(n2011), .ZN(n2812) );
  AOI22D1BWP12T U2353 ( .A1(b[10]), .A2(n2086), .B1(n2085), .B2(n2013), .ZN(
        n2015) );
  AOI22D1BWP12T U2354 ( .A1(b[9]), .A2(n2074), .B1(b[8]), .B2(n2112), .ZN(
        n2014) );
  ND2D1BWP12T U2355 ( .A1(n2015), .A2(n2014), .ZN(n2016) );
  MAOI22D0BWP12T U2356 ( .A1(a[2]), .A2(n2016), .B1(a[2]), .B2(n2016), .ZN(
        n2826) );
  AOI22D1BWP12T U2357 ( .A1(b[9]), .A2(n2086), .B1(n2085), .B2(n2017), .ZN(
        n2019) );
  AOI22D1BWP12T U2358 ( .A1(b[8]), .A2(n2074), .B1(b[7]), .B2(n2112), .ZN(
        n2018) );
  ND2D1BWP12T U2359 ( .A1(n2019), .A2(n2018), .ZN(n2020) );
  MAOI22D0BWP12T U2360 ( .A1(a[2]), .A2(n2020), .B1(a[2]), .B2(n2020), .ZN(
        n2828) );
  AOI22D1BWP12T U2361 ( .A1(b[5]), .A2(n2086), .B1(n2085), .B2(n2140), .ZN(
        n2023) );
  AOI22D1BWP12T U2362 ( .A1(b[4]), .A2(n2074), .B1(b[3]), .B2(n2112), .ZN(
        n2022) );
  ND2D1BWP12T U2363 ( .A1(n2023), .A2(n2022), .ZN(n2024) );
  MAOI22D0BWP12T U2364 ( .A1(a[2]), .A2(n2024), .B1(a[2]), .B2(n2024), .ZN(
        n2836) );
  NR2D1BWP12T U2365 ( .A1(n3170), .A2(n2025), .ZN(n2780) );
  AO222D1BWP12T U2366 ( .A1(b[3]), .A2(n2086), .B1(b[2]), .B2(n2074), .C1(
        n2085), .C2(n2026), .Z(n2030) );
  AOI21D1BWP12T U2367 ( .A1(b[1]), .A2(n2112), .B(n2030), .ZN(n2031) );
  ND2D1BWP12T U2368 ( .A1(b[0]), .A2(a[0]), .ZN(n3147) );
  INVD1BWP12T U2369 ( .I(n3147), .ZN(n2474) );
  AOI22D1BWP12T U2370 ( .A1(b[1]), .A2(n2086), .B1(n2085), .B2(n3881), .ZN(
        n3172) );
  OAI31D1BWP12T U2371 ( .A1(a[0]), .A2(n2470), .A3(n3170), .B(n3172), .ZN(
        n3173) );
  NR2D1BWP12T U2372 ( .A1(n2474), .A2(n3173), .ZN(n3952) );
  ND2D1BWP12T U2373 ( .A1(b[1]), .A2(a[1]), .ZN(n3163) );
  NR2D1BWP12T U2374 ( .A1(a[0]), .A2(n3163), .ZN(n2029) );
  OAI22D1BWP12T U2375 ( .A1(n2652), .A2(n2115), .B1(n2034), .B2(n2027), .ZN(
        n2028) );
  AOI211D1BWP12T U2376 ( .A1(n2112), .A2(b[0]), .B(n2029), .C(n2028), .ZN(
        n3954) );
  ND2D1BWP12T U2377 ( .A1(n3952), .A2(n3954), .ZN(n2846) );
  INVD1BWP12T U2378 ( .I(n2846), .ZN(n2032) );
  AN2D1BWP12T U2379 ( .A1(n2031), .A2(n2032), .Z(n2778) );
  OAI32D1BWP12T U2380 ( .A1(n3961), .A2(n2032), .A3(n2031), .B1(a[2]), .B2(
        n2030), .ZN(n2777) );
  RCIAO21D0BWP12T U2381 ( .A1(n2780), .A2(n2778), .B(n2777), .ZN(n2839) );
  OAI222D1BWP12T U2382 ( .A1(n2113), .A2(n2886), .B1(n2034), .B2(n2033), .C1(
        n3219), .C2(n2115), .ZN(n2036) );
  ND2D1BWP12T U2383 ( .A1(a[2]), .A2(n2652), .ZN(n3941) );
  ND2D1BWP12T U2384 ( .A1(a[2]), .A2(n2087), .ZN(n3944) );
  ND2D1BWP12T U2385 ( .A1(n3941), .A2(n3944), .ZN(n2035) );
  MAOI22D0BWP12T U2386 ( .A1(n2036), .A2(a[2]), .B1(n2036), .B2(n2035), .ZN(
        n2838) );
  AOI21D1BWP12T U2387 ( .A1(n2039), .A2(n2038), .B(n2037), .ZN(n2837) );
  AOI21D1BWP12T U2388 ( .A1(n2042), .A2(n2041), .B(n2040), .ZN(n2834) );
  AOI222D1BWP12T U2389 ( .A1(b[6]), .A2(n2086), .B1(b[5]), .B2(n2074), .C1(
        n2085), .C2(n2043), .ZN(n2045) );
  OAI211D1BWP12T U2390 ( .A1(n2087), .A2(n3219), .B(a[2]), .C(n2045), .ZN(
        n2044) );
  OAI21D1BWP12T U2391 ( .A1(n2045), .A2(a[2]), .B(n2044), .ZN(n2832) );
  INVD1BWP12T U2392 ( .I(b[0]), .ZN(n2534) );
  OAI32D1BWP12T U2393 ( .A1(n2048), .A2(n2047), .A3(n2534), .B1(n2046), .B2(
        n2048), .ZN(n2831) );
  FA1D0BWP12T U2394 ( .A(n2051), .B(n2050), .CI(n2049), .CO(n2055), .S(n2052)
         );
  FA1D0BWP12T U2395 ( .A(n2055), .B(n2054), .CI(n2053), .CO(n1897), .S(n2056)
         );
  AOI222D1BWP12T U2396 ( .A1(b[11]), .A2(n2086), .B1(b[10]), .B2(n2074), .C1(
        n2085), .C2(n2154), .ZN(n2058) );
  INVD1BWP12T U2397 ( .I(b[9]), .ZN(n3341) );
  OAI211D1BWP12T U2398 ( .A1(n2087), .A2(n3341), .B(a[2]), .C(n2058), .ZN(
        n2057) );
  OAI21D1BWP12T U2399 ( .A1(n2058), .A2(a[2]), .B(n2057), .ZN(n2823) );
  AOI222D1BWP12T U2400 ( .A1(b[12]), .A2(n2086), .B1(b[11]), .B2(n2074), .C1(
        n2085), .C2(n2059), .ZN(n2061) );
  INVD1BWP12T U2401 ( .I(b[10]), .ZN(n3370) );
  OAI211D1BWP12T U2402 ( .A1(n2087), .A2(n3370), .B(a[2]), .C(n2061), .ZN(
        n2060) );
  OAI21D1BWP12T U2403 ( .A1(n2061), .A2(a[2]), .B(n2060), .ZN(n2821) );
  AOI222D1BWP12T U2404 ( .A1(b[13]), .A2(n2086), .B1(b[12]), .B2(n2074), .C1(
        n2085), .C2(n2062), .ZN(n2064) );
  INVD1BWP12T U2405 ( .I(b[11]), .ZN(n2759) );
  OAI211D1BWP12T U2406 ( .A1(n2087), .A2(n2759), .B(a[2]), .C(n2064), .ZN(
        n2063) );
  OAI21D1BWP12T U2407 ( .A1(n2064), .A2(a[2]), .B(n2063), .ZN(n2819) );
  AOI222D1BWP12T U2408 ( .A1(b[14]), .A2(n2086), .B1(b[13]), .B2(n2074), .C1(
        n2085), .C2(n2174), .ZN(n2066) );
  INVD1BWP12T U2409 ( .I(b[12]), .ZN(n3416) );
  OAI211D1BWP12T U2410 ( .A1(n2087), .A2(n3416), .B(a[2]), .C(n2066), .ZN(
        n2065) );
  OAI21D1BWP12T U2411 ( .A1(n2066), .A2(a[2]), .B(n2065), .ZN(n2817) );
  AOI222D1BWP12T U2412 ( .A1(b[15]), .A2(n2086), .B1(b[14]), .B2(n2074), .C1(
        n2085), .C2(n2067), .ZN(n2069) );
  INVD1BWP12T U2413 ( .I(b[13]), .ZN(n2371) );
  OAI211D1BWP12T U2414 ( .A1(n2087), .A2(n2371), .B(a[2]), .C(n2069), .ZN(
        n2068) );
  OAI21D1BWP12T U2415 ( .A1(n2069), .A2(a[2]), .B(n2068), .ZN(n2815) );
  AOI222D1BWP12T U2416 ( .A1(b[16]), .A2(n2086), .B1(b[15]), .B2(n2074), .C1(
        n2085), .C2(n2070), .ZN(n2072) );
  INVD1BWP12T U2417 ( .I(b[14]), .ZN(n3465) );
  OAI211D1BWP12T U2418 ( .A1(n2087), .A2(n3465), .B(a[2]), .C(n2072), .ZN(
        n2071) );
  OAI21D1BWP12T U2419 ( .A1(n2072), .A2(a[2]), .B(n2071), .ZN(n2813) );
  AOI22D1BWP12T U2420 ( .A1(b[24]), .A2(n2086), .B1(n2085), .B2(n2073), .ZN(
        n2076) );
  AOI22D1BWP12T U2421 ( .A1(b[22]), .A2(n2112), .B1(b[23]), .B2(n2074), .ZN(
        n2075) );
  ND2D1BWP12T U2422 ( .A1(n2076), .A2(n2075), .ZN(n2077) );
  MAOI22D0BWP12T U2423 ( .A1(a[2]), .A2(n2077), .B1(a[2]), .B2(n2077), .ZN(
        n2794) );
  AOI22D1BWP12T U2424 ( .A1(b[26]), .A2(n2086), .B1(n2085), .B2(n2147), .ZN(
        n2079) );
  AOI22D1BWP12T U2425 ( .A1(b[25]), .A2(n2074), .B1(b[24]), .B2(n2112), .ZN(
        n2078) );
  ND2D1BWP12T U2426 ( .A1(n2079), .A2(n2078), .ZN(n2080) );
  MAOI22D0BWP12T U2427 ( .A1(a[2]), .A2(n2080), .B1(a[2]), .B2(n2080), .ZN(
        n2790) );
  AOI222D1BWP12T U2428 ( .A1(b[28]), .A2(n2086), .B1(b[27]), .B2(n2074), .C1(
        n2085), .C2(n2081), .ZN(n2083) );
  INVD1BWP12T U2429 ( .I(b[26]), .ZN(n2360) );
  OAI211D1BWP12T U2430 ( .A1(n2087), .A2(n2360), .B(a[2]), .C(n2083), .ZN(
        n2082) );
  OAI21D1BWP12T U2431 ( .A1(n2083), .A2(a[2]), .B(n2082), .ZN(n2785) );
  FA1D0BWP12T U2432 ( .A(b[28]), .B(b[29]), .CI(n2084), .CO(n1980), .S(n2199)
         );
  AOI222D1BWP12T U2433 ( .A1(b[29]), .A2(n2086), .B1(b[28]), .B2(n2074), .C1(
        n2085), .C2(n2199), .ZN(n2089) );
  INVD1BWP12T U2434 ( .I(b[27]), .ZN(n2361) );
  OAI211D1BWP12T U2435 ( .A1(n2087), .A2(n2361), .B(a[2]), .C(n2089), .ZN(
        n2088) );
  OAI21D1BWP12T U2436 ( .A1(n2089), .A2(a[2]), .B(n2088), .ZN(n2783) );
  INVD1BWP12T U2437 ( .I(n2787), .ZN(n2227) );
  NR2D1BWP12T U2438 ( .A1(n3958), .A2(n2227), .ZN(n3195) );
  AOI22D1BWP12T U2439 ( .A1(a[29]), .A2(a[26]), .B1(n3790), .B2(n3869), .ZN(
        n2109) );
  AOI22D1BWP12T U2440 ( .A1(b[2]), .A2(n2091), .B1(b[1]), .B2(n2090), .ZN(
        n2107) );
  AOI22D1BWP12T U2441 ( .A1(b[20]), .A2(n2093), .B1(b[19]), .B2(n2092), .ZN(
        n2098) );
  AOI22D1BWP12T U2442 ( .A1(b[18]), .A2(n2096), .B1(n2095), .B2(n2094), .ZN(
        n2097) );
  ND2D1BWP12T U2443 ( .A1(n2098), .A2(n2097), .ZN(n2105) );
  FA1D0BWP12T U2444 ( .A(n2101), .B(n2100), .CI(n2099), .CO(n2103), .S(n1951)
         );
  AOI22D1BWP12T U2445 ( .A1(a[11]), .A2(n3961), .B1(a[2]), .B2(n4005), .ZN(
        n2102) );
  MAOI22D0BWP12T U2446 ( .A1(n2103), .A2(n2102), .B1(n2103), .B2(n2102), .ZN(
        n2104) );
  MAOI22D0BWP12T U2447 ( .A1(n2105), .A2(n2104), .B1(n2105), .B2(n2104), .ZN(
        n2106) );
  MAOI22D0BWP12T U2448 ( .A1(n2107), .A2(n2106), .B1(n2107), .B2(n2106), .ZN(
        n2108) );
  MAOI22D0BWP12T U2449 ( .A1(n2109), .A2(n2108), .B1(n2109), .B2(n2108), .ZN(
        n2210) );
  FA1D0BWP12T U2450 ( .A(b[30]), .B(b[31]), .CI(n2110), .CO(n2111), .S(n1975)
         );
  AOI22D1BWP12T U2451 ( .A1(b[30]), .A2(n2112), .B1(n2111), .B2(n2085), .ZN(
        n2114) );
  AOI32D1BWP12T U2452 ( .A1(n2115), .A2(n2114), .A3(n2113), .B1(n3193), .B2(
        n2114), .ZN(n2136) );
  AOI22D1BWP12T U2453 ( .A1(a[8]), .A2(a[5]), .B1(n3247), .B2(n3321), .ZN(
        n2122) );
  AOI22D1BWP12T U2454 ( .A1(a[17]), .A2(a[14]), .B1(n3479), .B2(n3565), .ZN(
        n2120) );
  FA1D0BWP12T U2455 ( .A(mult_x_18_n231), .B(n2117), .CI(n2116), .CO(n2118), 
        .S(n2787) );
  MAOI22D0BWP12T U2456 ( .A1(mult_x_18_n239), .A2(n2118), .B1(mult_x_18_n239), 
        .B2(n2118), .ZN(n2119) );
  MAOI22D0BWP12T U2457 ( .A1(n2120), .A2(n2119), .B1(n2120), .B2(n2119), .ZN(
        n2121) );
  MAOI22D0BWP12T U2458 ( .A1(n2122), .A2(n2121), .B1(n2122), .B2(n2121), .ZN(
        n2126) );
  XOR3D1BWP12T U2459 ( .A1(n3632), .A2(n2126), .A3(n2125), .Z(n2134) );
  MAOI22D0BWP12T U2460 ( .A1(a[23]), .A2(mult_x_18_n230), .B1(a[23]), .B2(
        mult_x_18_n230), .ZN(n2132) );
  MAOI22D0BWP12T U2461 ( .A1(mult_x_18_n235), .A2(mult_x_18_n229), .B1(
        mult_x_18_n235), .B2(mult_x_18_n229), .ZN(n2130) );
  MAOI22D0BWP12T U2462 ( .A1(mult_x_18_n233), .A2(mult_x_18_n232), .B1(
        mult_x_18_n233), .B2(mult_x_18_n232), .ZN(n2128) );
  MOAI22D0BWP12T U2463 ( .A1(mult_x_18_n236), .A2(mult_x_18_n238), .B1(
        mult_x_18_n236), .B2(mult_x_18_n238), .ZN(n2127) );
  MAOI22D0BWP12T U2464 ( .A1(n2128), .A2(n2127), .B1(n2128), .B2(n2127), .ZN(
        n2129) );
  MAOI22D0BWP12T U2465 ( .A1(n2130), .A2(n2129), .B1(n2130), .B2(n2129), .ZN(
        n2131) );
  MAOI22D0BWP12T U2466 ( .A1(n2132), .A2(n2131), .B1(n2132), .B2(n2131), .ZN(
        n2133) );
  MAOI22D0BWP12T U2467 ( .A1(n2134), .A2(n2133), .B1(n2134), .B2(n2133), .ZN(
        n2135) );
  MAOI22D0BWP12T U2468 ( .A1(n2136), .A2(n2135), .B1(n2136), .B2(n2135), .ZN(
        n2208) );
  AOI22D1BWP12T U2469 ( .A1(b[5]), .A2(n2138), .B1(b[4]), .B2(n2137), .ZN(
        n2143) );
  AOI22D1BWP12T U2470 ( .A1(b[3]), .A2(n2141), .B1(n2140), .B2(n2139), .ZN(
        n2142) );
  ND2D1BWP12T U2471 ( .A1(n2143), .A2(n2142), .ZN(n2170) );
  AOI22D1BWP12T U2472 ( .A1(b[26]), .A2(n2145), .B1(b[25]), .B2(n2144), .ZN(
        n2150) );
  AOI22D1BWP12T U2473 ( .A1(b[24]), .A2(n2148), .B1(n2147), .B2(n2146), .ZN(
        n2149) );
  ND2D1BWP12T U2474 ( .A1(n2150), .A2(n2149), .ZN(n2159) );
  AOI22D1BWP12T U2475 ( .A1(b[11]), .A2(n2152), .B1(b[10]), .B2(n2151), .ZN(
        n2157) );
  AOI22D1BWP12T U2476 ( .A1(b[9]), .A2(n2155), .B1(n2154), .B2(n2153), .ZN(
        n2156) );
  ND2D1BWP12T U2477 ( .A1(n2157), .A2(n2156), .ZN(n2158) );
  MAOI22D0BWP12T U2478 ( .A1(n2159), .A2(n2158), .B1(n2159), .B2(n2158), .ZN(
        n2168) );
  AOI22D1BWP12T U2479 ( .A1(b[8]), .A2(n2161), .B1(b[7]), .B2(n2160), .ZN(
        n2166) );
  AOI22D1BWP12T U2480 ( .A1(b[6]), .A2(n2164), .B1(n2163), .B2(n2162), .ZN(
        n2165) );
  ND2D1BWP12T U2481 ( .A1(n2166), .A2(n2165), .ZN(n2167) );
  MAOI22D0BWP12T U2482 ( .A1(n2168), .A2(n2167), .B1(n2168), .B2(n2167), .ZN(
        n2169) );
  MAOI22D0BWP12T U2483 ( .A1(n2170), .A2(n2169), .B1(n2170), .B2(n2169), .ZN(
        n2206) );
  AOI22D1BWP12T U2484 ( .A1(b[14]), .A2(n2172), .B1(b[13]), .B2(n2171), .ZN(
        n2177) );
  AOI22D1BWP12T U2485 ( .A1(b[12]), .A2(n2175), .B1(n2174), .B2(n2173), .ZN(
        n2176) );
  ND2D1BWP12T U2486 ( .A1(n2177), .A2(n2176), .ZN(n2195) );
  AOI22D1BWP12T U2487 ( .A1(b[17]), .A2(n2179), .B1(b[16]), .B2(n2178), .ZN(
        n2184) );
  AOI22D1BWP12T U2488 ( .A1(b[15]), .A2(n2182), .B1(n2181), .B2(n2180), .ZN(
        n2183) );
  ND2D1BWP12T U2489 ( .A1(n2184), .A2(n2183), .ZN(n2193) );
  AOI22D1BWP12T U2490 ( .A1(b[22]), .A2(n2186), .B1(b[23]), .B2(n2185), .ZN(
        n2191) );
  AOI22D1BWP12T U2491 ( .A1(b[21]), .A2(n2189), .B1(n2188), .B2(n2187), .ZN(
        n2190) );
  ND2D1BWP12T U2492 ( .A1(n2191), .A2(n2190), .ZN(n2192) );
  MOAI22D0BWP12T U2493 ( .A1(n2193), .A2(n2192), .B1(n2193), .B2(n2192), .ZN(
        n2194) );
  MAOI22D0BWP12T U2494 ( .A1(n2195), .A2(n2194), .B1(n2195), .B2(n2194), .ZN(
        n2204) );
  AOI22D1BWP12T U2495 ( .A1(b[29]), .A2(n2197), .B1(b[28]), .B2(n2196), .ZN(
        n2202) );
  AOI22D1BWP12T U2496 ( .A1(b[27]), .A2(n2200), .B1(n2199), .B2(n2198), .ZN(
        n2201) );
  ND2D1BWP12T U2497 ( .A1(n2202), .A2(n2201), .ZN(n2203) );
  MAOI22D0BWP12T U2498 ( .A1(n2204), .A2(n2203), .B1(n2204), .B2(n2203), .ZN(
        n2205) );
  MAOI22D0BWP12T U2499 ( .A1(n2206), .A2(n2205), .B1(n2206), .B2(n2205), .ZN(
        n2207) );
  MAOI22D0BWP12T U2500 ( .A1(n2208), .A2(n2207), .B1(n2208), .B2(n2207), .ZN(
        n2209) );
  MAOI22D0BWP12T U2501 ( .A1(n2210), .A2(n2209), .B1(n2210), .B2(n2209), .ZN(
        n2212) );
  AOI22D1BWP12T U2502 ( .A1(n3143), .A2(n2211), .B1(n3195), .B2(n2212), .ZN(
        n2230) );
  NR2D1BWP12T U2503 ( .A1(n2212), .A2(n3958), .ZN(n3139) );
  NR2D1BWP12T U2504 ( .A1(n3194), .A2(b[31]), .ZN(n2773) );
  INVD1BWP12T U2505 ( .I(n2773), .ZN(n2226) );
  ND2D1BWP12T U2506 ( .A1(n3851), .A2(b[28]), .ZN(n2756) );
  INVD1BWP12T U2507 ( .I(n2756), .ZN(n3842) );
  NR2D1BWP12T U2508 ( .A1(a[26]), .A2(n2360), .ZN(n2753) );
  INVD1BWP12T U2509 ( .I(b[22]), .ZN(n2359) );
  NR2D1BWP12T U2510 ( .A1(a[22]), .A2(n2359), .ZN(n3678) );
  INVD1BWP12T U2511 ( .I(b[21]), .ZN(n2774) );
  OAI22D1BWP12T U2512 ( .A1(n2774), .A2(a[21]), .B1(n3628), .B2(a[20]), .ZN(
        n2764) );
  INVD1BWP12T U2513 ( .I(n2764), .ZN(n2213) );
  OAI22D1BWP12T U2514 ( .A1(n3578), .A2(b[18]), .B1(n3565), .B2(b[17]), .ZN(
        n2223) );
  INVD1BWP12T U2515 ( .I(n2223), .ZN(n2741) );
  INVD1BWP12T U2516 ( .I(b[17]), .ZN(n3544) );
  NR2D1BWP12T U2517 ( .A1(n3544), .A2(a[17]), .ZN(n2752) );
  NR2D1BWP12T U2518 ( .A1(a[16]), .A2(n2232), .ZN(n3522) );
  NR2D1BWP12T U2519 ( .A1(b[14]), .A2(n3479), .ZN(n3469) );
  NR2D1BWP12T U2520 ( .A1(b[13]), .A2(n3446), .ZN(n3443) );
  NR2D1BWP12T U2521 ( .A1(n3469), .A2(n3443), .ZN(n2742) );
  NR2D1BWP12T U2522 ( .A1(n2371), .A2(a[13]), .ZN(n3444) );
  ND2D1BWP12T U2523 ( .A1(n3341), .A2(a[9]), .ZN(n3343) );
  OAI21D1BWP12T U2524 ( .A1(n3380), .A2(b[10]), .B(n3343), .ZN(n2221) );
  INVD1BWP12T U2525 ( .I(n2221), .ZN(n2743) );
  NR2D1BWP12T U2526 ( .A1(n3341), .A2(a[9]), .ZN(n2757) );
  OAI22D1BWP12T U2527 ( .A1(n3321), .A2(b[8]), .B1(n3292), .B2(b[7]), .ZN(
        n2220) );
  INVD1BWP12T U2528 ( .I(n2220), .ZN(n2744) );
  INVD1BWP12T U2529 ( .I(b[7]), .ZN(n3291) );
  NR2D1BWP12T U2530 ( .A1(n3291), .A2(a[7]), .ZN(n3296) );
  INVD1BWP12T U2531 ( .I(b[6]), .ZN(n3277) );
  NR2D1BWP12T U2532 ( .A1(b[5]), .A2(n3247), .ZN(n2982) );
  AOI21D1BWP12T U2533 ( .A1(a[6]), .A2(n3277), .B(n2982), .ZN(n2745) );
  OAI22D1BWP12T U2534 ( .A1(n3218), .A2(b[4]), .B1(n2471), .B2(b[3]), .ZN(
        n2217) );
  INVD1BWP12T U2535 ( .I(n2217), .ZN(n2746) );
  ND2D1BWP12T U2536 ( .A1(b[3]), .A2(n2471), .ZN(n4000) );
  ND2D1BWP12T U2537 ( .A1(n3961), .A2(b[2]), .ZN(n2334) );
  ND2D1BWP12T U2538 ( .A1(n3941), .A2(n2334), .ZN(n3107) );
  INVD1BWP12T U2539 ( .I(n3107), .ZN(n2974) );
  INVD1BWP12T U2540 ( .I(b[1]), .ZN(n2593) );
  ND2D1BWP12T U2541 ( .A1(a[1]), .A2(n2593), .ZN(n2736) );
  NR2D1BWP12T U2542 ( .A1(b[1]), .A2(a[1]), .ZN(n3168) );
  INVD1BWP12T U2543 ( .I(n3168), .ZN(n2413) );
  ND2D1BWP12T U2544 ( .A1(n3163), .A2(n2413), .ZN(n2976) );
  ND2D1BWP12T U2545 ( .A1(n3169), .A2(b[0]), .ZN(n2769) );
  ND2D1BWP12T U2546 ( .A1(a[0]), .A2(n2534), .ZN(n3155) );
  IOA21D1BWP12T U2547 ( .A1(n2769), .A2(c_in), .B(n3155), .ZN(n2977) );
  ND2D1BWP12T U2548 ( .A1(n2976), .A2(n2977), .ZN(n2975) );
  ND2D1BWP12T U2549 ( .A1(n2736), .A2(n2975), .ZN(n2973) );
  ND2D1BWP12T U2550 ( .A1(n2974), .A2(n2973), .ZN(n2972) );
  ND2D1BWP12T U2551 ( .A1(n3941), .A2(n2972), .ZN(n2967) );
  ND2D1BWP12T U2552 ( .A1(n4000), .A2(n2967), .ZN(n2969) );
  AOI22D1BWP12T U2553 ( .A1(n2746), .A2(n2969), .B1(b[4]), .B2(n3218), .ZN(
        n2971) );
  ND2D1BWP12T U2554 ( .A1(b[5]), .A2(n3247), .ZN(n3240) );
  ND2D1BWP12T U2555 ( .A1(n2971), .A2(n3240), .ZN(n2983) );
  NR2D1BWP12T U2556 ( .A1(a[6]), .A2(n3277), .ZN(n3271) );
  AOI21D1BWP12T U2557 ( .A1(n2745), .A2(n2983), .B(n3271), .ZN(n2966) );
  IND2D1BWP12T U2558 ( .A1(n3296), .B1(n2966), .ZN(n2980) );
  ND2D1BWP12T U2559 ( .A1(n3321), .A2(b[8]), .ZN(n2219) );
  INVD1BWP12T U2560 ( .I(n2219), .ZN(n3328) );
  AOI21D1BWP12T U2561 ( .A1(n2744), .A2(n2980), .B(n3328), .ZN(n2965) );
  IND2D1BWP12T U2562 ( .A1(n2757), .B1(n2965), .ZN(n2962) );
  AOI22D1BWP12T U2563 ( .A1(n2743), .A2(n2962), .B1(b[10]), .B2(n3380), .ZN(
        n2964) );
  MAOI222D1BWP12T U2564 ( .A(a[11]), .B(n2964), .C(n2759), .ZN(n2961) );
  MAOI222D1BWP12T U2565 ( .A(b[12]), .B(n3428), .C(n2961), .ZN(n2960) );
  IND2D1BWP12T U2566 ( .A1(n3444), .B1(n2960), .ZN(n2987) );
  AOI22D1BWP12T U2567 ( .A1(n2742), .A2(n2987), .B1(b[14]), .B2(n3479), .ZN(
        n2959) );
  MAOI222D1BWP12T U2568 ( .A(a[15]), .B(n2959), .C(n2231), .ZN(n2958) );
  ND2D1BWP12T U2569 ( .A1(a[16]), .A2(n2232), .ZN(n3523) );
  OAI21D1BWP12T U2570 ( .A1(n3522), .A2(n2958), .B(n3523), .ZN(n2957) );
  IND2D1BWP12T U2571 ( .A1(n2752), .B1(n2957), .ZN(n2993) );
  AOI22D1BWP12T U2572 ( .A1(n2741), .A2(n2993), .B1(b[18]), .B2(n3578), .ZN(
        n2956) );
  INVD1BWP12T U2573 ( .I(b[19]), .ZN(n3598) );
  MAOI222D1BWP12T U2574 ( .A(a[19]), .B(n2956), .C(n3598), .ZN(n2991) );
  ND2D1BWP12T U2575 ( .A1(a[20]), .A2(n3628), .ZN(n2739) );
  ND2D1BWP12T U2576 ( .A1(n2991), .A2(n2739), .ZN(n2954) );
  AOI22D1BWP12T U2577 ( .A1(n2213), .A2(n2954), .B1(a[21]), .B2(n2774), .ZN(
        n2952) );
  NR2D1BWP12T U2578 ( .A1(n3678), .A2(n2952), .ZN(n2950) );
  INVD1BWP12T U2579 ( .I(b[23]), .ZN(n3697) );
  ND2D1BWP12T U2580 ( .A1(a[23]), .A2(n3697), .ZN(n3699) );
  ND2D1BWP12T U2581 ( .A1(a[22]), .A2(n2359), .ZN(n3675) );
  ND2D1BWP12T U2582 ( .A1(n3699), .A2(n3675), .ZN(n2216) );
  NR2D1BWP12T U2583 ( .A1(n2950), .A2(n2216), .ZN(n2948) );
  AOI22D1BWP12T U2584 ( .A1(n2518), .A2(b[24]), .B1(n3701), .B2(b[23]), .ZN(
        n2224) );
  INVD1BWP12T U2585 ( .I(n2224), .ZN(n2765) );
  OAI22D1BWP12T U2586 ( .A1(n2948), .A2(n2765), .B1(b[24]), .B2(n2518), .ZN(
        n2997) );
  MAOI222D1BWP12T U2587 ( .A(a[25]), .B(n3757), .C(n2997), .ZN(n2946) );
  NR2D1BWP12T U2588 ( .A1(n2753), .A2(n2946), .ZN(n2943) );
  ND2D1BWP12T U2589 ( .A1(a[27]), .A2(n2361), .ZN(n3821) );
  ND2D1BWP12T U2590 ( .A1(a[26]), .A2(n2360), .ZN(n3787) );
  ND2D1BWP12T U2591 ( .A1(n3821), .A2(n3787), .ZN(n2215) );
  OAI22D1BWP12T U2592 ( .A1(n2943), .A2(n2215), .B1(a[27]), .B2(n2361), .ZN(
        n2945) );
  NR2D1BWP12T U2593 ( .A1(n3842), .A2(n2945), .ZN(n2941) );
  INVD1BWP12T U2594 ( .I(b[29]), .ZN(n2363) );
  ND2D1BWP12T U2595 ( .A1(a[29]), .A2(n2363), .ZN(n3865) );
  NR2D1BWP12T U2596 ( .A1(n3851), .A2(b[28]), .ZN(n3841) );
  INVD1BWP12T U2597 ( .I(n3841), .ZN(n2304) );
  ND2D1BWP12T U2598 ( .A1(n3865), .A2(n2304), .ZN(n2214) );
  NR2D1BWP12T U2599 ( .A1(n2363), .A2(a[29]), .ZN(n2770) );
  INVD1BWP12T U2600 ( .I(n2770), .ZN(n3864) );
  OAI21D1BWP12T U2601 ( .A1(n2941), .A2(n2214), .B(n3864), .ZN(n2940) );
  MAOI222D1BWP12T U2602 ( .A(b[30]), .B(n3932), .C(n2940), .ZN(n2939) );
  AOI21D1BWP12T U2603 ( .A1(n2226), .A2(n2939), .B(n3949), .ZN(n2225) );
  INVD1BWP12T U2604 ( .I(n2214), .ZN(n2775) );
  INVD1BWP12T U2605 ( .I(n2215), .ZN(n2776) );
  INVD1BWP12T U2606 ( .I(n2216), .ZN(n2740) );
  ND2D1BWP12T U2607 ( .A1(a[15]), .A2(n2231), .ZN(n3491) );
  INVD1BWP12T U2608 ( .I(n3240), .ZN(n2768) );
  NR2D1BWP12T U2609 ( .A1(a[1]), .A2(n3165), .ZN(n2766) );
  INVD1BWP12T U2610 ( .I(n2976), .ZN(n3105) );
  NR2D1BWP12T U2611 ( .A1(n3105), .A2(n2769), .ZN(n2339) );
  NR2D1BWP12T U2612 ( .A1(n2766), .A2(n2339), .ZN(n2338) );
  NR2D1BWP12T U2613 ( .A1(n2338), .A2(n3107), .ZN(n2337) );
  ND2D1BWP12T U2614 ( .A1(n4000), .A2(n2334), .ZN(n2763) );
  NR2D1BWP12T U2615 ( .A1(n2337), .A2(n2763), .ZN(n2331) );
  OAI22D1BWP12T U2616 ( .A1(a[4]), .A2(n3219), .B1(n2331), .B2(n2217), .ZN(
        n2333) );
  NR2D1BWP12T U2617 ( .A1(n2768), .A2(n2333), .ZN(n2329) );
  INVD1BWP12T U2618 ( .I(n2329), .ZN(n2218) );
  AO21D1BWP12T U2619 ( .A1(n2218), .A2(n2745), .B(n3271), .Z(n2328) );
  NR2D1BWP12T U2620 ( .A1(n3296), .A2(n2328), .ZN(n2341) );
  OAI21D1BWP12T U2621 ( .A1(n2341), .A2(n2220), .B(n2219), .ZN(n2327) );
  NR2D1BWP12T U2622 ( .A1(n2757), .A2(n2327), .ZN(n2323) );
  OAI22D1BWP12T U2623 ( .A1(a[10]), .A2(n3370), .B1(n2323), .B2(n2221), .ZN(
        n2325) );
  MAOI222D1BWP12T U2624 ( .A(b[11]), .B(n4005), .C(n2325), .ZN(n2326) );
  MAOI222D1BWP12T U2625 ( .A(a[12]), .B(n2326), .C(n3416), .ZN(n2345) );
  NR2D1BWP12T U2626 ( .A1(n3444), .A2(n2345), .ZN(n2346) );
  INVD1BWP12T U2627 ( .I(n2742), .ZN(n2222) );
  OAI22D1BWP12T U2628 ( .A1(a[14]), .A2(n3465), .B1(n2346), .B2(n2222), .ZN(
        n2322) );
  NR2D1BWP12T U2629 ( .A1(a[15]), .A2(n2231), .ZN(n3494) );
  AOI21D1BWP12T U2630 ( .A1(n3491), .A2(n2322), .B(n3494), .ZN(n2321) );
  MAOI222D1BWP12T U2631 ( .A(a[16]), .B(n2321), .C(n2232), .ZN(n2320) );
  NR2D1BWP12T U2632 ( .A1(n2752), .A2(n2320), .ZN(n2318) );
  OAI22D1BWP12T U2633 ( .A1(a[18]), .A2(n2751), .B1(n2318), .B2(n2223), .ZN(
        n2317) );
  MAOI222D1BWP12T U2634 ( .A(b[19]), .B(n3618), .C(n2317), .ZN(n2316) );
  INR2D1BWP12T U2635 ( .A1(n2739), .B1(n2316), .ZN(n2314) );
  OAI22D1BWP12T U2636 ( .A1(b[21]), .A2(n3685), .B1(n2314), .B2(n2764), .ZN(
        n2309) );
  IND2D1BWP12T U2637 ( .A1(n3678), .B1(n2309), .ZN(n2310) );
  ND2D1BWP12T U2638 ( .A1(n2740), .A2(n2310), .ZN(n2312) );
  INVD1BWP12T U2639 ( .I(b[24]), .ZN(n3725) );
  AOI22D1BWP12T U2640 ( .A1(n2224), .A2(n2312), .B1(a[24]), .B2(n3725), .ZN(
        n2354) );
  MAOI222D1BWP12T U2641 ( .A(b[25]), .B(n2354), .C(n3768), .ZN(n2308) );
  IND2D1BWP12T U2642 ( .A1(n2753), .B1(n2308), .ZN(n2352) );
  AOI22D1BWP12T U2643 ( .A1(n2776), .A2(n2352), .B1(b[27]), .B2(n3824), .ZN(
        n2307) );
  ND2D1BWP12T U2644 ( .A1(n2307), .A2(n2756), .ZN(n2303) );
  AOI21D1BWP12T U2645 ( .A1(n2775), .A2(n2303), .B(n2770), .ZN(n2306) );
  MAOI222D1BWP12T U2646 ( .A(a[30]), .B(n2306), .C(n3912), .ZN(n2302) );
  INVD1BWP12T U2647 ( .I(n3976), .ZN(n3926) );
  OAI32D1BWP12T U2648 ( .A1(n2225), .A2(n2773), .A3(n2302), .B1(n3926), .B2(
        n2225), .ZN(n3142) );
  MAOI22D0BWP12T U2649 ( .A1(n3139), .A2(n2227), .B1(n3142), .B2(n2226), .ZN(
        n2229) );
  ND2D1BWP12T U2650 ( .A1(n3684), .A2(n3685), .ZN(n2715) );
  NR3D1BWP12T U2651 ( .A1(a[19]), .A2(a[18]), .A3(a[17]), .ZN(n2723) );
  ND2D1BWP12T U2652 ( .A1(n3174), .A2(n3961), .ZN(n3992) );
  NR3D1BWP12T U2653 ( .A1(a[4]), .A2(a[3]), .A3(n3992), .ZN(n3248) );
  ND2D1BWP12T U2654 ( .A1(n3248), .A2(n3247), .ZN(n3297) );
  ND2D1BWP12T U2655 ( .A1(n3292), .A2(n3276), .ZN(n2718) );
  NR2D1BWP12T U2656 ( .A1(n3297), .A2(n2718), .ZN(n3322) );
  ND2D1BWP12T U2657 ( .A1(n3322), .A2(n3321), .ZN(n3339) );
  NR2D1BWP12T U2658 ( .A1(a[9]), .A2(n3339), .ZN(n3381) );
  ND2D1BWP12T U2659 ( .A1(n4005), .A2(n3380), .ZN(n2717) );
  INR2D1BWP12T U2660 ( .A1(n3381), .B1(n2717), .ZN(n3429) );
  AN3XD1BWP12T U2661 ( .A1(n3429), .A2(n3446), .A3(n3428), .Z(n3480) );
  ND2D1BWP12T U2662 ( .A1(n3480), .A2(n3479), .ZN(n3504) );
  ND2D1BWP12T U2663 ( .A1(n3529), .A2(n2485), .ZN(n2716) );
  NR2D1BWP12T U2664 ( .A1(n3504), .A2(n2716), .ZN(n3566) );
  ND2D1BWP12T U2665 ( .A1(n2723), .A2(n3566), .ZN(n3625) );
  NR2D1BWP12T U2666 ( .A1(a[20]), .A2(n3625), .ZN(n3686) );
  IND2D1BWP12T U2667 ( .A1(n2715), .B1(n3686), .ZN(n3708) );
  NR2D1BWP12T U2668 ( .A1(a[23]), .A2(n3708), .ZN(n3722) );
  NR2D1BWP12T U2669 ( .A1(a[25]), .A2(a[24]), .ZN(n2720) );
  ND2D1BWP12T U2670 ( .A1(n3722), .A2(n2720), .ZN(n3781) );
  NR2D1BWP12T U2671 ( .A1(a[26]), .A2(n3781), .ZN(n3810) );
  NR2D1BWP12T U2672 ( .A1(a[28]), .A2(a[27]), .ZN(n2719) );
  ND2D1BWP12T U2673 ( .A1(n3810), .A2(n2719), .ZN(n3874) );
  NR2D1BWP12T U2674 ( .A1(a[29]), .A2(n3874), .ZN(n3933) );
  ND2D1BWP12T U2675 ( .A1(n3933), .A2(n3932), .ZN(n3931) );
  INVD1BWP12T U2676 ( .I(n3931), .ZN(n2938) );
  ND2D1BWP12T U2677 ( .A1(n2228), .A2(n3102), .ZN(n3990) );
  INVD1BWP12T U2678 ( .I(n3990), .ZN(n3945) );
  ND3D1BWP12T U2679 ( .A1(a[31]), .A2(n2938), .A3(n3945), .ZN(n3205) );
  ND3D1BWP12T U2680 ( .A1(n2230), .A2(n2229), .A3(n3205), .ZN(v) );
  NR2D1BWP12T U2681 ( .A1(a[29]), .A2(b[29]), .ZN(n3025) );
  NR2D1BWP12T U2682 ( .A1(a[28]), .A2(b[28]), .ZN(n3024) );
  NR2D1BWP12T U2683 ( .A1(a[27]), .A2(b[27]), .ZN(n3023) );
  NR2D1BWP12T U2684 ( .A1(a[26]), .A2(b[26]), .ZN(n3794) );
  NR2D1BWP12T U2685 ( .A1(a[25]), .A2(b[25]), .ZN(n3022) );
  ND2D1BWP12T U2686 ( .A1(n3725), .A2(n2518), .ZN(n3728) );
  INVD1BWP12T U2687 ( .I(n3728), .ZN(n3021) );
  NR2D1BWP12T U2688 ( .A1(b[23]), .A2(a[23]), .ZN(n3020) );
  NR2D1BWP12T U2689 ( .A1(a[22]), .A2(b[22]), .ZN(n3019) );
  NR2D1BWP12T U2690 ( .A1(b[21]), .A2(a[21]), .ZN(n3657) );
  NR2D1BWP12T U2691 ( .A1(b[20]), .A2(a[20]), .ZN(n3018) );
  NR2D1BWP12T U2692 ( .A1(b[19]), .A2(a[19]), .ZN(n3017) );
  NR2D1BWP12T U2693 ( .A1(a[18]), .A2(b[18]), .ZN(n3016) );
  NR2D1BWP12T U2694 ( .A1(a[17]), .A2(b[17]), .ZN(n3015) );
  NR2D1BWP12T U2695 ( .A1(b[16]), .A2(a[16]), .ZN(n3014) );
  ND2D1BWP12T U2696 ( .A1(n2485), .A2(n2231), .ZN(n3495) );
  INVD1BWP12T U2697 ( .I(n3495), .ZN(n3013) );
  NR2D1BWP12T U2698 ( .A1(a[14]), .A2(b[14]), .ZN(n3012) );
  ND2D1BWP12T U2699 ( .A1(n3446), .A2(n2371), .ZN(n2721) );
  INVD1BWP12T U2700 ( .I(n2721), .ZN(n3011) );
  NR2D1BWP12T U2701 ( .A1(a[12]), .A2(b[12]), .ZN(n3010) );
  NR2D1BWP12T U2702 ( .A1(a[11]), .A2(b[11]), .ZN(n3009) );
  ND2D1BWP12T U2703 ( .A1(n3380), .A2(n3370), .ZN(n3373) );
  INVD1BWP12T U2704 ( .I(n3373), .ZN(n3008) );
  NR2D1BWP12T U2705 ( .A1(a[9]), .A2(b[9]), .ZN(n3007) );
  NR2D1BWP12T U2706 ( .A1(a[8]), .A2(b[8]), .ZN(n3006) );
  NR2D1BWP12T U2707 ( .A1(a[7]), .A2(b[7]), .ZN(n3005) );
  NR2D1BWP12T U2708 ( .A1(a[6]), .A2(b[6]), .ZN(n3004) );
  NR2D1BWP12T U2709 ( .A1(a[5]), .A2(b[5]), .ZN(n3003) );
  NR2D1BWP12T U2710 ( .A1(a[4]), .A2(b[4]), .ZN(n3002) );
  ND2D1BWP12T U2711 ( .A1(a[4]), .A2(b[4]), .ZN(n2726) );
  IND2D1BWP12T U2712 ( .A1(n3002), .B1(n2726), .ZN(n3097) );
  ND2D1BWP12T U2713 ( .A1(a[3]), .A2(b[3]), .ZN(n3993) );
  NR2D1BWP12T U2714 ( .A1(a[3]), .A2(b[3]), .ZN(n3001) );
  IND2D1BWP12T U2715 ( .A1(n3001), .B1(n3993), .ZN(n3100) );
  INVD1BWP12T U2716 ( .I(n3100), .ZN(n2336) );
  ND2D1BWP12T U2717 ( .A1(b[2]), .A2(a[2]), .ZN(n3939) );
  INR2D1BWP12T U2718 ( .A1(n3163), .B1(n2474), .ZN(n2725) );
  NR2D1BWP12T U2719 ( .A1(n3168), .A2(n2725), .ZN(n2290) );
  ND2D1BWP12T U2720 ( .A1(n2290), .A2(n3107), .ZN(n2289) );
  ND2D1BWP12T U2721 ( .A1(n3939), .A2(n2289), .ZN(n2292) );
  ND2D1BWP12T U2722 ( .A1(n2336), .A2(n2292), .ZN(n2291) );
  ND2D1BWP12T U2723 ( .A1(n3993), .A2(n2291), .ZN(n2286) );
  NR2D1BWP12T U2724 ( .A1(n3097), .A2(n2286), .ZN(n2285) );
  NR2D1BWP12T U2725 ( .A1(n3002), .A2(n2285), .ZN(n2284) );
  INVD1BWP12T U2726 ( .I(n3003), .ZN(n3241) );
  ND2D1BWP12T U2727 ( .A1(a[5]), .A2(b[5]), .ZN(n3239) );
  ND2D1BWP12T U2728 ( .A1(n3241), .A2(n3239), .ZN(n3116) );
  NR2D1BWP12T U2729 ( .A1(n2284), .A2(n3116), .ZN(n2283) );
  NR2D1BWP12T U2730 ( .A1(n3003), .A2(n2283), .ZN(n2282) );
  ND2D1BWP12T U2731 ( .A1(a[6]), .A2(b[6]), .ZN(n3273) );
  IND2D1BWP12T U2732 ( .A1(n3004), .B1(n3273), .ZN(n3113) );
  NR2D1BWP12T U2733 ( .A1(n2282), .A2(n3113), .ZN(n2281) );
  NR2D1BWP12T U2734 ( .A1(n3004), .A2(n2281), .ZN(n2280) );
  ND2D1BWP12T U2735 ( .A1(a[7]), .A2(b[7]), .ZN(n3290) );
  IND2D1BWP12T U2736 ( .A1(n3005), .B1(n3290), .ZN(n3110) );
  NR2D1BWP12T U2737 ( .A1(n2280), .A2(n3110), .ZN(n2279) );
  NR2D1BWP12T U2738 ( .A1(n3005), .A2(n2279), .ZN(n2278) );
  ND2D1BWP12T U2739 ( .A1(a[8]), .A2(b[8]), .ZN(n3318) );
  IND2D1BWP12T U2740 ( .A1(n3006), .B1(n3318), .ZN(n3094) );
  NR2D1BWP12T U2741 ( .A1(n2278), .A2(n3094), .ZN(n2277) );
  NR2D1BWP12T U2742 ( .A1(n3006), .A2(n2277), .ZN(n2276) );
  ND2D1BWP12T U2743 ( .A1(a[9]), .A2(b[9]), .ZN(n3342) );
  IND2D1BWP12T U2744 ( .A1(n3007), .B1(n3342), .ZN(n3091) );
  NR2D1BWP12T U2745 ( .A1(n2276), .A2(n3091), .ZN(n2275) );
  NR2D1BWP12T U2746 ( .A1(n3007), .A2(n2275), .ZN(n2274) );
  ND2D1BWP12T U2747 ( .A1(a[10]), .A2(b[10]), .ZN(n3372) );
  ND2D1BWP12T U2748 ( .A1(n3373), .A2(n3372), .ZN(n3088) );
  NR2D1BWP12T U2749 ( .A1(n2274), .A2(n3088), .ZN(n2273) );
  NR2D1BWP12T U2750 ( .A1(n3008), .A2(n2273), .ZN(n2272) );
  ND2D1BWP12T U2751 ( .A1(a[11]), .A2(b[11]), .ZN(n3394) );
  IND2D1BWP12T U2752 ( .A1(n3009), .B1(n3394), .ZN(n3085) );
  NR2D1BWP12T U2753 ( .A1(n2272), .A2(n3085), .ZN(n2271) );
  NR2D1BWP12T U2754 ( .A1(n3009), .A2(n2271), .ZN(n2270) );
  ND2D1BWP12T U2755 ( .A1(a[12]), .A2(b[12]), .ZN(n3418) );
  IND2D1BWP12T U2756 ( .A1(n3010), .B1(n3418), .ZN(n3082) );
  NR2D1BWP12T U2757 ( .A1(n2270), .A2(n3082), .ZN(n2269) );
  NR2D1BWP12T U2758 ( .A1(n3010), .A2(n2269), .ZN(n2268) );
  ND2D1BWP12T U2759 ( .A1(a[13]), .A2(b[13]), .ZN(n3442) );
  ND2D1BWP12T U2760 ( .A1(n2721), .A2(n3442), .ZN(n3079) );
  NR2D1BWP12T U2761 ( .A1(n2268), .A2(n3079), .ZN(n2267) );
  NR2D1BWP12T U2762 ( .A1(n3011), .A2(n2267), .ZN(n2266) );
  ND2D1BWP12T U2763 ( .A1(a[14]), .A2(b[14]), .ZN(n3474) );
  IND2D1BWP12T U2764 ( .A1(n3012), .B1(n3474), .ZN(n3076) );
  NR2D1BWP12T U2765 ( .A1(n2266), .A2(n3076), .ZN(n2265) );
  NR2D1BWP12T U2766 ( .A1(n3012), .A2(n2265), .ZN(n2264) );
  ND2D1BWP12T U2767 ( .A1(a[15]), .A2(b[15]), .ZN(n3493) );
  ND2D1BWP12T U2768 ( .A1(n3495), .A2(n3493), .ZN(n3073) );
  NR2D1BWP12T U2769 ( .A1(n2264), .A2(n3073), .ZN(n2263) );
  NR2D1BWP12T U2770 ( .A1(n3013), .A2(n2263), .ZN(n2262) );
  AOI22D1BWP12T U2771 ( .A1(b[16]), .A2(n3529), .B1(a[16]), .B2(n2232), .ZN(
        n3070) );
  NR2D1BWP12T U2772 ( .A1(n2262), .A2(n3070), .ZN(n2261) );
  NR2D1BWP12T U2773 ( .A1(n3014), .A2(n2261), .ZN(n2260) );
  ND2D1BWP12T U2774 ( .A1(a[17]), .A2(b[17]), .ZN(n3556) );
  IND2D1BWP12T U2775 ( .A1(n3015), .B1(n3556), .ZN(n3067) );
  NR2D1BWP12T U2776 ( .A1(n2260), .A2(n3067), .ZN(n2259) );
  NR2D1BWP12T U2777 ( .A1(n3015), .A2(n2259), .ZN(n2258) );
  ND2D1BWP12T U2778 ( .A1(a[18]), .A2(b[18]), .ZN(n3574) );
  IND2D1BWP12T U2779 ( .A1(n3016), .B1(n3574), .ZN(n3064) );
  NR2D1BWP12T U2780 ( .A1(n2258), .A2(n3064), .ZN(n2257) );
  NR2D1BWP12T U2781 ( .A1(n3016), .A2(n2257), .ZN(n2256) );
  ND2D1BWP12T U2782 ( .A1(b[19]), .A2(a[19]), .ZN(n3608) );
  IND2D1BWP12T U2783 ( .A1(n3017), .B1(n3608), .ZN(n3061) );
  NR2D1BWP12T U2784 ( .A1(n2256), .A2(n3061), .ZN(n2255) );
  NR2D1BWP12T U2785 ( .A1(n3017), .A2(n2255), .ZN(n2254) );
  AOI22D1BWP12T U2786 ( .A1(b[20]), .A2(n3632), .B1(a[20]), .B2(n3628), .ZN(
        n3629) );
  NR2D1BWP12T U2787 ( .A1(n2254), .A2(n3629), .ZN(n2253) );
  NR2D1BWP12T U2788 ( .A1(n3018), .A2(n2253), .ZN(n2252) );
  ND2D1BWP12T U2789 ( .A1(b[21]), .A2(a[21]), .ZN(n3651) );
  IND2D1BWP12T U2790 ( .A1(n3657), .B1(n3651), .ZN(n3056) );
  NR2D1BWP12T U2791 ( .A1(n2252), .A2(n3056), .ZN(n2251) );
  NR2D1BWP12T U2792 ( .A1(n3657), .A2(n2251), .ZN(n2250) );
  ND2D1BWP12T U2793 ( .A1(a[22]), .A2(b[22]), .ZN(n3672) );
  IND2D1BWP12T U2794 ( .A1(n3019), .B1(n3672), .ZN(n3053) );
  NR2D1BWP12T U2795 ( .A1(n2250), .A2(n3053), .ZN(n2249) );
  NR2D1BWP12T U2796 ( .A1(n3019), .A2(n2249), .ZN(n2248) );
  ND2D1BWP12T U2797 ( .A1(b[23]), .A2(a[23]), .ZN(n3698) );
  IND2D1BWP12T U2798 ( .A1(n3020), .B1(n3698), .ZN(n3050) );
  NR2D1BWP12T U2799 ( .A1(n2248), .A2(n3050), .ZN(n2247) );
  NR2D1BWP12T U2800 ( .A1(n3020), .A2(n2247), .ZN(n2246) );
  ND2D1BWP12T U2801 ( .A1(b[24]), .A2(a[24]), .ZN(n3727) );
  ND2D1BWP12T U2802 ( .A1(n3728), .A2(n3727), .ZN(n3047) );
  NR2D1BWP12T U2803 ( .A1(n2246), .A2(n3047), .ZN(n2245) );
  NR2D1BWP12T U2804 ( .A1(n3021), .A2(n2245), .ZN(n2244) );
  ND2D1BWP12T U2805 ( .A1(a[25]), .A2(b[25]), .ZN(n3759) );
  IND2D1BWP12T U2806 ( .A1(n3022), .B1(n3759), .ZN(n3044) );
  NR2D1BWP12T U2807 ( .A1(n2244), .A2(n3044), .ZN(n2243) );
  NR2D1BWP12T U2808 ( .A1(n3022), .A2(n2243), .ZN(n2242) );
  ND2D1BWP12T U2809 ( .A1(a[26]), .A2(b[26]), .ZN(n3788) );
  IND2D1BWP12T U2810 ( .A1(n3794), .B1(n3788), .ZN(n3041) );
  NR2D1BWP12T U2811 ( .A1(n2242), .A2(n3041), .ZN(n2241) );
  NR2D1BWP12T U2812 ( .A1(n3794), .A2(n2241), .ZN(n2240) );
  AOI22D1BWP12T U2813 ( .A1(a[27]), .A2(n2361), .B1(b[27]), .B2(n3824), .ZN(
        n3038) );
  NR2D1BWP12T U2814 ( .A1(n2240), .A2(n3038), .ZN(n2239) );
  NR2D1BWP12T U2815 ( .A1(n3023), .A2(n2239), .ZN(n2238) );
  INVD1BWP12T U2816 ( .I(b[28]), .ZN(n2362) );
  AOI22D1BWP12T U2817 ( .A1(a[28]), .A2(n2362), .B1(b[28]), .B2(n3851), .ZN(
        n3035) );
  NR2D1BWP12T U2818 ( .A1(n2238), .A2(n3035), .ZN(n2237) );
  NR2D1BWP12T U2819 ( .A1(n3024), .A2(n2237), .ZN(n2236) );
  ND2D1BWP12T U2820 ( .A1(a[29]), .A2(b[29]), .ZN(n3866) );
  IND2D1BWP12T U2821 ( .A1(n3025), .B1(n3866), .ZN(n3032) );
  NR2D1BWP12T U2822 ( .A1(n2236), .A2(n3032), .ZN(n2235) );
  NR2D1BWP12T U2823 ( .A1(n3025), .A2(n2235), .ZN(n2233) );
  ND2D1BWP12T U2824 ( .A1(n3912), .A2(n3932), .ZN(n2722) );
  ND2D1BWP12T U2825 ( .A1(b[30]), .A2(a[30]), .ZN(n3918) );
  ND2D1BWP12T U2826 ( .A1(n2722), .A2(n3918), .ZN(n3029) );
  NR2D1BWP12T U2827 ( .A1(n2233), .A2(n3029), .ZN(n2234) );
  AOI21D1BWP12T U2828 ( .A1(n2233), .A2(n3029), .B(n2234), .ZN(n3928) );
  INVD1BWP12T U2829 ( .I(n2722), .ZN(n3026) );
  NR2D1BWP12T U2830 ( .A1(n3026), .A2(n2234), .ZN(n3137) );
  NR2D1BWP12T U2831 ( .A1(n3143), .A2(n2773), .ZN(n3027) );
  MOAI22D0BWP12T U2832 ( .A1(n3137), .A2(n3027), .B1(n3137), .B2(n3027), .ZN(
        n3211) );
  AO21D1BWP12T U2833 ( .A1(n2236), .A2(n3032), .B(n2235), .Z(n3905) );
  AO21D1BWP12T U2834 ( .A1(n2238), .A2(n3035), .B(n2237), .Z(n3859) );
  AOI21D1BWP12T U2835 ( .A1(n2240), .A2(n3038), .B(n2239), .ZN(n3827) );
  AOI21D1BWP12T U2836 ( .A1(n2242), .A2(n3041), .B(n2241), .ZN(n3809) );
  AOI21D1BWP12T U2837 ( .A1(n2244), .A2(n3044), .B(n2243), .ZN(n3780) );
  AO21D1BWP12T U2838 ( .A1(n2246), .A2(n3047), .B(n2245), .Z(n3751) );
  AO21D1BWP12T U2839 ( .A1(n2248), .A2(n3050), .B(n2247), .Z(n3717) );
  AO21D1BWP12T U2840 ( .A1(n2250), .A2(n3053), .B(n2249), .Z(n3692) );
  AOI21D1BWP12T U2841 ( .A1(n2252), .A2(n3056), .B(n2251), .ZN(n3668) );
  AOI21D1BWP12T U2842 ( .A1(n2254), .A2(n3629), .B(n2253), .ZN(n3645) );
  AOI21D1BWP12T U2843 ( .A1(n2256), .A2(n3061), .B(n2255), .ZN(n3619) );
  AO21D1BWP12T U2844 ( .A1(n2258), .A2(n3064), .B(n2257), .Z(n3593) );
  AO21D1BWP12T U2845 ( .A1(n2260), .A2(n3067), .B(n2259), .Z(n3572) );
  AO21D1BWP12T U2846 ( .A1(n2262), .A2(n3070), .B(n2261), .Z(n3539) );
  AOI21D1BWP12T U2847 ( .A1(n2264), .A2(n3073), .B(n2263), .ZN(n3515) );
  AOI21D1BWP12T U2848 ( .A1(n2266), .A2(n3076), .B(n2265), .ZN(n3490) );
  AOI21D1BWP12T U2849 ( .A1(n2268), .A2(n3079), .B(n2267), .ZN(n3461) );
  AO21D1BWP12T U2850 ( .A1(n2270), .A2(n3082), .B(n2269), .Z(n3436) );
  AO21D1BWP12T U2851 ( .A1(n2272), .A2(n3085), .B(n2271), .Z(n3409) );
  AO21D1BWP12T U2852 ( .A1(n2274), .A2(n3088), .B(n2273), .Z(n3388) );
  AOI21D1BWP12T U2853 ( .A1(n2276), .A2(n3091), .B(n2275), .ZN(n3361) );
  AOI21D1BWP12T U2854 ( .A1(n2278), .A2(n3094), .B(n2277), .ZN(n3338) );
  AOI21D1BWP12T U2855 ( .A1(n2280), .A2(n3110), .B(n2279), .ZN(n3313) );
  AO21D1BWP12T U2856 ( .A1(n2282), .A2(n3113), .B(n2281), .Z(n3263) );
  AO21D1BWP12T U2857 ( .A1(n2284), .A2(n3116), .B(n2283), .Z(n3238) );
  AO21D1BWP12T U2858 ( .A1(n3097), .A2(n2286), .B(n2285), .Z(n3228) );
  NR2D1BWP12T U2859 ( .A1(n2288), .A2(n2287), .ZN(n3906) );
  OAI21D1BWP12T U2860 ( .A1(n2290), .A2(n3107), .B(n2289), .ZN(n3964) );
  OAI21D1BWP12T U2861 ( .A1(n2336), .A2(n2292), .B(n2291), .ZN(n3974) );
  AOI22D1BWP12T U2862 ( .A1(n3105), .A2(n3147), .B1(n2474), .B2(n2976), .ZN(
        n3175) );
  ND4D1BWP12T U2863 ( .A1(n3906), .A2(n3964), .A3(n3974), .A4(n3175), .ZN(
        n2293) );
  NR4D0BWP12T U2864 ( .A1(n3263), .A2(n3238), .A3(n3228), .A4(n2293), .ZN(
        n2294) );
  ND4D1BWP12T U2865 ( .A1(n3361), .A2(n3338), .A3(n3313), .A4(n2294), .ZN(
        n2295) );
  NR4D0BWP12T U2866 ( .A1(n3436), .A2(n3409), .A3(n3388), .A4(n2295), .ZN(
        n2296) );
  ND4D1BWP12T U2867 ( .A1(n3515), .A2(n3490), .A3(n3461), .A4(n2296), .ZN(
        n2297) );
  NR4D0BWP12T U2868 ( .A1(n3593), .A2(n3572), .A3(n3539), .A4(n2297), .ZN(
        n2298) );
  ND4D1BWP12T U2869 ( .A1(n3668), .A2(n3645), .A3(n3619), .A4(n2298), .ZN(
        n2299) );
  NR4D0BWP12T U2870 ( .A1(n3751), .A2(n3717), .A3(n3692), .A4(n2299), .ZN(
        n2300) );
  ND4D1BWP12T U2871 ( .A1(n3827), .A2(n3809), .A3(n3780), .A4(n2300), .ZN(
        n2301) );
  NR4D0BWP12T U2872 ( .A1(n3211), .A2(n3905), .A3(n3859), .A4(n2301), .ZN(
        n2358) );
  MAOI22D0BWP12T U2873 ( .A1(n2302), .A2(n3027), .B1(n2302), .B2(n3027), .ZN(
        n3207) );
  ND2D1BWP12T U2874 ( .A1(n2304), .A2(n2303), .ZN(n2305) );
  MAOI22D0BWP12T U2875 ( .A1(n3032), .A2(n2305), .B1(n3032), .B2(n2305), .ZN(
        n3895) );
  MAOI22D0BWP12T U2876 ( .A1(n2306), .A2(n3029), .B1(n2306), .B2(n3029), .ZN(
        n3925) );
  MAOI22D0BWP12T U2877 ( .A1(n2307), .A2(n3035), .B1(n2307), .B2(n3035), .ZN(
        n3858) );
  MOAI22D0BWP12T U2878 ( .A1(n2308), .A2(n3041), .B1(n2308), .B2(n3041), .ZN(
        n3801) );
  MAOI22D0BWP12T U2879 ( .A1(n2309), .A2(n3053), .B1(n2309), .B2(n3053), .ZN(
        n3691) );
  ND2D1BWP12T U2880 ( .A1(n3675), .A2(n2310), .ZN(n2311) );
  MAOI22D0BWP12T U2881 ( .A1(n3050), .A2(n2311), .B1(n3050), .B2(n2311), .ZN(
        n3714) );
  NR2D1BWP12T U2882 ( .A1(n3697), .A2(a[23]), .ZN(n2947) );
  IND2D1BWP12T U2883 ( .A1(n2947), .B1(n2312), .ZN(n2313) );
  MOAI22D0BWP12T U2884 ( .A1(n3047), .A2(n2313), .B1(n3047), .B2(n2313), .ZN(
        n3750) );
  ND2D1BWP12T U2885 ( .A1(n3632), .A2(b[20]), .ZN(n2953) );
  INR2D1BWP12T U2886 ( .A1(n2953), .B1(n2314), .ZN(n2315) );
  MOAI22D0BWP12T U2887 ( .A1(n2315), .A2(n3056), .B1(n2315), .B2(n3056), .ZN(
        n3666) );
  MOAI22D0BWP12T U2888 ( .A1(n2316), .A2(n3629), .B1(n2316), .B2(n3629), .ZN(
        n3648) );
  MAOI22D0BWP12T U2889 ( .A1(n2317), .A2(n3061), .B1(n2317), .B2(n3061), .ZN(
        n3614) );
  ND2D1BWP12T U2890 ( .A1(n3544), .A2(a[17]), .ZN(n2992) );
  INR2D1BWP12T U2891 ( .A1(n2992), .B1(n2318), .ZN(n2319) );
  MOAI22D0BWP12T U2892 ( .A1(n2319), .A2(n3064), .B1(n2319), .B2(n3064), .ZN(
        n3592) );
  MOAI22D0BWP12T U2893 ( .A1(n2320), .A2(n3067), .B1(n2320), .B2(n3067), .ZN(
        n3561) );
  MAOI22D0BWP12T U2894 ( .A1(n2321), .A2(n3070), .B1(n2321), .B2(n3070), .ZN(
        n3538) );
  MAOI22D0BWP12T U2895 ( .A1(n2322), .A2(n3073), .B1(n2322), .B2(n3073), .ZN(
        n3513) );
  INR2D1BWP12T U2896 ( .A1(n3343), .B1(n2323), .ZN(n2324) );
  MOAI22D0BWP12T U2897 ( .A1(n2324), .A2(n3088), .B1(n2324), .B2(n3088), .ZN(
        n3387) );
  MOAI22D0BWP12T U2898 ( .A1(n2325), .A2(n3085), .B1(n2325), .B2(n3085), .ZN(
        n3408) );
  MAOI22D0BWP12T U2899 ( .A1(n2326), .A2(n3082), .B1(n2326), .B2(n3082), .ZN(
        n3435) );
  MAOI22D0BWP12T U2900 ( .A1(n2327), .A2(n3091), .B1(n2327), .B2(n3091), .ZN(
        n3359) );
  MAOI22D0BWP12T U2901 ( .A1(n2328), .A2(n3110), .B1(n2328), .B2(n3110), .ZN(
        n3305) );
  NR2D1BWP12T U2902 ( .A1(n2982), .A2(n2329), .ZN(n2330) );
  MOAI22D0BWP12T U2903 ( .A1(n2330), .A2(n3113), .B1(n2330), .B2(n3113), .ZN(
        n3285) );
  ND2D1BWP12T U2904 ( .A1(n2886), .A2(a[3]), .ZN(n2968) );
  INR2D1BWP12T U2905 ( .A1(n2968), .B1(n2331), .ZN(n2332) );
  MOAI22D0BWP12T U2906 ( .A1(n2332), .A2(n3097), .B1(n2332), .B2(n3097), .ZN(
        n3226) );
  MOAI22D0BWP12T U2907 ( .A1(n2333), .A2(n3116), .B1(n2333), .B2(n3116), .ZN(
        n3255) );
  INR2D1BWP12T U2908 ( .A1(n2334), .B1(n2337), .ZN(n2335) );
  MAOI22D0BWP12T U2909 ( .A1(n2336), .A2(n2335), .B1(n2336), .B2(n2335), .ZN(
        n3977) );
  AOI21D1BWP12T U2910 ( .A1(n2338), .A2(n3107), .B(n2337), .ZN(n3942) );
  AOI21D1BWP12T U2911 ( .A1(n3105), .A2(n2769), .B(n2339), .ZN(n3177) );
  ND4D1BWP12T U2912 ( .A1(n3926), .A2(n3977), .A3(n3942), .A4(n3177), .ZN(
        n2340) );
  NR4D0BWP12T U2913 ( .A1(n3285), .A2(n3226), .A3(n3255), .A4(n2340), .ZN(
        n2343) );
  ND2D1BWP12T U2914 ( .A1(n3291), .A2(a[7]), .ZN(n2979) );
  INR2D1BWP12T U2915 ( .A1(n2979), .B1(n2341), .ZN(n2342) );
  MAOI22D0BWP12T U2916 ( .A1(n2342), .A2(n3094), .B1(n2342), .B2(n3094), .ZN(
        n3331) );
  ND4D1BWP12T U2917 ( .A1(n3359), .A2(n3305), .A3(n2343), .A4(n3331), .ZN(
        n2344) );
  NR4D0BWP12T U2918 ( .A1(n3387), .A2(n3408), .A3(n3435), .A4(n2344), .ZN(
        n2348) );
  MAOI22D0BWP12T U2919 ( .A1(n2345), .A2(n3079), .B1(n2345), .B2(n3079), .ZN(
        n3459) );
  NR2D1BWP12T U2920 ( .A1(n3443), .A2(n2346), .ZN(n2347) );
  MAOI22D0BWP12T U2921 ( .A1(n2347), .A2(n3076), .B1(n2347), .B2(n3076), .ZN(
        n3483) );
  ND4D1BWP12T U2922 ( .A1(n3513), .A2(n2348), .A3(n3459), .A4(n3483), .ZN(
        n2349) );
  NR4D0BWP12T U2923 ( .A1(n3592), .A2(n3561), .A3(n3538), .A4(n2349), .ZN(
        n2350) );
  ND4D1BWP12T U2924 ( .A1(n3666), .A2(n3648), .A3(n3614), .A4(n2350), .ZN(
        n2351) );
  NR4D0BWP12T U2925 ( .A1(n3691), .A2(n3714), .A3(n3750), .A4(n2351), .ZN(
        n2355) );
  ND2D1BWP12T U2926 ( .A1(n3787), .A2(n2352), .ZN(n2353) );
  MOAI22D0BWP12T U2927 ( .A1(n3038), .A2(n2353), .B1(n3038), .B2(n2353), .ZN(
        n3829) );
  MAOI22D0BWP12T U2928 ( .A1(n2354), .A2(n3044), .B1(n2354), .B2(n3044), .ZN(
        n3772) );
  ND4D1BWP12T U2929 ( .A1(n3801), .A2(n2355), .A3(n3829), .A4(n3772), .ZN(
        n2356) );
  NR4D0BWP12T U2930 ( .A1(n3895), .A2(n3925), .A3(n3858), .A4(n2356), .ZN(
        n2357) );
  AOI22D1BWP12T U2931 ( .A1(n3928), .A2(n2358), .B1(n3207), .B2(n2357), .ZN(
        n3132) );
  ND2D1BWP12T U2932 ( .A1(n3155), .A2(n2769), .ZN(n3151) );
  NR2D1BWP12T U2933 ( .A1(a[31]), .A2(n3990), .ZN(n3140) );
  ND4D1BWP12T U2934 ( .A1(n3757), .A2(n3725), .A3(n2359), .A4(n2774), .ZN(
        n2370) );
  ND4D1BWP12T U2935 ( .A1(n2363), .A2(n2362), .A3(n2361), .A4(n2360), .ZN(
        n2369) );
  NR4D0BWP12T U2936 ( .A1(b[11]), .A2(b[10]), .A3(b[9]), .A4(b[8]), .ZN(n2367)
         );
  NR4D0BWP12T U2937 ( .A1(b[7]), .A2(b[6]), .A3(b[5]), .A4(b[23]), .ZN(n2366)
         );
  NR4D0BWP12T U2938 ( .A1(b[16]), .A2(b[15]), .A3(b[14]), .A4(b[12]), .ZN(
        n2365) );
  NR4D0BWP12T U2939 ( .A1(b[20]), .A2(b[19]), .A3(b[18]), .A4(b[17]), .ZN(
        n2364) );
  ND4D1BWP12T U2940 ( .A1(n2367), .A2(n2366), .A3(n2365), .A4(n2364), .ZN(
        n2368) );
  NR3D1BWP12T U2941 ( .A1(n2370), .A2(n2369), .A3(n2368), .ZN(n2735) );
  AN4XD1BWP12T U2942 ( .A1(n2735), .A2(n3193), .A3(n3912), .A4(n2371), .Z(
        n3144) );
  INVD1BWP12T U2943 ( .I(n3144), .ZN(n2626) );
  NR2D1BWP12T U2944 ( .A1(n2512), .A2(n2652), .ZN(n2508) );
  INVD1BWP12T U2945 ( .I(n2508), .ZN(n2469) );
  AOI22D1BWP12T U2946 ( .A1(b[0]), .A2(n3932), .B1(n3869), .B2(n2534), .ZN(
        n2881) );
  AOI22D1BWP12T U2947 ( .A1(b[0]), .A2(n3851), .B1(n3824), .B2(n2534), .ZN(
        n2373) );
  AOI22D1BWP12T U2948 ( .A1(b[1]), .A2(n2881), .B1(n2373), .B2(n3165), .ZN(
        n2438) );
  MOAI22D0BWP12T U2949 ( .A1(n2652), .A2(a[31]), .B1(n2438), .B2(n2652), .ZN(
        n2397) );
  NR2D1BWP12T U2950 ( .A1(b[3]), .A2(n2397), .ZN(n2856) );
  ND2D1BWP12T U2951 ( .A1(n2469), .A2(n2856), .ZN(n3825) );
  INVD1BWP12T U2952 ( .I(n3825), .ZN(n2547) );
  AOI22D1BWP12T U2953 ( .A1(b[0]), .A2(a[18]), .B1(a[17]), .B2(n2534), .ZN(
        n2376) );
  AOI22D1BWP12T U2954 ( .A1(b[0]), .A2(a[16]), .B1(a[15]), .B2(n3170), .ZN(
        n2379) );
  AOI22D1BWP12T U2955 ( .A1(b[1]), .A2(n2376), .B1(n2379), .B2(n3165), .ZN(
        n2435) );
  AOI22D1BWP12T U2956 ( .A1(b[0]), .A2(a[14]), .B1(a[13]), .B2(n3170), .ZN(
        n2378) );
  AOI22D1BWP12T U2957 ( .A1(b[0]), .A2(a[12]), .B1(a[11]), .B2(n3170), .ZN(
        n2380) );
  AOI22D1BWP12T U2958 ( .A1(b[1]), .A2(n2378), .B1(n2380), .B2(n3165), .ZN(
        n2457) );
  AOI22D1BWP12T U2959 ( .A1(b[2]), .A2(n2435), .B1(n2457), .B2(n2652), .ZN(
        n2568) );
  AOI22D1BWP12T U2960 ( .A1(b[0]), .A2(a[22]), .B1(a[21]), .B2(n3170), .ZN(
        n2374) );
  AOI22D1BWP12T U2961 ( .A1(b[0]), .A2(a[20]), .B1(a[19]), .B2(n3170), .ZN(
        n2377) );
  AOI22D1BWP12T U2962 ( .A1(b[1]), .A2(n2374), .B1(n2377), .B2(n3165), .ZN(
        n2436) );
  OAI22D1BWP12T U2963 ( .A1(n2534), .A2(n3790), .B1(n3768), .B2(b[0]), .ZN(
        n2372) );
  AOI22D1BWP12T U2964 ( .A1(b[0]), .A2(a[24]), .B1(a[23]), .B2(n3170), .ZN(
        n2375) );
  MOAI22D0BWP12T U2965 ( .A1(n3165), .A2(n2372), .B1(n2375), .B2(n2593), .ZN(
        n2437) );
  MAOI22D0BWP12T U2966 ( .A1(n2436), .A2(n2652), .B1(n2652), .B2(n2437), .ZN(
        n2496) );
  AOI22D1BWP12T U2967 ( .A1(n3784), .A2(n2568), .B1(n2912), .B2(n2496), .ZN(
        n2857) );
  OAI21D1BWP12T U2968 ( .A1(n2547), .A2(n3219), .B(n2857), .ZN(n3406) );
  NR2D1BWP12T U2969 ( .A1(n2626), .A2(n3406), .ZN(n3405) );
  NR2D1BWP12T U2970 ( .A1(b[1]), .A2(n2881), .ZN(n2383) );
  OAI21D1BWP12T U2971 ( .A1(a[31]), .A2(n2593), .B(b[2]), .ZN(n2869) );
  AOI22D1BWP12T U2972 ( .A1(b[1]), .A2(n2373), .B1(n2372), .B2(n3165), .ZN(
        n2426) );
  OAI22D1BWP12T U2973 ( .A1(n2383), .A2(n2869), .B1(b[2]), .B2(n2426), .ZN(
        n2444) );
  ND2D1BWP12T U2974 ( .A1(n2886), .A2(n2444), .ZN(n2873) );
  IND2D1BWP12T U2975 ( .A1(n2873), .B1(n2445), .ZN(n2564) );
  INVD1BWP12T U2976 ( .I(n2564), .ZN(n3767) );
  AOI22D1BWP12T U2977 ( .A1(b[1]), .A2(n2375), .B1(n2374), .B2(n3165), .ZN(
        n2425) );
  AOI22D1BWP12T U2978 ( .A1(b[1]), .A2(n2377), .B1(n2376), .B2(n3165), .ZN(
        n2428) );
  AOI22D1BWP12T U2979 ( .A1(b[2]), .A2(n2425), .B1(n2428), .B2(n2652), .ZN(
        n2890) );
  AOI22D1BWP12T U2980 ( .A1(b[1]), .A2(n2379), .B1(n2378), .B2(n3165), .ZN(
        n2427) );
  OAI22D1BWP12T U2981 ( .A1(n3170), .A2(n3380), .B1(n3346), .B2(b[0]), .ZN(
        n2398) );
  MAOI22D0BWP12T U2982 ( .A1(b[1]), .A2(n2380), .B1(n2398), .B2(b[1]), .ZN(
        n2431) );
  AOI22D1BWP12T U2983 ( .A1(b[2]), .A2(n2427), .B1(n2431), .B2(n2652), .ZN(
        n2891) );
  OAI22D1BWP12T U2984 ( .A1(n2890), .A2(n2662), .B1(n2891), .B2(n2914), .ZN(
        n2558) );
  AOI21D1BWP12T U2985 ( .A1(b[4]), .A2(n3767), .B(n2558), .ZN(n3353) );
  NR2D1BWP12T U2986 ( .A1(n3353), .A2(n2626), .ZN(n3356) );
  AOI22D1BWP12T U2987 ( .A1(b[0]), .A2(n3685), .B1(n3632), .B2(n3170), .ZN(
        n2395) );
  OAI22D1BWP12T U2988 ( .A1(n3170), .A2(a[19]), .B1(a[18]), .B2(b[0]), .ZN(
        n2385) );
  MAOI22D0BWP12T U2989 ( .A1(b[1]), .A2(n2395), .B1(n2385), .B2(b[1]), .ZN(
        n2401) );
  OAI22D1BWP12T U2990 ( .A1(n3170), .A2(a[17]), .B1(a[16]), .B2(b[0]), .ZN(
        n2384) );
  OAI22D1BWP12T U2991 ( .A1(n3170), .A2(a[15]), .B1(a[14]), .B2(b[0]), .ZN(
        n2387) );
  OA22D1BWP12T U2992 ( .A1(n2593), .A2(n2384), .B1(n2387), .B2(b[1]), .Z(n2405) );
  AOI22D1BWP12T U2993 ( .A1(b[2]), .A2(n2401), .B1(n2405), .B2(n2652), .ZN(
        n2434) );
  OAI22D1BWP12T U2994 ( .A1(n3170), .A2(a[13]), .B1(a[12]), .B2(b[0]), .ZN(
        n2386) );
  OAI22D1BWP12T U2995 ( .A1(n3170), .A2(a[11]), .B1(a[10]), .B2(b[0]), .ZN(
        n2389) );
  OA22D1BWP12T U2996 ( .A1(n2593), .A2(n2386), .B1(n2389), .B2(b[1]), .Z(n2404) );
  NR2D1BWP12T U2997 ( .A1(n2652), .A2(b[3]), .ZN(n2456) );
  INVD1BWP12T U2998 ( .I(n2456), .ZN(n2399) );
  NR2D1BWP12T U2999 ( .A1(b[3]), .A2(b[2]), .ZN(n2860) );
  OAI22D1BWP12T U3000 ( .A1(n3170), .A2(a[9]), .B1(a[8]), .B2(b[0]), .ZN(n2388) );
  OAI22D1BWP12T U3001 ( .A1(n3170), .A2(a[7]), .B1(a[6]), .B2(b[0]), .ZN(n2390) );
  OAI22D1BWP12T U3002 ( .A1(n2593), .A2(n2388), .B1(n2390), .B2(b[1]), .ZN(
        n2406) );
  MOAI22D0BWP12T U3003 ( .A1(n2404), .A2(n2399), .B1(n2860), .B2(n2406), .ZN(
        n2381) );
  AO211D1BWP12T U3004 ( .A1(b[3]), .A2(n2434), .B(b[4]), .C(n2381), .Z(n2850)
         );
  AOI22D1BWP12T U3005 ( .A1(b[0]), .A2(a[31]), .B1(a[30]), .B2(n2534), .ZN(
        n2870) );
  INVD1BWP12T U3006 ( .I(n2849), .ZN(n2878) );
  AOI22D1BWP12T U3007 ( .A1(b[0]), .A2(a[29]), .B1(a[28]), .B2(n3170), .ZN(
        n2392) );
  OAI22D1BWP12T U3008 ( .A1(n3170), .A2(n3824), .B1(n3790), .B2(b[0]), .ZN(
        n2394) );
  MAOI22D0BWP12T U3009 ( .A1(b[1]), .A2(n2392), .B1(n2394), .B2(b[1]), .ZN(
        n2400) );
  OAI22D1BWP12T U3010 ( .A1(n3170), .A2(n3768), .B1(n2518), .B2(b[0]), .ZN(
        n2393) );
  OAI22D1BWP12T U3011 ( .A1(n3170), .A2(n3701), .B1(n3684), .B2(b[0]), .ZN(
        n2396) );
  OAI22D1BWP12T U3012 ( .A1(n2593), .A2(n2393), .B1(n2396), .B2(b[1]), .ZN(
        n2402) );
  MAOI22D0BWP12T U3013 ( .A1(b[2]), .A2(n2400), .B1(n2402), .B2(b[2]), .ZN(
        n2433) );
  OAI32D1BWP12T U3014 ( .A1(n2886), .A2(n2870), .A3(n2878), .B1(b[3]), .B2(
        n2433), .ZN(n3679) );
  INVD1BWP12T U3015 ( .I(n3679), .ZN(n2443) );
  ND2D1BWP12T U3016 ( .A1(b[4]), .A2(n2443), .ZN(n2851) );
  ND2D1BWP12T U3017 ( .A1(n2850), .A2(n2851), .ZN(n2472) );
  IND2D1BWP12T U3018 ( .A1(n2472), .B1(n3144), .ZN(n3266) );
  AOI211D1BWP12T U3019 ( .A1(b[1]), .A2(n3194), .B(n2383), .C(n2382), .ZN(
        n2565) );
  ND2D1BWP12T U3020 ( .A1(n2565), .A2(n2886), .ZN(n2479) );
  NR2D1BWP12T U3021 ( .A1(n2626), .A2(b[4]), .ZN(n3199) );
  INVD1BWP12T U3022 ( .I(n3199), .ZN(n3908) );
  AOI32D1BWP12T U3023 ( .A1(n2564), .A2(n3266), .A3(n2479), .B1(n3908), .B2(
        n3266), .ZN(n2467) );
  AOI22D1BWP12T U3024 ( .A1(b[1]), .A2(n2385), .B1(n2384), .B2(n3165), .ZN(
        n2419) );
  AOI22D1BWP12T U3025 ( .A1(b[1]), .A2(n2387), .B1(n2386), .B2(n3165), .ZN(
        n2411) );
  AOI22D1BWP12T U3026 ( .A1(b[2]), .A2(n2419), .B1(n2411), .B2(n2652), .ZN(
        n2494) );
  AOI22D1BWP12T U3027 ( .A1(b[1]), .A2(n2389), .B1(n2388), .B2(n3165), .ZN(
        n2410) );
  OAI22D1BWP12T U3028 ( .A1(n3170), .A2(n3247), .B1(n3218), .B2(b[0]), .ZN(
        n2403) );
  MAOI22D0BWP12T U3029 ( .A1(b[1]), .A2(n2390), .B1(n2403), .B2(b[1]), .ZN(
        n2412) );
  AOI22D1BWP12T U3030 ( .A1(n2456), .A2(n2410), .B1(n2860), .B2(n2412), .ZN(
        n2391) );
  OA211D1BWP12T U3031 ( .A1(n2494), .A2(n2886), .B(n2391), .C(n3219), .Z(n2897) );
  OAI22D1BWP12T U3032 ( .A1(n3165), .A2(n2870), .B1(n2392), .B2(b[1]), .ZN(
        n2421) );
  AN2D1BWP12T U3033 ( .A1(n2421), .A2(n2652), .Z(n2862) );
  AOI22D1BWP12T U3034 ( .A1(b[1]), .A2(n2394), .B1(n2393), .B2(n3165), .ZN(
        n2417) );
  AOI22D1BWP12T U3035 ( .A1(b[1]), .A2(n2396), .B1(n2395), .B2(n3165), .ZN(
        n2418) );
  AOI22D1BWP12T U3036 ( .A1(b[2]), .A2(n2417), .B1(n2418), .B2(n2652), .ZN(
        n2493) );
  AOI22D1BWP12T U3037 ( .A1(b[3]), .A2(n2862), .B1(n2493), .B2(n2886), .ZN(
        n3637) );
  INVD1BWP12T U3038 ( .I(n3637), .ZN(n2441) );
  NR2D1BWP12T U3039 ( .A1(n3219), .A2(n2441), .ZN(n2899) );
  NR2D1BWP12T U3040 ( .A1(n2897), .A2(n2899), .ZN(n2478) );
  AN2D1BWP12T U3041 ( .A1(n2478), .A2(n3144), .Z(n3216) );
  AOI22D1BWP12T U3042 ( .A1(b[3]), .A2(n2397), .B1(n2496), .B2(n2886), .ZN(
        n2440) );
  ND2D1BWP12T U3043 ( .A1(n3165), .A2(n2860), .ZN(n2867) );
  INVD1BWP12T U3044 ( .I(n2867), .ZN(n2906) );
  AOI22D1BWP12T U3045 ( .A1(b[0]), .A2(n3218), .B1(n2471), .B2(n3170), .ZN(
        n2448) );
  AOI22D1BWP12T U3046 ( .A1(b[0]), .A2(a[6]), .B1(a[5]), .B2(n3170), .ZN(n2429) );
  INVD1BWP12T U3047 ( .I(n2860), .ZN(n2847) );
  OAI22D1BWP12T U3048 ( .A1(n3170), .A2(a[8]), .B1(a[7]), .B2(b[0]), .ZN(n2430) );
  MAOI22D0BWP12T U3049 ( .A1(b[1]), .A2(n2398), .B1(n2430), .B2(b[1]), .ZN(
        n2455) );
  NR2D1BWP12T U3050 ( .A1(n2626), .A2(n2500), .ZN(n3997) );
  ND2D1BWP12T U3051 ( .A1(n2508), .A2(n2625), .ZN(n3883) );
  AN2D1BWP12T U3052 ( .A1(n3997), .A2(n3883), .Z(n3983) );
  ND2D1BWP12T U3053 ( .A1(n2652), .A2(n2400), .ZN(n2871) );
  OAI31D1BWP12T U3054 ( .A1(n2652), .A2(n2870), .A3(b[1]), .B(n2871), .ZN(
        n3783) );
  AOI22D1BWP12T U3055 ( .A1(b[2]), .A2(n2402), .B1(n2401), .B2(n2652), .ZN(
        n2556) );
  INVD1BWP12T U3056 ( .I(n2556), .ZN(n2422) );
  ND2D1BWP12T U3057 ( .A1(n2886), .A2(n2422), .ZN(n2884) );
  OAI21D1BWP12T U3058 ( .A1(n2886), .A2(n3783), .B(n2884), .ZN(n3581) );
  OAI22D1BWP12T U3059 ( .A1(n3170), .A2(n2471), .B1(n3961), .B2(b[0]), .ZN(
        n2414) );
  INVD1BWP12T U3060 ( .I(n2414), .ZN(n2409) );
  AOI31D1BWP12T U3061 ( .A1(b[1]), .A2(n2860), .A3(n2403), .B(b[4]), .ZN(n2408) );
  AOI22D1BWP12T U3062 ( .A1(b[2]), .A2(n2405), .B1(n2404), .B2(n2652), .ZN(
        n2557) );
  AOI22D1BWP12T U3063 ( .A1(b[3]), .A2(n2557), .B1(n2456), .B2(n2406), .ZN(
        n2407) );
  OA211D1BWP12T U3064 ( .A1(n2409), .A2(n2867), .B(n2408), .C(n2407), .Z(n2887) );
  AOI21D1BWP12T U3065 ( .A1(n3581), .A2(b[4]), .B(n2887), .ZN(n3968) );
  AN2D1BWP12T U3066 ( .A1(n3968), .A2(n3144), .Z(n3967) );
  NR2D1BWP12T U3067 ( .A1(n3155), .A2(n2867), .ZN(n3158) );
  OAI22D1BWP12T U3068 ( .A1(n2652), .A2(n2411), .B1(n2410), .B2(b[2]), .ZN(
        n2566) );
  MAOI22D0BWP12T U3069 ( .A1(n2456), .A2(n2412), .B1(n2886), .B2(n2566), .ZN(
        n2416) );
  NR2D1BWP12T U3070 ( .A1(n2512), .A2(n2847), .ZN(n2447) );
  OAI211D1BWP12T U3071 ( .A1(n3165), .A2(n2414), .B(n2447), .C(n2413), .ZN(
        n2415) );
  ND2D1BWP12T U3072 ( .A1(n2416), .A2(n2415), .ZN(n2420) );
  MAOI22D0BWP12T U3073 ( .A1(b[2]), .A2(n2421), .B1(n2417), .B2(b[2]), .ZN(
        n2424) );
  MAOI22D0BWP12T U3074 ( .A1(n2419), .A2(n2652), .B1(n2652), .B2(n2418), .ZN(
        n2497) );
  AOI22D1BWP12T U3075 ( .A1(b[3]), .A2(n2424), .B1(n2497), .B2(n2886), .ZN(
        n2905) );
  OAI32D1BWP12T U3076 ( .A1(b[4]), .A2(n3158), .A3(n2420), .B1(n2905), .B2(
        n3219), .ZN(n3162) );
  NR2D1BWP12T U3077 ( .A1(n3162), .A2(n2626), .ZN(n2866) );
  NR4D0BWP12T U3078 ( .A1(n3216), .A2(n3983), .A3(n3967), .A4(n2866), .ZN(
        n2465) );
  MAOI22D0BWP12T U3079 ( .A1(n3784), .A2(n2494), .B1(n2662), .B2(n2493), .ZN(
        n2848) );
  ND2D1BWP12T U3080 ( .A1(n2860), .A2(n2421), .ZN(n3855) );
  ND2D1BWP12T U3081 ( .A1(b[4]), .A2(n3855), .ZN(n2483) );
  ND2D1BWP12T U3082 ( .A1(n2848), .A2(n2483), .ZN(n3421) );
  NR2D1BWP12T U3083 ( .A1(n2626), .A2(n3421), .ZN(n3427) );
  ND2D1BWP12T U3084 ( .A1(n2886), .A2(n3783), .ZN(n3791) );
  MAOI22D0BWP12T U3085 ( .A1(n2912), .A2(n2422), .B1(n2914), .B2(n2557), .ZN(
        n2423) );
  ND2D1BWP12T U3086 ( .A1(n3144), .A2(n2423), .ZN(n2888) );
  AOI21D1BWP12T U3087 ( .A1(b[4]), .A2(n3791), .B(n2888), .ZN(n3365) );
  NR2D1BWP12T U3088 ( .A1(b[3]), .A2(n2424), .ZN(n2875) );
  AOI22D1BWP12T U3089 ( .A1(n3784), .A2(n2566), .B1(n2912), .B2(n2497), .ZN(
        n2876) );
  OAI21D1BWP12T U3090 ( .A1(n2875), .A2(n3219), .B(n2876), .ZN(n3314) );
  NR2D1BWP12T U3091 ( .A1(n2626), .A2(n3314), .ZN(n3316) );
  MAOI22D0BWP12T U3092 ( .A1(b[2]), .A2(n2426), .B1(n2425), .B2(b[2]), .ZN(
        n2492) );
  AN2D1BWP12T U3093 ( .A1(n2492), .A2(n2886), .Z(n2879) );
  AOI21D1BWP12T U3094 ( .A1(n2565), .A2(b[3]), .B(n2879), .ZN(n3653) );
  INVD1BWP12T U3095 ( .I(n3653), .ZN(n2503) );
  NR2D1BWP12T U3096 ( .A1(n3219), .A2(n2503), .ZN(n2475) );
  AOI22D1BWP12T U3097 ( .A1(b[2]), .A2(n2428), .B1(n2427), .B2(n2652), .ZN(
        n2439) );
  AOI22D1BWP12T U3098 ( .A1(b[1]), .A2(n2430), .B1(n2429), .B2(n3165), .ZN(
        n2449) );
  AOI22D1BWP12T U3099 ( .A1(n2431), .A2(n2456), .B1(n2860), .B2(n2449), .ZN(
        n2432) );
  OAI211D1BWP12T U3100 ( .A1(n2439), .A2(n2886), .B(n2432), .C(n3219), .ZN(
        n2473) );
  ND2D1BWP12T U3101 ( .A1(n3144), .A2(n2473), .ZN(n2883) );
  NR2D1BWP12T U3102 ( .A1(n2475), .A2(n2883), .ZN(n3253) );
  NR4D0BWP12T U3103 ( .A1(n3427), .A2(n3365), .A3(n3316), .A4(n3253), .ZN(
        n2464) );
  NR2D1BWP12T U3104 ( .A1(n2870), .A2(n2867), .ZN(n2907) );
  INVD1BWP12T U3105 ( .I(n2907), .ZN(n3921) );
  MOAI22D0BWP12T U3106 ( .A1(n2914), .A2(n2434), .B1(n2912), .B2(n2433), .ZN(
        n2908) );
  AO21D1BWP12T U3107 ( .A1(n3921), .A2(b[4]), .B(n2908), .Z(n3475) );
  NR2D1BWP12T U3108 ( .A1(n2626), .A2(n3475), .ZN(n3478) );
  OAI22D1BWP12T U3109 ( .A1(n2652), .A2(n2436), .B1(n2435), .B2(b[2]), .ZN(
        n2915) );
  INVD1BWP12T U3110 ( .I(n2915), .ZN(n2458) );
  AOI22D1BWP12T U3111 ( .A1(b[2]), .A2(n2438), .B1(n2437), .B2(n2652), .ZN(
        n2911) );
  ND2D1BWP12T U3112 ( .A1(n2512), .A2(n2860), .ZN(n2486) );
  NR2D1BWP12T U3113 ( .A1(n3194), .A2(n2486), .ZN(n2442) );
  OAI222D1BWP12T U3114 ( .A1(n2458), .A2(n2914), .B1(n2662), .B2(n2911), .C1(
        n3219), .C2(n2442), .ZN(n3505) );
  NR2D1BWP12T U3115 ( .A1(n2626), .A2(n3505), .ZN(n3510) );
  INVD1BWP12T U3116 ( .I(n2439), .ZN(n2491) );
  OAI22D1BWP12T U3117 ( .A1(n2914), .A2(n2491), .B1(n2662), .B2(n2492), .ZN(
        n2909) );
  AO21D1BWP12T U3118 ( .A1(n2479), .A2(b[4]), .B(n2909), .Z(n3452) );
  NR2D1BWP12T U3119 ( .A1(n2626), .A2(n3452), .ZN(n3456) );
  ND2D1BWP12T U3120 ( .A1(op[0]), .A2(op[1]), .ZN(n2926) );
  INVD1BWP12T U3121 ( .I(n2926), .ZN(n2489) );
  NR2D1BWP12T U3122 ( .A1(op[3]), .A2(op[2]), .ZN(n2754) );
  ND2D1BWP12T U3123 ( .A1(n2489), .A2(n2754), .ZN(n3265) );
  NR4D0BWP12T U3124 ( .A1(n3478), .A2(n3510), .A3(n3456), .A4(n3265), .ZN(
        n2463) );
  INVD1BWP12T U3125 ( .I(n2440), .ZN(n2903) );
  AOI21D1BWP12T U3126 ( .A1(b[3]), .A2(n2508), .B(n2903), .ZN(n3610) );
  NR3D1BWP12T U3127 ( .A1(n2905), .A2(n3610), .A3(n2441), .ZN(n2577) );
  INVD1BWP12T U3128 ( .I(n2442), .ZN(n3201) );
  ND3D1BWP12T U3129 ( .A1(n3201), .A2(n3921), .A3(n3855), .ZN(n2567) );
  INVD1BWP12T U3130 ( .I(n2875), .ZN(n3732) );
  NR2D1BWP12T U3131 ( .A1(b[3]), .A2(n2890), .ZN(n2446) );
  AOI21D1BWP12T U3132 ( .A1(n2444), .A2(b[3]), .B(n2446), .ZN(n2852) );
  RCIAO21D0BWP12T U3133 ( .A1(n2446), .A2(n2445), .B(n2852), .ZN(n2454) );
  INVD1BWP12T U3134 ( .I(n2454), .ZN(n3558) );
  NR2D1BWP12T U3135 ( .A1(n3194), .A2(n2886), .ZN(n2874) );
  AOI21D1BWP12T U3136 ( .A1(n2886), .A2(n2911), .B(n2874), .ZN(n2459) );
  INVD1BWP12T U3137 ( .I(n2459), .ZN(n2854) );
  ND2D1BWP12T U3138 ( .A1(n2512), .A2(n2652), .ZN(n2468) );
  ND2D1BWP12T U3139 ( .A1(b[3]), .A2(n2468), .ZN(n2482) );
  ND2D1BWP12T U3140 ( .A1(n2854), .A2(n2482), .ZN(n3702) );
  INVD1BWP12T U3141 ( .I(n2891), .ZN(n2453) );
  OA221D1BWP12T U3142 ( .A1(n2448), .A2(n3165), .B1(a[2]), .B2(b[1]), .C(n2447), .Z(n2452) );
  ND2D1BWP12T U3143 ( .A1(a[1]), .A2(n2534), .ZN(n2450) );
  MOAI22D0BWP12T U3144 ( .A1(n2867), .A2(n2450), .B1(n2456), .B2(n2449), .ZN(
        n2451) );
  AOI211D1BWP12T U3145 ( .A1(b[3]), .A2(n2453), .B(n2452), .C(n2451), .ZN(
        n2490) );
  ND2D1BWP12T U3146 ( .A1(n2490), .A2(n3219), .ZN(n2853) );
  OAI21D1BWP12T U3147 ( .A1(n2454), .A2(n3219), .B(n2853), .ZN(n3186) );
  NR2D1BWP12T U3148 ( .A1(n2626), .A2(n3186), .ZN(n3189) );
  MAOI22D0BWP12T U3149 ( .A1(n2457), .A2(n2456), .B1(n2847), .B2(n2455), .ZN(
        n2461) );
  ND2D1BWP12T U3150 ( .A1(b[3]), .A2(n2458), .ZN(n2460) );
  AOI32D1BWP12T U3151 ( .A1(n2461), .A2(n3219), .A3(n2460), .B1(n2459), .B2(
        b[4]), .ZN(n2896) );
  ND2D1BWP12T U3152 ( .A1(n2625), .A2(n2468), .ZN(n3550) );
  ND2D1BWP12T U3153 ( .A1(n2896), .A2(n3550), .ZN(n2488) );
  NR2D1BWP12T U3154 ( .A1(n2626), .A2(n2488), .ZN(n3308) );
  ND4D1BWP12T U3155 ( .A1(n2465), .A2(n2464), .A3(n2463), .A4(n2462), .ZN(
        n2466) );
  NR4D0BWP12T U3156 ( .A1(n3405), .A2(n3356), .A3(n2467), .A4(n2466), .ZN(
        n2937) );
  ND2D1BWP12T U3157 ( .A1(n2469), .A2(n2468), .ZN(n2571) );
  OAI22D1BWP12T U3158 ( .A1(n3170), .A2(n2470), .B1(n3961), .B2(b[0]), .ZN(
        n2594) );
  MOAI22D0BWP12T U3159 ( .A1(n2593), .A2(n3155), .B1(n2594), .B2(n3878), .ZN(
        n3969) );
  INVD1BWP12T U3160 ( .I(n3969), .ZN(n2487) );
  OAI22D1BWP12T U3161 ( .A1(n3170), .A2(n2471), .B1(n3218), .B2(b[0]), .ZN(
        n2596) );
  OAI22D1BWP12T U3162 ( .A1(n3170), .A2(n3247), .B1(n3276), .B2(b[0]), .ZN(
        n2595) );
  OAI22D1BWP12T U3163 ( .A1(n3878), .A2(n2596), .B1(n2595), .B2(n2570), .ZN(
        n2507) );
  INVD1BWP12T U3164 ( .I(n2571), .ZN(n2573) );
  OAI22D1BWP12T U3165 ( .A1(n2571), .A2(n2487), .B1(n2507), .B2(n2573), .ZN(
        n2526) );
  INVD1BWP12T U3166 ( .I(n3550), .ZN(n2575) );
  IOA21D1BWP12T U3167 ( .A1(n2526), .A2(n2575), .B(n2472), .ZN(n3262) );
  INVD1BWP12T U3168 ( .I(n2473), .ZN(n2476) );
  OAI22D1BWP12T U3169 ( .A1(n3170), .A2(n3218), .B1(n3247), .B2(b[0]), .ZN(
        n2610) );
  AOI22D1BWP12T U3170 ( .A1(b[0]), .A2(a[2]), .B1(a[3]), .B2(n3170), .ZN(n2609) );
  MOAI22D0BWP12T U3171 ( .A1(n2610), .A2(n3881), .B1(n2570), .B2(n2609), .ZN(
        n2517) );
  AOI21D1BWP12T U3172 ( .A1(a[1]), .A2(n2534), .B(n2474), .ZN(n2620) );
  NR2D1BWP12T U3173 ( .A1(n2620), .A2(n3881), .ZN(n3187) );
  MOAI22D0BWP12T U3174 ( .A1(n2517), .A2(n2573), .B1(n2573), .B2(n3187), .ZN(
        n2543) );
  MOAI22D0BWP12T U3175 ( .A1(n2476), .A2(n2475), .B1(n2543), .B2(n2575), .ZN(
        n3237) );
  AOI22D1BWP12T U3176 ( .A1(n2570), .A2(n2594), .B1(n2596), .B2(n3878), .ZN(
        n2480) );
  ND2D1BWP12T U3177 ( .A1(b[2]), .A2(n2593), .ZN(n2477) );
  OAI22D1BWP12T U3178 ( .A1(n2573), .A2(n2480), .B1(n3155), .B2(n2477), .ZN(
        n2576) );
  AOI21D1BWP12T U3179 ( .A1(n2575), .A2(n2576), .B(n2478), .ZN(n3231) );
  INVD1BWP12T U3180 ( .I(n2479), .ZN(n3873) );
  OAI22D1BWP12T U3181 ( .A1(n3170), .A2(n3346), .B1(n3380), .B2(b[0]), .ZN(
        n2597) );
  AOI22D1BWP12T U3182 ( .A1(b[0]), .A2(a[11]), .B1(a[12]), .B2(n3170), .ZN(
        n2600) );
  MOAI22D0BWP12T U3183 ( .A1(n3878), .A2(n2597), .B1(n2600), .B2(n3878), .ZN(
        n2548) );
  AOI22D1BWP12T U3184 ( .A1(b[0]), .A2(a[13]), .B1(a[14]), .B2(n3170), .ZN(
        n2599) );
  AOI22D1BWP12T U3185 ( .A1(b[0]), .A2(a[15]), .B1(a[16]), .B2(n3170), .ZN(
        n2602) );
  AO22D1BWP12T U3186 ( .A1(n2570), .A2(n2599), .B1(n2602), .B2(n3878), .Z(
        n2572) );
  OA22D1BWP12T U3187 ( .A1(n2571), .A2(n2548), .B1(n2572), .B2(n2573), .Z(
        n3741) );
  ND2D1BWP12T U3188 ( .A1(n2486), .A2(n2482), .ZN(n2559) );
  INVD1BWP12T U3189 ( .I(n2559), .ZN(n2561) );
  AOI22D1BWP12T U3190 ( .A1(b[0]), .A2(n3292), .B1(n3321), .B2(n3170), .ZN(
        n2598) );
  AOI22D1BWP12T U3191 ( .A1(n2570), .A2(n2595), .B1(n2598), .B2(n3878), .ZN(
        n2549) );
  ND2D1BWP12T U3192 ( .A1(n2549), .A2(n2571), .ZN(n2562) );
  ND2D1BWP12T U3193 ( .A1(n2573), .A2(n2480), .ZN(n2560) );
  AOI31D1BWP12T U3194 ( .A1(n2561), .A2(n2562), .A3(n2560), .B(n3158), .ZN(
        n2481) );
  OAI21D1BWP12T U3195 ( .A1(n3741), .A2(n2482), .B(n2481), .ZN(n3525) );
  NR3D1BWP12T U3196 ( .A1(n3873), .A2(n2483), .A3(n3525), .ZN(n2484) );
  AOI32D1BWP12T U3197 ( .A1(n3219), .A2(n3231), .A3(n3581), .B1(n2484), .B2(
        n3231), .ZN(n2541) );
  AOI22D1BWP12T U3198 ( .A1(b[0]), .A2(a[10]), .B1(a[11]), .B2(n3170), .ZN(
        n2614) );
  OAI22D1BWP12T U3199 ( .A1(n3170), .A2(n3321), .B1(n3346), .B2(b[0]), .ZN(
        n2611) );
  MAOI22D0BWP12T U3200 ( .A1(n2614), .A2(n3878), .B1(n3878), .B2(n2611), .ZN(
        n2544) );
  OAI22D1BWP12T U3201 ( .A1(n3170), .A2(n3428), .B1(n3446), .B2(b[0]), .ZN(
        n2588) );
  OAI22D1BWP12T U3202 ( .A1(n3170), .A2(n3479), .B1(n2485), .B2(b[0]), .ZN(
        n2587) );
  OAI22D1BWP12T U3203 ( .A1(n3878), .A2(n2588), .B1(n2587), .B2(n2570), .ZN(
        n2554) );
  MAOI22D0BWP12T U3204 ( .A1(n2573), .A2(n2544), .B1(n2554), .B2(n2573), .ZN(
        n2531) );
  NR2D1BWP12T U3205 ( .A1(n3219), .A2(n2559), .ZN(n3889) );
  INVD1BWP12T U3206 ( .I(n3889), .ZN(n3814) );
  AOI22D1BWP12T U3207 ( .A1(n2570), .A2(n2725), .B1(n2609), .B2(n3878), .ZN(
        n3979) );
  OAI22D1BWP12T U3208 ( .A1(n3170), .A2(n3276), .B1(n3292), .B2(b[0]), .ZN(
        n2612) );
  OA22D1BWP12T U3209 ( .A1(n3878), .A2(n2610), .B1(n2612), .B2(n2570), .Z(
        n2545) );
  AOI22D1BWP12T U3210 ( .A1(n2573), .A2(n3979), .B1(n2545), .B2(n2571), .ZN(
        n2532) );
  ND2D1BWP12T U3211 ( .A1(b[4]), .A2(n2486), .ZN(n3506) );
  INVD1BWP12T U3212 ( .I(n3506), .ZN(n3818) );
  NR3D1BWP12T U3213 ( .A1(n3784), .A2(n2561), .A3(n3818), .ZN(n3585) );
  INVD1BWP12T U3214 ( .I(n3585), .ZN(n3603) );
  OAI22D1BWP12T U3215 ( .A1(n3170), .A2(n3529), .B1(n3565), .B2(b[0]), .ZN(
        n2589) );
  OAI22D1BWP12T U3216 ( .A1(n3170), .A2(n3578), .B1(n3618), .B2(b[0]), .ZN(
        n2608) );
  OAI22D1BWP12T U3217 ( .A1(n3878), .A2(n2589), .B1(n2608), .B2(n2570), .ZN(
        n2553) );
  OAI22D1BWP12T U3218 ( .A1(n2534), .A2(n3684), .B1(n3701), .B2(b[0]), .ZN(
        n2606) );
  INVD1BWP12T U3219 ( .I(n2606), .ZN(n2519) );
  OAI22D1BWP12T U3220 ( .A1(n2534), .A2(n3632), .B1(n3685), .B2(b[0]), .ZN(
        n2607) );
  MAOI22D0BWP12T U3221 ( .A1(n2519), .A2(n3878), .B1(n3878), .B2(n2607), .ZN(
        n3816) );
  MOAI22D0BWP12T U3222 ( .A1(n2571), .A2(n2553), .B1(n3816), .B2(n2571), .ZN(
        n2533) );
  NR2D1BWP12T U3223 ( .A1(n2573), .A2(n2487), .ZN(n3586) );
  OAI21D1BWP12T U3224 ( .A1(n3550), .A2(n2532), .B(n2488), .ZN(n3298) );
  ND2D1BWP12T U3225 ( .A1(n3268), .A2(n2489), .ZN(n3891) );
  INVD1BWP12T U3226 ( .I(n3891), .ZN(n3981) );
  ND2D1BWP12T U3227 ( .A1(n3187), .A2(n2571), .ZN(n3549) );
  ND4D1BWP12T U3228 ( .A1(n2490), .A2(n3981), .A3(n3791), .A4(n3549), .ZN(
        n2499) );
  INR4D0BWP12T U3229 ( .A1(n2494), .B1(n2493), .B2(n2492), .B3(n2491), .ZN(
        n2495) );
  ND4D1BWP12T U3230 ( .A1(n2497), .A2(n2496), .A3(n2495), .A4(n3732), .ZN(
        n2498) );
  NR4D0BWP12T U3231 ( .A1(n3586), .A2(n3298), .A3(n2499), .A4(n2498), .ZN(
        n2539) );
  INVD1BWP12T U3232 ( .I(n3883), .ZN(n3980) );
  NR2D1BWP12T U3233 ( .A1(n3980), .A2(n2500), .ZN(n3978) );
  AOI22D1BWP12T U3234 ( .A1(n2570), .A2(n2598), .B1(n2597), .B2(n3878), .ZN(
        n2506) );
  OAI22D1BWP12T U3235 ( .A1(n3878), .A2(n2600), .B1(n2599), .B2(n2570), .ZN(
        n2511) );
  MAOI22D0BWP12T U3236 ( .A1(n2573), .A2(n2506), .B1(n2511), .B2(n2573), .ZN(
        n2525) );
  AOI22D1BWP12T U3237 ( .A1(n3889), .A2(n2525), .B1(n3219), .B2(n3679), .ZN(
        n2502) );
  AOI22D1BWP12T U3238 ( .A1(b[0]), .A2(n3618), .B1(n3632), .B2(n2534), .ZN(
        n2592) );
  AOI22D1BWP12T U3239 ( .A1(b[0]), .A2(n3685), .B1(n3684), .B2(n2534), .ZN(
        n3740) );
  AOI22D1BWP12T U3240 ( .A1(n2570), .A2(n2592), .B1(n3740), .B2(n3878), .ZN(
        n2509) );
  OAI22D1BWP12T U3241 ( .A1(n2534), .A2(a[17]), .B1(a[18]), .B2(b[0]), .ZN(
        n2601) );
  OAI22D1BWP12T U3242 ( .A1(n3878), .A2(n2602), .B1(n2601), .B2(n2570), .ZN(
        n2510) );
  MAOI22D0BWP12T U3243 ( .A1(n2509), .A2(n2571), .B1(n2571), .B2(n2510), .ZN(
        n2528) );
  AOI22D1BWP12T U3244 ( .A1(n2575), .A2(n2528), .B1(n3585), .B2(n2526), .ZN(
        n2501) );
  ND2D1BWP12T U3245 ( .A1(n2502), .A2(n2501), .ZN(n3680) );
  AOI22D1BWP12T U3246 ( .A1(n2570), .A2(n2612), .B1(n2611), .B2(n3878), .ZN(
        n2516) );
  INVD1BWP12T U3247 ( .I(n2588), .ZN(n2613) );
  OAI22D1BWP12T U3248 ( .A1(n3878), .A2(n2614), .B1(n2613), .B2(n2570), .ZN(
        n2521) );
  MAOI22D0BWP12T U3249 ( .A1(n2573), .A2(n2516), .B1(n2521), .B2(n2573), .ZN(
        n2542) );
  AOI22D1BWP12T U3250 ( .A1(n3889), .A2(n2542), .B1(n3219), .B2(n2503), .ZN(
        n2505) );
  AOI22D1BWP12T U3251 ( .A1(n2570), .A2(n2608), .B1(n2607), .B2(n3878), .ZN(
        n2522) );
  INVD1BWP12T U3252 ( .I(n2587), .ZN(n2616) );
  INVD1BWP12T U3253 ( .I(n2589), .ZN(n2615) );
  OAI22D1BWP12T U3254 ( .A1(n3878), .A2(n2616), .B1(n2615), .B2(n2570), .ZN(
        n2520) );
  MAOI22D0BWP12T U3255 ( .A1(n2522), .A2(n2571), .B1(n2571), .B2(n2520), .ZN(
        n3888) );
  AOI22D1BWP12T U3256 ( .A1(n2575), .A2(n3888), .B1(n3585), .B2(n2543), .ZN(
        n2504) );
  ND2D1BWP12T U3257 ( .A1(n2505), .A2(n2504), .ZN(n3662) );
  NR4D0BWP12T U3258 ( .A1(n3968), .A2(n3978), .A3(n3680), .A4(n3662), .ZN(
        n2538) );
  AOI22D1BWP12T U3259 ( .A1(n2573), .A2(n2507), .B1(n2506), .B2(n2571), .ZN(
        n2551) );
  AOI22D1BWP12T U3260 ( .A1(n2561), .A2(n3586), .B1(n2551), .B2(n2559), .ZN(
        n3368) );
  NR2D1BWP12T U3261 ( .A1(n3550), .A2(n2508), .ZN(n3877) );
  INVD1BWP12T U3262 ( .I(n3877), .ZN(n3836) );
  INVD1BWP12T U3263 ( .I(n2509), .ZN(n2514) );
  AOI22D1BWP12T U3264 ( .A1(b[0]), .A2(n3701), .B1(n2518), .B2(n2534), .ZN(
        n3739) );
  AOI22D1BWP12T U3265 ( .A1(b[0]), .A2(n3768), .B1(n3790), .B2(n2534), .ZN(
        n3843) );
  AOI22D1BWP12T U3266 ( .A1(n2570), .A2(n3739), .B1(n3843), .B2(n3878), .ZN(
        n2527) );
  AOI22D1BWP12T U3267 ( .A1(n2573), .A2(n2511), .B1(n2510), .B2(n2571), .ZN(
        n2552) );
  AOI22D1BWP12T U3268 ( .A1(n3980), .A2(n2527), .B1(n3889), .B2(n2552), .ZN(
        n2513) );
  ND2D1BWP12T U3269 ( .A1(n2652), .A2(n3784), .ZN(n2679) );
  INVD1BWP12T U3270 ( .I(n2679), .ZN(n2635) );
  ND2D1BWP12T U3271 ( .A1(n2512), .A2(n2635), .ZN(n3737) );
  OAI211D1BWP12T U3272 ( .A1(n3836), .A2(n2514), .B(n2513), .C(n3737), .ZN(
        n2515) );
  AOI21D1BWP12T U3273 ( .A1(n3368), .A2(n3506), .B(n2515), .ZN(n3782) );
  AOI22D1BWP12T U3274 ( .A1(n2573), .A2(n2517), .B1(n2516), .B2(n2571), .ZN(
        n3553) );
  MAOI22D0BWP12T U3275 ( .A1(n3553), .A2(n2559), .B1(n2559), .B2(n3549), .ZN(
        n3354) );
  OAI22D1BWP12T U3276 ( .A1(n2534), .A2(n2518), .B1(n3768), .B2(b[0]), .ZN(
        n2605) );
  MAOI22D0BWP12T U3277 ( .A1(n2570), .A2(n2519), .B1(n2605), .B2(n2570), .ZN(
        n3876) );
  AOI22D1BWP12T U3278 ( .A1(n2573), .A2(n2521), .B1(n2520), .B2(n2571), .ZN(
        n3551) );
  AOI22D1BWP12T U3279 ( .A1(n3889), .A2(n3551), .B1(n3877), .B2(n2522), .ZN(
        n2523) );
  OAI211D1BWP12T U3280 ( .A1(n3883), .A2(n3876), .B(n2523), .C(n3737), .ZN(
        n2524) );
  AOI21D1BWP12T U3281 ( .A1(n3354), .A2(n3506), .B(n2524), .ZN(n3775) );
  AOI22D1BWP12T U3282 ( .A1(n2561), .A2(n2526), .B1(n2525), .B2(n2559), .ZN(
        n3476) );
  ND2D1BWP12T U3283 ( .A1(n3506), .A2(n3737), .ZN(n3884) );
  MAOI22D0BWP12T U3284 ( .A1(n3889), .A2(n2528), .B1(n3836), .B2(n2527), .ZN(
        n2530) );
  AOI22D1BWP12T U3285 ( .A1(b[0]), .A2(n3869), .B1(n3932), .B2(n2534), .ZN(
        n2672) );
  AOI22D1BWP12T U3286 ( .A1(b[0]), .A2(n3824), .B1(n3851), .B2(n2534), .ZN(
        n3844) );
  OAI221D1BWP12T U3287 ( .A1(n3881), .A2(n2672), .B1(n3878), .B2(n3844), .C(
        n3980), .ZN(n2529) );
  OAI211D1BWP12T U3288 ( .A1(n3476), .A2(n3884), .B(n2530), .C(n2529), .ZN(
        n3911) );
  AOI22D1BWP12T U3289 ( .A1(b[0]), .A2(n3790), .B1(n3824), .B2(n2534), .ZN(
        n3880) );
  AOI22D1BWP12T U3290 ( .A1(n2570), .A2(n2605), .B1(n3880), .B2(n3878), .ZN(
        n3813) );
  AOI22D1BWP12T U3291 ( .A1(n2561), .A2(n2532), .B1(n2531), .B2(n2559), .ZN(
        n2546) );
  INVD1BWP12T U3292 ( .I(n2546), .ZN(n3507) );
  MAOI22D0BWP12T U3293 ( .A1(n2533), .A2(n3889), .B1(n3884), .B2(n3507), .ZN(
        n2536) );
  AOI22D1BWP12T U3294 ( .A1(b[0]), .A2(n3932), .B1(n3194), .B2(n2534), .ZN(
        n2659) );
  AOI22D1BWP12T U3295 ( .A1(b[0]), .A2(n3851), .B1(n3869), .B2(n2534), .ZN(
        n3879) );
  OAI221D1BWP12T U3296 ( .A1(n3881), .A2(n2659), .B1(n3878), .B2(n3879), .C(
        n3980), .ZN(n2535) );
  OAI211D1BWP12T U3297 ( .A1(n3813), .A2(n3836), .B(n2536), .C(n2535), .ZN(
        n3210) );
  NR4D0BWP12T U3298 ( .A1(n3782), .A2(n3775), .A3(n3911), .A4(n3210), .ZN(
        n2537) );
  ND4D1BWP12T U3299 ( .A1(n3703), .A2(n2539), .A3(n2538), .A4(n2537), .ZN(
        n2540) );
  NR4D0BWP12T U3300 ( .A1(n3262), .A2(n3237), .A3(n2541), .A4(n2540), .ZN(
        n2714) );
  AOI22D1BWP12T U3301 ( .A1(n2561), .A2(n2543), .B1(n2542), .B2(n2559), .ZN(
        n3885) );
  ND2D1BWP12T U3302 ( .A1(n2571), .A2(n3979), .ZN(n3602) );
  AOI22D1BWP12T U3303 ( .A1(n2573), .A2(n2545), .B1(n2544), .B2(n2571), .ZN(
        n2555) );
  AOI22D1BWP12T U3304 ( .A1(n2561), .A2(n3602), .B1(n2555), .B2(n2559), .ZN(
        n3817) );
  INR4D0BWP12T U3305 ( .A1(n3476), .B1(n2547), .B2(n2546), .B3(n3817), .ZN(
        n2550) );
  AOI22D1BWP12T U3306 ( .A1(n2573), .A2(n2549), .B1(n2548), .B2(n2571), .ZN(
        n2574) );
  AOI22D1BWP12T U3307 ( .A1(n2561), .A2(n2576), .B1(n2574), .B2(n2559), .ZN(
        n3835) );
  ND4D1BWP12T U3308 ( .A1(n3885), .A2(n2550), .A3(n3475), .A4(n3835), .ZN(
        n2582) );
  MOAI22D0BWP12T U3309 ( .A1(n3550), .A2(n2552), .B1(n3889), .B2(n2551), .ZN(
        n3584) );
  AOI22D1BWP12T U3310 ( .A1(n2573), .A2(n2554), .B1(n2553), .B2(n2571), .ZN(
        n3815) );
  MAOI22D0BWP12T U3311 ( .A1(n2575), .A2(n3815), .B1(n3814), .B2(n2555), .ZN(
        n3601) );
  AOI22D1BWP12T U3312 ( .A1(n3784), .A2(n2557), .B1(n2912), .B2(n2556), .ZN(
        n3367) );
  IIND4D1BWP12T U3313 ( .A1(n2558), .A2(n3584), .B1(n3601), .B2(n3367), .ZN(
        n2581) );
  AN2D1BWP12T U3314 ( .A1(n2560), .A2(n2559), .Z(n2563) );
  NR2D1BWP12T U3315 ( .A1(n3155), .A2(n2878), .ZN(n2639) );
  OAI22D1BWP12T U3316 ( .A1(n2563), .A2(n2639), .B1(n2562), .B2(n2561), .ZN(
        n3736) );
  ND4D1BWP12T U3317 ( .A1(n3368), .A2(n3354), .A3(n2564), .A4(n3736), .ZN(
        n2580) );
  ND2D1BWP12T U3318 ( .A1(n3784), .A2(n2565), .ZN(n3875) );
  IND4D1BWP12T U3319 ( .A1(n2567), .B1(n2566), .B2(n3875), .B3(n3602), .ZN(
        n2569) );
  IND4D1BWP12T U3320 ( .A1(n2569), .B1(n2568), .B2(n3558), .B3(n3505), .ZN(
        n2578) );
  INVD1BWP12T U3321 ( .I(n2601), .ZN(n2583) );
  AOI22D1BWP12T U3322 ( .A1(n2570), .A2(n2583), .B1(n2592), .B2(n3878), .ZN(
        n3738) );
  AOI22D1BWP12T U3323 ( .A1(n2573), .A2(n2572), .B1(n3738), .B2(n2571), .ZN(
        n3839) );
  AOI222D1BWP12T U3324 ( .A1(n2576), .A2(n3585), .B1(n2575), .B2(n3839), .C1(
        n2574), .C2(n3889), .ZN(n3635) );
  IND4D1BWP12T U3325 ( .A1(n2578), .B1(n3162), .B2(n2577), .B3(n3635), .ZN(
        n2579) );
  NR4D0BWP12T U3326 ( .A1(n2582), .A2(n2581), .A3(n2580), .A4(n2579), .ZN(
        n2713) );
  AOI22D1BWP12T U3327 ( .A1(b[1]), .A2(n2594), .B1(n2596), .B2(n3165), .ZN(
        n2637) );
  OAI32D1BWP12T U3328 ( .A1(n2652), .A2(b[1]), .A3(n3155), .B1(b[2]), .B2(
        n2637), .ZN(n3227) );
  AOI22D1BWP12T U3329 ( .A1(b[1]), .A2(n2595), .B1(n2598), .B2(n3165), .ZN(
        n2638) );
  MOAI22D0BWP12T U3330 ( .A1(n2600), .A2(b[1]), .B1(b[1]), .B2(n2597), .ZN(
        n2642) );
  MAOI22D0BWP12T U3331 ( .A1(b[2]), .A2(n2638), .B1(n2642), .B2(b[2]), .ZN(
        n2687) );
  AOI22D1BWP12T U3332 ( .A1(b[3]), .A2(n3227), .B1(n2687), .B2(n2886), .ZN(
        n2704) );
  AOI22D1BWP12T U3333 ( .A1(b[1]), .A2(n2599), .B1(n2602), .B2(n3165), .ZN(
        n2641) );
  OAI22D1BWP12T U3334 ( .A1(n3165), .A2(n2583), .B1(n2592), .B2(b[1]), .ZN(
        n2636) );
  MAOI22D0BWP12T U3335 ( .A1(b[2]), .A2(n2641), .B1(n2636), .B2(b[2]), .ZN(
        n2688) );
  AOI22D1BWP12T U3336 ( .A1(b[4]), .A2(n2704), .B1(n2912), .B2(n2688), .ZN(
        n2586) );
  NR2D1BWP12T U3337 ( .A1(n2652), .A2(n2914), .ZN(n2684) );
  AOI22D1BWP12T U3338 ( .A1(b[1]), .A2(n3740), .B1(n3739), .B2(n3165), .ZN(
        n2634) );
  AOI221D1BWP12T U3339 ( .A1(n3844), .A2(n3165), .B1(n3843), .B2(b[1]), .C(
        n2679), .ZN(n2584) );
  AOI211D1BWP12T U3340 ( .A1(n2684), .A2(n2634), .B(n2584), .C(n2626), .ZN(
        n2585) );
  ND2D1BWP12T U3341 ( .A1(n2586), .A2(n2585), .ZN(n3830) );
  AOI22D1BWP12T U3342 ( .A1(b[1]), .A2(n2605), .B1(n3880), .B2(n3165), .ZN(
        n2665) );
  AOI22D1BWP12T U3343 ( .A1(b[1]), .A2(n2607), .B1(n2606), .B2(n3165), .ZN(
        n2629) );
  AOI22D1BWP12T U3344 ( .A1(n2635), .A2(n2665), .B1(n2684), .B2(n2629), .ZN(
        n2591) );
  OAI22D1BWP12T U3345 ( .A1(n3165), .A2(n2620), .B1(n2609), .B2(b[1]), .ZN(
        n2690) );
  INR2D1BWP12T U3346 ( .A1(n2690), .B1(b[2]), .ZN(n3985) );
  AOI22D1BWP12T U3347 ( .A1(b[1]), .A2(n2610), .B1(n2612), .B2(n3165), .ZN(
        n2623) );
  MAOI22D0BWP12T U3348 ( .A1(b[1]), .A2(n2611), .B1(n2614), .B2(b[1]), .ZN(
        n2628) );
  AOI22D1BWP12T U3349 ( .A1(b[2]), .A2(n2623), .B1(n2628), .B2(n2652), .ZN(
        n2691) );
  AOI22D1BWP12T U3350 ( .A1(b[3]), .A2(n3985), .B1(n2691), .B2(n2886), .ZN(
        n2705) );
  OAI22D1BWP12T U3351 ( .A1(n3165), .A2(n2588), .B1(n2587), .B2(b[1]), .ZN(
        n2627) );
  OAI22D1BWP12T U3352 ( .A1(n3165), .A2(n2589), .B1(n2608), .B2(b[1]), .ZN(
        n2630) );
  OA22D1BWP12T U3353 ( .A1(n2652), .A2(n2627), .B1(n2630), .B2(b[2]), .Z(n2692) );
  AOI22D1BWP12T U3354 ( .A1(b[4]), .A2(n2705), .B1(n2912), .B2(n2692), .ZN(
        n2590) );
  ND3D1BWP12T U3355 ( .A1(n3144), .A2(n2591), .A3(n2590), .ZN(n3819) );
  AOI22D1BWP12T U3356 ( .A1(b[1]), .A2(n3739), .B1(n3843), .B2(n3165), .ZN(
        n2677) );
  AOI22D1BWP12T U3357 ( .A1(b[1]), .A2(n2592), .B1(n3740), .B2(n3165), .ZN(
        n2647) );
  AOI22D1BWP12T U3358 ( .A1(n2635), .A2(n2677), .B1(n2684), .B2(n2647), .ZN(
        n2604) );
  NR2D1BWP12T U3359 ( .A1(b[2]), .A2(n2622), .ZN(n3951) );
  AOI22D1BWP12T U3360 ( .A1(b[1]), .A2(n2596), .B1(n2595), .B2(n3165), .ZN(
        n2621) );
  AOI22D1BWP12T U3361 ( .A1(b[1]), .A2(n2598), .B1(n2597), .B2(n3165), .ZN(
        n2645) );
  AOI22D1BWP12T U3362 ( .A1(b[2]), .A2(n2621), .B1(n2645), .B2(n2652), .ZN(
        n2693) );
  AOI22D1BWP12T U3363 ( .A1(b[3]), .A2(n3951), .B1(n2693), .B2(n2886), .ZN(
        n2706) );
  AOI22D1BWP12T U3364 ( .A1(b[1]), .A2(n2600), .B1(n2599), .B2(n3165), .ZN(
        n2646) );
  AOI22D1BWP12T U3365 ( .A1(b[1]), .A2(n2602), .B1(n2601), .B2(n3165), .ZN(
        n2648) );
  AOI22D1BWP12T U3366 ( .A1(b[2]), .A2(n2646), .B1(n2648), .B2(n2652), .ZN(
        n2694) );
  AOI22D1BWP12T U3367 ( .A1(b[4]), .A2(n2706), .B1(n2912), .B2(n2694), .ZN(
        n2603) );
  ND3D1BWP12T U3368 ( .A1(n3144), .A2(n2604), .A3(n2603), .ZN(n3785) );
  AOI22D1BWP12T U3369 ( .A1(b[1]), .A2(n2606), .B1(n2605), .B2(n3165), .ZN(
        n2685) );
  AOI22D1BWP12T U3370 ( .A1(b[1]), .A2(n2608), .B1(n2607), .B2(n3165), .ZN(
        n2654) );
  AOI22D1BWP12T U3371 ( .A1(n2635), .A2(n2685), .B1(n2684), .B2(n2654), .ZN(
        n2618) );
  NR2D1BWP12T U3372 ( .A1(n2620), .A2(n2878), .ZN(n3185) );
  MAOI22D0BWP12T U3373 ( .A1(n2610), .A2(n3165), .B1(n2593), .B2(n2609), .ZN(
        n2619) );
  AOI22D1BWP12T U3374 ( .A1(b[1]), .A2(n2612), .B1(n2611), .B2(n3165), .ZN(
        n2651) );
  AOI22D1BWP12T U3375 ( .A1(b[2]), .A2(n2619), .B1(n2651), .B2(n2652), .ZN(
        n2696) );
  AOI22D1BWP12T U3376 ( .A1(n3185), .A2(n2847), .B1(n2696), .B2(n2886), .ZN(
        n2707) );
  AOI22D1BWP12T U3377 ( .A1(b[1]), .A2(n2614), .B1(n2613), .B2(n3165), .ZN(
        n2653) );
  AOI22D1BWP12T U3378 ( .A1(b[1]), .A2(n2616), .B1(n2615), .B2(n3165), .ZN(
        n2655) );
  AOI22D1BWP12T U3379 ( .A1(b[2]), .A2(n2653), .B1(n2655), .B2(n2652), .ZN(
        n2697) );
  AOI22D1BWP12T U3380 ( .A1(b[4]), .A2(n2707), .B1(n2912), .B2(n2697), .ZN(
        n2617) );
  ND3D1BWP12T U3381 ( .A1(n3144), .A2(n2618), .A3(n2617), .ZN(n3763) );
  ND4D1BWP12T U3382 ( .A1(n3830), .A2(n3819), .A3(n3785), .A4(n3763), .ZN(
        n2703) );
  NR2D1BWP12T U3383 ( .A1(n2626), .A2(n2914), .ZN(n2863) );
  OAI32D1BWP12T U3384 ( .A1(b[1]), .A2(n2652), .A3(n2620), .B1(n2619), .B2(
        b[2]), .ZN(n2657) );
  INVD1BWP12T U3385 ( .I(n2657), .ZN(n3251) );
  NR4D0BWP12T U3386 ( .A1(n3185), .A2(n3951), .A3(n2639), .A4(n3227), .ZN(
        n2624) );
  OAI22D1BWP12T U3387 ( .A1(n2652), .A2(n2622), .B1(n2621), .B2(b[2]), .ZN(
        n2650) );
  INVD1BWP12T U3388 ( .I(n2650), .ZN(n3264) );
  MAOI22D0BWP12T U3389 ( .A1(b[2]), .A2(n2690), .B1(n2623), .B2(b[2]), .ZN(
        n3303) );
  ND4D1BWP12T U3390 ( .A1(n3251), .A2(n2624), .A3(n3264), .A4(n3303), .ZN(
        n2633) );
  NR2D1BWP12T U3391 ( .A1(n2626), .A2(n2625), .ZN(n2699) );
  INVD1BWP12T U3392 ( .I(n2699), .ZN(n2632) );
  AOI22D1BWP12T U3393 ( .A1(b[2]), .A2(n2628), .B1(n2627), .B2(n2652), .ZN(
        n2660) );
  AOI22D1BWP12T U3394 ( .A1(b[2]), .A2(n2630), .B1(n2629), .B2(n2652), .ZN(
        n2661) );
  OAI22D1BWP12T U3395 ( .A1(n2886), .A2(n2660), .B1(n2914), .B2(n2661), .ZN(
        n2631) );
  AOI211D1BWP12T U3396 ( .A1(b[4]), .A2(n3303), .B(n2632), .C(n2631), .ZN(
        n3709) );
  ND2D1BWP12T U3397 ( .A1(n2772), .A2(n2754), .ZN(n3920) );
  AOI211D1BWP12T U3398 ( .A1(n2863), .A2(n2633), .B(n3709), .C(n3920), .ZN(
        n2658) );
  AOI22D1BWP12T U3399 ( .A1(n2636), .A2(n2684), .B1(n2635), .B2(n2634), .ZN(
        n2644) );
  ND2D1BWP12T U3400 ( .A1(n2637), .A2(b[2]), .ZN(n2668) );
  AN2D1BWP12T U3401 ( .A1(n2668), .A2(n2886), .Z(n2640) );
  ND2D1BWP12T U3402 ( .A1(n2652), .A2(n2638), .ZN(n2667) );
  OAI22D1BWP12T U3403 ( .A1(n2640), .A2(n2639), .B1(n2667), .B2(b[3]), .ZN(
        n3324) );
  AOI22D1BWP12T U3404 ( .A1(b[2]), .A2(n2642), .B1(n2641), .B2(n2652), .ZN(
        n2669) );
  AOI22D1BWP12T U3405 ( .A1(b[4]), .A2(n3324), .B1(n2912), .B2(n2669), .ZN(
        n2643) );
  ND3D1BWP12T U3406 ( .A1(n3144), .A2(n2644), .A3(n2643), .ZN(n3747) );
  MAOI22D0BWP12T U3407 ( .A1(n2646), .A2(n2652), .B1(n2652), .B2(n2645), .ZN(
        n2673) );
  MAOI22D0BWP12T U3408 ( .A1(b[2]), .A2(n2648), .B1(n2647), .B2(b[2]), .ZN(
        n2674) );
  AOI22D1BWP12T U3409 ( .A1(b[3]), .A2(n2673), .B1(n3784), .B2(n2674), .ZN(
        n2649) );
  OAI211D1BWP12T U3410 ( .A1(n2650), .A2(n3219), .B(n2699), .C(n2649), .ZN(
        n3683) );
  MAOI22D0BWP12T U3411 ( .A1(n2653), .A2(n2652), .B1(n2652), .B2(n2651), .ZN(
        n2680) );
  MAOI22D0BWP12T U3412 ( .A1(b[2]), .A2(n2655), .B1(n2654), .B2(b[2]), .ZN(
        n2681) );
  AOI22D1BWP12T U3413 ( .A1(b[3]), .A2(n2680), .B1(n3784), .B2(n2681), .ZN(
        n2656) );
  OAI211D1BWP12T U3414 ( .A1(n3219), .A2(n2657), .B(n2699), .C(n2656), .ZN(
        n3652) );
  ND4D1BWP12T U3415 ( .A1(n2658), .A2(n3747), .A3(n3683), .A4(n3652), .ZN(
        n2702) );
  AOI221D1BWP12T U3416 ( .A1(b[1]), .A2(n3879), .B1(n3165), .B2(n2659), .C(
        n2679), .ZN(n2664) );
  MAOI22D0BWP12T U3417 ( .A1(b[3]), .A2(n3303), .B1(n2660), .B2(b[3]), .ZN(
        n3503) );
  OAI22D1BWP12T U3418 ( .A1(n3503), .A2(n3219), .B1(n2662), .B2(n2661), .ZN(
        n2663) );
  AOI211D1BWP12T U3419 ( .A1(n2665), .A2(n2684), .B(n2664), .C(n2663), .ZN(
        n2666) );
  ND2D1BWP12T U3420 ( .A1(n3144), .A2(n2666), .ZN(n3200) );
  ND2D1BWP12T U3421 ( .A1(n2668), .A2(n2667), .ZN(n2670) );
  AOI22D1BWP12T U3422 ( .A1(b[3]), .A2(n2670), .B1(n3784), .B2(n2669), .ZN(
        n2671) );
  OAI211D1BWP12T U3423 ( .A1(n3158), .A2(n3219), .B(n3144), .C(n2671), .ZN(
        n3519) );
  AOI221D1BWP12T U3424 ( .A1(n3844), .A2(b[1]), .B1(n2672), .B2(n3165), .C(
        n2679), .ZN(n2676) );
  AOI22D1BWP12T U3425 ( .A1(b[3]), .A2(n3264), .B1(n2673), .B2(n2886), .ZN(
        n3471) );
  MOAI22D0BWP12T U3426 ( .A1(n3471), .A2(n3219), .B1(n2674), .B2(n2912), .ZN(
        n2675) );
  AOI211D1BWP12T U3427 ( .A1(n2677), .A2(n2684), .B(n2676), .C(n2675), .ZN(
        n2678) );
  ND2D1BWP12T U3428 ( .A1(n3144), .A2(n2678), .ZN(n3919) );
  AOI221D1BWP12T U3429 ( .A1(n3880), .A2(b[1]), .B1(n3879), .B2(n3165), .C(
        n2679), .ZN(n2683) );
  AOI22D1BWP12T U3430 ( .A1(b[3]), .A2(n3251), .B1(n2680), .B2(n2886), .ZN(
        n3451) );
  MOAI22D0BWP12T U3431 ( .A1(n3451), .A2(n3219), .B1(n2912), .B2(n2681), .ZN(
        n2682) );
  AOI211D1BWP12T U3432 ( .A1(n2685), .A2(n2684), .B(n2683), .C(n2682), .ZN(
        n2686) );
  ND2D1BWP12T U3433 ( .A1(n3144), .A2(n2686), .ZN(n3890) );
  ND4D1BWP12T U3434 ( .A1(n3200), .A2(n3519), .A3(n3919), .A4(n3890), .ZN(
        n2701) );
  MAOI22D0BWP12T U3435 ( .A1(n3784), .A2(n2688), .B1(n2886), .B2(n2687), .ZN(
        n2689) );
  OAI211D1BWP12T U3436 ( .A1(n3219), .A2(n3227), .B(n2699), .C(n2689), .ZN(
        n3636) );
  ND2D1BWP12T U3437 ( .A1(n2860), .A2(n2690), .ZN(n2708) );
  MAOI22D0BWP12T U3438 ( .A1(n3784), .A2(n2694), .B1(n2886), .B2(n2693), .ZN(
        n2695) );
  OAI211D1BWP12T U3439 ( .A1(n3951), .A2(n3219), .B(n2699), .C(n2695), .ZN(
        n3589) );
  MAOI22D0BWP12T U3440 ( .A1(n3784), .A2(n2697), .B1(n2886), .B2(n2696), .ZN(
        n2698) );
  OAI211D1BWP12T U3441 ( .A1(n3185), .A2(n3219), .B(n2699), .C(n2698), .ZN(
        n3557) );
  ND4D1BWP12T U3442 ( .A1(n3636), .A2(n3609), .A3(n3589), .A4(n3557), .ZN(
        n2700) );
  NR4D0BWP12T U3443 ( .A1(n2703), .A2(n2702), .A3(n2701), .A4(n2700), .ZN(
        n2712) );
  INVD1BWP12T U3444 ( .I(n2704), .ZN(n3423) );
  INVD1BWP12T U3445 ( .I(n2705), .ZN(n3396) );
  INVD1BWP12T U3446 ( .I(n2706), .ZN(n3379) );
  INVD1BWP12T U3447 ( .I(n2707), .ZN(n3352) );
  NR4D0BWP12T U3448 ( .A1(n3423), .A2(n3396), .A3(n3379), .A4(n3352), .ZN(
        n2709) );
  IND4D1BWP12T U3449 ( .A1(n3503), .B1(n2709), .B2(n3324), .B3(n2708), .ZN(
        n2710) );
  OAI31D1BWP12T U3450 ( .A1(n3471), .A2(n3451), .A3(n2710), .B(n3199), .ZN(
        n2711) );
  AOI22D1BWP12T U3451 ( .A1(n2714), .A2(n2713), .B1(n2712), .B2(n2711), .ZN(
        n2935) );
  NR2D1BWP12T U3452 ( .A1(op[0]), .A2(op[1]), .ZN(n2859) );
  ND2D1BWP12T U3453 ( .A1(n2771), .A2(n2859), .ZN(n3988) );
  INVD1BWP12T U3454 ( .I(n3988), .ZN(n3940) );
  AN2D1BWP12T U3455 ( .A1(n3627), .A2(n2859), .Z(n3531) );
  ND4D1BWP12T U3456 ( .A1(n3239), .A2(n3273), .A3(n3290), .A4(n3318), .ZN(
        n2731) );
  ND2D1BWP12T U3457 ( .A1(a[31]), .A2(b[31]), .ZN(n3135) );
  ND4D1BWP12T U3458 ( .A1(n3135), .A2(n3939), .A3(n3993), .A4(n2726), .ZN(
        n2730) );
  ND2D1BWP12T U3459 ( .A1(b[16]), .A2(a[16]), .ZN(n2727) );
  ND4D1BWP12T U3460 ( .A1(n3442), .A2(n3474), .A3(n3493), .A4(n2727), .ZN(
        n2729) );
  ND4D1BWP12T U3461 ( .A1(n3342), .A2(n3372), .A3(n3394), .A4(n3418), .ZN(
        n2728) );
  NR4D0BWP12T U3462 ( .A1(n2731), .A2(n2730), .A3(n2729), .A4(n2728), .ZN(
        n2732) );
  AOI22D1BWP12T U3463 ( .A1(n2735), .A2(n2734), .B1(n2733), .B2(n2732), .ZN(
        n2934) );
  ND2D1BWP12T U3464 ( .A1(a[12]), .A2(n3416), .ZN(n3426) );
  ND2D1BWP12T U3465 ( .A1(a[11]), .A2(n2759), .ZN(n2737) );
  ND4D1BWP12T U3466 ( .A1(n3426), .A2(n2737), .A3(n3941), .A4(n2736), .ZN(
        n2750) );
  ND2D1BWP12T U3467 ( .A1(a[19]), .A2(n3598), .ZN(n2738) );
  ND4D1BWP12T U3468 ( .A1(n2739), .A2(n2738), .A3(n3523), .A4(n3491), .ZN(
        n2749) );
  ND4D1BWP12T U3469 ( .A1(n2743), .A2(n2742), .A3(n2741), .A4(n2740), .ZN(
        n2748) );
  ND4D1BWP12T U3470 ( .A1(n2746), .A2(n2745), .A3(n2744), .A4(n3155), .ZN(
        n2747) );
  NR4D0BWP12T U3471 ( .A1(n2750), .A2(n2749), .A3(n2748), .A4(n2747), .ZN(
        n2925) );
  NR2D1BWP12T U3472 ( .A1(b[25]), .A2(n3768), .ZN(n3758) );
  ND2D1BWP12T U3473 ( .A1(n3102), .A2(n2754), .ZN(n3724) );
  INVD1BWP12T U3474 ( .I(n3724), .ZN(n3823) );
  ND2D1BWP12T U3475 ( .A1(b[27]), .A2(n3824), .ZN(n2755) );
  NR2D1BWP12T U3476 ( .A1(a[10]), .A2(n3370), .ZN(n2758) );
  NR2D1BWP12T U3477 ( .A1(a[14]), .A2(n3465), .ZN(n2762) );
  NR2D1BWP12T U3478 ( .A1(a[12]), .A2(n3416), .ZN(n2761) );
  NR2D1BWP12T U3479 ( .A1(a[11]), .A2(n2759), .ZN(n2760) );
  NR2D1BWP12T U3480 ( .A1(a[4]), .A2(n3219), .ZN(n2767) );
  ND2D1BWP12T U3481 ( .A1(n2772), .A2(n2771), .ZN(n3650) );
  NR2D1BWP12T U3482 ( .A1(n2778), .A2(n2777), .ZN(n2779) );
  MAOI22D0BWP12T U3483 ( .A1(n2780), .A2(n2779), .B1(n2780), .B2(n2779), .ZN(
        n4004) );
  INVD1BWP12T U3484 ( .I(n3958), .ZN(n4003) );
  FA1D0BWP12T U3485 ( .A(mult_x_18_n247), .B(n2782), .CI(n2781), .CO(n2116), 
        .S(n3914) );
  FA1D0BWP12T U3486 ( .A(mult_x_18_n263), .B(n2784), .CI(n2783), .CO(n2781), 
        .S(n3867) );
  FA1D0BWP12T U3487 ( .A(mult_x_18_n277), .B(n2786), .CI(n2785), .CO(n2784), 
        .S(n3850) );
  NR4D0BWP12T U3488 ( .A1(n2787), .A2(n3914), .A3(n3867), .A4(n3850), .ZN(
        n2806) );
  FA1D0BWP12T U3489 ( .A(mult_x_18_n291), .B(n2789), .CI(n2788), .CO(n2786), 
        .S(n3822) );
  FA1D0BWP12T U3490 ( .A(mult_x_18_n305), .B(n2791), .CI(n2790), .CO(n2788), 
        .S(n3797) );
  FA1D0BWP12T U3491 ( .A(mult_x_18_n318), .B(n2793), .CI(n2792), .CO(n2791), 
        .S(n3760) );
  FA1D0BWP12T U3492 ( .A(mult_x_18_n331), .B(n2795), .CI(n2794), .CO(n2792), 
        .S(n3735) );
  NR4D0BWP12T U3493 ( .A1(n3822), .A2(n3797), .A3(n3760), .A4(n3735), .ZN(
        n2805) );
  FA1D0BWP12T U3494 ( .A(mult_x_18_n344), .B(n2797), .CI(n2796), .CO(n2795), 
        .S(n3700) );
  FA1D0BWP12T U3495 ( .A(mult_x_18_n355), .B(n2799), .CI(n2798), .CO(n2796), 
        .S(n3673) );
  FA1D0BWP12T U3496 ( .A(mult_x_18_n366), .B(n2801), .CI(n2800), .CO(n2798), 
        .S(n3656) );
  FA1D0BWP12T U3497 ( .A(mult_x_18_n377), .B(n2803), .CI(n2802), .CO(n2800), 
        .S(n3626) );
  NR4D0BWP12T U3498 ( .A1(n3700), .A2(n3673), .A3(n3656), .A4(n3626), .ZN(
        n2804) );
  ND4D1BWP12T U3499 ( .A1(n4003), .A2(n2806), .A3(n2805), .A4(n2804), .ZN(
        n2845) );
  FA1D0BWP12T U3500 ( .A(mult_x_18_n387), .B(n2808), .CI(n2807), .CO(n2802), 
        .S(n3599) );
  FA1D0BWP12T U3501 ( .A(mult_x_18_n397), .B(n2810), .CI(n2809), .CO(n2807), 
        .S(n3577) );
  FA1D0BWP12T U3502 ( .A(mult_x_18_n407), .B(n2812), .CI(n2811), .CO(n2809), 
        .S(n3548) );
  FA1D0BWP12T U3503 ( .A(mult_x_18_n415), .B(n2814), .CI(n2813), .CO(n2811), 
        .S(n3521) );
  NR4D0BWP12T U3504 ( .A1(n3599), .A2(n3577), .A3(n3548), .A4(n3521), .ZN(
        n2843) );
  FA1D0BWP12T U3505 ( .A(mult_x_18_n423), .B(n2816), .CI(n2815), .CO(n2814), 
        .S(n3496) );
  FA1D0BWP12T U3506 ( .A(mult_x_18_n431), .B(n2818), .CI(n2817), .CO(n2816), 
        .S(n3466) );
  FA1D0BWP12T U3507 ( .A(mult_x_18_n438), .B(n2820), .CI(n2819), .CO(n2818), 
        .S(n3441) );
  FA1D0BWP12T U3508 ( .A(mult_x_18_n445), .B(n2822), .CI(n2821), .CO(n2820), 
        .S(n3417) );
  NR4D0BWP12T U3509 ( .A1(n3496), .A2(n3466), .A3(n3441), .A4(n3417), .ZN(
        n2842) );
  FA1D0BWP12T U3510 ( .A(mult_x_18_n452), .B(n2824), .CI(n2823), .CO(n2822), 
        .S(n3395) );
  FA1D0BWP12T U3511 ( .A(mult_x_18_n457), .B(n2826), .CI(n2825), .CO(n2824), 
        .S(n3371) );
  FA1D0BWP12T U3512 ( .A(mult_x_18_n462), .B(n2828), .CI(n2827), .CO(n2825), 
        .S(n3340) );
  NR4D0BWP12T U3513 ( .A1(n3395), .A2(n3371), .A3(n3340), .A4(n3317), .ZN(
        n2841) );
  FA1D0BWP12T U3514 ( .A(n2833), .B(n2832), .CI(n2831), .CO(n2830), .S(n3270)
         );
  FA1D0BWP12T U3515 ( .A(n2836), .B(n2835), .CI(n2834), .CO(n2833), .S(n3246)
         );
  FA1D0BWP12T U3516 ( .A(n2839), .B(n2838), .CI(n2837), .CO(n2835), .S(n3220)
         );
  NR4D0BWP12T U3517 ( .A1(n3289), .A2(n3270), .A3(n3246), .A4(n3220), .ZN(
        n2840) );
  ND4D1BWP12T U3518 ( .A1(n2843), .A2(n2842), .A3(n2841), .A4(n2840), .ZN(
        n2844) );
  NR4D0BWP12T U3519 ( .A1(n4004), .A2(n2846), .A3(n2845), .A4(n2844), .ZN(
        n2923) );
  AOI31D1BWP12T U3520 ( .A1(a[31]), .A2(n2848), .A3(n2847), .B(n3427), .ZN(
        n3432) );
  INVD1BWP12T U3521 ( .I(n2874), .ZN(n2872) );
  NR2D1BWP12T U3522 ( .A1(n2849), .A2(n2872), .ZN(n2880) );
  OAI32D1BWP12T U3523 ( .A1(n3908), .A2(n2880), .A3(n3679), .B1(a[31]), .B2(
        n3199), .ZN(n3688) );
  OAI211D1BWP12T U3524 ( .A1(n2880), .A2(n2851), .B(n3144), .C(n2850), .ZN(
        n3288) );
  NR2D1BWP12T U3525 ( .A1(n2852), .A2(n2626), .ZN(n2855) );
  OAI21D1BWP12T U3526 ( .A1(n3199), .A2(n2855), .B(n2853), .ZN(n3192) );
  ND4D1BWP12T U3527 ( .A1(n3432), .A2(n3688), .A3(n3288), .A4(n3192), .ZN(
        n2921) );
  ND2D1BWP12T U3528 ( .A1(n3908), .A2(a[31]), .ZN(n3907) );
  INVD1BWP12T U3529 ( .I(n3907), .ZN(n3899) );
  AOI21D1BWP12T U3530 ( .A1(n3199), .A2(n2854), .B(n3899), .ZN(n3711) );
  AN2D1BWP12T U3531 ( .A1(n2855), .A2(n3219), .Z(n3564) );
  NR2D1BWP12T U3532 ( .A1(n2856), .A2(n2874), .ZN(n2868) );
  INVD1BWP12T U3533 ( .I(n2857), .ZN(n2858) );
  AOI211D1BWP12T U3534 ( .A1(b[4]), .A2(n2868), .B(n2626), .C(n2858), .ZN(
        n3397) );
  INVD1BWP12T U3535 ( .I(n2859), .ZN(n3269) );
  INVD1BWP12T U3536 ( .I(n3996), .ZN(n3831) );
  NR2D1BWP12T U3537 ( .A1(n2860), .A2(n3194), .ZN(n2861) );
  AOI211D1BWP12T U3538 ( .A1(n2863), .A2(n2862), .B(n3899), .C(n2861), .ZN(
        n3832) );
  OAI211D1BWP12T U3539 ( .A1(n3908), .A2(n3921), .B(n3832), .C(n3194), .ZN(
        n2864) );
  NR4D0BWP12T U3540 ( .A1(n3564), .A2(n3397), .A3(n3831), .A4(n2864), .ZN(
        n2865) );
  ND3D1BWP12T U3541 ( .A1(a[31]), .A2(b[3]), .A3(b[2]), .ZN(n2898) );
  IOA21D1BWP12T U3542 ( .A1(n2898), .A2(n3637), .B(n3199), .ZN(n3624) );
  IND4D1BWP12T U3543 ( .A1(n2866), .B1(n3711), .B2(n2865), .B3(n3624), .ZN(
        n2920) );
  AOI22D1BWP12T U3544 ( .A1(n2906), .A2(n2881), .B1(a[31]), .B2(n2867), .ZN(
        n2910) );
  NR2D1BWP12T U3545 ( .A1(n2910), .A2(n3908), .ZN(n3898) );
  NR2D1BWP12T U3546 ( .A1(n2868), .A2(n3908), .ZN(n3820) );
  AOI32D1BWP12T U3547 ( .A1(n3165), .A2(n2871), .A3(n2870), .B1(n2869), .B2(
        n2871), .ZN(n2885) );
  AOI21D1BWP12T U3548 ( .A1(n2886), .A2(n2885), .B(n2874), .ZN(n2889) );
  NR2D1BWP12T U3549 ( .A1(n2889), .A2(n3908), .ZN(n3798) );
  ND2D1BWP12T U3550 ( .A1(n2873), .A2(n2872), .ZN(n2893) );
  AN2D1BWP12T U3551 ( .A1(n2893), .A2(n3199), .Z(n3756) );
  NR4D0BWP12T U3552 ( .A1(n3898), .A2(n3820), .A3(n3798), .A4(n3756), .ZN(
        n2895) );
  NR2D1BWP12T U3553 ( .A1(n2875), .A2(n2874), .ZN(n2901) );
  INVD1BWP12T U3554 ( .I(n2876), .ZN(n2877) );
  AOI211D1BWP12T U3555 ( .A1(b[4]), .A2(n2901), .B(n2626), .C(n2877), .ZN(
        n3315) );
  NR2D1BWP12T U3556 ( .A1(n2886), .A2(n2878), .ZN(n2882) );
  AOI211D1BWP12T U3557 ( .A1(n2882), .A2(n2881), .B(n2880), .C(n2879), .ZN(
        n2902) );
  AOI21D1BWP12T U3558 ( .A1(b[4]), .A2(n2902), .B(n2883), .ZN(n3254) );
  OAI21D1BWP12T U3559 ( .A1(n2886), .A2(n2885), .B(n2884), .ZN(n2904) );
  AOI211D1BWP12T U3560 ( .A1(b[4]), .A2(n2904), .B(n2887), .C(n2626), .ZN(
        n3950) );
  NR4D0BWP12T U3561 ( .A1(n3997), .A2(n3315), .A3(n3254), .A4(n3950), .ZN(
        n2894) );
  AO21D1BWP12T U3562 ( .A1(b[4]), .A2(n2889), .B(n2888), .Z(n3366) );
  AOI22D1BWP12T U3563 ( .A1(n3784), .A2(n2891), .B1(n2912), .B2(n2890), .ZN(
        n2892) );
  OAI211D1BWP12T U3564 ( .A1(n3219), .A2(n2893), .B(n3144), .C(n2892), .ZN(
        n3349) );
  ND4D1BWP12T U3565 ( .A1(n2895), .A2(n2894), .A3(n3366), .A4(n3349), .ZN(
        n2919) );
  NR2D1BWP12T U3566 ( .A1(n3144), .A2(n3194), .ZN(n3159) );
  AOI21D1BWP12T U3567 ( .A1(n2896), .A2(n3144), .B(n3159), .ZN(n3304) );
  AOI211D1BWP12T U3568 ( .A1(n2899), .A2(n2898), .B(n2897), .C(n2626), .ZN(
        n2900) );
  NR2D1BWP12T U3569 ( .A1(n3159), .A2(n2900), .ZN(n3236) );
  NR2D1BWP12T U3570 ( .A1(n2901), .A2(n3908), .ZN(n3726) );
  NR2D1BWP12T U3571 ( .A1(n2902), .A2(n3908), .ZN(n3649) );
  NR2D1BWP12T U3572 ( .A1(n3908), .A2(n2903), .ZN(n3604) );
  NR2D1BWP12T U3573 ( .A1(n3908), .A2(n2904), .ZN(n3582) );
  NR4D0BWP12T U3574 ( .A1(n3726), .A2(n3649), .A3(n3604), .A4(n3582), .ZN(
        n2917) );
  INVD1BWP12T U3575 ( .I(n2905), .ZN(n3520) );
  NR2D1BWP12T U3576 ( .A1(n3908), .A2(n3520), .ZN(n3526) );
  AOI211D1BWP12T U3577 ( .A1(b[4]), .A2(n3909), .B(n2626), .C(n2908), .ZN(
        n3470) );
  AOI211D1BWP12T U3578 ( .A1(b[4]), .A2(n2910), .B(n2626), .C(n2909), .ZN(
        n3449) );
  ND2D1BWP12T U3579 ( .A1(n2912), .A2(n2911), .ZN(n2913) );
  OAI32D1BWP12T U3580 ( .A1(n2626), .A2(n2915), .A3(n2914), .B1(n2913), .B2(
        n2626), .ZN(n3492) );
  NR4D0BWP12T U3581 ( .A1(n3526), .A2(n3470), .A3(n3449), .A4(n3492), .ZN(
        n2916) );
  ND4D1BWP12T U3582 ( .A1(n3304), .A2(n3236), .A3(n2917), .A4(n2916), .ZN(
        n2918) );
  NR4D0BWP12T U3583 ( .A1(n2921), .A2(n2920), .A3(n2919), .A4(n2918), .ZN(
        n2922) );
  AOI211D1BWP12T U3584 ( .A1(n2925), .A2(n2924), .B(n2923), .C(n2922), .ZN(
        n2933) );
  NR2D1BWP12T U3585 ( .A1(n2927), .A2(n2926), .ZN(n3959) );
  INVD1BWP12T U3586 ( .I(n3959), .ZN(n3995) );
  ND4D1BWP12T U3587 ( .A1(n2931), .A2(n2930), .A3(n2929), .A4(n2928), .ZN(
        n2932) );
  ND4D1BWP12T U3588 ( .A1(n2935), .A2(n2934), .A3(n2933), .A4(n2932), .ZN(
        n2936) );
  AOI211D1BWP12T U3589 ( .A1(n3140), .A2(n2938), .B(n2937), .C(n2936), .ZN(
        n3131) );
  MOAI22D0BWP12T U3590 ( .A1(n3027), .A2(n2939), .B1(n3027), .B2(n2939), .ZN(
        n3215) );
  MAOI22D0BWP12T U3591 ( .A1(n2940), .A2(n3029), .B1(n2940), .B2(n3029), .ZN(
        n3927) );
  NR2D1BWP12T U3592 ( .A1(n2941), .A2(n3841), .ZN(n2942) );
  MOAI22D0BWP12T U3593 ( .A1(n2942), .A2(n3032), .B1(n2942), .B2(n3032), .ZN(
        n3897) );
  INR2D1BWP12T U3594 ( .A1(n3787), .B1(n2943), .ZN(n2944) );
  MOAI22D0BWP12T U3595 ( .A1(n2944), .A2(n3038), .B1(n2944), .B2(n3038), .ZN(
        n3828) );
  MOAI22D0BWP12T U3596 ( .A1(n2945), .A2(n3035), .B1(n2945), .B2(n3035), .ZN(
        n3860) );
  MAOI22D0BWP12T U3597 ( .A1(n2946), .A2(n3041), .B1(n2946), .B2(n3041), .ZN(
        n3802) );
  NR2D1BWP12T U3598 ( .A1(n2948), .A2(n2947), .ZN(n2949) );
  MOAI22D0BWP12T U3599 ( .A1(n2949), .A2(n3047), .B1(n2949), .B2(n3047), .ZN(
        n3755) );
  INR2D1BWP12T U3600 ( .A1(n3675), .B1(n2950), .ZN(n2951) );
  MOAI22D0BWP12T U3601 ( .A1(n2951), .A2(n3050), .B1(n2951), .B2(n3050), .ZN(
        n3716) );
  MOAI22D0BWP12T U3602 ( .A1(n2952), .A2(n3053), .B1(n2952), .B2(n3053), .ZN(
        n3693) );
  ND2D1BWP12T U3603 ( .A1(n2954), .A2(n2953), .ZN(n2955) );
  MOAI22D0BWP12T U3604 ( .A1(n3056), .A2(n2955), .B1(n3056), .B2(n2955), .ZN(
        n3671) );
  MOAI22D0BWP12T U3605 ( .A1(n2956), .A2(n3061), .B1(n2956), .B2(n3061), .ZN(
        n3623) );
  MAOI22D0BWP12T U3606 ( .A1(n2957), .A2(n3067), .B1(n2957), .B2(n3067), .ZN(
        n3563) );
  MOAI22D0BWP12T U3607 ( .A1(n2958), .A2(n3070), .B1(n2958), .B2(n3070), .ZN(
        n3540) );
  MAOI22D0BWP12T U3608 ( .A1(n2959), .A2(n3073), .B1(n2959), .B2(n3073), .ZN(
        n3518) );
  MOAI22D0BWP12T U3609 ( .A1(n2960), .A2(n3079), .B1(n2960), .B2(n3079), .ZN(
        n3460) );
  MAOI22D0BWP12T U3610 ( .A1(n2961), .A2(n3082), .B1(n2961), .B2(n3082), .ZN(
        n3440) );
  ND2D1BWP12T U3611 ( .A1(n2962), .A2(n3343), .ZN(n2963) );
  MAOI22D0BWP12T U3612 ( .A1(n3088), .A2(n2963), .B1(n3088), .B2(n2963), .ZN(
        n3389) );
  MAOI22D0BWP12T U3613 ( .A1(n2964), .A2(n3085), .B1(n2964), .B2(n3085), .ZN(
        n3411) );
  MAOI22D0BWP12T U3614 ( .A1(n2965), .A2(n3091), .B1(n2965), .B2(n3091), .ZN(
        n3364) );
  MOAI22D0BWP12T U3615 ( .A1(n2966), .A2(n3110), .B1(n2966), .B2(n3110), .ZN(
        n3309) );
  MAOI22D0BWP12T U3616 ( .A1(n2967), .A2(n3100), .B1(n2967), .B2(n3100), .ZN(
        n3998) );
  ND2D1BWP12T U3617 ( .A1(n2969), .A2(n2968), .ZN(n2970) );
  MAOI22D0BWP12T U3618 ( .A1(n3097), .A2(n2970), .B1(n3097), .B2(n2970), .ZN(
        n3217) );
  MAOI22D0BWP12T U3619 ( .A1(n2971), .A2(n3116), .B1(n2971), .B2(n3116), .ZN(
        n3257) );
  ND2D1BWP12T U3620 ( .A1(c_in), .A2(n3151), .ZN(n3000) );
  OAI21D1BWP12T U3621 ( .A1(c_in), .A2(n3151), .B(n3000), .ZN(n3145) );
  INVD1BWP12T U3622 ( .I(n3145), .ZN(n3148) );
  INVD1BWP12T U3623 ( .I(n3949), .ZN(n3999) );
  OAI21D1BWP12T U3624 ( .A1(n2974), .A2(n2973), .B(n2972), .ZN(n3948) );
  OAI21D1BWP12T U3625 ( .A1(n2977), .A2(n2976), .B(n2975), .ZN(n3176) );
  ND4D1BWP12T U3626 ( .A1(n3148), .A2(n3999), .A3(n3948), .A4(n3176), .ZN(
        n2978) );
  NR4D0BWP12T U3627 ( .A1(n3998), .A2(n3217), .A3(n3257), .A4(n2978), .ZN(
        n2985) );
  ND2D1BWP12T U3628 ( .A1(n2980), .A2(n2979), .ZN(n2981) );
  MOAI22D0BWP12T U3629 ( .A1(n3094), .A2(n2981), .B1(n3094), .B2(n2981), .ZN(
        n3332) );
  INVD1BWP12T U3630 ( .I(n2982), .ZN(n3243) );
  ND2D1BWP12T U3631 ( .A1(n2983), .A2(n3243), .ZN(n2984) );
  MOAI22D0BWP12T U3632 ( .A1(n3113), .A2(n2984), .B1(n3113), .B2(n2984), .ZN(
        n3281) );
  ND4D1BWP12T U3633 ( .A1(n3309), .A2(n2985), .A3(n3332), .A4(n3281), .ZN(
        n2986) );
  NR4D0BWP12T U3634 ( .A1(n3389), .A2(n3411), .A3(n3364), .A4(n2986), .ZN(
        n2989) );
  IND2D1BWP12T U3635 ( .A1(n3443), .B1(n2987), .ZN(n2988) );
  MOAI22D0BWP12T U3636 ( .A1(n3076), .A2(n2988), .B1(n3076), .B2(n2988), .ZN(
        n3484) );
  ND4D1BWP12T U3637 ( .A1(n3460), .A2(n3440), .A3(n2989), .A4(n3484), .ZN(
        n2990) );
  NR4D0BWP12T U3638 ( .A1(n3563), .A2(n3540), .A3(n3518), .A4(n2990), .ZN(
        n2995) );
  MAOI22D0BWP12T U3639 ( .A1(n2991), .A2(n3629), .B1(n2991), .B2(n3629), .ZN(
        n3642) );
  ND2D1BWP12T U3640 ( .A1(n2993), .A2(n2992), .ZN(n2994) );
  MOAI22D0BWP12T U3641 ( .A1(n3064), .A2(n2994), .B1(n3064), .B2(n2994), .ZN(
        n3597) );
  ND4D1BWP12T U3642 ( .A1(n3623), .A2(n2995), .A3(n3642), .A4(n3597), .ZN(
        n2996) );
  NR4D0BWP12T U3643 ( .A1(n3716), .A2(n3693), .A3(n3671), .A4(n2996), .ZN(
        n2998) );
  MOAI22D0BWP12T U3644 ( .A1(n2997), .A2(n3044), .B1(n2997), .B2(n3044), .ZN(
        n3776) );
  ND4D1BWP12T U3645 ( .A1(n3802), .A2(n3755), .A3(n2998), .A4(n3776), .ZN(
        n2999) );
  NR4D0BWP12T U3646 ( .A1(n3897), .A2(n3828), .A3(n3860), .A4(n2999), .ZN(
        n3129) );
  ND2D1BWP12T U3647 ( .A1(n3147), .A2(n3000), .ZN(n3104) );
  ND2D1BWP12T U3648 ( .A1(n3105), .A2(n3104), .ZN(n3103) );
  ND2D1BWP12T U3649 ( .A1(n3163), .A2(n3103), .ZN(n3108) );
  ND2D1BWP12T U3650 ( .A1(n3107), .A2(n3108), .ZN(n3106) );
  ND2D1BWP12T U3651 ( .A1(n3939), .A2(n3106), .ZN(n3101) );
  NR2D1BWP12T U3652 ( .A1(n3101), .A2(n3100), .ZN(n3099) );
  NR2D1BWP12T U3653 ( .A1(n3001), .A2(n3099), .ZN(n3098) );
  NR2D1BWP12T U3654 ( .A1(n3098), .A2(n3097), .ZN(n3096) );
  NR2D1BWP12T U3655 ( .A1(n3002), .A2(n3096), .ZN(n3117) );
  NR2D1BWP12T U3656 ( .A1(n3117), .A2(n3116), .ZN(n3115) );
  NR2D1BWP12T U3657 ( .A1(n3003), .A2(n3115), .ZN(n3114) );
  NR2D1BWP12T U3658 ( .A1(n3114), .A2(n3113), .ZN(n3112) );
  NR2D1BWP12T U3659 ( .A1(n3004), .A2(n3112), .ZN(n3111) );
  NR2D1BWP12T U3660 ( .A1(n3111), .A2(n3110), .ZN(n3109) );
  NR2D1BWP12T U3661 ( .A1(n3005), .A2(n3109), .ZN(n3095) );
  NR2D1BWP12T U3662 ( .A1(n3095), .A2(n3094), .ZN(n3093) );
  NR2D1BWP12T U3663 ( .A1(n3006), .A2(n3093), .ZN(n3092) );
  NR2D1BWP12T U3664 ( .A1(n3092), .A2(n3091), .ZN(n3090) );
  NR2D1BWP12T U3665 ( .A1(n3007), .A2(n3090), .ZN(n3089) );
  NR2D1BWP12T U3666 ( .A1(n3089), .A2(n3088), .ZN(n3087) );
  NR2D1BWP12T U3667 ( .A1(n3008), .A2(n3087), .ZN(n3086) );
  NR2D1BWP12T U3668 ( .A1(n3086), .A2(n3085), .ZN(n3084) );
  NR2D1BWP12T U3669 ( .A1(n3009), .A2(n3084), .ZN(n3083) );
  NR2D1BWP12T U3670 ( .A1(n3083), .A2(n3082), .ZN(n3081) );
  NR2D1BWP12T U3671 ( .A1(n3010), .A2(n3081), .ZN(n3080) );
  NR2D1BWP12T U3672 ( .A1(n3080), .A2(n3079), .ZN(n3078) );
  NR2D1BWP12T U3673 ( .A1(n3011), .A2(n3078), .ZN(n3077) );
  NR2D1BWP12T U3674 ( .A1(n3077), .A2(n3076), .ZN(n3075) );
  NR2D1BWP12T U3675 ( .A1(n3012), .A2(n3075), .ZN(n3074) );
  NR2D1BWP12T U3676 ( .A1(n3074), .A2(n3073), .ZN(n3072) );
  NR2D1BWP12T U3677 ( .A1(n3013), .A2(n3072), .ZN(n3071) );
  NR2D1BWP12T U3678 ( .A1(n3071), .A2(n3070), .ZN(n3069) );
  NR2D1BWP12T U3679 ( .A1(n3014), .A2(n3069), .ZN(n3068) );
  NR2D1BWP12T U3680 ( .A1(n3068), .A2(n3067), .ZN(n3066) );
  NR2D1BWP12T U3681 ( .A1(n3015), .A2(n3066), .ZN(n3065) );
  NR2D1BWP12T U3682 ( .A1(n3065), .A2(n3064), .ZN(n3063) );
  NR2D1BWP12T U3683 ( .A1(n3016), .A2(n3063), .ZN(n3062) );
  NR2D1BWP12T U3684 ( .A1(n3062), .A2(n3061), .ZN(n3060) );
  NR2D1BWP12T U3685 ( .A1(n3017), .A2(n3060), .ZN(n3059) );
  NR2D1BWP12T U3686 ( .A1(n3059), .A2(n3629), .ZN(n3058) );
  NR2D1BWP12T U3687 ( .A1(n3018), .A2(n3058), .ZN(n3057) );
  NR2D1BWP12T U3688 ( .A1(n3057), .A2(n3056), .ZN(n3055) );
  NR2D1BWP12T U3689 ( .A1(n3657), .A2(n3055), .ZN(n3054) );
  NR2D1BWP12T U3690 ( .A1(n3054), .A2(n3053), .ZN(n3052) );
  NR2D1BWP12T U3691 ( .A1(n3019), .A2(n3052), .ZN(n3051) );
  NR2D1BWP12T U3692 ( .A1(n3051), .A2(n3050), .ZN(n3049) );
  NR2D1BWP12T U3693 ( .A1(n3020), .A2(n3049), .ZN(n3048) );
  NR2D1BWP12T U3694 ( .A1(n3048), .A2(n3047), .ZN(n3046) );
  NR2D1BWP12T U3695 ( .A1(n3021), .A2(n3046), .ZN(n3045) );
  NR2D1BWP12T U3696 ( .A1(n3045), .A2(n3044), .ZN(n3043) );
  NR2D1BWP12T U3697 ( .A1(n3022), .A2(n3043), .ZN(n3042) );
  NR2D1BWP12T U3698 ( .A1(n3042), .A2(n3041), .ZN(n3040) );
  NR2D1BWP12T U3699 ( .A1(n3794), .A2(n3040), .ZN(n3039) );
  NR2D1BWP12T U3700 ( .A1(n3039), .A2(n3038), .ZN(n3037) );
  NR2D1BWP12T U3701 ( .A1(n3023), .A2(n3037), .ZN(n3036) );
  NR2D1BWP12T U3702 ( .A1(n3036), .A2(n3035), .ZN(n3034) );
  NR2D1BWP12T U3703 ( .A1(n3024), .A2(n3034), .ZN(n3033) );
  NR2D1BWP12T U3704 ( .A1(n3033), .A2(n3032), .ZN(n3031) );
  NR2D1BWP12T U3705 ( .A1(n3025), .A2(n3031), .ZN(n3030) );
  NR2D1BWP12T U3706 ( .A1(n3030), .A2(n3029), .ZN(n3028) );
  NR2D1BWP12T U3707 ( .A1(n3026), .A2(n3028), .ZN(n3133) );
  MOAI22D0BWP12T U3708 ( .A1(n3133), .A2(n3027), .B1(n3133), .B2(n3027), .ZN(
        n3212) );
  AO21D1BWP12T U3709 ( .A1(n3030), .A2(n3029), .B(n3028), .Z(n3930) );
  AO21D1BWP12T U3710 ( .A1(n3033), .A2(n3032), .B(n3031), .Z(n3896) );
  AOI21D1BWP12T U3711 ( .A1(n3036), .A2(n3035), .B(n3034), .ZN(n3863) );
  AOI21D1BWP12T U3712 ( .A1(n3039), .A2(n3038), .B(n3037), .ZN(n3826) );
  AOI21D1BWP12T U3713 ( .A1(n3042), .A2(n3041), .B(n3040), .ZN(n3803) );
  AO21D1BWP12T U3714 ( .A1(n3045), .A2(n3044), .B(n3043), .Z(n3777) );
  AO21D1BWP12T U3715 ( .A1(n3048), .A2(n3047), .B(n3046), .Z(n3752) );
  AO21D1BWP12T U3716 ( .A1(n3051), .A2(n3050), .B(n3049), .Z(n3715) );
  AOI21D1BWP12T U3717 ( .A1(n3054), .A2(n3053), .B(n3052), .ZN(n3696) );
  AOI21D1BWP12T U3718 ( .A1(n3057), .A2(n3056), .B(n3055), .ZN(n3667) );
  AOI21D1BWP12T U3719 ( .A1(n3059), .A2(n3629), .B(n3058), .ZN(n3643) );
  AO21D1BWP12T U3720 ( .A1(n3062), .A2(n3061), .B(n3060), .Z(n3620) );
  AO21D1BWP12T U3721 ( .A1(n3065), .A2(n3064), .B(n3063), .Z(n3594) );
  AO21D1BWP12T U3722 ( .A1(n3068), .A2(n3067), .B(n3066), .Z(n3562) );
  AOI21D1BWP12T U3723 ( .A1(n3071), .A2(n3070), .B(n3069), .ZN(n3543) );
  AOI21D1BWP12T U3724 ( .A1(n3074), .A2(n3073), .B(n3072), .ZN(n3514) );
  AOI21D1BWP12T U3725 ( .A1(n3077), .A2(n3076), .B(n3075), .ZN(n3485) );
  AO21D1BWP12T U3726 ( .A1(n3080), .A2(n3079), .B(n3078), .Z(n3464) );
  AO21D1BWP12T U3727 ( .A1(n3083), .A2(n3082), .B(n3081), .Z(n3437) );
  AO21D1BWP12T U3728 ( .A1(n3086), .A2(n3085), .B(n3084), .Z(n3410) );
  AOI21D1BWP12T U3729 ( .A1(n3089), .A2(n3088), .B(n3087), .ZN(n3392) );
  AOI21D1BWP12T U3730 ( .A1(n3092), .A2(n3091), .B(n3090), .ZN(n3360) );
  AOI21D1BWP12T U3731 ( .A1(n3095), .A2(n3094), .B(n3093), .ZN(n3333) );
  AO21D1BWP12T U3732 ( .A1(n3098), .A2(n3097), .B(n3096), .Z(n3233) );
  AO21D1BWP12T U3733 ( .A1(n3101), .A2(n3100), .B(n3099), .Z(n3986) );
  ND2D1BWP12T U3734 ( .A1(n3268), .A2(n3102), .ZN(n3956) );
  INVD1BWP12T U3735 ( .I(n3956), .ZN(n3987) );
  OAI21D1BWP12T U3736 ( .A1(n3105), .A2(n3104), .B(n3103), .ZN(n3166) );
  OAI21D1BWP12T U3737 ( .A1(n3108), .A2(n3107), .B(n3106), .ZN(n3955) );
  ND4D1BWP12T U3738 ( .A1(n3987), .A2(n3166), .A3(n3955), .A4(n3145), .ZN(
        n3119) );
  AOI21D1BWP12T U3739 ( .A1(n3111), .A2(n3110), .B(n3109), .ZN(n3310) );
  AOI21D1BWP12T U3740 ( .A1(n3114), .A2(n3113), .B(n3112), .ZN(n3282) );
  AOI21D1BWP12T U3741 ( .A1(n3117), .A2(n3116), .B(n3115), .ZN(n3256) );
  ND3D1BWP12T U3742 ( .A1(n3310), .A2(n3282), .A3(n3256), .ZN(n3118) );
  NR4D0BWP12T U3743 ( .A1(n3233), .A2(n3986), .A3(n3119), .A4(n3118), .ZN(
        n3120) );
  ND4D1BWP12T U3744 ( .A1(n3392), .A2(n3360), .A3(n3333), .A4(n3120), .ZN(
        n3121) );
  NR4D0BWP12T U3745 ( .A1(n3464), .A2(n3437), .A3(n3410), .A4(n3121), .ZN(
        n3122) );
  ND4D1BWP12T U3746 ( .A1(n3543), .A2(n3514), .A3(n3485), .A4(n3122), .ZN(
        n3123) );
  NR4D0BWP12T U3747 ( .A1(n3620), .A2(n3594), .A3(n3562), .A4(n3123), .ZN(
        n3124) );
  ND4D1BWP12T U3748 ( .A1(n3696), .A2(n3667), .A3(n3643), .A4(n3124), .ZN(
        n3125) );
  NR4D0BWP12T U3749 ( .A1(n3777), .A2(n3752), .A3(n3715), .A4(n3125), .ZN(
        n3126) );
  ND4D1BWP12T U3750 ( .A1(n3863), .A2(n3826), .A3(n3803), .A4(n3126), .ZN(
        n3127) );
  NR4D0BWP12T U3751 ( .A1(n3212), .A2(n3930), .A3(n3896), .A4(n3127), .ZN(
        n3128) );
  AOI31D1BWP12T U3752 ( .A1(n3215), .A2(n3927), .A3(n3129), .B(n3128), .ZN(
        n3130) );
  OAI211D1BWP12T U3753 ( .A1(n3132), .A2(n3151), .B(n3131), .C(n3130), .ZN(z)
         );
  INVD1BWP12T U3754 ( .I(n3135), .ZN(n3134) );
  OAI21D1BWP12T U3755 ( .A1(n3134), .A2(n3133), .B(n3987), .ZN(n3136) );
  INVD1BWP12T U3756 ( .I(n3906), .ZN(n3975) );
  AOI32D1BWP12T U3757 ( .A1(n3137), .A2(n3136), .A3(n3135), .B1(n3975), .B2(
        n3136), .ZN(n3138) );
  OAI32D1BWP12T U3758 ( .A1(n3139), .A2(a[31]), .A3(b[31]), .B1(n3138), .B2(
        n3139), .ZN(n3141) );
  ND2D1BWP12T U3759 ( .A1(n3140), .A2(n3931), .ZN(n3206) );
  OAI211D1BWP12T U3760 ( .A1(n3143), .A2(n3142), .B(n3141), .C(n3206), .ZN(
        c_out) );
  INVD1BWP12T U3761 ( .I(n3265), .ZN(n3982) );
  OAI32D1BWP12T U3762 ( .A1(n3981), .A2(n3982), .A3(n3996), .B1(n3144), .B2(
        n3981), .ZN(n3161) );
  NR2D1BWP12T U3763 ( .A1(n3908), .A2(n3920), .ZN(n3502) );
  OAI32D1BWP12T U3764 ( .A1(n3170), .A2(a[0]), .A3(n3724), .B1(n3988), .B2(
        n3170), .ZN(n3157) );
  ND2D1BWP12T U3765 ( .A1(n3650), .A2(n3724), .ZN(n3840) );
  INVD1BWP12T U3766 ( .I(n3840), .ZN(n3989) );
  AOI211D1BWP12T U3767 ( .A1(b[0]), .A2(n4003), .B(n3945), .C(n3940), .ZN(
        n3146) );
  OAI22D1BWP12T U3768 ( .A1(n3146), .A2(n3169), .B1(n3956), .B2(n3145), .ZN(
        n3150) );
  INVD1BWP12T U3769 ( .I(n3531), .ZN(n3938) );
  OAI22D1BWP12T U3770 ( .A1(n3148), .A2(n3949), .B1(n3147), .B2(n3938), .ZN(
        n3149) );
  AOI211D1BWP12T U3771 ( .A1(n3959), .A2(n3169), .B(n3150), .C(n3149), .ZN(
        n3154) );
  ND2D1BWP12T U3772 ( .A1(n3152), .A2(n3151), .ZN(n3153) );
  OAI211D1BWP12T U3773 ( .A1(n3989), .A2(n3155), .B(n3154), .C(n3153), .ZN(
        n3156) );
  AOI211D1BWP12T U3774 ( .A1(n3502), .A2(n3158), .B(n3157), .C(n3156), .ZN(
        n3160) );
  ND2D1BWP12T U3775 ( .A1(n3996), .A2(n3159), .ZN(n3963) );
  OAI211D1BWP12T U3776 ( .A1(n3162), .A2(n3161), .B(n3160), .C(n3963), .ZN(
        result[0]) );
  INVD1BWP12T U3777 ( .I(n3502), .ZN(n3325) );
  NR2D1BWP12T U3778 ( .A1(n3325), .A2(b[3]), .ZN(n3984) );
  OAI22D1BWP12T U3779 ( .A1(a[1]), .A2(n3724), .B1(n3938), .B2(n3163), .ZN(
        n3164) );
  AOI211D1BWP12T U3780 ( .A1(n3165), .A2(n3840), .B(n3940), .C(n3164), .ZN(
        n3167) );
  OAI22D1BWP12T U3781 ( .A1(n3168), .A2(n3167), .B1(n3166), .B2(n3956), .ZN(
        n3184) );
  NR3D1BWP12T U3782 ( .A1(n3961), .A2(n3170), .A3(n3169), .ZN(n3171) );
  MUX2ND0BWP12T U3783 ( .I0(n3173), .I1(n3172), .S(n3171), .ZN(n3182) );
  INVD1BWP12T U3784 ( .I(n3963), .ZN(n4002) );
  AOI211D1BWP12T U3785 ( .A1(a[0]), .A2(a[1]), .B(n3174), .C(n3990), .ZN(n3180) );
  OAI22D1BWP12T U3786 ( .A1(a[1]), .A2(n3995), .B1(n3175), .B2(n3975), .ZN(
        n3179) );
  OAI22D1BWP12T U3787 ( .A1(n3177), .A2(n3976), .B1(n3949), .B2(n3176), .ZN(
        n3178) );
  NR4D0BWP12T U3788 ( .A1(n4002), .A2(n3180), .A3(n3179), .A4(n3178), .ZN(
        n3181) );
  OAI21D1BWP12T U3789 ( .A1(n3958), .A2(n3182), .B(n3181), .ZN(n3183) );
  AOI211D1BWP12T U3790 ( .A1(n3185), .A2(n3984), .B(n3184), .C(n3183), .ZN(
        n3191) );
  IOA21D1BWP12T U3791 ( .A1(n3980), .A2(n3187), .B(n3186), .ZN(n3188) );
  AOI22D1BWP12T U3792 ( .A1(n3982), .A2(n3189), .B1(n3981), .B2(n3188), .ZN(
        n3190) );
  OAI211D1BWP12T U3793 ( .A1(n3192), .A2(n3831), .B(n3191), .C(n3190), .ZN(
        result[1]) );
  OAI221D1BWP12T U3794 ( .A1(b[31]), .A2(n3989), .B1(n3193), .B2(n3938), .C(
        n3831), .ZN(n3204) );
  NR2D1BWP12T U3795 ( .A1(a[31]), .A2(b[31]), .ZN(n3198) );
  AOI32D1BWP12T U3796 ( .A1(b[31]), .A2(n3194), .A3(n3823), .B1(n3959), .B2(
        n3194), .ZN(n3197) );
  INVD1BWP12T U3797 ( .I(n3195), .ZN(n3196) );
  OAI211D1BWP12T U3798 ( .A1(n3198), .A2(n3988), .B(n3197), .C(n3196), .ZN(
        n3203) );
  ND2D1BWP12T U3799 ( .A1(n3199), .A2(n3982), .ZN(n3792) );
  OAI21D1BWP12T U3800 ( .A1(n3891), .A2(b[4]), .B(n3792), .ZN(n3766) );
  INVD1BWP12T U3801 ( .I(n3766), .ZN(n3922) );
  OAI22D1BWP12T U3802 ( .A1(n3922), .A2(n3201), .B1(n3920), .B2(n3200), .ZN(
        n3202) );
  AO211D1BWP12T U3803 ( .A1(a[31]), .A2(n3204), .B(n3203), .C(n3202), .Z(n3209) );
  OAI211D1BWP12T U3804 ( .A1(n3207), .A2(n3976), .B(n3206), .C(n3205), .ZN(
        n3208) );
  AOI211D1BWP12T U3805 ( .A1(n3981), .A2(n3210), .B(n3209), .C(n3208), .ZN(
        n3214) );
  AOI22D1BWP12T U3806 ( .A1(n3987), .A2(n3212), .B1(n3906), .B2(n3211), .ZN(
        n3213) );
  OAI211D1BWP12T U3807 ( .A1(n3215), .A2(n3949), .B(n3214), .C(n3213), .ZN(
        result[31]) );
  CKBD1BWP12T U3808 ( .I(result[31]), .Z(n) );
  AOI22D1BWP12T U3809 ( .A1(n3999), .A2(n3217), .B1(n3216), .B2(n3982), .ZN(
        n3235) );
  ND2D1BWP12T U3810 ( .A1(n3724), .A2(n3988), .ZN(n3960) );
  INVD1BWP12T U3811 ( .I(n3960), .ZN(n4001) );
  OAI32D1BWP12T U3812 ( .A1(a[4]), .A2(n4001), .A3(n3219), .B1(n3995), .B2(
        a[4]), .ZN(n3225) );
  NR2D1BWP12T U3813 ( .A1(a[3]), .A2(n3992), .ZN(n3991) );
  OAI21D1BWP12T U3814 ( .A1(n3991), .A2(n3218), .B(n3945), .ZN(n3223) );
  OAI221D1BWP12T U3815 ( .A1(b[4]), .A2(n3840), .B1(n3219), .B2(n3531), .C(
        a[4]), .ZN(n3222) );
  AOI22D1BWP12T U3816 ( .A1(a[4]), .A2(n3940), .B1(n4003), .B2(n3220), .ZN(
        n3221) );
  OAI211D1BWP12T U3817 ( .A1(n3248), .A2(n3223), .B(n3222), .C(n3221), .ZN(
        n3224) );
  AOI211D1BWP12T U3818 ( .A1(n3226), .A2(n3926), .B(n3225), .C(n3224), .ZN(
        n3230) );
  AOI22D1BWP12T U3819 ( .A1(n3906), .A2(n3228), .B1(n3984), .B2(n3227), .ZN(
        n3229) );
  OAI211D1BWP12T U3820 ( .A1(n3231), .A2(n3891), .B(n3230), .C(n3229), .ZN(
        n3232) );
  AOI21D1BWP12T U3821 ( .A1(n3987), .A2(n3233), .B(n3232), .ZN(n3234) );
  OAI211D1BWP12T U3822 ( .A1(n3236), .A2(n3831), .B(n3235), .C(n3234), .ZN(
        result[4]) );
  AOI22D1BWP12T U3823 ( .A1(n3906), .A2(n3238), .B1(n3981), .B2(n3237), .ZN(
        n3261) );
  INVD1BWP12T U3824 ( .I(n3984), .ZN(n3302) );
  OAI22D1BWP12T U3825 ( .A1(n3240), .A2(n3724), .B1(n3239), .B2(n3938), .ZN(
        n3245) );
  AOI22D1BWP12T U3826 ( .A1(n3940), .A2(n3241), .B1(n3959), .B2(n3247), .ZN(
        n3242) );
  OAI21D1BWP12T U3827 ( .A1(n3989), .A2(n3243), .B(n3242), .ZN(n3244) );
  AOI211D1BWP12T U3828 ( .A1(n4003), .A2(n3246), .B(n3245), .C(n3244), .ZN(
        n3250) );
  OAI211D1BWP12T U3829 ( .A1(n3248), .A2(n3247), .B(n3945), .C(n3297), .ZN(
        n3249) );
  OAI211D1BWP12T U3830 ( .A1(n3251), .A2(n3302), .B(n3250), .C(n3249), .ZN(
        n3252) );
  AOI211D1BWP12T U3831 ( .A1(n3253), .A2(n3982), .B(n4002), .C(n3252), .ZN(
        n3260) );
  AOI22D1BWP12T U3832 ( .A1(n3926), .A2(n3255), .B1(n3996), .B2(n3254), .ZN(
        n3259) );
  MAOI22D0BWP12T U3833 ( .A1(n3999), .A2(n3257), .B1(n3256), .B2(n3956), .ZN(
        n3258) );
  ND4D1BWP12T U3834 ( .A1(n3261), .A2(n3260), .A3(n3259), .A4(n3258), .ZN(
        result[5]) );
  AOI22D1BWP12T U3835 ( .A1(n3906), .A2(n3263), .B1(n3981), .B2(n3262), .ZN(
        n3287) );
  OAI22D1BWP12T U3836 ( .A1(n3266), .A2(n3265), .B1(n3264), .B2(n3302), .ZN(
        n3280) );
  NR2D1BWP12T U3837 ( .A1(a[6]), .A2(n3297), .ZN(n3267) );
  AOI211D1BWP12T U3838 ( .A1(a[6]), .A2(n3297), .B(n3267), .C(n3990), .ZN(
        n3275) );
  NR2D1BWP12T U3839 ( .A1(n3269), .A2(n3268), .ZN(n3833) );
  INVD1BWP12T U3840 ( .I(n3833), .ZN(n3994) );
  AOI22D1BWP12T U3841 ( .A1(n3271), .A2(n3960), .B1(n4003), .B2(n3270), .ZN(
        n3272) );
  OAI21D1BWP12T U3842 ( .A1(n3273), .A2(n3994), .B(n3272), .ZN(n3274) );
  AOI211D1BWP12T U3843 ( .A1(n3959), .A2(n3276), .B(n3275), .C(n3274), .ZN(
        n3279) );
  AOI32D1BWP12T U3844 ( .A1(n3840), .A2(a[6]), .A3(n3277), .B1(n3940), .B2(
        a[6]), .ZN(n3278) );
  IND4D1BWP12T U3845 ( .A1(n3280), .B1(n3279), .B2(n3963), .B3(n3278), .ZN(
        n3284) );
  OAI22D1BWP12T U3846 ( .A1(n3282), .A2(n3956), .B1(n3949), .B2(n3281), .ZN(
        n3283) );
  AOI211D1BWP12T U3847 ( .A1(n3926), .A2(n3285), .B(n3284), .C(n3283), .ZN(
        n3286) );
  OAI211D1BWP12T U3848 ( .A1(n3288), .A2(n3831), .B(n3287), .C(n3286), .ZN(
        result[6]) );
  MOAI22D0BWP12T U3849 ( .A1(n3290), .A2(n3994), .B1(n4003), .B2(n3289), .ZN(
        n3295) );
  ND2D1BWP12T U3850 ( .A1(n3291), .A2(n3840), .ZN(n3293) );
  AOI32D1BWP12T U3851 ( .A1(n3988), .A2(a[7]), .A3(n3293), .B1(n3995), .B2(
        n3292), .ZN(n3294) );
  AOI211D1BWP12T U3852 ( .A1(n3296), .A2(n3960), .B(n3295), .C(n3294), .ZN(
        n3301) );
  OAI32D1BWP12T U3853 ( .A1(n3322), .A2(a[6]), .A3(n3297), .B1(a[7]), .B2(
        n3322), .ZN(n3299) );
  AOI22D1BWP12T U3854 ( .A1(n3945), .A2(n3299), .B1(n3981), .B2(n3298), .ZN(
        n3300) );
  OAI211D1BWP12T U3855 ( .A1(n3303), .A2(n3302), .B(n3301), .C(n3300), .ZN(
        n3307) );
  OAI22D1BWP12T U3856 ( .A1(n3305), .A2(n3976), .B1(n3304), .B2(n3831), .ZN(
        n3306) );
  AOI211D1BWP12T U3857 ( .A1(n3982), .A2(n3308), .B(n3307), .C(n3306), .ZN(
        n3312) );
  OA22D1BWP12T U3858 ( .A1(n3310), .A2(n3956), .B1(n3309), .B2(n3949), .Z(
        n3311) );
  OAI211D1BWP12T U3859 ( .A1(n3313), .A2(n3975), .B(n3312), .C(n3311), .ZN(
        result[7]) );
  OAI21D1BWP12T U3860 ( .A1(n3506), .A2(n3736), .B(n3314), .ZN(n3336) );
  AOI22D1BWP12T U3861 ( .A1(n3982), .A2(n3316), .B1(n3996), .B2(n3315), .ZN(
        n3330) );
  MOAI22D0BWP12T U3862 ( .A1(n3318), .A2(n3938), .B1(n4003), .B2(n3317), .ZN(
        n3319) );
  AOI221D1BWP12T U3863 ( .A1(n3940), .A2(a[8]), .B1(n3959), .B2(n3321), .C(
        n3319), .ZN(n3320) );
  OAI31D1BWP12T U3864 ( .A1(b[8]), .A2(n3989), .A3(n3321), .B(n3320), .ZN(
        n3327) );
  OAI211D1BWP12T U3865 ( .A1(n3322), .A2(n3321), .B(n3945), .C(n3339), .ZN(
        n3323) );
  OAI211D1BWP12T U3866 ( .A1(n3325), .A2(n3324), .B(n3963), .C(n3323), .ZN(
        n3326) );
  AOI211D1BWP12T U3867 ( .A1(n3328), .A2(n3960), .B(n3327), .C(n3326), .ZN(
        n3329) );
  OAI211D1BWP12T U3868 ( .A1(n3976), .A2(n3331), .B(n3330), .C(n3329), .ZN(
        n3335) );
  OAI22D1BWP12T U3869 ( .A1(n3333), .A2(n3956), .B1(n3949), .B2(n3332), .ZN(
        n3334) );
  AOI211D1BWP12T U3870 ( .A1(n3981), .A2(n3336), .B(n3335), .C(n3334), .ZN(
        n3337) );
  OAI21D1BWP12T U3871 ( .A1(n3338), .A2(n3975), .B(n3337), .ZN(result[8]) );
  AOI211D1BWP12T U3872 ( .A1(a[9]), .A2(n3339), .B(n3381), .C(n3990), .ZN(
        n3351) );
  AOI22D1BWP12T U3873 ( .A1(a[9]), .A2(n3940), .B1(n4003), .B2(n3340), .ZN(
        n3348) );
  OAI21D1BWP12T U3874 ( .A1(n4001), .A2(n3341), .B(n3995), .ZN(n3345) );
  OAI22D1BWP12T U3875 ( .A1(n3989), .A2(n3343), .B1(n3342), .B2(n3938), .ZN(
        n3344) );
  AOI211D1BWP12T U3876 ( .A1(n3346), .A2(n3345), .B(n4002), .C(n3344), .ZN(
        n3347) );
  OAI211D1BWP12T U3877 ( .A1(n3831), .A2(n3349), .B(n3348), .C(n3347), .ZN(
        n3350) );
  AOI211D1BWP12T U3878 ( .A1(n3502), .A2(n3352), .B(n3351), .C(n3350), .ZN(
        n3358) );
  OAI21D1BWP12T U3879 ( .A1(n3354), .A2(n3506), .B(n3353), .ZN(n3355) );
  AOI22D1BWP12T U3880 ( .A1(n3356), .A2(n3982), .B1(n3981), .B2(n3355), .ZN(
        n3357) );
  OAI211D1BWP12T U3881 ( .A1(n3359), .A2(n3976), .B(n3358), .C(n3357), .ZN(
        n3363) );
  OAI22D1BWP12T U3882 ( .A1(n3361), .A2(n3975), .B1(n3360), .B2(n3956), .ZN(
        n3362) );
  AO211D1BWP12T U3883 ( .A1(n3999), .A2(n3364), .B(n3363), .C(n3362), .Z(
        result[9]) );
  MOAI22D0BWP12T U3884 ( .A1(n3831), .A2(n3366), .B1(n3982), .B2(n3365), .ZN(
        n3386) );
  OAI21D1BWP12T U3885 ( .A1(n3368), .A2(n3506), .B(n3367), .ZN(n3369) );
  AOI31D1BWP12T U3886 ( .A1(b[4]), .A2(n2886), .A3(n3783), .B(n3369), .ZN(
        n3384) );
  ND2D1BWP12T U3887 ( .A1(a[10]), .A2(n3370), .ZN(n3377) );
  AOI22D1BWP12T U3888 ( .A1(n3371), .A2(n4003), .B1(n3959), .B2(n3380), .ZN(
        n3376) );
  OAI22D1BWP12T U3889 ( .A1(a[10]), .A2(n3724), .B1(n3938), .B2(n3372), .ZN(
        n3374) );
  OAI21D1BWP12T U3890 ( .A1(n3940), .A2(n3374), .B(n3373), .ZN(n3375) );
  OAI211D1BWP12T U3891 ( .A1(n3989), .A2(n3377), .B(n3376), .C(n3375), .ZN(
        n3378) );
  AOI211D1BWP12T U3892 ( .A1(n3502), .A2(n3379), .B(n4002), .C(n3378), .ZN(
        n3383) );
  ND2D1BWP12T U3893 ( .A1(n3381), .A2(n3380), .ZN(n3393) );
  OAI211D1BWP12T U3894 ( .A1(n3381), .A2(n3380), .B(n3945), .C(n3393), .ZN(
        n3382) );
  OAI211D1BWP12T U3895 ( .A1(n3384), .A2(n3891), .B(n3383), .C(n3382), .ZN(
        n3385) );
  AOI211D1BWP12T U3896 ( .A1(n3926), .A2(n3387), .B(n3386), .C(n3385), .ZN(
        n3391) );
  AOI22D1BWP12T U3897 ( .A1(n3999), .A2(n3389), .B1(n3906), .B2(n3388), .ZN(
        n3390) );
  OAI211D1BWP12T U3898 ( .A1(n3392), .A2(n3956), .B(n3391), .C(n3390), .ZN(
        result[10]) );
  AOI211D1BWP12T U3899 ( .A1(a[11]), .A2(n3393), .B(n3429), .C(n3990), .ZN(
        n3404) );
  MAOI22D0BWP12T U3900 ( .A1(n4003), .A2(n3395), .B1(n3394), .B2(n3938), .ZN(
        n3402) );
  AOI31D1BWP12T U3901 ( .A1(b[11]), .A2(n3960), .A3(n4005), .B(n4002), .ZN(
        n3401) );
  AOI22D1BWP12T U3902 ( .A1(n3996), .A2(n3397), .B1(n3502), .B2(n3396), .ZN(
        n3400) );
  NR2D1BWP12T U3903 ( .A1(b[11]), .A2(n3989), .ZN(n3398) );
  OAI32D1BWP12T U3904 ( .A1(n4005), .A2(n3940), .A3(n3398), .B1(a[11]), .B2(
        n3959), .ZN(n3399) );
  ND4D1BWP12T U3905 ( .A1(n3402), .A2(n3401), .A3(n3400), .A4(n3399), .ZN(
        n3403) );
  AOI211D1BWP12T U3906 ( .A1(n3982), .A2(n3405), .B(n3404), .C(n3403), .ZN(
        n3415) );
  IOA21D1BWP12T U3907 ( .A1(n3818), .A2(n3817), .B(n3406), .ZN(n3407) );
  AOI22D1BWP12T U3908 ( .A1(n3926), .A2(n3408), .B1(n3981), .B2(n3407), .ZN(
        n3414) );
  AOI22D1BWP12T U3909 ( .A1(n3987), .A2(n3410), .B1(n3906), .B2(n3409), .ZN(
        n3413) );
  ND2D1BWP12T U3910 ( .A1(n3999), .A2(n3411), .ZN(n3412) );
  ND4D1BWP12T U3911 ( .A1(n3415), .A2(n3414), .A3(n3413), .A4(n3412), .ZN(
        result[11]) );
  OAI21D1BWP12T U3912 ( .A1(n4001), .A2(n3416), .B(n3995), .ZN(n3420) );
  MOAI22D0BWP12T U3913 ( .A1(n3418), .A2(n3938), .B1(n4003), .B2(n3417), .ZN(
        n3419) );
  AOI221D1BWP12T U3914 ( .A1(n3940), .A2(a[12]), .B1(n3420), .B2(n3428), .C(
        n3419), .ZN(n3425) );
  OAI32D1BWP12T U3915 ( .A1(n3891), .A2(n3506), .A3(n3835), .B1(n3421), .B2(
        n3891), .ZN(n3422) );
  AOI211D1BWP12T U3916 ( .A1(n3502), .A2(n3423), .B(n4002), .C(n3422), .ZN(
        n3424) );
  OAI211D1BWP12T U3917 ( .A1(n3989), .A2(n3426), .B(n3425), .C(n3424), .ZN(
        n3434) );
  ND2D1BWP12T U3918 ( .A1(n3982), .A2(n3427), .ZN(n3431) );
  ND2D1BWP12T U3919 ( .A1(n3429), .A2(n3428), .ZN(n3453) );
  OAI211D1BWP12T U3920 ( .A1(n3429), .A2(n3428), .B(n3945), .C(n3453), .ZN(
        n3430) );
  OAI211D1BWP12T U3921 ( .A1(n3432), .A2(n3831), .B(n3431), .C(n3430), .ZN(
        n3433) );
  AOI211D1BWP12T U3922 ( .A1(n3926), .A2(n3435), .B(n3434), .C(n3433), .ZN(
        n3439) );
  AOI22D1BWP12T U3923 ( .A1(n3987), .A2(n3437), .B1(n3906), .B2(n3436), .ZN(
        n3438) );
  OAI211D1BWP12T U3924 ( .A1(n3440), .A2(n3949), .B(n3439), .C(n3438), .ZN(
        result[12]) );
  MOAI22D0BWP12T U3925 ( .A1(n3442), .A2(n3938), .B1(n4003), .B2(n3441), .ZN(
        n3448) );
  AOI22D1BWP12T U3926 ( .A1(n3444), .A2(n3960), .B1(n3443), .B2(n3840), .ZN(
        n3445) );
  OAI221D1BWP12T U3927 ( .A1(a[13]), .A2(n3995), .B1(n3446), .B2(n3988), .C(
        n3445), .ZN(n3447) );
  AO211D1BWP12T U3928 ( .A1(n3996), .A2(n3449), .B(n3448), .C(n3447), .Z(n3450) );
  AOI211D1BWP12T U3929 ( .A1(n3502), .A2(n3451), .B(n4002), .C(n3450), .ZN(
        n3458) );
  OAI32D1BWP12T U3930 ( .A1(n3891), .A2(n3885), .A3(n3506), .B1(n3452), .B2(
        n3891), .ZN(n3455) );
  AOI211D1BWP12T U3931 ( .A1(a[13]), .A2(n3453), .B(n3480), .C(n3990), .ZN(
        n3454) );
  AOI211D1BWP12T U3932 ( .A1(n3456), .A2(n3982), .B(n3455), .C(n3454), .ZN(
        n3457) );
  OAI211D1BWP12T U3933 ( .A1(n3976), .A2(n3459), .B(n3458), .C(n3457), .ZN(
        n3463) );
  OAI22D1BWP12T U3934 ( .A1(n3461), .A2(n3975), .B1(n3460), .B2(n3949), .ZN(
        n3462) );
  AO211D1BWP12T U3935 ( .A1(n3987), .A2(n3464), .B(n3463), .C(n3462), .Z(
        result[13]) );
  OAI32D1BWP12T U3936 ( .A1(a[14]), .A2(n4001), .A3(n3465), .B1(n3995), .B2(
        a[14]), .ZN(n3468) );
  MOAI22D0BWP12T U3937 ( .A1(n3479), .A2(n3988), .B1(n4003), .B2(n3466), .ZN(
        n3467) );
  AOI211D1BWP12T U3938 ( .A1(n3469), .A2(n3840), .B(n3468), .C(n3467), .ZN(
        n3473) );
  AOI22D1BWP12T U3939 ( .A1(n3471), .A2(n3502), .B1(n3996), .B2(n3470), .ZN(
        n3472) );
  OAI211D1BWP12T U3940 ( .A1(n3474), .A2(n3938), .B(n3473), .C(n3472), .ZN(
        n3488) );
  OAI21D1BWP12T U3941 ( .A1(n3476), .A2(n3506), .B(n3475), .ZN(n3477) );
  AOI22D1BWP12T U3942 ( .A1(n3982), .A2(n3478), .B1(n3981), .B2(n3477), .ZN(
        n3482) );
  OAI211D1BWP12T U3943 ( .A1(n3480), .A2(n3479), .B(n3945), .C(n3504), .ZN(
        n3481) );
  OAI211D1BWP12T U3944 ( .A1(n3483), .A2(n3976), .B(n3482), .C(n3481), .ZN(
        n3487) );
  OAI22D1BWP12T U3945 ( .A1(n3485), .A2(n3956), .B1(n3949), .B2(n3484), .ZN(
        n3486) );
  NR4D0BWP12T U3946 ( .A1(n4002), .A2(n3488), .A3(n3487), .A4(n3486), .ZN(
        n3489) );
  OAI21D1BWP12T U3947 ( .A1(n3490), .A2(n3975), .B(n3489), .ZN(result[14]) );
  OAI22D1BWP12T U3948 ( .A1(a[15]), .A2(n3995), .B1(n3989), .B2(n3491), .ZN(
        n3501) );
  NR2D1BWP12T U3949 ( .A1(n3899), .A2(n3492), .ZN(n3499) );
  MAOI22D0BWP12T U3950 ( .A1(n3494), .A2(n3823), .B1(n3493), .B2(n3938), .ZN(
        n3498) );
  AOI22D1BWP12T U3951 ( .A1(n4003), .A2(n3496), .B1(n3940), .B2(n3495), .ZN(
        n3497) );
  OAI211D1BWP12T U3952 ( .A1(n3499), .A2(n3831), .B(n3498), .C(n3497), .ZN(
        n3500) );
  AOI211D1BWP12T U3953 ( .A1(n3503), .A2(n3502), .B(n3501), .C(n3500), .ZN(
        n3512) );
  NR2D1BWP12T U3954 ( .A1(a[15]), .A2(n3504), .ZN(n3530) );
  AOI211D1BWP12T U3955 ( .A1(a[15]), .A2(n3504), .B(n3530), .C(n3990), .ZN(
        n3509) );
  OAI32D1BWP12T U3956 ( .A1(n3891), .A2(n3507), .A3(n3506), .B1(n3505), .B2(
        n3891), .ZN(n3508) );
  AOI211D1BWP12T U3957 ( .A1(n3510), .A2(n3982), .B(n3509), .C(n3508), .ZN(
        n3511) );
  OAI211D1BWP12T U3958 ( .A1(n3513), .A2(n3976), .B(n3512), .C(n3511), .ZN(
        n3517) );
  OAI22D1BWP12T U3959 ( .A1(n3515), .A2(n3975), .B1(n3514), .B2(n3956), .ZN(
        n3516) );
  AO211D1BWP12T U3960 ( .A1(n3999), .A2(n3518), .B(n3517), .C(n3516), .Z(
        result[15]) );
  OAI22D1BWP12T U3961 ( .A1(n3922), .A2(n3520), .B1(n3920), .B2(n3519), .ZN(
        n3537) );
  AOI22D1BWP12T U3962 ( .A1(n3521), .A2(n4003), .B1(n3959), .B2(n3529), .ZN(
        n3535) );
  MOAI22D0BWP12T U3963 ( .A1(n3989), .A2(n3523), .B1(n3960), .B2(n3522), .ZN(
        n3524) );
  AO31D1BWP12T U3964 ( .A1(b[4]), .A2(n3981), .A3(n3525), .B(n3524), .Z(n3527)
         );
  OAI32D1BWP12T U3965 ( .A1(n3527), .A2(n3899), .A3(n3526), .B1(n3996), .B2(
        n3527), .ZN(n3534) );
  INVD1BWP12T U3966 ( .I(n3566), .ZN(n3528) );
  OAI211D1BWP12T U3967 ( .A1(n3530), .A2(n3529), .B(n3945), .C(n3528), .ZN(
        n3533) );
  AOI32D1BWP12T U3968 ( .A1(b[16]), .A2(a[16]), .A3(n3531), .B1(n3940), .B2(
        a[16]), .ZN(n3532) );
  ND4D1BWP12T U3969 ( .A1(n3535), .A2(n3534), .A3(n3533), .A4(n3532), .ZN(
        n3536) );
  AOI211D1BWP12T U3970 ( .A1(n3926), .A2(n3538), .B(n3537), .C(n3536), .ZN(
        n3542) );
  AOI22D1BWP12T U3971 ( .A1(n3999), .A2(n3540), .B1(n3906), .B2(n3539), .ZN(
        n3541) );
  OAI211D1BWP12T U3972 ( .A1(n3543), .A2(n3956), .B(n3542), .C(n3541), .ZN(
        result[16]) );
  NR3D1BWP12T U3973 ( .A1(n3544), .A2(a[17]), .A3(n4001), .ZN(n3547) );
  ND2D1BWP12T U3974 ( .A1(n3544), .A2(n3840), .ZN(n3545) );
  AOI32D1BWP12T U3975 ( .A1(n3988), .A2(a[17]), .A3(n3545), .B1(n3565), .B2(
        n3995), .ZN(n3546) );
  AOI211D1BWP12T U3976 ( .A1(n3548), .A2(n4003), .B(n3547), .C(n3546), .ZN(
        n3555) );
  OAI22D1BWP12T U3977 ( .A1(n3551), .A2(n3550), .B1(n3603), .B2(n3549), .ZN(
        n3552) );
  AOI32D1BWP12T U3978 ( .A1(n3889), .A2(n3981), .A3(n3553), .B1(n3552), .B2(
        n3981), .ZN(n3554) );
  OAI211D1BWP12T U3979 ( .A1(n3938), .A2(n3556), .B(n3555), .C(n3554), .ZN(
        n3560) );
  OAI22D1BWP12T U3980 ( .A1(n3922), .A2(n3558), .B1(n3920), .B2(n3557), .ZN(
        n3559) );
  AOI211D1BWP12T U3981 ( .A1(n3926), .A2(n3561), .B(n3560), .C(n3559), .ZN(
        n3570) );
  AOI22D1BWP12T U3982 ( .A1(n3999), .A2(n3563), .B1(n3987), .B2(n3562), .ZN(
        n3569) );
  OAI21D1BWP12T U3983 ( .A1(n3899), .A2(n3564), .B(n3996), .ZN(n3568) );
  ND2D1BWP12T U3984 ( .A1(n3566), .A2(n3565), .ZN(n3573) );
  OAI211D1BWP12T U3985 ( .A1(n3566), .A2(n3565), .B(n3945), .C(n3573), .ZN(
        n3567) );
  ND4D1BWP12T U3986 ( .A1(n3570), .A2(n3569), .A3(n3568), .A4(n3567), .ZN(
        n3571) );
  AO21D1BWP12T U3987 ( .A1(n3906), .A2(n3572), .B(n3571), .Z(result[17]) );
  NR2D1BWP12T U3988 ( .A1(a[18]), .A2(n3573), .ZN(n3611) );
  AOI211D1BWP12T U3989 ( .A1(a[18]), .A2(n3573), .B(n3611), .C(n3990), .ZN(
        n3591) );
  NR2D1BWP12T U3990 ( .A1(n3574), .A2(n3938), .ZN(n3576) );
  OAI32D1BWP12T U3991 ( .A1(n3578), .A2(b[18]), .A3(n3989), .B1(n3988), .B2(
        n3578), .ZN(n3575) );
  AOI211D1BWP12T U3992 ( .A1(n3577), .A2(n4003), .B(n3576), .C(n3575), .ZN(
        n3580) );
  AOI32D1BWP12T U3993 ( .A1(b[18]), .A2(n3578), .A3(n3960), .B1(n3959), .B2(
        n3578), .ZN(n3579) );
  OAI211D1BWP12T U3994 ( .A1(n3922), .A2(n3581), .B(n3580), .C(n3579), .ZN(
        n3583) );
  OAI32D1BWP12T U3995 ( .A1(n3583), .A2(n3899), .A3(n3582), .B1(n3996), .B2(
        n3583), .ZN(n3588) );
  AOI32D1BWP12T U3996 ( .A1(n3586), .A2(n3981), .A3(n3585), .B1(n3584), .B2(
        n3981), .ZN(n3587) );
  OAI211D1BWP12T U3997 ( .A1(n3589), .A2(n3920), .B(n3588), .C(n3587), .ZN(
        n3590) );
  AOI211D1BWP12T U3998 ( .A1(n3592), .A2(n3926), .B(n3591), .C(n3590), .ZN(
        n3596) );
  AOI22D1BWP12T U3999 ( .A1(n3987), .A2(n3594), .B1(n3906), .B2(n3593), .ZN(
        n3595) );
  OAI211D1BWP12T U4000 ( .A1(n3949), .A2(n3597), .B(n3596), .C(n3595), .ZN(
        result[18]) );
  OAI21D1BWP12T U4001 ( .A1(n4001), .A2(n3598), .B(n3995), .ZN(n3617) );
  OAI21D1BWP12T U4002 ( .A1(b[19]), .A2(n3989), .B(n3988), .ZN(n3600) );
  AOI22D1BWP12T U4003 ( .A1(a[19]), .A2(n3600), .B1(n4003), .B2(n3599), .ZN(
        n3607) );
  OAI32D1BWP12T U4004 ( .A1(n3891), .A2(n3603), .A3(n3602), .B1(n3601), .B2(
        n3891), .ZN(n3605) );
  OAI32D1BWP12T U4005 ( .A1(n3605), .A2(n3899), .A3(n3604), .B1(n3996), .B2(
        n3605), .ZN(n3606) );
  OAI211D1BWP12T U4006 ( .A1(n3608), .A2(n3938), .B(n3607), .C(n3606), .ZN(
        n3616) );
  MAOI22D0BWP12T U4007 ( .A1(n3610), .A2(n3766), .B1(n3920), .B2(n3609), .ZN(
        n3613) );
  OAI211D1BWP12T U4008 ( .A1(n3611), .A2(n3618), .B(n3945), .C(n3625), .ZN(
        n3612) );
  OAI211D1BWP12T U4009 ( .A1(n3614), .A2(n3976), .B(n3613), .C(n3612), .ZN(
        n3615) );
  AOI211D1BWP12T U4010 ( .A1(n3618), .A2(n3617), .B(n3616), .C(n3615), .ZN(
        n3622) );
  MAOI22D0BWP12T U4011 ( .A1(n3987), .A2(n3620), .B1(n3619), .B2(n3975), .ZN(
        n3621) );
  OAI211D1BWP12T U4012 ( .A1(n3623), .A2(n3949), .B(n3622), .C(n3621), .ZN(
        result[19]) );
  AOI21D1BWP12T U4013 ( .A1(n3907), .A2(n3624), .B(n3831), .ZN(n3641) );
  AOI211D1BWP12T U4014 ( .A1(a[20]), .A2(n3625), .B(n3686), .C(n3990), .ZN(
        n3640) );
  AOI22D1BWP12T U4015 ( .A1(b[20]), .A2(n3940), .B1(n4003), .B2(n3626), .ZN(
        n3634) );
  AOI211D1BWP12T U4016 ( .A1(n3628), .A2(n3627), .B(n3632), .C(n3994), .ZN(
        n3631) );
  AOI211D1BWP12T U4017 ( .A1(n3632), .A2(n3724), .B(n3989), .C(n3629), .ZN(
        n3630) );
  AOI211D1BWP12T U4018 ( .A1(n3959), .A2(n3632), .B(n3631), .C(n3630), .ZN(
        n3633) );
  OAI211D1BWP12T U4019 ( .A1(n3635), .A2(n3891), .B(n3634), .C(n3633), .ZN(
        n3639) );
  OAI22D1BWP12T U4020 ( .A1(n3637), .A2(n3922), .B1(n3636), .B2(n3920), .ZN(
        n3638) );
  NR4D0BWP12T U4021 ( .A1(n3641), .A2(n3640), .A3(n3639), .A4(n3638), .ZN(
        n3647) );
  OAI22D1BWP12T U4022 ( .A1(n3643), .A2(n3956), .B1(n3949), .B2(n3642), .ZN(
        n3644) );
  RCIAO21D0BWP12T U4023 ( .A1(n3645), .A2(n3975), .B(n3644), .ZN(n3646) );
  OAI211D1BWP12T U4024 ( .A1(n3648), .A2(n3976), .B(n3647), .C(n3646), .ZN(
        result[20]) );
  RCIAO21D0BWP12T U4025 ( .A1(n3899), .A2(n3649), .B(n3831), .ZN(n3661) );
  MAOI22D0BWP12T U4026 ( .A1(n3823), .A2(n3651), .B1(n3650), .B2(b[21]), .ZN(
        n3659) );
  OAI22D1BWP12T U4027 ( .A1(a[21]), .A2(n3995), .B1(n3938), .B2(n3651), .ZN(
        n3655) );
  OAI22D1BWP12T U4028 ( .A1(n3653), .A2(n3792), .B1(n3652), .B2(n3920), .ZN(
        n3654) );
  AOI211D1BWP12T U4029 ( .A1(n4003), .A2(n3656), .B(n3655), .C(n3654), .ZN(
        n3658) );
  AOI32D1BWP12T U4030 ( .A1(n3659), .A2(n3658), .A3(n3988), .B1(n3657), .B2(
        n3658), .ZN(n3660) );
  AOI211D1BWP12T U4031 ( .A1(n3981), .A2(n3662), .B(n3661), .C(n3660), .ZN(
        n3665) );
  ND2D1BWP12T U4032 ( .A1(n3686), .A2(n3685), .ZN(n3663) );
  OAI211D1BWP12T U4033 ( .A1(n3686), .A2(n3685), .B(n3945), .C(n3663), .ZN(
        n3664) );
  OAI211D1BWP12T U4034 ( .A1(n3666), .A2(n3976), .B(n3665), .C(n3664), .ZN(
        n3670) );
  OAI22D1BWP12T U4035 ( .A1(n3668), .A2(n3975), .B1(n3667), .B2(n3956), .ZN(
        n3669) );
  AO211D1BWP12T U4036 ( .A1(n3999), .A2(n3671), .B(n3670), .C(n3669), .Z(
        result[21]) );
  OAI22D1BWP12T U4037 ( .A1(a[22]), .A2(n3995), .B1(n3938), .B2(n3672), .ZN(
        n3677) );
  AOI22D1BWP12T U4038 ( .A1(a[22]), .A2(n3940), .B1(n4003), .B2(n3673), .ZN(
        n3674) );
  OAI21D1BWP12T U4039 ( .A1(n3989), .A2(n3675), .B(n3674), .ZN(n3676) );
  AOI211D1BWP12T U4040 ( .A1(n3678), .A2(n3960), .B(n3677), .C(n3676), .ZN(
        n3682) );
  INVD1BWP12T U4041 ( .I(n3792), .ZN(n3872) );
  AOI22D1BWP12T U4042 ( .A1(n3981), .A2(n3680), .B1(n3872), .B2(n3679), .ZN(
        n3681) );
  OAI211D1BWP12T U4043 ( .A1(n3920), .A2(n3683), .B(n3682), .C(n3681), .ZN(
        n3690) );
  AOI32D1BWP12T U4044 ( .A1(n3686), .A2(n3708), .A3(n3685), .B1(n3684), .B2(
        n3708), .ZN(n3687) );
  OAI22D1BWP12T U4045 ( .A1(n3688), .A2(n3831), .B1(n3990), .B2(n3687), .ZN(
        n3689) );
  AOI211D1BWP12T U4046 ( .A1(n3926), .A2(n3691), .B(n3690), .C(n3689), .ZN(
        n3695) );
  AOI22D1BWP12T U4047 ( .A1(n3999), .A2(n3693), .B1(n3906), .B2(n3692), .ZN(
        n3694) );
  OAI211D1BWP12T U4048 ( .A1(n3696), .A2(n3956), .B(n3695), .C(n3694), .ZN(
        result[22]) );
  OAI32D1BWP12T U4049 ( .A1(a[23]), .A2(n4001), .A3(n3697), .B1(n3995), .B2(
        a[23]), .ZN(n3707) );
  OAI22D1BWP12T U4050 ( .A1(n3989), .A2(n3699), .B1(n3698), .B2(n3938), .ZN(
        n3706) );
  MOAI22D0BWP12T U4051 ( .A1(n3701), .A2(n3988), .B1(n4003), .B2(n3700), .ZN(
        n3705) );
  OAI22D1BWP12T U4052 ( .A1(n3703), .A2(n3891), .B1(n3702), .B2(n3792), .ZN(
        n3704) );
  NR4D0BWP12T U4053 ( .A1(n3707), .A2(n3706), .A3(n3705), .A4(n3704), .ZN(
        n3721) );
  AOI211D1BWP12T U4054 ( .A1(a[23]), .A2(n3708), .B(n3722), .C(n3990), .ZN(
        n3713) );
  INVD1BWP12T U4055 ( .I(n3709), .ZN(n3710) );
  OAI22D1BWP12T U4056 ( .A1(n3711), .A2(n3831), .B1(n3920), .B2(n3710), .ZN(
        n3712) );
  AOI211D1BWP12T U4057 ( .A1(n3714), .A2(n3926), .B(n3713), .C(n3712), .ZN(
        n3720) );
  AOI22D1BWP12T U4058 ( .A1(n3999), .A2(n3716), .B1(n3987), .B2(n3715), .ZN(
        n3719) );
  ND2D1BWP12T U4059 ( .A1(n3906), .A2(n3717), .ZN(n3718) );
  ND4D1BWP12T U4060 ( .A1(n3721), .A2(n3720), .A3(n3719), .A4(n3718), .ZN(
        result[23]) );
  INVD1BWP12T U4061 ( .I(n3722), .ZN(n3723) );
  NR2D1BWP12T U4062 ( .A1(a[24]), .A2(n3723), .ZN(n3769) );
  AOI211D1BWP12T U4063 ( .A1(a[24]), .A2(n3723), .B(n3769), .C(n3990), .ZN(
        n3749) );
  OAI32D1BWP12T U4064 ( .A1(a[24]), .A2(n3725), .A3(n3724), .B1(n3995), .B2(
        a[24]), .ZN(n3734) );
  OAI21D1BWP12T U4065 ( .A1(n3899), .A2(n3726), .B(n3996), .ZN(n3731) );
  OAI22D1BWP12T U4066 ( .A1(b[24]), .A2(n3989), .B1(n3938), .B2(n3727), .ZN(
        n3729) );
  OAI21D1BWP12T U4067 ( .A1(n3940), .A2(n3729), .B(n3728), .ZN(n3730) );
  OAI211D1BWP12T U4068 ( .A1(n3922), .A2(n3732), .B(n3731), .C(n3730), .ZN(
        n3733) );
  AOI211D1BWP12T U4069 ( .A1(n4003), .A2(n3735), .B(n3734), .C(n3733), .ZN(
        n3746) );
  INVD1BWP12T U4070 ( .I(n3736), .ZN(n3744) );
  INVD1BWP12T U4071 ( .I(n3737), .ZN(n3812) );
  AOI211D1BWP12T U4072 ( .A1(n3877), .A2(n3738), .B(n3812), .C(n3891), .ZN(
        n3743) );
  AOI22D1BWP12T U4073 ( .A1(n3881), .A2(n3740), .B1(n3739), .B2(n3878), .ZN(
        n3837) );
  AOI22D1BWP12T U4074 ( .A1(n3980), .A2(n3837), .B1(n3889), .B2(n3741), .ZN(
        n3742) );
  OAI211D1BWP12T U4075 ( .A1(n3818), .A2(n3744), .B(n3743), .C(n3742), .ZN(
        n3745) );
  OAI211D1BWP12T U4076 ( .A1(n3920), .A2(n3747), .B(n3746), .C(n3745), .ZN(
        n3748) );
  AOI211D1BWP12T U4077 ( .A1(n3926), .A2(n3750), .B(n3749), .C(n3748), .ZN(
        n3754) );
  AOI22D1BWP12T U4078 ( .A1(n3987), .A2(n3752), .B1(n3906), .B2(n3751), .ZN(
        n3753) );
  OAI211D1BWP12T U4079 ( .A1(n3755), .A2(n3949), .B(n3754), .C(n3753), .ZN(
        result[24]) );
  RCIAO21D0BWP12T U4080 ( .A1(n3899), .A2(n3756), .B(n3831), .ZN(n3774) );
  OAI32D1BWP12T U4081 ( .A1(a[25]), .A2(n4001), .A3(n3757), .B1(n3995), .B2(
        a[25]), .ZN(n3765) );
  AOI22D1BWP12T U4082 ( .A1(a[25]), .A2(n3940), .B1(n3758), .B2(n3840), .ZN(
        n3762) );
  MAOI22D0BWP12T U4083 ( .A1(n4003), .A2(n3760), .B1(n3759), .B2(n3938), .ZN(
        n3761) );
  OAI211D1BWP12T U4084 ( .A1(n3763), .A2(n3920), .B(n3762), .C(n3761), .ZN(
        n3764) );
  AOI211D1BWP12T U4085 ( .A1(n3767), .A2(n3766), .B(n3765), .C(n3764), .ZN(
        n3771) );
  OAI211D1BWP12T U4086 ( .A1(n3769), .A2(n3768), .B(n3945), .C(n3781), .ZN(
        n3770) );
  OAI211D1BWP12T U4087 ( .A1(n3772), .A2(n3976), .B(n3771), .C(n3770), .ZN(
        n3773) );
  AOI211D1BWP12T U4088 ( .A1(n3775), .A2(n3981), .B(n3774), .C(n3773), .ZN(
        n3779) );
  MAOI22D0BWP12T U4089 ( .A1(n3987), .A2(n3777), .B1(n3949), .B2(n3776), .ZN(
        n3778) );
  OAI211D1BWP12T U4090 ( .A1(n3780), .A2(n3975), .B(n3779), .C(n3778), .ZN(
        result[25]) );
  AOI211D1BWP12T U4091 ( .A1(a[26]), .A2(n3781), .B(n3810), .C(n3990), .ZN(
        n3807) );
  AOI21D1BWP12T U4092 ( .A1(n3784), .A2(n3783), .B(n3782), .ZN(n3786) );
  OAI22D1BWP12T U4093 ( .A1(n3786), .A2(n3891), .B1(n3785), .B2(n3920), .ZN(
        n3806) );
  OAI22D1BWP12T U4094 ( .A1(a[26]), .A2(n3995), .B1(n3989), .B2(n3787), .ZN(
        n3796) );
  NR2D1BWP12T U4095 ( .A1(n3788), .A2(n3938), .ZN(n3789) );
  AOI211D1BWP12T U4096 ( .A1(n3823), .A2(n3790), .B(n3789), .C(n3940), .ZN(
        n3793) );
  OAI22D1BWP12T U4097 ( .A1(n3794), .A2(n3793), .B1(n3792), .B2(n3791), .ZN(
        n3795) );
  AOI211D1BWP12T U4098 ( .A1(n4003), .A2(n3797), .B(n3796), .C(n3795), .ZN(
        n3800) );
  OAI21D1BWP12T U4099 ( .A1(n3899), .A2(n3798), .B(n3996), .ZN(n3799) );
  OAI211D1BWP12T U4100 ( .A1(n3801), .A2(n3976), .B(n3800), .C(n3799), .ZN(
        n3805) );
  OAI22D1BWP12T U4101 ( .A1(n3803), .A2(n3956), .B1(n3802), .B2(n3949), .ZN(
        n3804) );
  NR4D0BWP12T U4102 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(
        n3808) );
  OAI21D1BWP12T U4103 ( .A1(n3809), .A2(n3975), .B(n3808), .ZN(result[26]) );
  INVD1BWP12T U4104 ( .I(n3810), .ZN(n3811) );
  NR2D1BWP12T U4105 ( .A1(a[27]), .A2(n3811), .ZN(n3852) );
  OAI22D1BWP12T U4106 ( .A1(n3832), .A2(n3831), .B1(n3830), .B2(n3920), .ZN(
        n3857) );
  ND2D1BWP12T U4107 ( .A1(b[28]), .A2(n3833), .ZN(n3834) );
  AOI32D1BWP12T U4108 ( .A1(n3988), .A2(a[28]), .A3(n3834), .B1(n3995), .B2(
        n3851), .ZN(n3849) );
  OAI22D1BWP12T U4109 ( .A1(n3837), .A2(n3836), .B1(n3884), .B2(n3835), .ZN(
        n3838) );
  AOI21D1BWP12T U4110 ( .A1(n3889), .A2(n3839), .B(n3838), .ZN(n3847) );
  AOI22D1BWP12T U4111 ( .A1(n3842), .A2(n3960), .B1(n3841), .B2(n3840), .ZN(
        n3846) );
  OAI221D1BWP12T U4112 ( .A1(n3881), .A2(n3844), .B1(n3878), .B2(n3843), .C(
        n3980), .ZN(n3845) );
  AOI32D1BWP12T U4113 ( .A1(n3847), .A2(n3846), .A3(n3845), .B1(n3891), .B2(
        n3846), .ZN(n3848) );
  AOI211D1BWP12T U4114 ( .A1(n4003), .A2(n3850), .B(n3849), .C(n3848), .ZN(
        n3854) );
  OAI211D1BWP12T U4115 ( .A1(n3852), .A2(n3851), .B(n3945), .C(n3874), .ZN(
        n3853) );
  OAI211D1BWP12T U4116 ( .A1(n3922), .A2(n3855), .B(n3854), .C(n3853), .ZN(
        n3856) );
  AOI211D1BWP12T U4117 ( .A1(n3926), .A2(n3858), .B(n3857), .C(n3856), .ZN(
        n3862) );
  AOI22D1BWP12T U4118 ( .A1(n3999), .A2(n3860), .B1(n3906), .B2(n3859), .ZN(
        n3861) );
  OAI211D1BWP12T U4119 ( .A1(n3863), .A2(n3956), .B(n3862), .C(n3861), .ZN(
        result[28]) );
  OAI22D1BWP12T U4120 ( .A1(n3989), .A2(n3865), .B1(n4001), .B2(n3864), .ZN(
        n3871) );
  MAOI22D0BWP12T U4121 ( .A1(n4003), .A2(n3867), .B1(n3866), .B2(n3994), .ZN(
        n3868) );
  OAI221D1BWP12T U4122 ( .A1(a[29]), .A2(n3995), .B1(n3869), .B2(n3988), .C(
        n3868), .ZN(n3870) );
  AOI211D1BWP12T U4123 ( .A1(n3873), .A2(n3872), .B(n3871), .C(n3870), .ZN(
        n3903) );
  AOI211D1BWP12T U4124 ( .A1(a[29]), .A2(n3874), .B(n3933), .C(n3990), .ZN(
        n3894) );
  IOA21D1BWP12T U4125 ( .A1(n3877), .A2(n3876), .B(n3875), .ZN(n3887) );
  AOI22D1BWP12T U4126 ( .A1(n3881), .A2(n3880), .B1(n3879), .B2(n3878), .ZN(
        n3882) );
  OAI22D1BWP12T U4127 ( .A1(n3885), .A2(n3884), .B1(n3883), .B2(n3882), .ZN(
        n3886) );
  AOI211D1BWP12T U4128 ( .A1(n3889), .A2(n3888), .B(n3887), .C(n3886), .ZN(
        n3892) );
  OAI22D1BWP12T U4129 ( .A1(n3892), .A2(n3891), .B1(n3920), .B2(n3890), .ZN(
        n3893) );
  AOI211D1BWP12T U4130 ( .A1(n3895), .A2(n3926), .B(n3894), .C(n3893), .ZN(
        n3902) );
  AOI22D1BWP12T U4131 ( .A1(n3999), .A2(n3897), .B1(n3987), .B2(n3896), .ZN(
        n3901) );
  OAI21D1BWP12T U4132 ( .A1(n3899), .A2(n3898), .B(n3996), .ZN(n3900) );
  ND4D1BWP12T U4133 ( .A1(n3903), .A2(n3902), .A3(n3901), .A4(n3900), .ZN(
        n3904) );
  AO21D1BWP12T U4134 ( .A1(n3906), .A2(n3905), .B(n3904), .Z(result[29]) );
  OAI21D1BWP12T U4135 ( .A1(n3909), .A2(n3908), .B(n3907), .ZN(n3910) );
  AOI22D1BWP12T U4136 ( .A1(n3981), .A2(n3911), .B1(n3996), .B2(n3910), .ZN(
        n3937) );
  NR3D1BWP12T U4137 ( .A1(n3912), .A2(a[30]), .A3(n4001), .ZN(n3913) );
  AOI21D1BWP12T U4138 ( .A1(n3914), .A2(n4003), .B(n3913), .ZN(n3917) );
  NR2D1BWP12T U4139 ( .A1(b[30]), .A2(n3989), .ZN(n3915) );
  OAI32D1BWP12T U4140 ( .A1(n3932), .A2(n3940), .A3(n3915), .B1(a[30]), .B2(
        n3959), .ZN(n3916) );
  OAI211D1BWP12T U4141 ( .A1(n3938), .A2(n3918), .B(n3917), .C(n3916), .ZN(
        n3924) );
  OAI22D1BWP12T U4142 ( .A1(n3922), .A2(n3921), .B1(n3920), .B2(n3919), .ZN(
        n3923) );
  AOI211D1BWP12T U4143 ( .A1(n3926), .A2(n3925), .B(n3924), .C(n3923), .ZN(
        n3936) );
  OAI22D1BWP12T U4144 ( .A1(n3928), .A2(n3975), .B1(n3927), .B2(n3949), .ZN(
        n3929) );
  AOI21D1BWP12T U4145 ( .A1(n3987), .A2(n3930), .B(n3929), .ZN(n3935) );
  OAI211D1BWP12T U4146 ( .A1(n3933), .A2(n3932), .B(n3945), .C(n3931), .ZN(
        n3934) );
  ND4D1BWP12T U4147 ( .A1(n3937), .A2(n3936), .A3(n3935), .A4(n3934), .ZN(
        result[30]) );
  MAOI22D0BWP12T U4148 ( .A1(a[2]), .A2(n3940), .B1(n3939), .B2(n3938), .ZN(
        n3947) );
  OAI22D1BWP12T U4149 ( .A1(n3942), .A2(n3976), .B1(n3989), .B2(n3941), .ZN(
        n3943) );
  AOI31D1BWP12T U4150 ( .A1(n3945), .A2(n3992), .A3(n3944), .B(n3943), .ZN(
        n3946) );
  OA211D1BWP12T U4151 ( .A1(n3949), .A2(n3948), .B(n3947), .C(n3946), .Z(n3973) );
  AOI22D1BWP12T U4152 ( .A1(n3951), .A2(n3984), .B1(n3996), .B2(n3950), .ZN(
        n3972) );
  NR2D1BWP12T U4153 ( .A1(n3952), .A2(n3961), .ZN(n3953) );
  MAOI22D0BWP12T U4154 ( .A1(n3954), .A2(n3953), .B1(n3954), .B2(n3953), .ZN(
        n3957) );
  OAI22D1BWP12T U4155 ( .A1(n3958), .A2(n3957), .B1(n3956), .B2(n3955), .ZN(
        n3966) );
  AOI32D1BWP12T U4156 ( .A1(b[2]), .A2(n3961), .A3(n3960), .B1(n3959), .B2(
        n3961), .ZN(n3962) );
  OAI211D1BWP12T U4157 ( .A1(n3964), .A2(n3975), .B(n3963), .C(n3962), .ZN(
        n3965) );
  AOI211D1BWP12T U4158 ( .A1(n3967), .A2(n3982), .B(n3966), .C(n3965), .ZN(
        n3971) );
  AOI32D1BWP12T U4159 ( .A1(n3980), .A2(n3981), .A3(n3969), .B1(n3968), .B2(
        n3981), .ZN(n3970) );
  ND4D1BWP12T U4160 ( .A1(n3973), .A2(n3972), .A3(n3971), .A4(n3970), .ZN(
        result[2]) );
  NR2D1BWP12T U4161 ( .A1(n4006), .A2(n4005), .ZN(n4007) );
  MOAI22D0BWP12T U4162 ( .A1(n4008), .A2(n4007), .B1(n4008), .B2(n4007), .ZN(
        mult_x_18_n454) );
endmodule

