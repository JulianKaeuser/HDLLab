
module register_file_v2 ( readA_sel, readB_sel, readC_sel, readD_sel, 
        write1_sel, write2_sel, write1_en, write2_en, write1_in, write2_in, 
        immediate1_in, immediate2_in, next_pc_in, next_cpsr_in, next_sp_in, 
        clk, reset, regA_out, regB_out, regC_out, regD_out, pc_out, cpsr_out, 
        sp_out, next_pc_en_BAR );
  input [4:0] readA_sel;
  input [4:0] readB_sel;
  input [4:0] readC_sel;
  input [4:0] readD_sel;
  input [4:0] write1_sel;
  input [4:0] write2_sel;
  input [31:0] write1_in;
  input [31:0] write2_in;
  input [31:0] immediate1_in;
  input [31:0] immediate2_in;
  input [31:0] next_pc_in;
  input [3:0] next_cpsr_in;
  input [31:0] next_sp_in;
  output [31:0] regA_out;
  output [31:0] regB_out;
  output [31:0] regC_out;
  output [31:0] regD_out;
  output [31:0] pc_out;
  output [3:0] cpsr_out;
  output [31:0] sp_out;
  input write1_en, write2_en, clk, reset, next_pc_en_BAR;
  wire   n2135, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2326, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2646, n2647, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2136, n2261, n2293, n2325, n2327,
         n2389, n2517, n2549, n2581, n2645, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548;
  wire   [3549:3580] n;
  wire   [31:0] r0;
  wire   [31:0] r1;
  wire   [31:0] r2;
  wire   [31:0] r3;
  wire   [31:0] r4;
  wire   [31:0] r5;
  wire   [31:0] r6;
  wire   [31:0] r7;
  wire   [31:0] r8;
  wire   [31:0] r9;
  wire   [31:0] r10;
  wire   [31:0] r11;
  wire   [31:0] r12;
  wire   [31:0] lr;
  wire   [31:0] tmp1;
  wire   [31:0] spin;
  wire   [3:2] cpsrin;

  DFQD1BWP12T r0_reg_30_ ( .D(n2646), .CP(clk), .Q(r0[30]) );
  DFQD1BWP12T r0_reg_28_ ( .D(n2644), .CP(clk), .Q(r0[28]) );
  DFQD1BWP12T r0_reg_27_ ( .D(n2643), .CP(clk), .Q(r0[27]) );
  DFQD1BWP12T r0_reg_26_ ( .D(n2642), .CP(clk), .Q(r0[26]) );
  DFQD1BWP12T r0_reg_25_ ( .D(n2641), .CP(clk), .Q(r0[25]) );
  DFQD1BWP12T r0_reg_24_ ( .D(n2640), .CP(clk), .Q(r0[24]) );
  DFQD1BWP12T r0_reg_23_ ( .D(n2639), .CP(clk), .Q(r0[23]) );
  DFQD1BWP12T r0_reg_22_ ( .D(n2638), .CP(clk), .Q(r0[22]) );
  DFQD1BWP12T r0_reg_21_ ( .D(n2637), .CP(clk), .Q(r0[21]) );
  DFQD1BWP12T r0_reg_20_ ( .D(n2636), .CP(clk), .Q(r0[20]) );
  DFQD1BWP12T r0_reg_19_ ( .D(n2635), .CP(clk), .Q(r0[19]) );
  DFQD1BWP12T r0_reg_18_ ( .D(n2634), .CP(clk), .Q(r0[18]) );
  DFQD1BWP12T r0_reg_17_ ( .D(n2633), .CP(clk), .Q(r0[17]) );
  DFQD1BWP12T r0_reg_16_ ( .D(n2632), .CP(clk), .Q(r0[16]) );
  DFQD1BWP12T r0_reg_15_ ( .D(n2631), .CP(clk), .Q(r0[15]) );
  DFQD1BWP12T r0_reg_14_ ( .D(n2630), .CP(clk), .Q(r0[14]) );
  DFQD1BWP12T r0_reg_13_ ( .D(n2629), .CP(clk), .Q(r0[13]) );
  DFQD1BWP12T r0_reg_11_ ( .D(n2627), .CP(clk), .Q(r0[11]) );
  DFQD1BWP12T r0_reg_10_ ( .D(n2626), .CP(clk), .Q(r0[10]) );
  DFQD1BWP12T r0_reg_9_ ( .D(n2625), .CP(clk), .Q(r0[9]) );
  DFQD1BWP12T r0_reg_8_ ( .D(n2624), .CP(clk), .Q(r0[8]) );
  DFQD1BWP12T r0_reg_6_ ( .D(n2622), .CP(clk), .Q(r0[6]) );
  DFQD1BWP12T r0_reg_5_ ( .D(n2621), .CP(clk), .Q(r0[5]) );
  DFQD1BWP12T r0_reg_4_ ( .D(n2620), .CP(clk), .Q(r0[4]) );
  DFQD1BWP12T r0_reg_3_ ( .D(n2619), .CP(clk), .Q(r0[3]) );
  DFQD1BWP12T r0_reg_2_ ( .D(n2618), .CP(clk), .Q(r0[2]) );
  DFQD1BWP12T r0_reg_0_ ( .D(n2616), .CP(clk), .Q(r0[0]) );
  DFQD1BWP12T r1_reg_30_ ( .D(n2614), .CP(clk), .Q(r1[30]) );
  DFQD1BWP12T r1_reg_29_ ( .D(n2613), .CP(clk), .Q(r1[29]) );
  DFQD1BWP12T r1_reg_28_ ( .D(n2612), .CP(clk), .Q(r1[28]) );
  DFQD1BWP12T r1_reg_27_ ( .D(n2611), .CP(clk), .Q(r1[27]) );
  DFQD1BWP12T r1_reg_26_ ( .D(n2610), .CP(clk), .Q(r1[26]) );
  DFQD1BWP12T r1_reg_25_ ( .D(n2609), .CP(clk), .Q(r1[25]) );
  DFQD1BWP12T r1_reg_24_ ( .D(n2608), .CP(clk), .Q(r1[24]) );
  DFQD1BWP12T r1_reg_23_ ( .D(n2607), .CP(clk), .Q(r1[23]) );
  DFQD1BWP12T r1_reg_22_ ( .D(n2606), .CP(clk), .Q(r1[22]) );
  DFQD1BWP12T r1_reg_21_ ( .D(n2605), .CP(clk), .Q(r1[21]) );
  DFQD1BWP12T r1_reg_20_ ( .D(n2604), .CP(clk), .Q(r1[20]) );
  DFQD1BWP12T r1_reg_19_ ( .D(n2603), .CP(clk), .Q(r1[19]) );
  DFQD1BWP12T r1_reg_17_ ( .D(n2601), .CP(clk), .Q(r1[17]) );
  DFQD1BWP12T r1_reg_16_ ( .D(n2600), .CP(clk), .Q(r1[16]) );
  DFQD1BWP12T r1_reg_15_ ( .D(n2599), .CP(clk), .Q(r1[15]) );
  DFQD1BWP12T r1_reg_14_ ( .D(n2598), .CP(clk), .Q(r1[14]) );
  DFQD1BWP12T r1_reg_13_ ( .D(n2597), .CP(clk), .Q(r1[13]) );
  DFQD1BWP12T r1_reg_12_ ( .D(n2596), .CP(clk), .Q(r1[12]) );
  DFQD1BWP12T r1_reg_11_ ( .D(n2595), .CP(clk), .Q(r1[11]) );
  DFQD1BWP12T r1_reg_10_ ( .D(n2594), .CP(clk), .Q(r1[10]) );
  DFQD1BWP12T r1_reg_9_ ( .D(n2593), .CP(clk), .Q(r1[9]) );
  DFQD1BWP12T r1_reg_8_ ( .D(n2592), .CP(clk), .Q(r1[8]) );
  DFQD1BWP12T r1_reg_7_ ( .D(n2591), .CP(clk), .Q(r1[7]) );
  DFQD1BWP12T r1_reg_6_ ( .D(n2590), .CP(clk), .Q(r1[6]) );
  DFQD1BWP12T r1_reg_5_ ( .D(n2589), .CP(clk), .Q(r1[5]) );
  DFQD1BWP12T r1_reg_4_ ( .D(n2588), .CP(clk), .Q(r1[4]) );
  DFQD1BWP12T r1_reg_3_ ( .D(n2587), .CP(clk), .Q(r1[3]) );
  DFQD1BWP12T r1_reg_2_ ( .D(n2586), .CP(clk), .Q(r1[2]) );
  DFQD1BWP12T r1_reg_1_ ( .D(n2585), .CP(clk), .Q(r1[1]) );
  DFQD1BWP12T r1_reg_0_ ( .D(n2584), .CP(clk), .Q(r1[0]) );
  DFQD1BWP12T r2_reg_31_ ( .D(n2583), .CP(clk), .Q(r2[31]) );
  DFQD1BWP12T r2_reg_30_ ( .D(n2582), .CP(clk), .Q(r2[30]) );
  DFQD1BWP12T r2_reg_28_ ( .D(n2580), .CP(clk), .Q(r2[28]) );
  DFQD1BWP12T r2_reg_27_ ( .D(n2579), .CP(clk), .Q(r2[27]) );
  DFQD1BWP12T r2_reg_26_ ( .D(n2578), .CP(clk), .Q(r2[26]) );
  DFQD1BWP12T r2_reg_25_ ( .D(n2577), .CP(clk), .Q(r2[25]) );
  DFQD1BWP12T r2_reg_24_ ( .D(n2576), .CP(clk), .Q(r2[24]) );
  DFQD1BWP12T r2_reg_23_ ( .D(n2575), .CP(clk), .Q(r2[23]) );
  DFQD1BWP12T r2_reg_22_ ( .D(n2574), .CP(clk), .Q(r2[22]) );
  DFQD1BWP12T r2_reg_21_ ( .D(n2573), .CP(clk), .Q(r2[21]) );
  DFQD1BWP12T r2_reg_20_ ( .D(n2572), .CP(clk), .Q(r2[20]) );
  DFQD1BWP12T r2_reg_19_ ( .D(n2571), .CP(clk), .Q(r2[19]) );
  DFQD1BWP12T r2_reg_18_ ( .D(n2570), .CP(clk), .Q(r2[18]) );
  DFQD1BWP12T r2_reg_17_ ( .D(n2569), .CP(clk), .Q(r2[17]) );
  DFQD1BWP12T r2_reg_16_ ( .D(n2568), .CP(clk), .Q(r2[16]) );
  DFQD1BWP12T r2_reg_15_ ( .D(n2567), .CP(clk), .Q(r2[15]) );
  DFQD1BWP12T r2_reg_14_ ( .D(n2566), .CP(clk), .Q(r2[14]) );
  DFQD1BWP12T r2_reg_13_ ( .D(n2565), .CP(clk), .Q(r2[13]) );
  DFQD1BWP12T r2_reg_12_ ( .D(n2564), .CP(clk), .Q(r2[12]) );
  DFQD1BWP12T r2_reg_11_ ( .D(n2563), .CP(clk), .Q(r2[11]) );
  DFQD1BWP12T r2_reg_10_ ( .D(n2562), .CP(clk), .Q(r2[10]) );
  DFQD1BWP12T r2_reg_9_ ( .D(n2561), .CP(clk), .Q(r2[9]) );
  DFQD1BWP12T r2_reg_8_ ( .D(n2560), .CP(clk), .Q(r2[8]) );
  DFQD1BWP12T r2_reg_7_ ( .D(n2559), .CP(clk), .Q(r2[7]) );
  DFQD1BWP12T r2_reg_6_ ( .D(n2558), .CP(clk), .Q(r2[6]) );
  DFQD1BWP12T r2_reg_5_ ( .D(n2557), .CP(clk), .Q(r2[5]) );
  DFQD1BWP12T r2_reg_4_ ( .D(n2556), .CP(clk), .Q(r2[4]) );
  DFQD1BWP12T r2_reg_3_ ( .D(n2555), .CP(clk), .Q(r2[3]) );
  DFQD1BWP12T r2_reg_2_ ( .D(n2554), .CP(clk), .Q(r2[2]) );
  DFQD1BWP12T r2_reg_1_ ( .D(n2553), .CP(clk), .Q(r2[1]) );
  DFQD1BWP12T r2_reg_0_ ( .D(n2552), .CP(clk), .Q(r2[0]) );
  DFQD1BWP12T r3_reg_31_ ( .D(n2551), .CP(clk), .Q(r3[31]) );
  DFQD1BWP12T r3_reg_30_ ( .D(n2550), .CP(clk), .Q(r3[30]) );
  DFQD1BWP12T r3_reg_28_ ( .D(n2548), .CP(clk), .Q(r3[28]) );
  DFQD1BWP12T r3_reg_27_ ( .D(n2547), .CP(clk), .Q(r3[27]) );
  DFQD1BWP12T r3_reg_26_ ( .D(n2546), .CP(clk), .Q(r3[26]) );
  DFQD1BWP12T r3_reg_25_ ( .D(n2545), .CP(clk), .Q(r3[25]) );
  DFQD1BWP12T r3_reg_24_ ( .D(n2544), .CP(clk), .Q(r3[24]) );
  DFQD1BWP12T r3_reg_23_ ( .D(n2543), .CP(clk), .Q(r3[23]) );
  DFQD1BWP12T r3_reg_22_ ( .D(n2542), .CP(clk), .Q(r3[22]) );
  DFQD1BWP12T r3_reg_21_ ( .D(n2541), .CP(clk), .Q(r3[21]) );
  DFQD1BWP12T r3_reg_20_ ( .D(n2540), .CP(clk), .Q(r3[20]) );
  DFQD1BWP12T r3_reg_19_ ( .D(n2539), .CP(clk), .Q(r3[19]) );
  DFQD1BWP12T r3_reg_18_ ( .D(n2538), .CP(clk), .Q(r3[18]) );
  DFQD1BWP12T r3_reg_17_ ( .D(n2537), .CP(clk), .Q(r3[17]) );
  DFQD1BWP12T r3_reg_16_ ( .D(n2536), .CP(clk), .Q(r3[16]) );
  DFQD1BWP12T r3_reg_15_ ( .D(n2535), .CP(clk), .Q(r3[15]) );
  DFQD1BWP12T r3_reg_14_ ( .D(n2534), .CP(clk), .Q(r3[14]) );
  DFQD1BWP12T r3_reg_13_ ( .D(n2533), .CP(clk), .Q(r3[13]) );
  DFQD1BWP12T r3_reg_12_ ( .D(n2532), .CP(clk), .Q(r3[12]) );
  DFQD1BWP12T r3_reg_11_ ( .D(n2531), .CP(clk), .Q(r3[11]) );
  DFQD1BWP12T r3_reg_10_ ( .D(n2530), .CP(clk), .Q(r3[10]) );
  DFQD1BWP12T r3_reg_9_ ( .D(n2529), .CP(clk), .Q(r3[9]) );
  DFQD1BWP12T r3_reg_8_ ( .D(n2528), .CP(clk), .Q(r3[8]) );
  DFQD1BWP12T r3_reg_7_ ( .D(n2527), .CP(clk), .Q(r3[7]) );
  DFQD1BWP12T r3_reg_6_ ( .D(n2526), .CP(clk), .Q(r3[6]) );
  DFQD1BWP12T r3_reg_5_ ( .D(n2525), .CP(clk), .Q(r3[5]) );
  DFQD1BWP12T r3_reg_4_ ( .D(n2524), .CP(clk), .Q(r3[4]) );
  DFQD1BWP12T r3_reg_3_ ( .D(n2523), .CP(clk), .Q(r3[3]) );
  DFQD1BWP12T r3_reg_2_ ( .D(n2522), .CP(clk), .Q(r3[2]) );
  DFQD1BWP12T r3_reg_1_ ( .D(n2521), .CP(clk), .Q(r3[1]) );
  DFQD1BWP12T r3_reg_0_ ( .D(n2520), .CP(clk), .Q(r3[0]) );
  DFQD1BWP12T r4_reg_30_ ( .D(n2518), .CP(clk), .Q(r4[30]) );
  DFQD1BWP12T r4_reg_28_ ( .D(n2516), .CP(clk), .Q(r4[28]) );
  DFQD1BWP12T r4_reg_27_ ( .D(n2515), .CP(clk), .Q(r4[27]) );
  DFQD1BWP12T r4_reg_26_ ( .D(n2514), .CP(clk), .Q(r4[26]) );
  DFQD1BWP12T r4_reg_25_ ( .D(n2513), .CP(clk), .Q(r4[25]) );
  DFQD1BWP12T r4_reg_24_ ( .D(n2512), .CP(clk), .Q(r4[24]) );
  DFQD1BWP12T r4_reg_23_ ( .D(n2511), .CP(clk), .Q(r4[23]) );
  DFQD1BWP12T r4_reg_22_ ( .D(n2510), .CP(clk), .Q(r4[22]) );
  DFQD1BWP12T r4_reg_21_ ( .D(n2509), .CP(clk), .Q(r4[21]) );
  DFQD1BWP12T r4_reg_20_ ( .D(n2508), .CP(clk), .Q(r4[20]) );
  DFQD1BWP12T r4_reg_19_ ( .D(n2507), .CP(clk), .Q(r4[19]) );
  DFQD1BWP12T r4_reg_18_ ( .D(n2506), .CP(clk), .Q(r4[18]) );
  DFQD1BWP12T r4_reg_17_ ( .D(n2505), .CP(clk), .Q(r4[17]) );
  DFQD1BWP12T r4_reg_16_ ( .D(n2504), .CP(clk), .Q(r4[16]) );
  DFQD1BWP12T r4_reg_15_ ( .D(n2503), .CP(clk), .Q(r4[15]) );
  DFQD1BWP12T r4_reg_14_ ( .D(n2502), .CP(clk), .Q(r4[14]) );
  DFQD1BWP12T r4_reg_13_ ( .D(n2501), .CP(clk), .Q(r4[13]) );
  DFQD1BWP12T r4_reg_12_ ( .D(n2500), .CP(clk), .Q(r4[12]) );
  DFQD1BWP12T r4_reg_11_ ( .D(n2499), .CP(clk), .Q(r4[11]) );
  DFQD1BWP12T r4_reg_10_ ( .D(n2498), .CP(clk), .Q(r4[10]) );
  DFQD1BWP12T r4_reg_9_ ( .D(n2497), .CP(clk), .Q(r4[9]) );
  DFQD1BWP12T r4_reg_8_ ( .D(n2496), .CP(clk), .Q(r4[8]) );
  DFQD1BWP12T r4_reg_6_ ( .D(n2494), .CP(clk), .Q(r4[6]) );
  DFQD1BWP12T r4_reg_5_ ( .D(n2493), .CP(clk), .Q(r4[5]) );
  DFQD1BWP12T r4_reg_4_ ( .D(n2492), .CP(clk), .Q(r4[4]) );
  DFQD1BWP12T r4_reg_3_ ( .D(n2491), .CP(clk), .Q(r4[3]) );
  DFQD1BWP12T r4_reg_2_ ( .D(n2490), .CP(clk), .Q(r4[2]) );
  DFQD1BWP12T r4_reg_1_ ( .D(n2489), .CP(clk), .Q(r4[1]) );
  DFQD1BWP12T r4_reg_0_ ( .D(n2488), .CP(clk), .Q(r4[0]) );
  DFQD1BWP12T r5_reg_31_ ( .D(n2487), .CP(clk), .Q(r5[31]) );
  DFQD1BWP12T r5_reg_30_ ( .D(n2486), .CP(clk), .Q(r5[30]) );
  DFQD1BWP12T r5_reg_29_ ( .D(n2485), .CP(clk), .Q(r5[29]) );
  DFQD1BWP12T r5_reg_28_ ( .D(n2484), .CP(clk), .Q(r5[28]) );
  DFQD1BWP12T r5_reg_27_ ( .D(n2483), .CP(clk), .Q(r5[27]) );
  DFQD1BWP12T r5_reg_26_ ( .D(n2482), .CP(clk), .Q(r5[26]) );
  DFQD1BWP12T r5_reg_25_ ( .D(n2481), .CP(clk), .Q(r5[25]) );
  DFQD1BWP12T r5_reg_24_ ( .D(n2480), .CP(clk), .Q(r5[24]) );
  DFQD1BWP12T r5_reg_23_ ( .D(n2479), .CP(clk), .Q(r5[23]) );
  DFQD1BWP12T r5_reg_22_ ( .D(n2478), .CP(clk), .Q(r5[22]) );
  DFQD1BWP12T r5_reg_20_ ( .D(n2476), .CP(clk), .Q(r5[20]) );
  DFQD1BWP12T r5_reg_19_ ( .D(n2475), .CP(clk), .Q(r5[19]) );
  DFQD1BWP12T r5_reg_18_ ( .D(n2474), .CP(clk), .Q(r5[18]) );
  DFQD1BWP12T r5_reg_17_ ( .D(n2473), .CP(clk), .Q(r5[17]) );
  DFQD1BWP12T r5_reg_16_ ( .D(n2472), .CP(clk), .Q(r5[16]) );
  DFQD1BWP12T r5_reg_14_ ( .D(n2470), .CP(clk), .Q(r5[14]) );
  DFQD1BWP12T r5_reg_13_ ( .D(n2469), .CP(clk), .Q(r5[13]) );
  DFQD1BWP12T r5_reg_12_ ( .D(n2468), .CP(clk), .Q(r5[12]) );
  DFQD1BWP12T r5_reg_11_ ( .D(n2467), .CP(clk), .Q(r5[11]) );
  DFQD1BWP12T r5_reg_10_ ( .D(n2466), .CP(clk), .Q(r5[10]) );
  DFQD1BWP12T r5_reg_9_ ( .D(n2465), .CP(clk), .Q(r5[9]) );
  DFQD1BWP12T r5_reg_8_ ( .D(n2464), .CP(clk), .Q(r5[8]) );
  DFQD1BWP12T r5_reg_7_ ( .D(n2463), .CP(clk), .Q(r5[7]) );
  DFQD1BWP12T r5_reg_6_ ( .D(n2462), .CP(clk), .Q(r5[6]) );
  DFQD1BWP12T r5_reg_5_ ( .D(n2461), .CP(clk), .Q(r5[5]) );
  DFQD1BWP12T r5_reg_4_ ( .D(n2460), .CP(clk), .Q(r5[4]) );
  DFQD1BWP12T r5_reg_3_ ( .D(n2459), .CP(clk), .Q(r5[3]) );
  DFQD1BWP12T r5_reg_1_ ( .D(n2457), .CP(clk), .Q(r5[1]) );
  DFQD1BWP12T r5_reg_0_ ( .D(n2456), .CP(clk), .Q(r5[0]) );
  DFQD1BWP12T r6_reg_31_ ( .D(n2455), .CP(clk), .Q(r6[31]) );
  DFQD1BWP12T r6_reg_30_ ( .D(n2454), .CP(clk), .Q(r6[30]) );
  DFQD1BWP12T r6_reg_29_ ( .D(n2453), .CP(clk), .Q(r6[29]) );
  DFQD1BWP12T r6_reg_28_ ( .D(n2452), .CP(clk), .Q(r6[28]) );
  DFQD1BWP12T r6_reg_27_ ( .D(n2451), .CP(clk), .Q(r6[27]) );
  DFQD1BWP12T r6_reg_25_ ( .D(n2449), .CP(clk), .Q(r6[25]) );
  DFQD1BWP12T r6_reg_24_ ( .D(n2448), .CP(clk), .Q(r6[24]) );
  DFQD1BWP12T r6_reg_23_ ( .D(n2447), .CP(clk), .Q(r6[23]) );
  DFQD1BWP12T r6_reg_22_ ( .D(n2446), .CP(clk), .Q(r6[22]) );
  DFQD1BWP12T r6_reg_21_ ( .D(n2445), .CP(clk), .Q(r6[21]) );
  DFQD1BWP12T r6_reg_20_ ( .D(n2444), .CP(clk), .Q(r6[20]) );
  DFQD1BWP12T r6_reg_19_ ( .D(n2443), .CP(clk), .Q(r6[19]) );
  DFQD1BWP12T r6_reg_18_ ( .D(n2442), .CP(clk), .Q(r6[18]) );
  DFQD1BWP12T r6_reg_17_ ( .D(n2441), .CP(clk), .Q(r6[17]) );
  DFQD1BWP12T r6_reg_16_ ( .D(n2440), .CP(clk), .Q(r6[16]) );
  DFQD1BWP12T r6_reg_15_ ( .D(n2439), .CP(clk), .Q(r6[15]) );
  DFQD1BWP12T r6_reg_14_ ( .D(n2438), .CP(clk), .Q(r6[14]) );
  DFQD1BWP12T r6_reg_13_ ( .D(n2437), .CP(clk), .Q(r6[13]) );
  DFQD1BWP12T r6_reg_12_ ( .D(n2436), .CP(clk), .Q(r6[12]) );
  DFQD1BWP12T r6_reg_11_ ( .D(n2435), .CP(clk), .Q(r6[11]) );
  DFQD1BWP12T r6_reg_10_ ( .D(n2434), .CP(clk), .Q(r6[10]) );
  DFQD1BWP12T r6_reg_9_ ( .D(n2433), .CP(clk), .Q(r6[9]) );
  DFQD1BWP12T r6_reg_8_ ( .D(n2432), .CP(clk), .Q(r6[8]) );
  DFQD1BWP12T r6_reg_6_ ( .D(n2430), .CP(clk), .Q(r6[6]) );
  DFQD1BWP12T r6_reg_4_ ( .D(n2428), .CP(clk), .Q(r6[4]) );
  DFQD1BWP12T r6_reg_3_ ( .D(n2427), .CP(clk), .Q(r6[3]) );
  DFQD1BWP12T r6_reg_2_ ( .D(n2426), .CP(clk), .Q(r6[2]) );
  DFQD1BWP12T r6_reg_1_ ( .D(n2425), .CP(clk), .Q(r6[1]) );
  DFQD1BWP12T r6_reg_0_ ( .D(n2424), .CP(clk), .Q(r6[0]) );
  DFQD1BWP12T r7_reg_31_ ( .D(n2423), .CP(clk), .Q(r7[31]) );
  DFQD1BWP12T r7_reg_30_ ( .D(n2422), .CP(clk), .Q(r7[30]) );
  DFQD1BWP12T r7_reg_29_ ( .D(n2421), .CP(clk), .Q(r7[29]) );
  DFQD1BWP12T r7_reg_28_ ( .D(n2420), .CP(clk), .Q(r7[28]) );
  DFQD1BWP12T r7_reg_27_ ( .D(n2419), .CP(clk), .Q(r7[27]) );
  DFQD1BWP12T r7_reg_26_ ( .D(n2418), .CP(clk), .Q(r7[26]) );
  DFQD1BWP12T r7_reg_25_ ( .D(n2417), .CP(clk), .Q(r7[25]) );
  DFQD1BWP12T r7_reg_24_ ( .D(n2416), .CP(clk), .Q(r7[24]) );
  DFQD1BWP12T r7_reg_23_ ( .D(n2415), .CP(clk), .Q(r7[23]) );
  DFQD1BWP12T r7_reg_22_ ( .D(n2414), .CP(clk), .Q(r7[22]) );
  DFQD1BWP12T r7_reg_21_ ( .D(n2413), .CP(clk), .Q(r7[21]) );
  DFQD1BWP12T r7_reg_20_ ( .D(n2412), .CP(clk), .Q(r7[20]) );
  DFQD1BWP12T r7_reg_19_ ( .D(n2411), .CP(clk), .Q(r7[19]) );
  DFQD1BWP12T r7_reg_18_ ( .D(n2410), .CP(clk), .Q(r7[18]) );
  DFQD1BWP12T r7_reg_16_ ( .D(n2408), .CP(clk), .Q(r7[16]) );
  DFQD1BWP12T r7_reg_15_ ( .D(n2407), .CP(clk), .Q(r7[15]) );
  DFQD1BWP12T r7_reg_14_ ( .D(n2406), .CP(clk), .Q(r7[14]) );
  DFQD1BWP12T r7_reg_13_ ( .D(n2405), .CP(clk), .Q(r7[13]) );
  DFQD1BWP12T r7_reg_12_ ( .D(n2404), .CP(clk), .Q(r7[12]) );
  DFQD1BWP12T r7_reg_11_ ( .D(n2403), .CP(clk), .Q(r7[11]) );
  DFQD1BWP12T r7_reg_10_ ( .D(n2402), .CP(clk), .Q(r7[10]) );
  DFQD1BWP12T r7_reg_9_ ( .D(n2401), .CP(clk), .Q(r7[9]) );
  DFQD1BWP12T r7_reg_8_ ( .D(n2400), .CP(clk), .Q(r7[8]) );
  DFQD1BWP12T r7_reg_7_ ( .D(n2399), .CP(clk), .Q(r7[7]) );
  DFQD1BWP12T r7_reg_6_ ( .D(n2398), .CP(clk), .Q(r7[6]) );
  DFQD1BWP12T r7_reg_5_ ( .D(n2397), .CP(clk), .Q(r7[5]) );
  DFQD1BWP12T r7_reg_4_ ( .D(n2396), .CP(clk), .Q(r7[4]) );
  DFQD1BWP12T r7_reg_3_ ( .D(n2395), .CP(clk), .Q(r7[3]) );
  DFQD1BWP12T r7_reg_2_ ( .D(n2394), .CP(clk), .Q(r7[2]) );
  DFQD1BWP12T r7_reg_1_ ( .D(n2393), .CP(clk), .Q(r7[1]) );
  DFQD1BWP12T r7_reg_0_ ( .D(n2392), .CP(clk), .Q(r7[0]) );
  DFQD1BWP12T r8_reg_30_ ( .D(n2390), .CP(clk), .Q(r8[30]) );
  DFQD1BWP12T r8_reg_28_ ( .D(n2388), .CP(clk), .Q(r8[28]) );
  DFQD1BWP12T r8_reg_27_ ( .D(n2387), .CP(clk), .Q(r8[27]) );
  DFQD1BWP12T r8_reg_26_ ( .D(n2386), .CP(clk), .Q(r8[26]) );
  DFQD1BWP12T r8_reg_25_ ( .D(n2385), .CP(clk), .Q(r8[25]) );
  DFQD1BWP12T r8_reg_24_ ( .D(n2384), .CP(clk), .Q(r8[24]) );
  DFQD1BWP12T r8_reg_23_ ( .D(n2383), .CP(clk), .Q(r8[23]) );
  DFQD1BWP12T r8_reg_22_ ( .D(n2382), .CP(clk), .Q(r8[22]) );
  DFQD1BWP12T r8_reg_21_ ( .D(n2381), .CP(clk), .Q(r8[21]) );
  DFQD1BWP12T r8_reg_20_ ( .D(n2380), .CP(clk), .Q(r8[20]) );
  DFQD1BWP12T r8_reg_19_ ( .D(n2379), .CP(clk), .Q(r8[19]) );
  DFQD1BWP12T r8_reg_18_ ( .D(n2378), .CP(clk), .Q(r8[18]) );
  DFQD1BWP12T r8_reg_17_ ( .D(n2377), .CP(clk), .Q(r8[17]) );
  DFQD1BWP12T r8_reg_16_ ( .D(n2376), .CP(clk), .Q(r8[16]) );
  DFQD1BWP12T r8_reg_15_ ( .D(n2375), .CP(clk), .Q(r8[15]) );
  DFQD1BWP12T r8_reg_14_ ( .D(n2374), .CP(clk), .Q(r8[14]) );
  DFQD1BWP12T r8_reg_13_ ( .D(n2373), .CP(clk), .Q(r8[13]) );
  DFQD1BWP12T r8_reg_12_ ( .D(n2372), .CP(clk), .Q(r8[12]) );
  DFQD1BWP12T r8_reg_11_ ( .D(n2371), .CP(clk), .Q(r8[11]) );
  DFQD1BWP12T r8_reg_10_ ( .D(n2370), .CP(clk), .Q(r8[10]) );
  DFQD1BWP12T r8_reg_9_ ( .D(n2369), .CP(clk), .Q(r8[9]) );
  DFQD1BWP12T r8_reg_8_ ( .D(n2368), .CP(clk), .Q(r8[8]) );
  DFQD1BWP12T r8_reg_7_ ( .D(n2367), .CP(clk), .Q(r8[7]) );
  DFQD1BWP12T r8_reg_6_ ( .D(n2366), .CP(clk), .Q(r8[6]) );
  DFQD1BWP12T r8_reg_5_ ( .D(n2365), .CP(clk), .Q(r8[5]) );
  DFQD1BWP12T r8_reg_4_ ( .D(n2364), .CP(clk), .Q(r8[4]) );
  DFQD1BWP12T r8_reg_3_ ( .D(n2363), .CP(clk), .Q(r8[3]) );
  DFQD1BWP12T r8_reg_2_ ( .D(n2362), .CP(clk), .Q(r8[2]) );
  DFQD1BWP12T r8_reg_1_ ( .D(n2361), .CP(clk), .Q(r8[1]) );
  DFQD1BWP12T r8_reg_0_ ( .D(n2360), .CP(clk), .Q(r8[0]) );
  DFQD1BWP12T r9_reg_31_ ( .D(n2359), .CP(clk), .Q(r9[31]) );
  DFQD1BWP12T r9_reg_30_ ( .D(n2358), .CP(clk), .Q(r9[30]) );
  DFQD1BWP12T r9_reg_29_ ( .D(n2357), .CP(clk), .Q(r9[29]) );
  DFQD1BWP12T r9_reg_28_ ( .D(n2356), .CP(clk), .Q(r9[28]) );
  DFQD1BWP12T r9_reg_27_ ( .D(n2355), .CP(clk), .Q(r9[27]) );
  DFQD1BWP12T r9_reg_26_ ( .D(n2354), .CP(clk), .Q(r9[26]) );
  DFQD1BWP12T r9_reg_25_ ( .D(n2353), .CP(clk), .Q(r9[25]) );
  DFQD1BWP12T r9_reg_24_ ( .D(n2352), .CP(clk), .Q(r9[24]) );
  DFQD1BWP12T r9_reg_23_ ( .D(n2351), .CP(clk), .Q(r9[23]) );
  DFQD1BWP12T r9_reg_22_ ( .D(n2350), .CP(clk), .Q(r9[22]) );
  DFQD1BWP12T r9_reg_21_ ( .D(n2349), .CP(clk), .Q(r9[21]) );
  DFQD1BWP12T r9_reg_20_ ( .D(n2348), .CP(clk), .Q(r9[20]) );
  DFQD1BWP12T r9_reg_19_ ( .D(n2347), .CP(clk), .Q(r9[19]) );
  DFQD1BWP12T r9_reg_18_ ( .D(n2346), .CP(clk), .Q(r9[18]) );
  DFQD1BWP12T r9_reg_17_ ( .D(n2345), .CP(clk), .Q(r9[17]) );
  DFQD1BWP12T r9_reg_16_ ( .D(n2344), .CP(clk), .Q(r9[16]) );
  DFQD1BWP12T r9_reg_15_ ( .D(n2343), .CP(clk), .Q(r9[15]) );
  DFQD1BWP12T r9_reg_14_ ( .D(n2342), .CP(clk), .Q(r9[14]) );
  DFQD1BWP12T r9_reg_13_ ( .D(n2341), .CP(clk), .Q(r9[13]) );
  DFQD1BWP12T r9_reg_12_ ( .D(n2340), .CP(clk), .Q(r9[12]) );
  DFQD1BWP12T r9_reg_11_ ( .D(n2339), .CP(clk), .Q(r9[11]) );
  DFQD1BWP12T r9_reg_10_ ( .D(n2338), .CP(clk), .Q(r9[10]) );
  DFQD1BWP12T r9_reg_9_ ( .D(n2337), .CP(clk), .Q(r9[9]) );
  DFQD1BWP12T r9_reg_8_ ( .D(n2336), .CP(clk), .Q(r9[8]) );
  DFQD1BWP12T r9_reg_6_ ( .D(n2334), .CP(clk), .Q(r9[6]) );
  DFQD1BWP12T r9_reg_5_ ( .D(n2333), .CP(clk), .Q(r9[5]) );
  DFQD1BWP12T r9_reg_4_ ( .D(n2332), .CP(clk), .Q(r9[4]) );
  DFQD1BWP12T r9_reg_3_ ( .D(n2331), .CP(clk), .Q(r9[3]) );
  DFQD1BWP12T r9_reg_2_ ( .D(n2330), .CP(clk), .Q(r9[2]) );
  DFQD1BWP12T r9_reg_1_ ( .D(n2329), .CP(clk), .Q(r9[1]) );
  DFQD1BWP12T r9_reg_0_ ( .D(n2328), .CP(clk), .Q(r9[0]) );
  DFQD1BWP12T r10_reg_30_ ( .D(n2326), .CP(clk), .Q(r10[30]) );
  DFQD1BWP12T r10_reg_28_ ( .D(n2324), .CP(clk), .Q(r10[28]) );
  DFQD1BWP12T r10_reg_27_ ( .D(n2323), .CP(clk), .Q(r10[27]) );
  DFQD1BWP12T r10_reg_26_ ( .D(n2322), .CP(clk), .Q(r10[26]) );
  DFQD1BWP12T r10_reg_25_ ( .D(n2321), .CP(clk), .Q(r10[25]) );
  DFQD1BWP12T r10_reg_24_ ( .D(n2320), .CP(clk), .Q(r10[24]) );
  DFQD1BWP12T r10_reg_23_ ( .D(n2319), .CP(clk), .Q(r10[23]) );
  DFQD1BWP12T r10_reg_22_ ( .D(n2318), .CP(clk), .Q(r10[22]) );
  DFQD1BWP12T r10_reg_21_ ( .D(n2317), .CP(clk), .Q(r10[21]) );
  DFQD1BWP12T r10_reg_20_ ( .D(n2316), .CP(clk), .Q(r10[20]) );
  DFQD1BWP12T r10_reg_19_ ( .D(n2315), .CP(clk), .Q(r10[19]) );
  DFQD1BWP12T r10_reg_18_ ( .D(n2314), .CP(clk), .Q(r10[18]) );
  DFQD1BWP12T r10_reg_16_ ( .D(n2312), .CP(clk), .Q(r10[16]) );
  DFQD1BWP12T r10_reg_15_ ( .D(n2311), .CP(clk), .Q(r10[15]) );
  DFQD1BWP12T r10_reg_14_ ( .D(n2310), .CP(clk), .Q(r10[14]) );
  DFQD1BWP12T r10_reg_12_ ( .D(n2308), .CP(clk), .Q(r10[12]) );
  DFQD1BWP12T r10_reg_11_ ( .D(n2307), .CP(clk), .Q(r10[11]) );
  DFQD1BWP12T r10_reg_10_ ( .D(n2306), .CP(clk), .Q(r10[10]) );
  DFQD1BWP12T r10_reg_9_ ( .D(n2305), .CP(clk), .Q(r10[9]) );
  DFQD1BWP12T r10_reg_8_ ( .D(n2304), .CP(clk), .Q(r10[8]) );
  DFQD1BWP12T r10_reg_7_ ( .D(n2303), .CP(clk), .Q(r10[7]) );
  DFQD1BWP12T r10_reg_6_ ( .D(n2302), .CP(clk), .Q(r10[6]) );
  DFQD1BWP12T r10_reg_5_ ( .D(n2301), .CP(clk), .Q(r10[5]) );
  DFQD1BWP12T r10_reg_4_ ( .D(n2300), .CP(clk), .Q(r10[4]) );
  DFQD1BWP12T r10_reg_3_ ( .D(n2299), .CP(clk), .Q(r10[3]) );
  DFQD1BWP12T r10_reg_2_ ( .D(n2298), .CP(clk), .Q(r10[2]) );
  DFQD1BWP12T r10_reg_1_ ( .D(n2297), .CP(clk), .Q(r10[1]) );
  DFQD1BWP12T r10_reg_0_ ( .D(n2296), .CP(clk), .Q(r10[0]) );
  DFQD1BWP12T r11_reg_30_ ( .D(n2294), .CP(clk), .Q(r11[30]) );
  DFQD1BWP12T r11_reg_28_ ( .D(n2292), .CP(clk), .Q(r11[28]) );
  DFQD1BWP12T r11_reg_27_ ( .D(n2291), .CP(clk), .Q(r11[27]) );
  DFQD1BWP12T r11_reg_26_ ( .D(n2290), .CP(clk), .Q(r11[26]) );
  DFQD1BWP12T r11_reg_25_ ( .D(n2289), .CP(clk), .Q(r11[25]) );
  DFQD1BWP12T r11_reg_24_ ( .D(n2288), .CP(clk), .Q(r11[24]) );
  DFQD1BWP12T r11_reg_23_ ( .D(n2287), .CP(clk), .Q(r11[23]) );
  DFQD1BWP12T r11_reg_22_ ( .D(n2286), .CP(clk), .Q(r11[22]) );
  DFQD1BWP12T r11_reg_21_ ( .D(n2285), .CP(clk), .Q(r11[21]) );
  DFQD1BWP12T r11_reg_20_ ( .D(n2284), .CP(clk), .Q(r11[20]) );
  DFQD1BWP12T r11_reg_19_ ( .D(n2283), .CP(clk), .Q(r11[19]) );
  DFQD1BWP12T r11_reg_18_ ( .D(n2282), .CP(clk), .Q(r11[18]) );
  DFQD1BWP12T r11_reg_16_ ( .D(n2280), .CP(clk), .Q(r11[16]) );
  DFQD1BWP12T r11_reg_15_ ( .D(n2279), .CP(clk), .Q(r11[15]) );
  DFQD1BWP12T r11_reg_14_ ( .D(n2278), .CP(clk), .Q(r11[14]) );
  DFQD1BWP12T r11_reg_13_ ( .D(n2277), .CP(clk), .Q(r11[13]) );
  DFQD1BWP12T r11_reg_12_ ( .D(n2276), .CP(clk), .Q(r11[12]) );
  DFQD1BWP12T r11_reg_11_ ( .D(n2275), .CP(clk), .Q(r11[11]) );
  DFQD1BWP12T r11_reg_10_ ( .D(n2274), .CP(clk), .Q(r11[10]) );
  DFQD1BWP12T r11_reg_9_ ( .D(n2273), .CP(clk), .Q(r11[9]) );
  DFQD1BWP12T r11_reg_8_ ( .D(n2272), .CP(clk), .Q(r11[8]) );
  DFQD1BWP12T r11_reg_7_ ( .D(n2271), .CP(clk), .Q(r11[7]) );
  DFQD1BWP12T r11_reg_6_ ( .D(n2270), .CP(clk), .Q(r11[6]) );
  DFQD1BWP12T r11_reg_5_ ( .D(n2269), .CP(clk), .Q(r11[5]) );
  DFQD1BWP12T r11_reg_4_ ( .D(n2268), .CP(clk), .Q(r11[4]) );
  DFQD1BWP12T r11_reg_3_ ( .D(n2267), .CP(clk), .Q(r11[3]) );
  DFQD1BWP12T r11_reg_2_ ( .D(n2266), .CP(clk), .Q(r11[2]) );
  DFQD1BWP12T r11_reg_1_ ( .D(n2265), .CP(clk), .Q(r11[1]) );
  DFQD1BWP12T r11_reg_0_ ( .D(n2264), .CP(clk), .Q(r11[0]) );
  DFQD1BWP12T r12_reg_30_ ( .D(n2262), .CP(clk), .Q(r12[30]) );
  DFQD1BWP12T r12_reg_28_ ( .D(n2260), .CP(clk), .Q(r12[28]) );
  DFQD1BWP12T r12_reg_27_ ( .D(n2259), .CP(clk), .Q(r12[27]) );
  DFQD1BWP12T r12_reg_26_ ( .D(n2258), .CP(clk), .Q(r12[26]) );
  DFQD1BWP12T r12_reg_25_ ( .D(n2257), .CP(clk), .Q(r12[25]) );
  DFQD1BWP12T r12_reg_24_ ( .D(n2256), .CP(clk), .Q(r12[24]) );
  DFQD1BWP12T r12_reg_23_ ( .D(n2255), .CP(clk), .Q(r12[23]) );
  DFQD1BWP12T r12_reg_22_ ( .D(n2254), .CP(clk), .Q(r12[22]) );
  DFQD1BWP12T r12_reg_21_ ( .D(n2253), .CP(clk), .Q(r12[21]) );
  DFQD1BWP12T r12_reg_20_ ( .D(n2252), .CP(clk), .Q(r12[20]) );
  DFQD1BWP12T r12_reg_19_ ( .D(n2251), .CP(clk), .Q(r12[19]) );
  DFQD1BWP12T r12_reg_17_ ( .D(n2249), .CP(clk), .Q(r12[17]) );
  DFQD1BWP12T r12_reg_16_ ( .D(n2248), .CP(clk), .Q(r12[16]) );
  DFQD1BWP12T r12_reg_15_ ( .D(n2247), .CP(clk), .Q(r12[15]) );
  DFQD1BWP12T r12_reg_14_ ( .D(n2246), .CP(clk), .Q(r12[14]) );
  DFQD1BWP12T r12_reg_13_ ( .D(n2245), .CP(clk), .Q(r12[13]) );
  DFQD1BWP12T r12_reg_11_ ( .D(n2243), .CP(clk), .Q(r12[11]) );
  DFQD1BWP12T r12_reg_10_ ( .D(n2242), .CP(clk), .Q(r12[10]) );
  DFQD1BWP12T r12_reg_9_ ( .D(n2241), .CP(clk), .Q(r12[9]) );
  DFQD1BWP12T r12_reg_8_ ( .D(n2240), .CP(clk), .Q(r12[8]) );
  DFQD1BWP12T r12_reg_7_ ( .D(n2239), .CP(clk), .Q(r12[7]) );
  DFQD1BWP12T r12_reg_6_ ( .D(n2238), .CP(clk), .Q(r12[6]) );
  DFQD1BWP12T r12_reg_5_ ( .D(n2237), .CP(clk), .Q(r12[5]) );
  DFQD1BWP12T r12_reg_4_ ( .D(n2236), .CP(clk), .Q(r12[4]) );
  DFQD1BWP12T r12_reg_3_ ( .D(n2235), .CP(clk), .Q(r12[3]) );
  DFQD1BWP12T r12_reg_2_ ( .D(n2234), .CP(clk), .Q(r12[2]) );
  DFQD1BWP12T r12_reg_1_ ( .D(n2233), .CP(clk), .Q(r12[1]) );
  DFQD1BWP12T r12_reg_0_ ( .D(n2232), .CP(clk), .Q(r12[0]) );
  DFQD1BWP12T lr_reg_31_ ( .D(n2231), .CP(clk), .Q(lr[31]) );
  DFQD1BWP12T lr_reg_30_ ( .D(n2230), .CP(clk), .Q(lr[30]) );
  DFQD1BWP12T lr_reg_29_ ( .D(n2229), .CP(clk), .Q(lr[29]) );
  DFQD1BWP12T lr_reg_28_ ( .D(n2228), .CP(clk), .Q(lr[28]) );
  DFQD1BWP12T lr_reg_27_ ( .D(n2227), .CP(clk), .Q(lr[27]) );
  DFQD1BWP12T lr_reg_26_ ( .D(n2226), .CP(clk), .Q(lr[26]) );
  DFQD1BWP12T lr_reg_25_ ( .D(n2225), .CP(clk), .Q(lr[25]) );
  DFQD1BWP12T lr_reg_24_ ( .D(n2224), .CP(clk), .Q(lr[24]) );
  DFQD1BWP12T lr_reg_23_ ( .D(n2223), .CP(clk), .Q(lr[23]) );
  DFQD1BWP12T lr_reg_22_ ( .D(n2222), .CP(clk), .Q(lr[22]) );
  DFQD1BWP12T lr_reg_20_ ( .D(n2220), .CP(clk), .Q(lr[20]) );
  DFQD1BWP12T lr_reg_19_ ( .D(n2219), .CP(clk), .Q(lr[19]) );
  DFQD1BWP12T lr_reg_16_ ( .D(n2216), .CP(clk), .Q(lr[16]) );
  DFQD1BWP12T lr_reg_15_ ( .D(n2215), .CP(clk), .Q(lr[15]) );
  DFQD1BWP12T lr_reg_14_ ( .D(n2214), .CP(clk), .Q(lr[14]) );
  DFQD1BWP12T lr_reg_13_ ( .D(n2213), .CP(clk), .Q(lr[13]) );
  DFQD1BWP12T lr_reg_12_ ( .D(n2212), .CP(clk), .Q(lr[12]) );
  DFQD1BWP12T lr_reg_11_ ( .D(n2211), .CP(clk), .Q(lr[11]) );
  DFQD1BWP12T lr_reg_10_ ( .D(n2210), .CP(clk), .Q(lr[10]) );
  DFQD1BWP12T lr_reg_9_ ( .D(n2209), .CP(clk), .Q(lr[9]) );
  DFQD1BWP12T lr_reg_8_ ( .D(n2208), .CP(clk), .Q(lr[8]) );
  DFQD1BWP12T lr_reg_7_ ( .D(n2207), .CP(clk), .Q(lr[7]) );
  DFQD1BWP12T lr_reg_6_ ( .D(n2206), .CP(clk), .Q(lr[6]) );
  DFQD1BWP12T lr_reg_5_ ( .D(n2205), .CP(clk), .Q(lr[5]) );
  DFQD1BWP12T lr_reg_4_ ( .D(n2204), .CP(clk), .Q(lr[4]) );
  DFQD1BWP12T lr_reg_3_ ( .D(n2203), .CP(clk), .Q(lr[3]) );
  DFQD1BWP12T lr_reg_2_ ( .D(n2202), .CP(clk), .Q(lr[2]) );
  DFQD1BWP12T lr_reg_1_ ( .D(n2201), .CP(clk), .Q(lr[1]) );
  DFQD1BWP12T lr_reg_0_ ( .D(n2200), .CP(clk), .Q(lr[0]) );
  DFQD1BWP12T sp_reg_30_ ( .D(spin[30]), .CP(clk), .Q(n[3550]) );
  DFQD1BWP12T sp_reg_29_ ( .D(spin[29]), .CP(clk), .Q(n[3551]) );
  DFQD1BWP12T sp_reg_28_ ( .D(spin[28]), .CP(clk), .Q(n[3552]) );
  DFQD1BWP12T sp_reg_27_ ( .D(spin[27]), .CP(clk), .Q(n[3553]) );
  DFQD1BWP12T sp_reg_26_ ( .D(spin[26]), .CP(clk), .Q(n[3554]) );
  DFQD1BWP12T sp_reg_25_ ( .D(spin[25]), .CP(clk), .Q(n[3555]) );
  DFQD1BWP12T sp_reg_24_ ( .D(spin[24]), .CP(clk), .Q(n[3556]) );
  DFQD1BWP12T sp_reg_23_ ( .D(spin[23]), .CP(clk), .Q(n[3557]) );
  DFQD1BWP12T sp_reg_22_ ( .D(spin[22]), .CP(clk), .Q(n[3558]) );
  DFQD1BWP12T sp_reg_21_ ( .D(spin[21]), .CP(clk), .Q(n[3559]) );
  DFQD1BWP12T sp_reg_20_ ( .D(spin[20]), .CP(clk), .Q(n[3560]) );
  DFQD1BWP12T sp_reg_19_ ( .D(spin[19]), .CP(clk), .Q(n[3561]) );
  DFQD1BWP12T sp_reg_18_ ( .D(spin[18]), .CP(clk), .Q(n[3562]) );
  DFQD1BWP12T sp_reg_17_ ( .D(spin[17]), .CP(clk), .Q(n[3563]) );
  DFQD1BWP12T sp_reg_16_ ( .D(spin[16]), .CP(clk), .Q(n[3564]) );
  DFQD1BWP12T sp_reg_15_ ( .D(spin[15]), .CP(clk), .Q(n[3565]) );
  DFQD1BWP12T sp_reg_13_ ( .D(spin[13]), .CP(clk), .Q(n[3567]) );
  DFQD1BWP12T sp_reg_12_ ( .D(spin[12]), .CP(clk), .Q(n[3568]) );
  DFQD1BWP12T sp_reg_11_ ( .D(spin[11]), .CP(clk), .Q(n[3569]) );
  DFQD1BWP12T sp_reg_10_ ( .D(spin[10]), .CP(clk), .Q(n[3570]) );
  DFQD1BWP12T sp_reg_9_ ( .D(spin[9]), .CP(clk), .Q(n[3571]) );
  DFQD1BWP12T sp_reg_8_ ( .D(spin[8]), .CP(clk), .Q(n[3572]) );
  DFQD1BWP12T sp_reg_7_ ( .D(spin[7]), .CP(clk), .Q(n[3573]) );
  DFQD1BWP12T sp_reg_6_ ( .D(spin[6]), .CP(clk), .Q(n[3574]) );
  DFQD1BWP12T sp_reg_5_ ( .D(spin[5]), .CP(clk), .Q(n[3575]) );
  DFQD1BWP12T sp_reg_4_ ( .D(spin[4]), .CP(clk), .Q(n[3576]) );
  DFQD1BWP12T sp_reg_3_ ( .D(spin[3]), .CP(clk), .Q(n[3577]) );
  DFQD1BWP12T sp_reg_2_ ( .D(spin[2]), .CP(clk), .Q(n[3578]) );
  DFQD1BWP12T sp_reg_1_ ( .D(spin[1]), .CP(clk), .Q(n[3579]) );
  DFQD1BWP12T sp_reg_0_ ( .D(spin[0]), .CP(clk), .Q(n[3580]) );
  DFQD1BWP12T pc_reg_24_ ( .D(n2192), .CP(clk), .Q(pc_out[24]) );
  DFQD1BWP12T pc_reg_20_ ( .D(n2188), .CP(clk), .Q(pc_out[20]) );
  DFQD1BWP12T pc_reg_19_ ( .D(n2187), .CP(clk), .Q(pc_out[19]) );
  DFQD1BWP12T pc_reg_18_ ( .D(n2186), .CP(clk), .Q(pc_out[18]) );
  DFQD1BWP12T pc_reg_17_ ( .D(n2185), .CP(clk), .Q(pc_out[17]) );
  DFQD1BWP12T pc_reg_16_ ( .D(n2184), .CP(clk), .Q(pc_out[16]) );
  DFQD1BWP12T pc_reg_14_ ( .D(n2182), .CP(clk), .Q(pc_out[14]) );
  DFQD1BWP12T pc_reg_13_ ( .D(n2181), .CP(clk), .Q(pc_out[13]) );
  DFQD1BWP12T pc_reg_12_ ( .D(n2180), .CP(clk), .Q(pc_out[12]) );
  DFQD1BWP12T pc_reg_10_ ( .D(n2178), .CP(clk), .Q(pc_out[10]) );
  DFQD1BWP12T pc_reg_9_ ( .D(n2177), .CP(clk), .Q(pc_out[9]) );
  DFQD1BWP12T pc_reg_8_ ( .D(n2176), .CP(clk), .Q(pc_out[8]) );
  DFQD1BWP12T pc_reg_5_ ( .D(n2173), .CP(clk), .Q(pc_out[5]) );
  DFQD1BWP12T pc_reg_4_ ( .D(n2172), .CP(clk), .Q(pc_out[4]) );
  DFQD1BWP12T pc_reg_2_ ( .D(n2170), .CP(clk), .Q(pc_out[2]) );
  DFQD1BWP12T pc_reg_0_ ( .D(n2168), .CP(clk), .Q(pc_out[0]) );
  DFQD1BWP12T cpsr_reg_3_ ( .D(cpsrin[3]), .CP(clk), .Q(cpsr_out[3]) );
  DFQD1BWP12T cpsr_reg_2_ ( .D(cpsrin[2]), .CP(clk), .Q(cpsr_out[2]) );
  DFQD1BWP12T tmp1_reg_30_ ( .D(n2166), .CP(clk), .Q(tmp1[30]) );
  DFQD1BWP12T tmp1_reg_29_ ( .D(n2165), .CP(clk), .Q(tmp1[29]) );
  DFQD1BWP12T tmp1_reg_28_ ( .D(n2164), .CP(clk), .Q(tmp1[28]) );
  DFQD1BWP12T tmp1_reg_27_ ( .D(n2163), .CP(clk), .Q(tmp1[27]) );
  DFQD1BWP12T tmp1_reg_26_ ( .D(n2162), .CP(clk), .Q(tmp1[26]) );
  DFQD1BWP12T tmp1_reg_25_ ( .D(n2161), .CP(clk), .Q(tmp1[25]) );
  DFQD1BWP12T tmp1_reg_24_ ( .D(n2160), .CP(clk), .Q(tmp1[24]) );
  DFQD1BWP12T tmp1_reg_23_ ( .D(n2159), .CP(clk), .Q(tmp1[23]) );
  DFQD1BWP12T tmp1_reg_22_ ( .D(n2158), .CP(clk), .Q(tmp1[22]) );
  DFQD1BWP12T tmp1_reg_21_ ( .D(n2157), .CP(clk), .Q(tmp1[21]) );
  DFQD1BWP12T tmp1_reg_20_ ( .D(n2156), .CP(clk), .Q(tmp1[20]) );
  DFQD1BWP12T tmp1_reg_19_ ( .D(n2155), .CP(clk), .Q(tmp1[19]) );
  DFQD1BWP12T tmp1_reg_18_ ( .D(n2154), .CP(clk), .Q(tmp1[18]) );
  DFQD1BWP12T tmp1_reg_17_ ( .D(n2153), .CP(clk), .Q(tmp1[17]) );
  DFQD1BWP12T tmp1_reg_16_ ( .D(n2152), .CP(clk), .Q(tmp1[16]) );
  DFQD1BWP12T tmp1_reg_15_ ( .D(n2151), .CP(clk), .Q(tmp1[15]) );
  DFQD1BWP12T tmp1_reg_14_ ( .D(n2150), .CP(clk), .Q(tmp1[14]) );
  DFQD1BWP12T tmp1_reg_13_ ( .D(n2149), .CP(clk), .Q(tmp1[13]) );
  DFQD1BWP12T tmp1_reg_12_ ( .D(n2148), .CP(clk), .Q(tmp1[12]) );
  DFQD1BWP12T tmp1_reg_11_ ( .D(n2147), .CP(clk), .Q(tmp1[11]) );
  DFQD1BWP12T tmp1_reg_10_ ( .D(n2146), .CP(clk), .Q(tmp1[10]) );
  DFQD1BWP12T tmp1_reg_9_ ( .D(n2145), .CP(clk), .Q(tmp1[9]) );
  DFQD1BWP12T tmp1_reg_8_ ( .D(n2144), .CP(clk), .Q(tmp1[8]) );
  DFQD1BWP12T tmp1_reg_7_ ( .D(n2143), .CP(clk), .Q(tmp1[7]) );
  DFQD1BWP12T tmp1_reg_6_ ( .D(n2142), .CP(clk), .Q(tmp1[6]) );
  DFQD1BWP12T tmp1_reg_5_ ( .D(n2141), .CP(clk), .Q(tmp1[5]) );
  DFQD1BWP12T tmp1_reg_4_ ( .D(n2140), .CP(clk), .Q(tmp1[4]) );
  DFQD1BWP12T tmp1_reg_3_ ( .D(n2139), .CP(clk), .Q(tmp1[3]) );
  DFQD1BWP12T tmp1_reg_2_ ( .D(n2138), .CP(clk), .Q(tmp1[2]) );
  DFQD1BWP12T tmp1_reg_1_ ( .D(n2137), .CP(clk), .Q(tmp1[1]) );
  DFQD1BWP12T tmp1_reg_0_ ( .D(n2135), .CP(clk), .Q(tmp1[0]) );
  DFQD4BWP12T pc_reg_1_ ( .D(n2169), .CP(clk), .Q(pc_out[1]) );
  DFQD2BWP12T pc_reg_23_ ( .D(n2191), .CP(clk), .Q(pc_out[23]) );
  DFQD1BWP12T sp_reg_31_ ( .D(spin[31]), .CP(clk), .Q(n[3549]) );
  DFKCNXD1BWP12T cpsr_reg_0_ ( .CN(n3532), .D(next_cpsr_in[0]), .CP(clk), .Q(
        cpsr_out[0]) );
  DFXD1BWP12T pc_reg_31_ ( .D(n2199), .CP(clk), .Q(pc_out[31]), .QN(n3548) );
  DFXD1BWP12T pc_reg_27_ ( .D(n2195), .CP(clk), .Q(pc_out[27]), .QN(n3538) );
  DFXD1BWP12T pc_reg_29_ ( .D(n2197), .CP(clk), .Q(pc_out[29]), .QN(n3533) );
  DFKCSND1BWP12T r2_reg_29_ ( .D(n3512), .SN(n3516), .CN(n3524), .CP(clk), .Q(
        n3540), .QN(r2[29]) );
  DFKCSND1BWP12T r3_reg_29_ ( .D(n3512), .SN(n3515), .CN(n3523), .CP(clk), .Q(
        n3534), .QN(r3[29]) );
  DFKCSND1BWP12T r10_reg_29_ ( .D(n3512), .SN(n3520), .CN(n3528), .CP(clk), 
        .Q(n3544), .QN(r10[29]) );
  DFXD1BWP12T pc_reg_22_ ( .D(n2190), .CP(clk), .Q(pc_out[22]), .QN(n3535) );
  DFXD1BWP12T pc_reg_21_ ( .D(n2189), .CP(clk), .Q(pc_out[21]), .QN(n3514) );
  DFXD1BWP12T pc_reg_25_ ( .D(n2193), .CP(clk), .Q(pc_out[25]), .QN(n3536) );
  DFKCSND1BWP12T r12_reg_29_ ( .D(n3512), .SN(n3521), .CN(n3529), .CP(clk), 
        .Q(n3541), .QN(r12[29]) );
  DFKCSND1BWP12T r4_reg_29_ ( .D(n3512), .SN(n3518), .CN(n3526), .CP(clk), .Q(
        n3543), .QN(r4[29]) );
  DFXD1BWP12T pc_reg_30_ ( .D(n2198), .CP(clk), .Q(pc_out[30]), .QN(n3547) );
  DFKCSND1BWP12T r8_reg_29_ ( .D(n3512), .SN(n3519), .CN(n3527), .CP(clk), .Q(
        n3542), .QN(r8[29]) );
  DFKCSND1BWP12T r0_reg_29_ ( .D(n3512), .SN(n3517), .CN(n3525), .CP(clk), .Q(
        n3546), .QN(r0[29]) );
  DFXD1BWP12T pc_reg_28_ ( .D(n2196), .CP(clk), .Q(pc_out[28]), .QN(n3539) );
  DFQD1BWP12T r11_reg_31_ ( .D(n2295), .CP(clk), .Q(r11[31]) );
  DFQD1BWP12T r1_reg_31_ ( .D(n2615), .CP(clk), .Q(r1[31]) );
  DFQD1BWP12T tmp1_reg_31_ ( .D(n2167), .CP(clk), .Q(tmp1[31]) );
  DFKCSND1BWP12T r10_reg_31_ ( .D(n3511), .SN(n3520), .CN(n3531), .CP(clk), 
        .Q(n3510), .QN(r10[31]) );
  DFKCSND1BWP12T r11_reg_29_ ( .D(n3513), .SN(n3522), .CN(n3530), .CP(clk), 
        .Q(n3545), .QN(r11[29]) );
  DFXD1BWP12T pc_reg_26_ ( .D(n2194), .CP(clk), .Q(pc_out[26]), .QN(n3537) );
  DFKCNQD1BWP12T cpsr_reg_1_ ( .CN(n3532), .D(next_cpsr_in[1]), .CP(clk), .Q(
        cpsr_out[1]) );
  DFQD1BWP12T pc_reg_11_ ( .D(n2179), .CP(clk), .Q(pc_out[11]) );
  DFQD1BWP12T pc_reg_3_ ( .D(n2171), .CP(clk), .Q(pc_out[3]) );
  DFQD1BWP12T r5_reg_2_ ( .D(n2458), .CP(clk), .Q(r5[2]) );
  DFQD1BWP12T r0_reg_1_ ( .D(n2617), .CP(clk), .Q(r0[1]) );
  DFQD1BWP12T pc_reg_7_ ( .D(n2175), .CP(clk), .Q(pc_out[7]) );
  DFQD1BWP12T r6_reg_7_ ( .D(n2431), .CP(clk), .Q(r6[7]) );
  DFQD1BWP12T r9_reg_7_ ( .D(n2335), .CP(clk), .Q(r9[7]) );
  DFQD1BWP12T sp_reg_14_ ( .D(spin[14]), .CP(clk), .Q(n[3566]) );
  DFQD1BWP12T r0_reg_7_ ( .D(n2623), .CP(clk), .Q(r0[7]) );
  DFQD1BWP12T r12_reg_18_ ( .D(n2250), .CP(clk), .Q(r12[18]) );
  DFQD1BWP12T r10_reg_13_ ( .D(n2309), .CP(clk), .Q(r10[13]) );
  DFQD1BWP12T r12_reg_12_ ( .D(n2244), .CP(clk), .Q(r12[12]) );
  DFQD1BWP12T r1_reg_18_ ( .D(n2602), .CP(clk), .Q(r1[18]) );
  DFQD1BWP12T r5_reg_21_ ( .D(n2477), .CP(clk), .Q(r5[21]) );
  DFQD1BWP12T lr_reg_18_ ( .D(n2218), .CP(clk), .Q(lr[18]) );
  DFQD1BWP12T lr_reg_21_ ( .D(n2221), .CP(clk), .Q(lr[21]) );
  DFQD1BWP12T r6_reg_5_ ( .D(n2429), .CP(clk), .Q(r6[5]) );
  DFQD1BWP12T r0_reg_12_ ( .D(n2628), .CP(clk), .Q(r0[12]) );
  DFQD1BWP12T r4_reg_7_ ( .D(n2495), .CP(clk), .Q(r4[7]) );
  DFQD1BWP12T r5_reg_15_ ( .D(n2471), .CP(clk), .Q(r5[15]) );
  DFQD1BWP12T pc_reg_6_ ( .D(n2174), .CP(clk), .Q(pc_out[6]) );
  DFQD1BWP12T r7_reg_17_ ( .D(n2409), .CP(clk), .Q(r7[17]) );
  DFQD1BWP12T r10_reg_17_ ( .D(n2313), .CP(clk), .Q(r10[17]) );
  DFQD1BWP12T r11_reg_17_ ( .D(n2281), .CP(clk), .Q(r11[17]) );
  DFQD1BWP12T lr_reg_17_ ( .D(n2217), .CP(clk), .Q(lr[17]) );
  DFQD1BWP12T r6_reg_26_ ( .D(n2450), .CP(clk), .Q(r6[26]) );
  DFQD1BWP12T r12_reg_31_ ( .D(n2263), .CP(clk), .Q(r12[31]) );
  DFQD1BWP12T r4_reg_31_ ( .D(n2519), .CP(clk), .Q(r4[31]) );
  DFQD1BWP12T r0_reg_31_ ( .D(n2647), .CP(clk), .Q(r0[31]) );
  DFQD1BWP12T r8_reg_31_ ( .D(n2391), .CP(clk), .Q(r8[31]) );
  DFQD1BWP12T pc_reg_15_ ( .D(n2183), .CP(clk), .Q(pc_out[15]) );
  TPNR3D1BWP12T U3 ( .A1(n849), .A2(n848), .A3(n847), .ZN(n850) );
  NR2D1BWP12T U4 ( .A1(n1246), .A2(n181), .ZN(n1253) );
  NR2D1BWP12T U5 ( .A1(n243), .A2(n242), .ZN(n248) );
  TPNR2D1BWP12T U6 ( .A1(n1251), .A2(n1250), .ZN(n1252) );
  TPNR2D2BWP12T U7 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  IOA21D1BWP12T U8 ( .A1(n846), .A2(lr[8]), .B(n845), .ZN(n849) );
  TPNR2D1BWP12T U9 ( .A1(n1425), .A2(n1424), .ZN(n1439) );
  OAI22D1BWP12T U10 ( .A1(n3396), .A2(n1752), .B1(n3442), .B2(n1751), .ZN(
        n1753) );
  OAI22D1BWP12T U11 ( .A1(n3396), .A2(n1830), .B1(n3442), .B2(n1829), .ZN(
        n1831) );
  OAI22D1BWP12T U12 ( .A1(n3452), .A2(n1828), .B1(n3393), .B2(n1827), .ZN(
        n1832) );
  IND2D1BWP12T U13 ( .A1(n1475), .B1(n1474), .ZN(n1476) );
  ND2D1BWP12T U14 ( .A1(n1200), .A2(r11[16]), .ZN(n1201) );
  ND2D1BWP12T U15 ( .A1(n1853), .A2(r4[16]), .ZN(n1221) );
  NR2D1BWP12T U16 ( .A1(n3442), .A2(n1223), .ZN(n1224) );
  IOA21D1BWP12T U17 ( .A1(n621), .A2(r12[16]), .B(n1208), .ZN(n1217) );
  ND3D1BWP12T U18 ( .A1(n632), .A2(n631), .A3(n630), .ZN(n633) );
  OAI22D1BWP12T U19 ( .A1(n3393), .A2(n604), .B1(n603), .B2(n3452), .ZN(n608)
         );
  OAI21D1BWP12T U20 ( .A1(n3414), .A2(n606), .B(n605), .ZN(n607) );
  INR2D1BWP12T U21 ( .A1(r12[11]), .B1(n3436), .ZN(n1298) );
  NR2D1BWP12T U22 ( .A1(n3396), .A2(n2880), .ZN(n1290) );
  NR2D1BWP12T U23 ( .A1(n3442), .A2(n2893), .ZN(n1291) );
  NR2D1BWP12T U24 ( .A1(n1920), .A2(n3541), .ZN(n754) );
  INR2D1BWP12T U25 ( .A1(pc_out[11]), .B1(n1917), .ZN(n259) );
  OAI22D1BWP12T U26 ( .A1(n1652), .A2(n2549), .B1(n1847), .B2(n1896), .ZN(
        n1556) );
  ND2D1BWP12T U27 ( .A1(next_pc_en_BAR), .A2(n536), .ZN(n3343) );
  INVD1BWP12T U28 ( .I(n535), .ZN(n536) );
  NR2D1BWP12T U29 ( .A1(n544), .A2(n561), .ZN(n547) );
  INR2D1BWP12T U30 ( .A1(n355), .B1(n361), .ZN(n531) );
  INVD1BWP12T U31 ( .I(n531), .ZN(n545) );
  INR2D1BWP12T U32 ( .A1(write2_sel[2]), .B1(n546), .ZN(n532) );
  ND2D1BWP12T U33 ( .A1(n594), .A2(n3532), .ZN(n595) );
  INR2D1BWP12T U34 ( .A1(write2_sel[2]), .B1(write2_sel[1]), .ZN(n594) );
  ND2D1BWP12T U35 ( .A1(n584), .A2(n3532), .ZN(n421) );
  INVD1BWP12T U36 ( .I(n1742), .ZN(n1739) );
  IND3D1BWP12T U37 ( .A1(write1_sel[0]), .B1(write1_sel[3]), .B2(n360), .ZN(
        n591) );
  IND3D1BWP12T U38 ( .A1(write1_sel[0]), .B1(n358), .B2(n360), .ZN(n585) );
  AOI21D1BWP12T U39 ( .A1(write1_in[20]), .A2(n530), .B(n1737), .ZN(n3506) );
  OR2XD1BWP12T U40 ( .A1(n421), .A2(n544), .Z(n2872) );
  AOI211D1BWP12T U41 ( .A1(n532), .A2(n593), .B(n3259), .C(reset), .ZN(n3261)
         );
  NR3D1BWP12T U42 ( .A1(n3259), .A2(n363), .A3(n596), .ZN(n3260) );
  INVD1BWP12T U43 ( .I(n3020), .ZN(n3259) );
  INR3D0BWP12T U44 ( .A1(n550), .B1(reset), .B2(n551), .ZN(n3198) );
  NR2D1BWP12T U45 ( .A1(n551), .A2(n550), .ZN(n3197) );
  OR2XD1BWP12T U46 ( .A1(n544), .A2(n422), .Z(n3015) );
  AOI211D1BWP12T U47 ( .A1(n531), .A2(n579), .B(n3269), .C(reset), .ZN(n3271)
         );
  NR3D1BWP12T U48 ( .A1(n3269), .A2(n580), .A3(n545), .ZN(n3270) );
  INVD1BWP12T U49 ( .I(n3015), .ZN(n3269) );
  NR3D1BWP12T U50 ( .A1(n3264), .A2(n364), .A3(n363), .ZN(n3265) );
  AOI211D1BWP12T U51 ( .A1(n532), .A2(n554), .B(n3264), .C(reset), .ZN(n3266)
         );
  INVD1BWP12T U52 ( .I(n2999), .ZN(n3264) );
  AOI211D1BWP12T U53 ( .A1(n532), .A2(n586), .B(n3274), .C(reset), .ZN(n3277)
         );
  NR3D1BWP12T U54 ( .A1(n3274), .A2(n363), .A3(n587), .ZN(n3276) );
  INVD1BWP12T U55 ( .I(n3007), .ZN(n3274) );
  NR3D1BWP12T U56 ( .A1(n3254), .A2(n364), .A3(n595), .ZN(n3255) );
  AOI211D1BWP12T U57 ( .A1(n594), .A2(n554), .B(n3254), .C(reset), .ZN(n3256)
         );
  INVD1BWP12T U58 ( .I(n3003), .ZN(n3254) );
  INR3D0BWP12T U59 ( .A1(n562), .B1(reset), .B2(n563), .ZN(n3194) );
  NR2D1BWP12T U60 ( .A1(n563), .A2(n562), .ZN(n3193) );
  INVD2BWP12T U61 ( .I(n3512), .ZN(n3247) );
  NR3D1BWP12T U62 ( .A1(n3231), .A2(n580), .A3(n364), .ZN(n3232) );
  INVD1BWP12T U63 ( .I(n3011), .ZN(n3231) );
  NR2D1BWP12T U64 ( .A1(n585), .A2(n421), .ZN(n3518) );
  NR2D1BWP12T U65 ( .A1(n591), .A2(n421), .ZN(n3521) );
  NR2D1BWP12T U66 ( .A1(n591), .A2(n420), .ZN(n3520) );
  NR2D1BWP12T U67 ( .A1(n555), .A2(n420), .ZN(n3515) );
  ND3D1BWP12T U68 ( .A1(n795), .A2(n794), .A3(n793), .ZN(regA_out[24]) );
  ND3D1BWP12T U69 ( .A1(n230), .A2(n229), .A3(n228), .ZN(regA_out[22]) );
  OAI22D1BWP12T U70 ( .A1(n3416), .A2(n1974), .B1(n3436), .B2(n1747), .ZN(
        n1756) );
  OAI22D1BWP12T U71 ( .A1(n3452), .A2(n1975), .B1(n3393), .B2(n1750), .ZN(
        n1754) );
  ND2D1BWP12T U72 ( .A1(n1886), .A2(n1885), .ZN(regA_out[20]) );
  ND3D1BWP12T U73 ( .A1(n352), .A2(n351), .A3(n350), .ZN(regA_out[26]) );
  INVD1BWP12T U74 ( .I(n1842), .ZN(n1843) );
  ND2D1BWP12T U75 ( .A1(n3384), .A2(r1[25]), .ZN(n1842) );
  AOI21D1BWP12T U76 ( .A1(n1839), .A2(r7[25]), .B(n1838), .ZN(n1845) );
  INR2D1BWP12T U77 ( .A1(r5[25]), .B1(n1837), .ZN(n1838) );
  OAI22D1BWP12T U78 ( .A1(n3416), .A2(n1824), .B1(n3436), .B2(n1823), .ZN(
        n1834) );
  OAI22D1BWP12T U79 ( .A1(n3436), .A2(n3541), .B1(n3416), .B2(n2656), .ZN(
        n1644) );
  NR3D2BWP12T U80 ( .A1(n1793), .A2(n1792), .A3(n1791), .ZN(n1801) );
  AN2D1BWP12T U81 ( .A1(n1853), .A2(r4[21]), .Z(n1792) );
  NR3D1BWP12T U82 ( .A1(n1799), .A2(n1798), .A3(n1797), .ZN(n1800) );
  NR2D1BWP12T U83 ( .A1(n3442), .A2(n1796), .ZN(n1798) );
  NR2D1BWP12T U84 ( .A1(n3432), .A2(n2824), .ZN(n456) );
  INR2D1BWP12T U85 ( .A1(r12[12]), .B1(n3436), .ZN(n1471) );
  OAI22D1BWP12T U86 ( .A1(n3402), .A2(n1816), .B1(n1959), .B2(n3452), .ZN(
        n1817) );
  OAI22D1BWP12T U87 ( .A1(n3390), .A2(n1957), .B1(n1956), .B2(n3442), .ZN(
        n1819) );
  CKND2D2BWP12T U88 ( .A1(n1622), .A2(r2[1]), .ZN(n1624) );
  ND2D1BWP12T U89 ( .A1(n1804), .A2(immediate1_in[1]), .ZN(n1623) );
  AOI21D1BWP12T U90 ( .A1(n1862), .A2(n[3563]), .B(n617), .ZN(n620) );
  NR2D1BWP12T U91 ( .A1(n616), .A2(n615), .ZN(n617) );
  INVD1BWP12T U92 ( .I(n3442), .ZN(n629) );
  INVD1BWP12T U93 ( .I(n876), .ZN(n878) );
  INR2D1BWP12T U94 ( .A1(n880), .B1(write1_in[18]), .ZN(n876) );
  ND2D1BWP12T U95 ( .A1(n657), .A2(n656), .ZN(n658) );
  NR2D1BWP12T U96 ( .A1(n655), .A2(n654), .ZN(n656) );
  ND3D1BWP12T U97 ( .A1(n1383), .A2(n1382), .A3(n1381), .ZN(n1384) );
  NR2D1BWP12T U98 ( .A1(n3432), .A2(n2943), .ZN(n1189) );
  INR2D1BWP12T U99 ( .A1(r5[5]), .B1(n3414), .ZN(n690) );
  ND2D1BWP12T U100 ( .A1(n1839), .A2(r7[5]), .ZN(n707) );
  NR2D1BWP12T U101 ( .A1(n1630), .A2(n1629), .ZN(n1631) );
  OAI22D1BWP12T U102 ( .A1(n2801), .A2(n3387), .B1(n3436), .B2(n1948), .ZN(
        n1630) );
  OAI22D1BWP12T U103 ( .A1(n3402), .A2(n2804), .B1(n2829), .B2(n3452), .ZN(
        n1629) );
  NR2D1BWP12T U104 ( .A1(n1616), .A2(n1615), .ZN(n1634) );
  OAI22D1BWP12T U105 ( .A1(n3414), .A2(n1614), .B1(n1810), .B2(n1613), .ZN(
        n1615) );
  OAI22D1BWP12T U106 ( .A1(n3406), .A2(n2807), .B1(n1612), .B2(n3444), .ZN(
        n1616) );
  NR2D1BWP12T U107 ( .A1(n1619), .A2(n1618), .ZN(n1633) );
  OAI22D1BWP12T U108 ( .A1(n3434), .A2(n1951), .B1(n3446), .B2(n2832), .ZN(
        n1618) );
  INR2D1BWP12T U109 ( .A1(r8[19]), .B1(n3387), .ZN(n665) );
  ND2D1BWP12T U110 ( .A1(n1853), .A2(r4[19]), .ZN(n666) );
  ND2D1BWP12T U111 ( .A1(n1859), .A2(lr[19]), .ZN(n669) );
  ND2D1BWP12T U112 ( .A1(n1788), .A2(pc_out[19]), .ZN(n678) );
  ND2D1BWP12T U113 ( .A1(n1380), .A2(tmp1[19]), .ZN(n679) );
  INVD1BWP12T U114 ( .I(write1_sel[1]), .ZN(n359) );
  INVD1BWP12T U115 ( .I(write2_sel[3]), .ZN(n361) );
  INVD1BWP12T U116 ( .I(n543), .ZN(n561) );
  AN2D1BWP12T U117 ( .A1(write2_sel[0]), .A2(n362), .Z(n355) );
  INR2D1BWP12T U118 ( .A1(write2_en), .B1(write2_sel[4]), .ZN(n362) );
  AOI21D1BWP12T U119 ( .A1(n3412), .A2(r6[7]), .B(n854), .ZN(n857) );
  INR3D0BWP12T U120 ( .A1(n1481), .B1(n1480), .B2(n1479), .ZN(n1482) );
  INR3D0BWP12T U121 ( .A1(n1468), .B1(n1467), .B2(n1466), .ZN(n1484) );
  ND2D1BWP12T U122 ( .A1(n645), .A2(n644), .ZN(n646) );
  ND2D1BWP12T U123 ( .A1(n642), .A2(n641), .ZN(n648) );
  NR2D1BWP12T U124 ( .A1(n640), .A2(n639), .ZN(n641) );
  ND2D1BWP12T U125 ( .A1(n3418), .A2(r11[14]), .ZN(n643) );
  ND2D1BWP12T U126 ( .A1(n3418), .A2(r11[15]), .ZN(n1371) );
  OAI21D1BWP12T U127 ( .A1(n3444), .A2(n1391), .B(n1390), .ZN(n1392) );
  ND2D1BWP12T U128 ( .A1(n1859), .A2(lr[15]), .ZN(n1390) );
  OAI22D1BWP12T U129 ( .A1(n3390), .A2(n2944), .B1(n2945), .B2(n3442), .ZN(
        n1187) );
  OAI22D1BWP12T U130 ( .A1(n3416), .A2(n2990), .B1(n3393), .B2(n2947), .ZN(
        n1188) );
  ND2D1BWP12T U131 ( .A1(n751), .A2(n750), .ZN(regA_out[4]) );
  NR3D1BWP12T U132 ( .A1(n1226), .A2(n1225), .A3(n1224), .ZN(n1227) );
  ND2D3BWP12T U133 ( .A1(n636), .A2(n635), .ZN(regA_out[17]) );
  INR2D2BWP12T U134 ( .A1(n634), .B1(n633), .ZN(n635) );
  ND2D1BWP12T U135 ( .A1(n1300), .A2(n1299), .ZN(n1301) );
  INVD1BWP12T U136 ( .I(n1298), .ZN(n1300) );
  ND2D1BWP12T U137 ( .A1(n1645), .A2(r9[11]), .ZN(n1306) );
  NR2D1BWP12T U138 ( .A1(n3435), .A2(n3025), .ZN(n1304) );
  ND2D1BWP12T U139 ( .A1(n1293), .A2(n1292), .ZN(n1294) );
  ND2D1BWP12T U140 ( .A1(n1411), .A2(n1410), .ZN(regA_out[10]) );
  INVD1BWP12T U141 ( .I(n1676), .ZN(n1677) );
  INR2D1BWP12T U142 ( .A1(r9[21]), .B1(n1553), .ZN(n329) );
  INR2D1BWP12T U143 ( .A1(r10[21]), .B1(n1899), .ZN(n328) );
  NR2D1BWP12T U144 ( .A1(n1895), .A2(n957), .ZN(n958) );
  INR2D1BWP12T U145 ( .A1(r10[5]), .B1(n1592), .ZN(n951) );
  ND2D1BWP12T U146 ( .A1(n1567), .A2(immediate2_in[16]), .ZN(n300) );
  NR2D1BWP12T U147 ( .A1(n1669), .A2(n2656), .ZN(n757) );
  NR2D1BWP12T U148 ( .A1(n1519), .A2(n3540), .ZN(n759) );
  ND2D1BWP12T U149 ( .A1(n1915), .A2(r6[10]), .ZN(n984) );
  INR2D1BWP12T U150 ( .A1(lr[10]), .B1(n1669), .ZN(n986) );
  INVD1BWP12T U151 ( .I(n1578), .ZN(n1580) );
  ND2D1BWP12T U152 ( .A1(n1907), .A2(immediate2_in[14]), .ZN(n1528) );
  NR2D1BWP12T U153 ( .A1(n1669), .A2(n1992), .ZN(n1535) );
  MOAI22D0BWP12T U154 ( .A1(n2851), .A2(n1669), .B1(n1713), .B2(
        immediate2_in[3]), .ZN(n1255) );
  INVD1BWP12T U155 ( .I(r12[4]), .ZN(n176) );
  ND2D1BWP12T U156 ( .A1(n1713), .A2(immediate2_in[7]), .ZN(n1716) );
  OR3XD1BWP12T U157 ( .A1(readC_sel[2]), .A2(n405), .A3(readC_sel[4]), .Z(n403) );
  NR2D1BWP12T U158 ( .A1(write1_in[28]), .A2(n3331), .ZN(n1033) );
  INR2D1BWP12T U159 ( .A1(write1_en), .B1(write1_sel[4]), .ZN(n360) );
  INVD1BWP12T U160 ( .I(write1_sel[3]), .ZN(n358) );
  NR2D1BWP12T U161 ( .A1(n359), .A2(write1_sel[2]), .ZN(n543) );
  NR2D1BWP12T U162 ( .A1(n530), .A2(n529), .ZN(n3318) );
  INR2D1BWP12T U163 ( .A1(write1_sel[2]), .B1(n359), .ZN(n482) );
  ND2D1BWP12T U164 ( .A1(n602), .A2(n3532), .ZN(n535) );
  INVD1BWP12T U165 ( .I(write2_sel[1]), .ZN(n546) );
  NR3D1BWP12T U166 ( .A1(n546), .A2(reset), .A3(write2_sel[2]), .ZN(n560) );
  INVD1BWP12T U167 ( .I(n593), .ZN(n596) );
  INR3D0BWP12T U168 ( .A1(n362), .B1(write2_sel[0]), .B2(n361), .ZN(n593) );
  ND2D1BWP12T U169 ( .A1(n482), .A2(n3532), .ZN(n366) );
  ND2D1BWP12T U170 ( .A1(n532), .A2(n3532), .ZN(n363) );
  NR2D1BWP12T U171 ( .A1(n555), .A2(n561), .ZN(n557) );
  ND2D1BWP12T U172 ( .A1(n419), .A2(n3532), .ZN(n422) );
  INVD1BWP12T U173 ( .I(n554), .ZN(n364) );
  INR2D1BWP12T U174 ( .A1(n355), .B1(write2_sel[3]), .ZN(n554) );
  INR3D0BWP12T U175 ( .A1(n362), .B1(write2_sel[3]), .B2(write2_sel[0]), .ZN(
        n586) );
  NR2D1BWP12T U176 ( .A1(write2_sel[1]), .A2(write2_sel[2]), .ZN(n579) );
  INVD1BWP12T U177 ( .I(n586), .ZN(n587) );
  ND2D1BWP12T U178 ( .A1(n579), .A2(n3532), .ZN(n580) );
  INR3D0BWP12T U179 ( .A1(n871), .B1(n870), .B2(n869), .ZN(n872) );
  ND2D1BWP12T U180 ( .A1(n1200), .A2(r11[7]), .ZN(n871) );
  INR2D1BWP12T U181 ( .A1(r8[7]), .B1(n3435), .ZN(n853) );
  NR2D2BWP12T U182 ( .A1(n165), .A2(n275), .ZN(n270) );
  OAI22D1BWP12T U183 ( .A1(n1887), .A2(n2062), .B1(n1889), .B2(n390), .ZN(n393) );
  ND3D1BWP12T U184 ( .A1(n381), .A2(n380), .A3(n379), .ZN(n382) );
  OR2XD1BWP12T U185 ( .A1(n1714), .A2(n378), .Z(n380) );
  ND2D1BWP12T U186 ( .A1(n1907), .A2(immediate2_in[22]), .ZN(n379) );
  IND3D1BWP12T U187 ( .A1(n720), .B1(n719), .B2(n718), .ZN(n728) );
  INVD1BWP12T U188 ( .I(n717), .ZN(n719) );
  IND2D1BWP12T U189 ( .A1(n1111), .B1(n1110), .ZN(n1116) );
  ND3D1BWP12T U190 ( .A1(n1114), .A2(n1113), .A3(n1112), .ZN(n1115) );
  ND2D1BWP12T U191 ( .A1(n1907), .A2(immediate2_in[18]), .ZN(n1112) );
  OAI22D1BWP12T U192 ( .A1(n1887), .A2(n2098), .B1(n160), .B2(n3413), .ZN(
        n1119) );
  IOA21D1BWP12T U193 ( .A1(n1921), .A2(tmp1[2]), .B(n1655), .ZN(n1656) );
  IND2D1BWP12T U194 ( .A1(n317), .B1(n316), .ZN(n325) );
  ND3D1BWP12T U195 ( .A1(n323), .A2(n322), .A3(n321), .ZN(n324) );
  ND2D1BWP12T U196 ( .A1(n1907), .A2(immediate2_in[21]), .ZN(n321) );
  IOA21D1BWP12T U197 ( .A1(n1909), .A2(lr[5]), .B(n974), .ZN(n979) );
  ND2D1BWP12T U198 ( .A1(n1907), .A2(immediate2_in[5]), .ZN(n974) );
  IOA21D1BWP12T U199 ( .A1(n1571), .A2(r8[5]), .B(n970), .ZN(n971) );
  OAI22D1BWP12T U200 ( .A1(n1587), .A2(n1223), .B1(n1222), .B2(n1895), .ZN(
        n311) );
  ND2D1BWP12T U201 ( .A1(n1907), .A2(immediate2_in[28]), .ZN(n1325) );
  AN3XD2BWP12T U202 ( .A1(n1328), .A2(n1327), .A3(n1326), .Z(n1329) );
  AOI22D1BWP12T U203 ( .A1(n1921), .A2(tmp1[28]), .B1(r8[28]), .B2(n1571), 
        .ZN(n1327) );
  AOI21D1BWP12T U204 ( .A1(n1918), .A2(r4[29]), .B(n754), .ZN(n755) );
  ND3D1BWP12T U205 ( .A1(n989), .A2(n988), .A3(n987), .ZN(n993) );
  AOI21D1BWP12T U206 ( .A1(immediate2_in[10]), .A2(n1567), .B(n986), .ZN(n987)
         );
  INR2D1BWP12T U207 ( .A1(n984), .B1(n983), .ZN(n989) );
  CKND2D2BWP12T U208 ( .A1(n1095), .A2(n182), .ZN(n1102) );
  TPOAI22D1BWP12T U209 ( .A1(n1663), .A2(n2662), .B1(n1367), .B2(n1592), .ZN(
        n1106) );
  OAI22D1BWP12T U210 ( .A1(n1887), .A2(n3392), .B1(n161), .B2(n3380), .ZN(n807) );
  OAI22D1BWP12T U211 ( .A1(n1519), .A2(n3376), .B1(n1911), .B2(n796), .ZN(n798) );
  INVD1BWP12T U212 ( .I(n259), .ZN(n264) );
  INR2D1BWP12T U213 ( .A1(n255), .B1(n254), .ZN(n265) );
  ND2D1BWP12T U214 ( .A1(n272), .A2(n271), .ZN(n273) );
  OAI22D1BWP12T U215 ( .A1(n1587), .A2(n2893), .B1(n2878), .B2(n1724), .ZN(
        n292) );
  ND3D1BWP12T U216 ( .A1(n1581), .A2(n1580), .A3(n1579), .ZN(n1582) );
  AOI22D1BWP12T U217 ( .A1(n1575), .A2(pc_out[24]), .B1(r6[24]), .B2(n1915), 
        .ZN(n1581) );
  ND2D1BWP12T U218 ( .A1(n1907), .A2(immediate2_in[24]), .ZN(n1579) );
  OAI22D1BWP12T U219 ( .A1(n1592), .A2(n1591), .B1(n1590), .B2(n1589), .ZN(
        n1593) );
  OAI21D1BWP12T U220 ( .A1(n1663), .A2(n1542), .B(n1541), .ZN(n1543) );
  INVD1BWP12T U221 ( .I(n1540), .ZN(n1541) );
  INR2D1BWP12T U222 ( .A1(r10[14]), .B1(n1899), .ZN(n1540) );
  NR2D1BWP12T U223 ( .A1(n1911), .A2(n1910), .ZN(n1912) );
  OAI21D1BWP12T U224 ( .A1(n1917), .A2(n2874), .B(n1916), .ZN(n1928) );
  ND2D1BWP12T U225 ( .A1(n1918), .A2(r4[6]), .ZN(n1919) );
  OAI22D1BWP12T U226 ( .A1(n1587), .A2(n1956), .B1(n1807), .B2(n1724), .ZN(
        n1269) );
  OAI22D1BWP12T U227 ( .A1(n1553), .A2(n1816), .B1(n1899), .B2(n1959), .ZN(
        n1270) );
  IND2D1BWP12T U228 ( .A1(n917), .B1(n916), .ZN(n922) );
  ND2D1BWP12T U229 ( .A1(n1907), .A2(immediate2_in[20]), .ZN(n918) );
  AOI22D1BWP12T U230 ( .A1(n1575), .A2(pc_out[25]), .B1(r6[25]), .B2(n1915), 
        .ZN(n1561) );
  OAI22D1BWP12T U231 ( .A1(n1519), .A2(n1841), .B1(n1911), .B2(n1563), .ZN(
        n1566) );
  NR2D2BWP12T U232 ( .A1(n1559), .A2(n1558), .ZN(n1570) );
  OR2XD2BWP12T U233 ( .A1(n1557), .A2(n1556), .Z(n1558) );
  INVD1BWP12T U234 ( .I(n3478), .ZN(n2810) );
  NR2D1BWP12T U235 ( .A1(n406), .A2(n403), .ZN(n3475) );
  NR2D1BWP12T U236 ( .A1(n407), .A2(n400), .ZN(n3473) );
  NR2D1BWP12T U237 ( .A1(n410), .A2(n404), .ZN(n3482) );
  NR2D1BWP12T U238 ( .A1(n406), .A2(n404), .ZN(n3481) );
  NR2D1BWP12T U239 ( .A1(n410), .A2(n409), .ZN(n3485) );
  NR2D1BWP12T U240 ( .A1(n409), .A2(n408), .ZN(n3486) );
  NR2D1BWP12T U241 ( .A1(n409), .A2(n406), .ZN(n3484) );
  NR2D1BWP12T U242 ( .A1(n409), .A2(n407), .ZN(n3483) );
  INVD1BWP12T U243 ( .I(readC_sel[4]), .ZN(n3492) );
  INVD1BWP12T U244 ( .I(n2800), .ZN(n3493) );
  INVD1BWP12T U245 ( .I(n2806), .ZN(n3480) );
  INVD1BWP12T U246 ( .I(n2744), .ZN(n3479) );
  NR3D1BWP12T U247 ( .A1(n1033), .A2(n1029), .A3(n3497), .ZN(n1035) );
  ND3D1BWP12T U248 ( .A1(n360), .A2(write1_sel[0]), .A3(n358), .ZN(n555) );
  ND2D1BWP12T U249 ( .A1(n543), .A2(n3532), .ZN(n420) );
  AOI21D1BWP12T U250 ( .A1(write1_in[28]), .A2(n530), .B(n1037), .ZN(n1605) );
  NR2D1BWP12T U251 ( .A1(n1602), .A2(n1601), .ZN(n1604) );
  NR2D1BWP12T U252 ( .A1(write1_in[29]), .A2(n3324), .ZN(n1602) );
  NR2D1BWP12T U253 ( .A1(n1038), .A2(n3497), .ZN(n533) );
  INVD1BWP12T U254 ( .I(r4[7]), .ZN(n2865) );
  CKBD1BWP12T U255 ( .I(write1_in[8]), .Z(n166) );
  IOA21D1BWP12T U256 ( .A1(write1_in[1]), .A2(n530), .B(n507), .ZN(n2844) );
  AOI21D1BWP12T U257 ( .A1(write1_in[3]), .A2(n530), .B(n508), .ZN(n2949) );
  RCOAI21D1BWP12T U258 ( .A1(n500), .A2(n3331), .B(n499), .ZN(n3058) );
  INVD1BWP12T U259 ( .I(write1_in[8]), .ZN(n500) );
  ND2D1BWP12T U260 ( .A1(n1936), .A2(n1935), .ZN(n3111) );
  CKBD1BWP12T U261 ( .I(n3250), .Z(n163) );
  INVD1BWP12T U262 ( .I(n3343), .ZN(n3498) );
  OAI21D1BWP12T U263 ( .A1(n3094), .A2(n3331), .B(n1160), .ZN(n3502) );
  OR2XD1BWP12T U264 ( .A1(n3506), .A2(n3497), .Z(n3501) );
  AN2D1BWP12T U265 ( .A1(n3307), .A2(n3505), .Z(n3298) );
  AOI211D1BWP12T U266 ( .A1(n531), .A2(n594), .B(n3184), .C(reset), .ZN(n3186)
         );
  NR3D1BWP12T U267 ( .A1(n3184), .A2(n545), .A3(n595), .ZN(n3185) );
  OR2XD1BWP12T U268 ( .A1(n366), .A2(n591), .Z(n3020) );
  INVD1BWP12T U269 ( .I(n3261), .ZN(n3022) );
  INVD1BWP12T U270 ( .I(n3260), .ZN(n3018) );
  INVD1BWP12T U271 ( .I(r12[7]), .ZN(n2846) );
  INVD1BWP12T U272 ( .I(n3521), .ZN(n2957) );
  INVD1BWP12T U273 ( .I(n3227), .ZN(n2958) );
  INVD1BWP12T U274 ( .I(n3228), .ZN(n2956) );
  INVD1BWP12T U275 ( .I(r11[0]), .ZN(n3067) );
  INVD1BWP12T U276 ( .I(r11[3]), .ZN(n2852) );
  INVD1BWP12T U277 ( .I(n3522), .ZN(n2965) );
  INVD1BWP12T U278 ( .I(n3201), .ZN(n2964) );
  INVD1BWP12T U279 ( .I(n3202), .ZN(n2966) );
  INVD1BWP12T U280 ( .I(n3520), .ZN(n2977) );
  INVD1BWP12T U281 ( .I(n3198), .ZN(n2976) );
  INVD1BWP12T U282 ( .I(n3197), .ZN(n2978) );
  INVD1BWP12T U283 ( .I(r9[0]), .ZN(n2711) );
  INVD1BWP12T U284 ( .I(r9[3]), .ZN(n1816) );
  INVD1BWP12T U285 ( .I(n3271), .ZN(n3016) );
  INVD1BWP12T U286 ( .I(n3270), .ZN(n3014) );
  INVD1BWP12T U287 ( .I(n3519), .ZN(n2961) );
  INVD1BWP12T U288 ( .I(n3214), .ZN(n2962) );
  INVD1BWP12T U289 ( .I(n3215), .ZN(n2960) );
  INVD1BWP12T U290 ( .I(r7[7]), .ZN(n1723) );
  OR2XD1BWP12T U291 ( .A1(n555), .A2(n366), .Z(n2999) );
  INVD1BWP12T U292 ( .I(n3265), .ZN(n2998) );
  INVD1BWP12T U293 ( .I(n3266), .ZN(n3000) );
  OR2XD1BWP12T U294 ( .A1(n366), .A2(n585), .Z(n3007) );
  INVD1BWP12T U295 ( .I(n3277), .ZN(n3008) );
  INVD1BWP12T U296 ( .I(n3276), .ZN(n3006) );
  INVD1BWP12T U297 ( .I(r5[0]), .ZN(n730) );
  OR2XD1BWP12T U298 ( .A1(n555), .A2(n421), .Z(n3003) );
  INVD1BWP12T U299 ( .I(n3255), .ZN(n3002) );
  INVD1BWP12T U300 ( .I(n3256), .ZN(n3004) );
  INVD1BWP12T U301 ( .I(n3518), .ZN(n2953) );
  INVD1BWP12T U302 ( .I(n3222), .ZN(n2954) );
  INVD1BWP12T U303 ( .I(n3223), .ZN(n2952) );
  INVD1BWP12T U304 ( .I(n3515), .ZN(n2969) );
  INVD1BWP12T U305 ( .I(r3[11]), .ZN(n2888) );
  INVD1BWP12T U306 ( .I(n3189), .ZN(n2970) );
  INVD1BWP12T U307 ( .I(n3190), .ZN(n2968) );
  INVD1BWP12T U308 ( .I(r2[3]), .ZN(n1960) );
  INVD1BWP12T U309 ( .I(r2[9]), .ZN(n2943) );
  INVD1BWP12T U310 ( .I(n3516), .ZN(n2973) );
  INVD1BWP12T U311 ( .I(r2[11]), .ZN(n2896) );
  INVD1BWP12T U312 ( .I(n3194), .ZN(n2972) );
  INVD1BWP12T U313 ( .I(n3193), .ZN(n2974) );
  INVD1BWP12T U314 ( .I(write1_in[1]), .ZN(n1953) );
  INVD1BWP12T U315 ( .I(write2_in[1]), .ZN(n1954) );
  INVD1BWP12T U316 ( .I(r1[3]), .ZN(n1809) );
  INVD1BWP12T U317 ( .I(write1_in[7]), .ZN(n2866) );
  INVD1BWP12T U318 ( .I(write2_in[7]), .ZN(n2867) );
  OR2XD1BWP12T U319 ( .A1(n555), .A2(n422), .Z(n3011) );
  INVD1BWP12T U320 ( .I(n3232), .ZN(n3010) );
  INVD1BWP12T U321 ( .I(n3233), .ZN(n3012) );
  CKBD1BWP12T U322 ( .I(write1_in[15]), .Z(n177) );
  INVD1BWP12T U323 ( .I(write1_in[0]), .ZN(n2825) );
  INVD1BWP12T U324 ( .I(write2_in[0]), .ZN(n2826) );
  INVD1BWP12T U325 ( .I(write1_in[2]), .ZN(n2003) );
  INVD1BWP12T U326 ( .I(write2_in[2]), .ZN(n2004) );
  INVD1BWP12T U327 ( .I(r0[3]), .ZN(n1956) );
  INVD1BWP12T U328 ( .I(write1_in[3]), .ZN(n1961) );
  INVD1BWP12T U329 ( .I(write2_in[3]), .ZN(n1962) );
  INVD1BWP12T U330 ( .I(write1_in[4]), .ZN(n2014) );
  INVD1BWP12T U331 ( .I(write2_in[4]), .ZN(n2015) );
  INVD1BWP12T U332 ( .I(write1_in[5]), .ZN(n2022) );
  INVD1BWP12T U333 ( .I(write2_in[5]), .ZN(n2023) );
  INVD1BWP12T U334 ( .I(write1_in[6]), .ZN(n2031) );
  INVD1BWP12T U335 ( .I(write2_in[6]), .ZN(n2032) );
  INVD1BWP12T U336 ( .I(n166), .ZN(n2934) );
  INVD1BWP12T U337 ( .I(write2_in[8]), .ZN(n2933) );
  INVD1BWP12T U338 ( .I(write1_in[9]), .ZN(n2989) );
  INVD1BWP12T U339 ( .I(write2_in[9]), .ZN(n2988) );
  INVD1BWP12T U340 ( .I(write1_in[10]), .ZN(n3021) );
  INVD1BWP12T U341 ( .I(n3517), .ZN(n2981) );
  INVD1BWP12T U342 ( .I(write2_in[10]), .ZN(n3019) );
  INVD1BWP12T U343 ( .I(r0[11]), .ZN(n2893) );
  INVD1BWP12T U344 ( .I(write2_in[11]), .ZN(n2902) );
  INVD1BWP12T U345 ( .I(n3218), .ZN(n2982) );
  INVD1BWP12T U346 ( .I(n3219), .ZN(n2980) );
  INVD1BWP12T U347 ( .I(n3050), .ZN(n3055) );
  CKBD1BWP12T U348 ( .I(write1_in[17]), .Z(n3054) );
  CKBD1BWP12T U349 ( .I(write1_in[18]), .Z(n3060) );
  INVD1BWP12T U350 ( .I(n3094), .ZN(n3096) );
  CKBD1BWP12T U351 ( .I(write1_in[21]), .Z(n3098) );
  BUFFD2BWP12T U352 ( .I(n172), .Z(n3150) );
  INVD2BWP12T U353 ( .I(n3153), .ZN(n3211) );
  INVD1BWP12T U354 ( .I(r5[1]), .ZN(n1614) );
  INVD1BWP12T U355 ( .I(r11[1]), .ZN(n2802) );
  INVD1BWP12T U356 ( .I(r9[2]), .ZN(n2855) );
  INVD1BWP12T U357 ( .I(r7[2]), .ZN(n1672) );
  INVD1BWP12T U358 ( .I(r9[10]), .ZN(n3017) );
  INVD2BWP12T U359 ( .I(n1837), .ZN(n1873) );
  INVD2BWP12T U360 ( .I(n618), .ZN(n3417) );
  ND2D8BWP12T U361 ( .A1(n193), .A2(n861), .ZN(n3436) );
  ND2D1BWP12T U362 ( .A1(n577), .A2(n576), .ZN(n2167) );
  ND2D1BWP12T U363 ( .A1(n3275), .A2(n3246), .ZN(n577) );
  ND2D1BWP12T U364 ( .A1(n3275), .A2(n3231), .ZN(n354) );
  ND2D1BWP12T U365 ( .A1(n583), .A2(n582), .ZN(n2391) );
  ND2D1BWP12T U366 ( .A1(n3275), .A2(n3519), .ZN(n583) );
  ND2D1BWP12T U367 ( .A1(n573), .A2(n572), .ZN(n2647) );
  ND2D1BWP12T U368 ( .A1(n3275), .A2(n3517), .ZN(n573) );
  ND2D1BWP12T U369 ( .A1(n590), .A2(n589), .ZN(n2519) );
  ND2D1BWP12T U370 ( .A1(n3275), .A2(n3518), .ZN(n590) );
  ND2D1BWP12T U371 ( .A1(n575), .A2(n574), .ZN(n2295) );
  ND2D1BWP12T U372 ( .A1(n3275), .A2(n3522), .ZN(n575) );
  NR2D1BWP12T U373 ( .A1(n570), .A2(reset), .ZN(n3517) );
  NR2D1BWP12T U374 ( .A1(n578), .A2(reset), .ZN(n3519) );
  ND3D1BWP12T U375 ( .A1(n1746), .A2(n1745), .A3(n1744), .ZN(n2189) );
  ND3D1BWP12T U376 ( .A1(n1739), .A2(n3289), .A3(n1738), .ZN(n1746) );
  ND2D1BWP12T U377 ( .A1(n599), .A2(n598), .ZN(n2263) );
  ND2D1BWP12T U378 ( .A1(n3275), .A2(n3521), .ZN(n599) );
  ND2D1BWP12T U379 ( .A1(n3275), .A2(n3184), .ZN(n357) );
  AN2D1BWP12T U380 ( .A1(next_cpsr_in[3]), .A2(n3532), .Z(cpsrin[3]) );
  ND2D1BWP12T U381 ( .A1(n3247), .A2(n3184), .ZN(n1126) );
  ND2D1BWP12T U382 ( .A1(n3275), .A2(n3259), .ZN(n3263) );
  ND2D1BWP12T U383 ( .A1(n549), .A2(n548), .ZN(n2294) );
  ND2D1BWP12T U384 ( .A1(n553), .A2(n552), .ZN(n2326) );
  ND2D1BWP12T U385 ( .A1(n3275), .A2(n3269), .ZN(n3273) );
  ND2D1BWP12T U386 ( .A1(n3275), .A2(n3264), .ZN(n3268) );
  ND2D1BWP12T U387 ( .A1(n3275), .A2(n3274), .ZN(n3279) );
  ND2D1BWP12T U388 ( .A1(n3275), .A2(n3254), .ZN(n3258) );
  ND2D1BWP12T U389 ( .A1(n3226), .A2(n3518), .ZN(n3225) );
  ND2D1BWP12T U390 ( .A1(n559), .A2(n558), .ZN(n2550) );
  ND2D1BWP12T U391 ( .A1(n567), .A2(n566), .ZN(n2551) );
  ND2D1BWP12T U392 ( .A1(n3275), .A2(n3515), .ZN(n567) );
  ND2D1BWP12T U393 ( .A1(n565), .A2(n564), .ZN(n2582) );
  ND2D1BWP12T U394 ( .A1(n569), .A2(n568), .ZN(n2583) );
  ND2D1BWP12T U395 ( .A1(n3275), .A2(n3516), .ZN(n569) );
  ND2D1BWP12T U396 ( .A1(n3247), .A2(n3231), .ZN(n3235) );
  OAI22D1BWP12T U397 ( .A1(n3406), .A2(n2997), .B1(n2931), .B2(n3444), .ZN(
        n1358) );
  OAI22D1BWP12T U398 ( .A1(n1587), .A2(n1233), .B1(n1232), .B2(n1895), .ZN(
        n1234) );
  ND2D1BWP12T U399 ( .A1(n1907), .A2(immediate2_in[8]), .ZN(n845) );
  AOI211D1BWP12T U400 ( .A1(n1668), .A2(immediate2_in[31]), .B(n1090), .C(
        n1089), .ZN(n1091) );
  OAI22D1BWP12T U401 ( .A1(n1787), .A2(n1577), .B1(n1621), .B2(n784), .ZN(n789) );
  CKBD1BWP12T U402 ( .I(write1_in[27]), .Z(n172) );
  OAI22D1BWP12T U403 ( .A1(n3390), .A2(n2903), .B1(n2904), .B2(n3442), .ZN(
        n1363) );
  OAI22D1BWP12T U404 ( .A1(n1887), .A2(n2722), .B1(n161), .B2(n1446), .ZN(
        n1450) );
  ND2D1BWP12T U405 ( .A1(n1907), .A2(immediate2_in[23]), .ZN(n813) );
  ND2D1BWP12T U406 ( .A1(n1907), .A2(immediate2_in[26]), .ZN(n1244) );
  ND2D1BWP12T U407 ( .A1(n1907), .A2(immediate2_in[17]), .ZN(n448) );
  NR2D1BWP12T U408 ( .A1(n1564), .A2(n3357), .ZN(n1089) );
  OAI22D1BWP12T U409 ( .A1(n1911), .A2(n815), .B1(n1519), .B2(n1757), .ZN(n817) );
  OAI22D1BWP12T U410 ( .A1(n3452), .A2(n1447), .B1(n3393), .B2(n2722), .ZN(
        n236) );
  OAI22D1BWP12T U411 ( .A1(n3416), .A2(n378), .B1(n3436), .B2(n194), .ZN(n211)
         );
  OAI22D1BWP12T U412 ( .A1(n3452), .A2(n384), .B1(n3393), .B2(n2062), .ZN(n209) );
  OAI22D1BWP12T U413 ( .A1(n3416), .A2(n1453), .B1(n3436), .B2(n231), .ZN(n238) );
  OAI22D1BWP12T U414 ( .A1(n3444), .A2(n1444), .B1(n1837), .B2(n1446), .ZN(
        n241) );
  OAI22D1BWP12T U415 ( .A1(n3416), .A2(n1243), .B1(n3436), .B2(n339), .ZN(n346) );
  OAI22D1BWP12T U416 ( .A1(n1887), .A2(n604), .B1(n161), .B2(n606), .ZN(n436)
         );
  OR2XD1BWP12T U417 ( .A1(n1564), .A2(n610), .Z(n443) );
  INR2D1BWP12T U418 ( .A1(r2[4]), .B1(n3432), .ZN(n737) );
  OAI22D1BWP12T U419 ( .A1(n3416), .A2(n2697), .B1(n3436), .B2(n2696), .ZN(
        n783) );
  OAI22D1BWP12T U420 ( .A1(n3452), .A2(n1591), .B1(n3393), .B2(n1588), .ZN(
        n781) );
  ND2D1BWP12T U421 ( .A1(n1839), .A2(r7[24]), .ZN(n787) );
  INR2D1BWP12T U422 ( .A1(r5[24]), .B1(n1837), .ZN(n785) );
  OAI22D1BWP12T U423 ( .A1(n1663), .A2(n1762), .B1(n1975), .B2(n1592), .ZN(
        n821) );
  AOI21D1BWP12T U424 ( .A1(n1892), .A2(r0[8]), .B(n827), .ZN(n837) );
  ND2D1BWP12T U425 ( .A1(n1900), .A2(r9[8]), .ZN(n829) );
  INR2D1BWP12T U426 ( .A1(r3[8]), .B1(n1896), .ZN(n832) );
  ND2D1BWP12T U427 ( .A1(n1526), .A2(tmp1[8]), .ZN(n840) );
  OAI22D1BWP12T U428 ( .A1(n3436), .A2(n934), .B1(n3416), .B2(n1320), .ZN(n941) );
  OR2XD1BWP12T U429 ( .A1(n1564), .A2(n2050), .Z(n1003) );
  OAI22D1BWP12T U430 ( .A1(n1587), .A2(n1046), .B1(n1724), .B2(n1016), .ZN(
        n1017) );
  ND2D1BWP12T U431 ( .A1(n1853), .A2(r4[13]), .ZN(n1060) );
  OAI21D1BWP12T U432 ( .A1(n3442), .A2(n1046), .B(n1045), .ZN(n1059) );
  NR2D1BWP12T U433 ( .A1(n1428), .A2(n1053), .ZN(n1054) );
  AOI22D1BWP12T U434 ( .A1(n1575), .A2(pc_out[26]), .B1(n1915), .B2(r6[26]), 
        .ZN(n1248) );
  AOI22D1BWP12T U435 ( .A1(n1532), .A2(pc_out[19]), .B1(r6[19]), .B2(n1915), 
        .ZN(n1337) );
  NR2D1BWP12T U436 ( .A1(n3432), .A2(n2908), .ZN(n1353) );
  OAI22D1BWP12T U437 ( .A1(n2905), .A2(n3387), .B1(n3436), .B2(n2906), .ZN(
        n1362) );
  OAI22D1BWP12T U438 ( .A1(n3402), .A2(n3017), .B1(n2975), .B2(n3452), .ZN(
        n1406) );
  INR2D1BWP12T U439 ( .A1(r9[6]), .B1(n3402), .ZN(n1423) );
  OAI22D1BWP12T U440 ( .A1(n1553), .A2(n1448), .B1(n1447), .B2(n1592), .ZN(
        n1449) );
  ND2D1BWP12T U441 ( .A1(n1567), .A2(immediate2_in[27]), .ZN(n1458) );
  OAI21D1BWP12T U442 ( .A1(n1663), .A2(n1493), .B(n1492), .ZN(n1494) );
  AOI22D1BWP12T U443 ( .A1(n1571), .A2(r8[1]), .B1(tmp1[1]), .B2(n1526), .ZN(
        n1521) );
  INR2D1BWP12T U444 ( .A1(r7[20]), .B1(n3444), .ZN(n1854) );
  ND2D1BWP12T U445 ( .A1(n3418), .A2(r11[20]), .ZN(n1879) );
  NR2D1BWP12T U446 ( .A1(n3442), .A2(n3441), .ZN(n3457) );
  NR3D1BWP12T U447 ( .A1(n1868), .A2(n1867), .A3(n1866), .ZN(n1886) );
  TPNR3D2BWP12T U448 ( .A1(n1496), .A2(n1495), .A3(n1494), .ZN(n1506) );
  OAI21D1BWP12T U449 ( .A1(n841), .A2(n2905), .B(n840), .ZN(n842) );
  ND2D1BWP12T U450 ( .A1(n1355), .A2(n1354), .ZN(n1360) );
  ND3D1BWP12T U451 ( .A1(n1004), .A2(n1003), .A3(n1002), .ZN(n1012) );
  ND3D1BWP12T U452 ( .A1(n445), .A2(n444), .A3(n443), .ZN(n452) );
  INVD1BWP12T U453 ( .I(r6[10]), .ZN(n158) );
  ND3D1BWP12T U454 ( .A1(n1337), .A2(n1336), .A3(n185), .ZN(n1338) );
  ND2D1BWP12T U455 ( .A1(n1085), .A2(n1084), .ZN(n1086) );
  ND3D1BWP12T U456 ( .A1(n814), .A2(n179), .A3(n813), .ZN(n819) );
  NR2D1BWP12T U457 ( .A1(n1419), .A2(n1418), .ZN(n1420) );
  NR2D1BWP12T U458 ( .A1(n437), .A2(n436), .ZN(n438) );
  IND2D1BWP12T U459 ( .A1(n817), .B1(n816), .ZN(n818) );
  ND2D1BWP12T U460 ( .A1(n1399), .A2(n1398), .ZN(n1405) );
  TPNR2D1BWP12T U461 ( .A1(n1081), .A2(n1080), .ZN(n1093) );
  TPNR2D1BWP12T U462 ( .A1(n1052), .A2(n1051), .ZN(n1057) );
  NR2D1BWP12T U463 ( .A1(n1280), .A2(n1279), .ZN(n1287) );
  IND2D1BWP12T U464 ( .A1(n1455), .B1(n1454), .ZN(n1461) );
  ND2D1BWP12T U465 ( .A1(n1144), .A2(n1143), .ZN(n1151) );
  NR2D1BWP12T U466 ( .A1(n1285), .A2(n1284), .ZN(n1286) );
  NR2D2BWP12T U467 ( .A1(n1242), .A2(n1241), .ZN(n1254) );
  NR2D1BWP12T U468 ( .A1(n1872), .A2(n1871), .ZN(n1875) );
  NR2D1BWP12T U469 ( .A1(n831), .A2(n830), .ZN(n834) );
  NR2D1BWP12T U470 ( .A1(n1855), .A2(n1854), .ZN(n1856) );
  OR2XD1BWP12T U471 ( .A1(n1488), .A2(n1487), .Z(n1496) );
  IND2D1BWP12T U472 ( .A1(n1249), .B1(n1248), .ZN(n1251) );
  INVD1BWP12T U473 ( .I(n1020), .ZN(n1021) );
  IND2D1BWP12T U474 ( .A1(n439), .B1(n438), .ZN(n442) );
  OR2XD1BWP12T U475 ( .A1(n1078), .A2(n1077), .Z(n1081) );
  ND2D1BWP12T U476 ( .A1(n1532), .A2(pc_out[1]), .ZN(n1515) );
  INVD1BWP12T U477 ( .I(n155), .ZN(n156) );
  AN2XD2BWP12T U478 ( .A1(n169), .A2(n170), .Z(n1009) );
  INVD1BWP12T U479 ( .I(n829), .ZN(n830) );
  INVD1BWP12T U480 ( .I(n785), .ZN(n786) );
  INVD1BWP12T U481 ( .I(n1152), .ZN(n1153) );
  INVD1BWP12T U482 ( .I(n1013), .ZN(n1014) );
  INVD1BWP12T U483 ( .I(n737), .ZN(n738) );
  AOI22D0BWP12T U484 ( .A1(r9[1]), .A2(n3063), .B1(n3064), .B2(r12[1]), .ZN(n1) );
  AOI22D0BWP12T U485 ( .A1(pc_out[1]), .A2(n3061), .B1(r11[1]), .B2(n2994), 
        .ZN(n2) );
  AOI22D0BWP12T U486 ( .A1(r1[1]), .A2(n3074), .B1(n3075), .B2(r5[1]), .ZN(n3)
         );
  AOI22D0BWP12T U487 ( .A1(r7[1]), .A2(n3076), .B1(n3077), .B2(r6[1]), .ZN(n4)
         );
  AOI22D0BWP12T U488 ( .A1(r3[1]), .A2(n3078), .B1(n3079), .B2(r2[1]), .ZN(n5)
         );
  AOI22D0BWP12T U489 ( .A1(r4[1]), .A2(n3080), .B1(n3081), .B2(r0[1]), .ZN(n6)
         );
  ND4D0BWP12T U490 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(n7) );
  OAI22D0BWP12T U491 ( .A1(n3042), .A2(n2831), .B1(n2832), .B2(n3069), .ZN(n8)
         );
  MOAI22D0BWP12T U492 ( .A1(n3066), .A2(n2829), .B1(n3073), .B2(r8[1]), .ZN(n9) );
  AOI211D0BWP12T U493 ( .A1(n3086), .A2(n7), .B(n8), .C(n9), .ZN(n10) );
  ND3D0BWP12T U494 ( .A1(n1), .A2(n2), .A3(n10), .ZN(regD_out[1]) );
  AOI22D0BWP12T U495 ( .A1(n[3560]), .A2(n3464), .B1(lr[20]), .B2(n3473), .ZN(
        n11) );
  AOI22D0BWP12T U496 ( .A1(r6[20]), .A2(n2770), .B1(r5[20]), .B2(n3481), .ZN(
        n12) );
  AOI22D0BWP12T U497 ( .A1(r7[20]), .A2(n3482), .B1(r4[20]), .B2(n2757), .ZN(
        n13) );
  AOI22D0BWP12T U498 ( .A1(r2[20]), .A2(n3483), .B1(r1[20]), .B2(n3484), .ZN(
        n14) );
  AOI22D0BWP12T U499 ( .A1(r0[20]), .A2(n3486), .B1(r3[20]), .B2(n3485), .ZN(
        n15) );
  ND4D0BWP12T U500 ( .A1(n12), .A2(n13), .A3(n14), .A4(n15), .ZN(n16) );
  AOI22D0BWP12T U501 ( .A1(r12[20]), .A2(n3479), .B1(n3492), .B2(n16), .ZN(n17) );
  CKND0BWP12T U502 ( .I(pc_out[20]), .ZN(n18) );
  MOAI22D0BWP12T U503 ( .A1(n2806), .A2(n18), .B1(r9[20]), .B2(n3475), .ZN(n19) );
  OAI22D0BWP12T U504 ( .A1(n2710), .A2(n2803), .B1(n2709), .B2(n2800), .ZN(n20) );
  AOI211D0BWP12T U505 ( .A1(r10[20]), .A2(n2810), .B(n19), .C(n20), .ZN(n21)
         );
  ND3D0BWP12T U506 ( .A1(n11), .A2(n17), .A3(n21), .ZN(regC_out[20]) );
  AO222D0BWP12T U507 ( .A1(n3274), .A2(n3108), .B1(n3276), .B2(write2_in[26]), 
        .C1(r6[26]), .C2(n3277), .Z(n2450) );
  AO222D0BWP12T U508 ( .A1(n3259), .A2(n3054), .B1(n3260), .B2(write2_in[17]), 
        .C1(lr[17]), .C2(n3261), .Z(n2217) );
  AO222D0BWP12T U509 ( .A1(n3254), .A2(write1_in[15]), .B1(n3255), .B2(
        write2_in[15]), .C1(r5[15]), .C2(n3256), .Z(n2471) );
  AO222D0BWP12T U510 ( .A1(n3517), .A2(write1_in[12]), .B1(write2_in[12]), 
        .B2(n3218), .C1(r0[12]), .C2(n3219), .Z(n2628) );
  AO222D0BWP12T U511 ( .A1(n3259), .A2(n3098), .B1(n3260), .B2(write2_in[21]), 
        .C1(lr[21]), .C2(n3261), .Z(n2221) );
  AO222D0BWP12T U512 ( .A1(n3259), .A2(n3060), .B1(write2_in[18]), .B2(n3260), 
        .C1(lr[18]), .C2(n3261), .Z(n2218) );
  AO222D0BWP12T U513 ( .A1(n3184), .A2(write1_in[14]), .B1(n3185), .B2(
        write2_in[14]), .C1(n[3566]), .C2(n3186), .Z(spin[14]) );
  AO222D0BWP12T U514 ( .A1(n3246), .A2(n3055), .B1(write2_in[16]), .B2(n1947), 
        .C1(tmp1[16]), .C2(n1946), .Z(n2152) );
  AO222D0BWP12T U515 ( .A1(n3246), .A2(n3096), .B1(tmp1[19]), .B2(n1946), .C1(
        n1947), .C2(write2_in[19]), .Z(n2155) );
  AO222D0BWP12T U516 ( .A1(n3246), .A2(n3095), .B1(tmp1[20]), .B2(n1946), .C1(
        n1947), .C2(write2_in[20]), .Z(n2156) );
  AO222D0BWP12T U517 ( .A1(n3246), .A2(n3282), .B1(tmp1[22]), .B2(n1946), .C1(
        n1947), .C2(write2_in[22]), .Z(n2158) );
  AO222D0BWP12T U518 ( .A1(n3246), .A2(write1_in[23]), .B1(tmp1[23]), .B2(
        n1946), .C1(n1947), .C2(write2_in[23]), .Z(n2159) );
  AO222D0BWP12T U519 ( .A1(n3246), .A2(n3097), .B1(tmp1[24]), .B2(n1946), .C1(
        n1947), .C2(write2_in[24]), .Z(n2160) );
  AO222D0BWP12T U520 ( .A1(n3246), .A2(n3113), .B1(tmp1[25]), .B2(n1946), .C1(
        n1947), .C2(write2_in[25]), .Z(n2161) );
  AOI22D0BWP12T U521 ( .A1(r12[2]), .A2(n3064), .B1(n2994), .B2(r11[2]), .ZN(
        n22) );
  AOI22D0BWP12T U522 ( .A1(pc_out[2]), .A2(n3061), .B1(n3062), .B2(lr[2]), 
        .ZN(n23) );
  AOI22D0BWP12T U523 ( .A1(r1[2]), .A2(n3074), .B1(n3075), .B2(r5[2]), .ZN(n24) );
  AOI22D0BWP12T U524 ( .A1(r7[2]), .A2(n3076), .B1(n3077), .B2(r6[2]), .ZN(n25) );
  AOI22D0BWP12T U525 ( .A1(r3[2]), .A2(n3078), .B1(n3079), .B2(r2[2]), .ZN(n26) );
  AOI22D0BWP12T U526 ( .A1(r4[2]), .A2(n3080), .B1(n3081), .B2(r0[2]), .ZN(n27) );
  ND4D0BWP12T U527 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(n28) );
  OAI22D0BWP12T U528 ( .A1(n2886), .A2(n2855), .B1(n2856), .B2(n3069), .ZN(n29) );
  MOAI22D0BWP12T U529 ( .A1(n3066), .A2(n2854), .B1(n3073), .B2(r8[2]), .ZN(
        n30) );
  AOI211D0BWP12T U530 ( .A1(n3086), .A2(n28), .B(n29), .C(n30), .ZN(n31) );
  ND3D0BWP12T U531 ( .A1(n22), .A2(n23), .A3(n31), .ZN(regD_out[2]) );
  AO222D0BWP12T U532 ( .A1(n3522), .A2(n3054), .B1(r11[17]), .B2(n3201), .C1(
        n3202), .C2(write2_in[17]), .Z(n2281) );
  AO222D0BWP12T U533 ( .A1(n3254), .A2(n3098), .B1(n3255), .B2(write2_in[21]), 
        .C1(r5[21]), .C2(n3256), .Z(n2477) );
  AO222D0BWP12T U534 ( .A1(n3231), .A2(n3060), .B1(write2_in[18]), .B2(n3232), 
        .C1(r1[18]), .C2(n3233), .Z(n2602) );
  AO222D0BWP12T U535 ( .A1(n3521), .A2(write1_in[12]), .B1(write2_in[12]), 
        .B2(n3227), .C1(r12[12]), .C2(n3228), .Z(n2244) );
  AO222D0BWP12T U536 ( .A1(n3246), .A2(write1_in[14]), .B1(tmp1[14]), .B2(
        n1946), .C1(n1947), .C2(write2_in[14]), .Z(n2150) );
  AO222D0BWP12T U537 ( .A1(n3246), .A2(write1_in[15]), .B1(tmp1[15]), .B2(
        n1946), .C1(n1947), .C2(write2_in[15]), .Z(n2151) );
  AO222D0BWP12T U538 ( .A1(n3246), .A2(n3108), .B1(tmp1[26]), .B2(n1946), .C1(
        n1947), .C2(write2_in[26]), .Z(n2162) );
  AO222D0BWP12T U539 ( .A1(n3184), .A2(n3055), .B1(write2_in[16]), .B2(n3185), 
        .C1(n[3564]), .C2(n3186), .Z(spin[16]) );
  AO222D0BWP12T U540 ( .A1(n3184), .A2(n3096), .B1(n3185), .B2(write2_in[19]), 
        .C1(n[3561]), .C2(n3186), .Z(spin[19]) );
  AO222D0BWP12T U541 ( .A1(n3184), .A2(n3095), .B1(n3185), .B2(write2_in[20]), 
        .C1(n[3560]), .C2(n3186), .Z(spin[20]) );
  AO222D0BWP12T U542 ( .A1(n3184), .A2(n3282), .B1(n3185), .B2(write2_in[22]), 
        .C1(n[3558]), .C2(n3186), .Z(spin[22]) );
  AO222D0BWP12T U543 ( .A1(n3184), .A2(write1_in[23]), .B1(n3185), .B2(
        write2_in[23]), .C1(n[3557]), .C2(n3186), .Z(spin[23]) );
  AO222D0BWP12T U544 ( .A1(n3184), .A2(n3097), .B1(n3185), .B2(write2_in[24]), 
        .C1(n[3556]), .C2(n3186), .Z(spin[24]) );
  AO222D0BWP12T U545 ( .A1(n3184), .A2(n3113), .B1(n3185), .B2(write2_in[25]), 
        .C1(n[3555]), .C2(n3186), .Z(spin[25]) );
  OAI22D0BWP12T U546 ( .A1(n2850), .A2(n2920), .B1(n3042), .B2(n2851), .ZN(n32) );
  OAI22D0BWP12T U547 ( .A1(n3068), .A2(n2852), .B1(n2853), .B2(n3069), .ZN(n33) );
  AOI211D0BWP12T U548 ( .A1(n3029), .A2(r10[3]), .B(n32), .C(n33), .ZN(n34) );
  AOI22D0BWP12T U549 ( .A1(pc_out[3]), .A2(n3061), .B1(r9[3]), .B2(n3063), 
        .ZN(n35) );
  AOI22D0BWP12T U550 ( .A1(r1[3]), .A2(n3074), .B1(n3075), .B2(r5[3]), .ZN(n36) );
  AOI22D0BWP12T U551 ( .A1(r7[3]), .A2(n3076), .B1(n3077), .B2(r6[3]), .ZN(n37) );
  AOI22D0BWP12T U552 ( .A1(r3[3]), .A2(n3078), .B1(n3079), .B2(r2[3]), .ZN(n38) );
  AOI22D0BWP12T U553 ( .A1(r4[3]), .A2(n3080), .B1(n3081), .B2(r0[3]), .ZN(n39) );
  ND4D0BWP12T U554 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n40) );
  AOI22D0BWP12T U555 ( .A1(r8[3]), .A2(n3073), .B1(n3086), .B2(n40), .ZN(n41)
         );
  ND3D0BWP12T U556 ( .A1(n34), .A2(n35), .A3(n41), .ZN(regD_out[3]) );
  AO222D0BWP12T U557 ( .A1(n3520), .A2(n3054), .B1(write2_in[17]), .B2(n3197), 
        .C1(r10[17]), .C2(n3198), .Z(n2313) );
  AO222D0BWP12T U558 ( .A1(n3521), .A2(n3060), .B1(write2_in[18]), .B2(n3227), 
        .C1(r12[18]), .C2(n3228), .Z(n2250) );
  AO222D0BWP12T U559 ( .A1(n3246), .A2(write1_in[12]), .B1(write2_in[12]), 
        .B2(n1947), .C1(tmp1[12]), .C2(n1946), .Z(n2148) );
  AO222D0BWP12T U560 ( .A1(n3246), .A2(n3098), .B1(tmp1[21]), .B2(n1946), .C1(
        n1947), .C2(write2_in[21]), .Z(n2157) );
  AO222D0BWP12T U561 ( .A1(n3184), .A2(n177), .B1(n3185), .B2(write2_in[15]), 
        .C1(n[3565]), .C2(n3186), .Z(spin[15]) );
  AO222D0BWP12T U562 ( .A1(n3184), .A2(n3108), .B1(n3185), .B2(write2_in[26]), 
        .C1(n[3554]), .C2(n3186), .Z(spin[26]) );
  AO222D0BWP12T U563 ( .A1(n3259), .A2(write1_in[14]), .B1(n3260), .B2(
        write2_in[14]), .C1(lr[14]), .C2(n3261), .Z(n2214) );
  AO222D0BWP12T U564 ( .A1(n3259), .A2(n3055), .B1(write2_in[16]), .B2(n3260), 
        .C1(lr[16]), .C2(n3261), .Z(n2216) );
  AO222D0BWP12T U565 ( .A1(n3259), .A2(n3096), .B1(n3260), .B2(write2_in[19]), 
        .C1(lr[19]), .C2(n3261), .Z(n2219) );
  AO222D0BWP12T U566 ( .A1(n3259), .A2(n3095), .B1(n3260), .B2(write2_in[20]), 
        .C1(lr[20]), .C2(n3261), .Z(n2220) );
  AO222D0BWP12T U567 ( .A1(n3259), .A2(n3282), .B1(n3260), .B2(write2_in[22]), 
        .C1(lr[22]), .C2(n3261), .Z(n2222) );
  AO222D0BWP12T U568 ( .A1(n3259), .A2(write1_in[23]), .B1(n3260), .B2(
        write2_in[23]), .C1(lr[23]), .C2(n3261), .Z(n2223) );
  AO222D0BWP12T U569 ( .A1(n3259), .A2(n3097), .B1(n3260), .B2(write2_in[24]), 
        .C1(lr[24]), .C2(n3261), .Z(n2224) );
  AO222D0BWP12T U570 ( .A1(n3259), .A2(n3113), .B1(n3260), .B2(write2_in[25]), 
        .C1(lr[25]), .C2(n3261), .Z(n2225) );
  AOI22D0BWP12T U571 ( .A1(r12[4]), .A2(n3064), .B1(n2994), .B2(r11[4]), .ZN(
        n42) );
  AOI22D0BWP12T U572 ( .A1(pc_out[4]), .A2(n3061), .B1(n3037), .B2(n[3576]), 
        .ZN(n43) );
  AOI22D0BWP12T U573 ( .A1(r1[4]), .A2(n3074), .B1(n3075), .B2(r5[4]), .ZN(n44) );
  AOI22D0BWP12T U574 ( .A1(r7[4]), .A2(n3076), .B1(n3077), .B2(r6[4]), .ZN(n45) );
  AOI22D0BWP12T U575 ( .A1(r3[4]), .A2(n3078), .B1(n3079), .B2(r2[4]), .ZN(n46) );
  AOI22D0BWP12T U576 ( .A1(r4[4]), .A2(n3080), .B1(n3081), .B2(r0[4]), .ZN(n47) );
  ND4D0BWP12T U577 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(n48) );
  OAI22D0BWP12T U578 ( .A1(n2842), .A2(n2886), .B1(n3042), .B2(n2843), .ZN(n49) );
  MOAI22D0BWP12T U579 ( .A1(n3066), .A2(n2841), .B1(n3073), .B2(r8[4]), .ZN(
        n50) );
  AOI211D0BWP12T U580 ( .A1(n3086), .A2(n48), .B(n49), .C(n50), .ZN(n51) );
  ND3D0BWP12T U581 ( .A1(n42), .A2(n43), .A3(n51), .ZN(regD_out[4]) );
  AO222D0BWP12T U582 ( .A1(n3264), .A2(n3054), .B1(n3265), .B2(write2_in[17]), 
        .C1(r7[17]), .C2(n3266), .Z(n2409) );
  AO222D0BWP12T U583 ( .A1(n3246), .A2(n3060), .B1(write2_in[18]), .B2(n1947), 
        .C1(tmp1[18]), .C2(n1946), .Z(n2154) );
  CKND0BWP12T U584 ( .I(write2_in[12]), .ZN(n52) );
  AOI21D0BWP12T U585 ( .A1(n[3568]), .A2(n3186), .B(reset), .ZN(n53) );
  CKND2D0BWP12T U586 ( .A1(n3184), .A2(write1_in[12]), .ZN(n54) );
  OAI211D0BWP12T U587 ( .A1(n2993), .A2(n52), .B(n53), .C(n54), .ZN(spin[12])
         );
  AO222D0BWP12T U588 ( .A1(n3184), .A2(n3098), .B1(n3185), .B2(write2_in[21]), 
        .C1(n[3559]), .C2(n3186), .Z(spin[21]) );
  AO222D0BWP12T U589 ( .A1(n3259), .A2(n177), .B1(n3260), .B2(write2_in[15]), 
        .C1(lr[15]), .C2(n3261), .Z(n2215) );
  AO222D0BWP12T U590 ( .A1(n3259), .A2(n3108), .B1(n3260), .B2(write2_in[26]), 
        .C1(lr[26]), .C2(n3261), .Z(n2226) );
  AO222D0BWP12T U591 ( .A1(n3521), .A2(write1_in[14]), .B1(n3227), .B2(
        write2_in[14]), .C1(r12[14]), .C2(n3228), .Z(n2246) );
  AO222D0BWP12T U592 ( .A1(n3521), .A2(n3055), .B1(write2_in[16]), .B2(n3227), 
        .C1(r12[16]), .C2(n3228), .Z(n2248) );
  AO222D0BWP12T U593 ( .A1(n3521), .A2(n3096), .B1(n3227), .B2(write2_in[19]), 
        .C1(r12[19]), .C2(n3228), .Z(n2251) );
  AO222D0BWP12T U594 ( .A1(n3521), .A2(n3095), .B1(n3227), .B2(write2_in[20]), 
        .C1(r12[20]), .C2(n3228), .Z(n2252) );
  AO222D0BWP12T U595 ( .A1(n3521), .A2(n3282), .B1(n3227), .B2(write2_in[22]), 
        .C1(r12[22]), .C2(n3228), .Z(n2254) );
  AO222D0BWP12T U596 ( .A1(n3521), .A2(write1_in[23]), .B1(n3227), .B2(
        write2_in[23]), .C1(r12[23]), .C2(n3228), .Z(n2255) );
  AO222D0BWP12T U597 ( .A1(n3521), .A2(n3097), .B1(n3227), .B2(write2_in[24]), 
        .C1(r12[24]), .C2(n3228), .Z(n2256) );
  AO222D0BWP12T U598 ( .A1(n3521), .A2(n3113), .B1(n3227), .B2(write2_in[25]), 
        .C1(r12[25]), .C2(n3228), .Z(n2257) );
  AOI22D0BWP12T U599 ( .A1(r9[5]), .A2(n3063), .B1(n3064), .B2(r12[5]), .ZN(
        n55) );
  AOI22D0BWP12T U600 ( .A1(pc_out[5]), .A2(n3061), .B1(n3062), .B2(lr[5]), 
        .ZN(n56) );
  AOI22D0BWP12T U601 ( .A1(r1[5]), .A2(n3074), .B1(n3075), .B2(r5[5]), .ZN(n57) );
  AOI22D0BWP12T U602 ( .A1(r7[5]), .A2(n3076), .B1(n3077), .B2(r6[5]), .ZN(n58) );
  AOI22D0BWP12T U603 ( .A1(r3[5]), .A2(n3078), .B1(n3079), .B2(r2[5]), .ZN(n59) );
  AOI22D0BWP12T U604 ( .A1(r4[5]), .A2(n3080), .B1(n3081), .B2(r0[5]), .ZN(n60) );
  ND4D0BWP12T U605 ( .A1(n57), .A2(n58), .A3(n59), .A4(n60), .ZN(n61) );
  CKND0BWP12T U606 ( .I(n[3575]), .ZN(n62) );
  OAI22D0BWP12T U607 ( .A1(n3069), .A2(n62), .B1(n3068), .B2(n2869), .ZN(n63)
         );
  MOAI22D0BWP12T U608 ( .A1(n3066), .A2(n2868), .B1(n3073), .B2(r8[5]), .ZN(
        n64) );
  AOI211D0BWP12T U609 ( .A1(n3086), .A2(n61), .B(n63), .C(n64), .ZN(n65) );
  ND3D0BWP12T U610 ( .A1(n55), .A2(n56), .A3(n65), .ZN(regD_out[5]) );
  AO222D0BWP12T U611 ( .A1(n3246), .A2(n3054), .B1(tmp1[17]), .B2(n1946), .C1(
        n1947), .C2(write2_in[17]), .Z(n2153) );
  MOAI22D0BWP12T U612 ( .A1(n3112), .A2(n3111), .B1(n3112), .B2(n3111), .ZN(
        n66) );
  AOI22D0BWP12T U613 ( .A1(pc_out[14]), .A2(n3498), .B1(n3499), .B2(
        next_pc_in[14]), .ZN(n67) );
  OAI21D0BWP12T U614 ( .A1(n3497), .A2(n66), .B(n67), .ZN(n2182) );
  AO222D0BWP12T U615 ( .A1(n3184), .A2(n3060), .B1(write2_in[18]), .B2(n3185), 
        .C1(n[3562]), .C2(n3186), .Z(spin[18]) );
  AO222D0BWP12T U616 ( .A1(n3259), .A2(write1_in[12]), .B1(write2_in[12]), 
        .B2(n3260), .C1(lr[12]), .C2(n3261), .Z(n2212) );
  AO222D0BWP12T U617 ( .A1(n3521), .A2(write1_in[15]), .B1(n3227), .B2(
        write2_in[15]), .C1(r12[15]), .C2(n3228), .Z(n2247) );
  AO222D0BWP12T U618 ( .A1(n3521), .A2(n3098), .B1(n3227), .B2(write2_in[21]), 
        .C1(r12[21]), .C2(n3228), .Z(n2253) );
  AO222D0BWP12T U619 ( .A1(n3521), .A2(n3108), .B1(n3227), .B2(write2_in[26]), 
        .C1(r12[26]), .C2(n3228), .Z(n2258) );
  AO222D0BWP12T U620 ( .A1(n3522), .A2(write1_in[14]), .B1(r11[14]), .B2(n3201), .C1(n3202), .C2(write2_in[14]), .Z(n2278) );
  AO222D0BWP12T U621 ( .A1(n3522), .A2(n3055), .B1(r11[16]), .B2(n3201), .C1(
        write2_in[16]), .C2(n3202), .Z(n2280) );
  AO222D0BWP12T U622 ( .A1(n3522), .A2(n3096), .B1(r11[19]), .B2(n3201), .C1(
        n3202), .C2(write2_in[19]), .Z(n2283) );
  AO222D0BWP12T U623 ( .A1(n3522), .A2(n3095), .B1(r11[20]), .B2(n3201), .C1(
        n3202), .C2(write2_in[20]), .Z(n2284) );
  AO222D0BWP12T U624 ( .A1(n3522), .A2(n3099), .B1(r11[22]), .B2(n3201), .C1(
        n3202), .C2(write2_in[22]), .Z(n2286) );
  AO222D0BWP12T U625 ( .A1(n3522), .A2(write1_in[23]), .B1(r11[23]), .B2(n3201), .C1(n3202), .C2(write2_in[23]), .Z(n2287) );
  AO222D0BWP12T U626 ( .A1(n3522), .A2(n3097), .B1(r11[24]), .B2(n3201), .C1(
        n3202), .C2(write2_in[24]), .Z(n2288) );
  AO222D0BWP12T U627 ( .A1(n3522), .A2(n3113), .B1(r11[25]), .B2(n3201), .C1(
        n3202), .C2(write2_in[25]), .Z(n2289) );
  AOI22D0BWP12T U628 ( .A1(r12[6]), .A2(n3064), .B1(n2994), .B2(r11[6]), .ZN(
        n68) );
  AOI22D0BWP12T U629 ( .A1(lr[6]), .A2(n3062), .B1(n3037), .B2(n[3574]), .ZN(
        n69) );
  AOI22D0BWP12T U630 ( .A1(r1[6]), .A2(n3074), .B1(n3075), .B2(r5[6]), .ZN(n70) );
  AOI22D0BWP12T U631 ( .A1(r7[6]), .A2(n3076), .B1(n3077), .B2(r6[6]), .ZN(n71) );
  AOI22D0BWP12T U632 ( .A1(r3[6]), .A2(n3078), .B1(n3079), .B2(r2[6]), .ZN(n72) );
  AOI22D0BWP12T U633 ( .A1(r4[6]), .A2(n3080), .B1(n3081), .B2(r0[6]), .ZN(n73) );
  ND4D0BWP12T U634 ( .A1(n70), .A2(n71), .A3(n72), .A4(n73), .ZN(n74) );
  OAI22D0BWP12T U635 ( .A1(n2886), .A2(n2873), .B1(n2874), .B2(n3028), .ZN(n75) );
  MOAI22D0BWP12T U636 ( .A1(n3066), .A2(n1412), .B1(n3073), .B2(r8[6]), .ZN(
        n76) );
  AOI211D0BWP12T U637 ( .A1(n3086), .A2(n74), .B(n75), .C(n76), .ZN(n77) );
  ND3D0BWP12T U638 ( .A1(n68), .A2(n69), .A3(n77), .ZN(regD_out[6]) );
  AO222D0BWP12T U639 ( .A1(n3184), .A2(n3054), .B1(n3185), .B2(write2_in[17]), 
        .C1(n[3563]), .C2(n3186), .Z(spin[17]) );
  AO222D0BWP12T U640 ( .A1(n3522), .A2(write1_in[12]), .B1(r11[12]), .B2(n3201), .C1(write2_in[12]), .C2(n3202), .Z(n2276) );
  AO222D0BWP12T U641 ( .A1(n3522), .A2(write1_in[15]), .B1(r11[15]), .B2(n3201), .C1(n3202), .C2(write2_in[15]), .Z(n2279) );
  AO222D0BWP12T U642 ( .A1(n3522), .A2(n3060), .B1(r11[18]), .B2(n3201), .C1(
        write2_in[18]), .C2(n3202), .Z(n2282) );
  AO222D0BWP12T U643 ( .A1(n3522), .A2(n3098), .B1(r11[21]), .B2(n3201), .C1(
        n3202), .C2(write2_in[21]), .Z(n2285) );
  AO222D0BWP12T U644 ( .A1(n3522), .A2(n3108), .B1(r11[26]), .B2(n3201), .C1(
        n3202), .C2(write2_in[26]), .Z(n2290) );
  AO222D0BWP12T U645 ( .A1(n3520), .A2(write1_in[14]), .B1(write2_in[14]), 
        .B2(n3197), .C1(r10[14]), .C2(n3198), .Z(n2310) );
  AO222D0BWP12T U646 ( .A1(n3520), .A2(n3055), .B1(write2_in[16]), .B2(n3197), 
        .C1(r10[16]), .C2(n3198), .Z(n2312) );
  AO222D0BWP12T U647 ( .A1(n3520), .A2(n3096), .B1(write2_in[19]), .B2(n3197), 
        .C1(r10[19]), .C2(n3198), .Z(n2315) );
  AO222D0BWP12T U648 ( .A1(n3520), .A2(n3095), .B1(write2_in[20]), .B2(n3197), 
        .C1(r10[20]), .C2(n3198), .Z(n2316) );
  AO222D0BWP12T U649 ( .A1(n3520), .A2(n3099), .B1(write2_in[22]), .B2(n3197), 
        .C1(r10[22]), .C2(n3198), .Z(n2318) );
  AO222D0BWP12T U650 ( .A1(n3520), .A2(write1_in[23]), .B1(write2_in[23]), 
        .B2(n3197), .C1(r10[23]), .C2(n3198), .Z(n2319) );
  AO222D0BWP12T U651 ( .A1(n3520), .A2(n3097), .B1(write2_in[24]), .B2(n3197), 
        .C1(r10[24]), .C2(n3198), .Z(n2320) );
  AO222D0BWP12T U652 ( .A1(n3520), .A2(n3113), .B1(write2_in[25]), .B2(n3197), 
        .C1(r10[25]), .C2(n3198), .Z(n2321) );
  AOI22D0BWP12T U653 ( .A1(r12[7]), .A2(n3064), .B1(n2994), .B2(r11[7]), .ZN(
        n78) );
  AOI22D0BWP12T U654 ( .A1(pc_out[7]), .A2(n3061), .B1(n3062), .B2(lr[7]), 
        .ZN(n79) );
  AOI22D0BWP12T U655 ( .A1(r1[7]), .A2(n3074), .B1(n3075), .B2(r5[7]), .ZN(n80) );
  AOI22D0BWP12T U656 ( .A1(r7[7]), .A2(n3076), .B1(n3077), .B2(r6[7]), .ZN(n81) );
  AOI22D0BWP12T U657 ( .A1(r3[7]), .A2(n3078), .B1(n3079), .B2(r2[7]), .ZN(n82) );
  AOI22D0BWP12T U658 ( .A1(r4[7]), .A2(n3080), .B1(n3081), .B2(r0[7]), .ZN(n83) );
  ND4D0BWP12T U659 ( .A1(n80), .A2(n81), .A3(n82), .A4(n83), .ZN(n84) );
  OAI22D0BWP12T U660 ( .A1(n3024), .A2(n2860), .B1(n2861), .B2(n3069), .ZN(n85) );
  MOAI22D0BWP12T U661 ( .A1(n3066), .A2(n2859), .B1(n3063), .B2(r9[7]), .ZN(
        n86) );
  AOI211D0BWP12T U662 ( .A1(n3086), .A2(n84), .B(n85), .C(n86), .ZN(n87) );
  ND3D0BWP12T U663 ( .A1(n78), .A2(n79), .A3(n87), .ZN(regD_out[7]) );
  AO222D0BWP12T U664 ( .A1(n3521), .A2(n3054), .B1(n3227), .B2(write2_in[17]), 
        .C1(r12[17]), .C2(n3228), .Z(n2249) );
  AO222D0BWP12T U665 ( .A1(n3520), .A2(write1_in[12]), .B1(write2_in[12]), 
        .B2(n3197), .C1(r10[12]), .C2(n3198), .Z(n2308) );
  AO222D0BWP12T U666 ( .A1(n3520), .A2(write1_in[15]), .B1(write2_in[15]), 
        .B2(n3197), .C1(r10[15]), .C2(n3198), .Z(n2311) );
  AO222D0BWP12T U667 ( .A1(n3520), .A2(n3060), .B1(write2_in[18]), .B2(n3197), 
        .C1(r10[18]), .C2(n3198), .Z(n2314) );
  AO222D0BWP12T U668 ( .A1(n3520), .A2(n3098), .B1(write2_in[21]), .B2(n3197), 
        .C1(r10[21]), .C2(n3198), .Z(n2317) );
  AO222D0BWP12T U669 ( .A1(n3520), .A2(n3108), .B1(write2_in[26]), .B2(n3197), 
        .C1(r10[26]), .C2(n3198), .Z(n2322) );
  AO222D0BWP12T U670 ( .A1(n3269), .A2(write1_in[14]), .B1(n3270), .B2(
        write2_in[14]), .C1(r9[14]), .C2(n3271), .Z(n2342) );
  AO222D0BWP12T U671 ( .A1(n3269), .A2(n3055), .B1(write2_in[16]), .B2(n3270), 
        .C1(r9[16]), .C2(n3271), .Z(n2344) );
  AO222D0BWP12T U672 ( .A1(n3269), .A2(n3096), .B1(n3270), .B2(write2_in[19]), 
        .C1(r9[19]), .C2(n3271), .Z(n2347) );
  AO222D0BWP12T U673 ( .A1(n3269), .A2(n3095), .B1(n3270), .B2(write2_in[20]), 
        .C1(r9[20]), .C2(n3271), .Z(n2348) );
  AO222D0BWP12T U674 ( .A1(n3269), .A2(n3099), .B1(n3270), .B2(write2_in[22]), 
        .C1(r9[22]), .C2(n3271), .Z(n2350) );
  AO222D0BWP12T U675 ( .A1(n3269), .A2(write1_in[23]), .B1(n3270), .B2(
        write2_in[23]), .C1(r9[23]), .C2(n3271), .Z(n2351) );
  AO222D0BWP12T U676 ( .A1(n3269), .A2(n3097), .B1(n3270), .B2(write2_in[24]), 
        .C1(r9[24]), .C2(n3271), .Z(n2352) );
  AO222D0BWP12T U677 ( .A1(n3269), .A2(n3113), .B1(n3270), .B2(write2_in[25]), 
        .C1(r9[25]), .C2(n3271), .Z(n2353) );
  AOI22D0BWP12T U678 ( .A1(r9[8]), .A2(n3063), .B1(n3064), .B2(r12[8]), .ZN(
        n88) );
  AOI22D0BWP12T U679 ( .A1(r11[8]), .A2(n2994), .B1(n3037), .B2(n[3572]), .ZN(
        n89) );
  AOI22D0BWP12T U680 ( .A1(r1[8]), .A2(n3074), .B1(n3075), .B2(r5[8]), .ZN(n90) );
  AOI22D0BWP12T U681 ( .A1(r7[8]), .A2(n3076), .B1(n3077), .B2(r6[8]), .ZN(n91) );
  AOI22D0BWP12T U682 ( .A1(r3[8]), .A2(n3078), .B1(n3079), .B2(r2[8]), .ZN(n92) );
  AOI22D0BWP12T U683 ( .A1(r4[8]), .A2(n3080), .B1(n3081), .B2(r0[8]), .ZN(n93) );
  ND4D0BWP12T U684 ( .A1(n90), .A2(n91), .A3(n92), .A4(n93), .ZN(n94) );
  OAI22D0BWP12T U685 ( .A1(n3042), .A2(n2996), .B1(n2997), .B2(n3028), .ZN(n95) );
  MOAI22D0BWP12T U686 ( .A1(n3066), .A2(n2995), .B1(n3073), .B2(r8[8]), .ZN(
        n96) );
  AOI211D0BWP12T U687 ( .A1(n3086), .A2(n94), .B(n95), .C(n96), .ZN(n97) );
  ND3D0BWP12T U688 ( .A1(n88), .A2(n89), .A3(n97), .ZN(regD_out[8]) );
  MOAI22D0BWP12T U689 ( .A1(n3137), .A2(n3136), .B1(n3137), .B2(n3136), .ZN(
        n98) );
  AOI22D0BWP12T U690 ( .A1(pc_out[15]), .A2(n3498), .B1(n3499), .B2(
        next_pc_in[15]), .ZN(n99) );
  OAI21D0BWP12T U691 ( .A1(n3497), .A2(n98), .B(n99), .ZN(n2183) );
  AO222D0BWP12T U692 ( .A1(n3269), .A2(write1_in[12]), .B1(write2_in[12]), 
        .B2(n3270), .C1(r9[12]), .C2(n3271), .Z(n2340) );
  AO222D0BWP12T U693 ( .A1(n3269), .A2(n177), .B1(n3270), .B2(write2_in[15]), 
        .C1(r9[15]), .C2(n3271), .Z(n2343) );
  AO222D0BWP12T U694 ( .A1(n3269), .A2(n3054), .B1(n3270), .B2(write2_in[17]), 
        .C1(r9[17]), .C2(n3271), .Z(n2345) );
  AO222D0BWP12T U695 ( .A1(n3269), .A2(n3060), .B1(write2_in[18]), .B2(n3270), 
        .C1(r9[18]), .C2(n3271), .Z(n2346) );
  AO222D0BWP12T U696 ( .A1(n3269), .A2(n3098), .B1(n3270), .B2(write2_in[21]), 
        .C1(r9[21]), .C2(n3271), .Z(n2349) );
  AO222D0BWP12T U697 ( .A1(n3269), .A2(n3108), .B1(n3270), .B2(write2_in[26]), 
        .C1(r9[26]), .C2(n3271), .Z(n2354) );
  AO222D0BWP12T U698 ( .A1(n3519), .A2(write1_in[14]), .B1(n3214), .B2(
        write2_in[14]), .C1(r8[14]), .C2(n3215), .Z(n2374) );
  AO222D0BWP12T U699 ( .A1(n3519), .A2(n3055), .B1(write2_in[16]), .B2(n3214), 
        .C1(r8[16]), .C2(n3215), .Z(n2376) );
  AO222D0BWP12T U700 ( .A1(n3519), .A2(n3096), .B1(n3214), .B2(write2_in[19]), 
        .C1(r8[19]), .C2(n3215), .Z(n2379) );
  AO222D0BWP12T U701 ( .A1(n3519), .A2(n3095), .B1(n3214), .B2(write2_in[20]), 
        .C1(r8[20]), .C2(n3215), .Z(n2380) );
  AO222D0BWP12T U702 ( .A1(n3519), .A2(n3099), .B1(n3214), .B2(write2_in[22]), 
        .C1(r8[22]), .C2(n3215), .Z(n2382) );
  AO222D0BWP12T U703 ( .A1(n3519), .A2(write1_in[23]), .B1(n3214), .B2(
        write2_in[23]), .C1(r8[23]), .C2(n3215), .Z(n2383) );
  AO222D0BWP12T U704 ( .A1(n3519), .A2(n3097), .B1(n3214), .B2(write2_in[24]), 
        .C1(r8[24]), .C2(n3215), .Z(n2384) );
  AO222D0BWP12T U705 ( .A1(n3519), .A2(n3113), .B1(n3214), .B2(write2_in[25]), 
        .C1(r8[25]), .C2(n3215), .Z(n2385) );
  AOI22D0BWP12T U706 ( .A1(r12[9]), .A2(n3064), .B1(n2994), .B2(r11[9]), .ZN(
        n100) );
  AOI22D0BWP12T U707 ( .A1(pc_out[9]), .A2(n3061), .B1(n3062), .B2(lr[9]), 
        .ZN(n101) );
  AOI22D0BWP12T U708 ( .A1(r1[9]), .A2(n3074), .B1(n3075), .B2(r5[9]), .ZN(
        n102) );
  AOI22D0BWP12T U709 ( .A1(r7[9]), .A2(n3076), .B1(n3077), .B2(r6[9]), .ZN(
        n103) );
  AOI22D0BWP12T U710 ( .A1(r3[9]), .A2(n3078), .B1(n3079), .B2(r2[9]), .ZN(
        n104) );
  AOI22D0BWP12T U711 ( .A1(r4[9]), .A2(n3080), .B1(n3081), .B2(r0[9]), .ZN(
        n105) );
  ND4D0BWP12T U712 ( .A1(n102), .A2(n103), .A3(n104), .A4(n105), .ZN(n106) );
  OAI22D0BWP12T U713 ( .A1(n2886), .A2(n2984), .B1(n2887), .B2(n3069), .ZN(
        n107) );
  MOAI22D0BWP12T U714 ( .A1(n3066), .A2(n2941), .B1(n3073), .B2(r8[9]), .ZN(
        n108) );
  AOI211D0BWP12T U715 ( .A1(n3086), .A2(n106), .B(n107), .C(n108), .ZN(n109)
         );
  ND3D0BWP12T U716 ( .A1(n100), .A2(n101), .A3(n109), .ZN(regD_out[9]) );
  AO222D0BWP12T U717 ( .A1(n3519), .A2(write1_in[12]), .B1(write2_in[12]), 
        .B2(n3214), .C1(r8[12]), .C2(n3215), .Z(n2372) );
  AO222D0BWP12T U718 ( .A1(n3519), .A2(write1_in[15]), .B1(n3214), .B2(
        write2_in[15]), .C1(r8[15]), .C2(n3215), .Z(n2375) );
  AO222D0BWP12T U719 ( .A1(n3519), .A2(n3054), .B1(n3214), .B2(write2_in[17]), 
        .C1(r8[17]), .C2(n3215), .Z(n2377) );
  AO222D0BWP12T U720 ( .A1(n3519), .A2(n3060), .B1(write2_in[18]), .B2(n3214), 
        .C1(r8[18]), .C2(n3215), .Z(n2378) );
  AO222D0BWP12T U721 ( .A1(n3519), .A2(n3098), .B1(n3214), .B2(write2_in[21]), 
        .C1(r8[21]), .C2(n3215), .Z(n2381) );
  AO222D0BWP12T U722 ( .A1(n3519), .A2(n3108), .B1(n3214), .B2(write2_in[26]), 
        .C1(r8[26]), .C2(n3215), .Z(n2386) );
  AO222D0BWP12T U723 ( .A1(n3264), .A2(write1_in[14]), .B1(n3265), .B2(
        write2_in[14]), .C1(r7[14]), .C2(n3266), .Z(n2406) );
  AO222D0BWP12T U724 ( .A1(n3264), .A2(n3055), .B1(write2_in[16]), .B2(n3265), 
        .C1(r7[16]), .C2(n3266), .Z(n2408) );
  AO222D0BWP12T U725 ( .A1(n3264), .A2(n3096), .B1(n3265), .B2(write2_in[19]), 
        .C1(r7[19]), .C2(n3266), .Z(n2411) );
  AO222D0BWP12T U726 ( .A1(n3264), .A2(n3095), .B1(n3265), .B2(write2_in[20]), 
        .C1(r7[20]), .C2(n3266), .Z(n2412) );
  AO222D0BWP12T U727 ( .A1(n3264), .A2(n3099), .B1(n3265), .B2(write2_in[22]), 
        .C1(r7[22]), .C2(n3266), .Z(n2414) );
  AO222D0BWP12T U728 ( .A1(n3264), .A2(write1_in[23]), .B1(n3265), .B2(
        write2_in[23]), .C1(r7[23]), .C2(n3266), .Z(n2415) );
  AO222D0BWP12T U729 ( .A1(n3264), .A2(n3097), .B1(n3265), .B2(write2_in[24]), 
        .C1(r7[24]), .C2(n3266), .Z(n2416) );
  AO222D0BWP12T U730 ( .A1(n3264), .A2(n3113), .B1(n3265), .B2(write2_in[25]), 
        .C1(r7[25]), .C2(n3266), .Z(n2417) );
  MOAI22D0BWP12T U731 ( .A1(n3434), .A2(n1387), .B1(n3445), .B2(pc_out[15]), 
        .ZN(n1389) );
  AOI22D0BWP12T U732 ( .A1(pc_out[10]), .A2(n3061), .B1(r9[10]), .B2(n3063), 
        .ZN(n110) );
  AOI22D0BWP12T U733 ( .A1(lr[10]), .A2(n3062), .B1(n[3570]), .B2(n3037), .ZN(
        n111) );
  AOI22D0BWP12T U734 ( .A1(r1[10]), .A2(n3074), .B1(r5[10]), .B2(n3075), .ZN(
        n112) );
  AOI22D0BWP12T U735 ( .A1(r6[10]), .A2(n3077), .B1(r7[10]), .B2(n3076), .ZN(
        n113) );
  AOI22D0BWP12T U736 ( .A1(r2[10]), .A2(n3079), .B1(r3[10]), .B2(n3078), .ZN(
        n114) );
  AOI22D0BWP12T U737 ( .A1(r0[10]), .A2(n3081), .B1(r4[10]), .B2(n3080), .ZN(
        n115) );
  ND4D0BWP12T U738 ( .A1(n112), .A2(n113), .A3(n114), .A4(n115), .ZN(n116) );
  OAI22D0BWP12T U739 ( .A1(n2955), .A2(n2920), .B1(n2963), .B2(n3068), .ZN(
        n117) );
  MOAI22D0BWP12T U740 ( .A1(n2975), .A2(n3066), .B1(n3073), .B2(r8[10]), .ZN(
        n118) );
  AOI211D0BWP12T U741 ( .A1(n3086), .A2(n116), .B(n117), .C(n118), .ZN(n119)
         );
  ND3D0BWP12T U742 ( .A1(n110), .A2(n111), .A3(n119), .ZN(regD_out[10]) );
  AO222D0BWP12T U743 ( .A1(n3264), .A2(write1_in[12]), .B1(write2_in[12]), 
        .B2(n3265), .C1(r7[12]), .C2(n3266), .Z(n2404) );
  AO222D0BWP12T U744 ( .A1(n3264), .A2(n177), .B1(n3265), .B2(write2_in[15]), 
        .C1(r7[15]), .C2(n3266), .Z(n2407) );
  AO222D0BWP12T U745 ( .A1(n3264), .A2(n3060), .B1(write2_in[18]), .B2(n3265), 
        .C1(r7[18]), .C2(n3266), .Z(n2410) );
  AO222D0BWP12T U746 ( .A1(n3264), .A2(n3098), .B1(n3265), .B2(write2_in[21]), 
        .C1(r7[21]), .C2(n3266), .Z(n2413) );
  AO222D0BWP12T U747 ( .A1(n3264), .A2(n3108), .B1(n3265), .B2(write2_in[26]), 
        .C1(r7[26]), .C2(n3266), .Z(n2418) );
  AO222D0BWP12T U748 ( .A1(n3274), .A2(write1_in[14]), .B1(n3276), .B2(
        write2_in[14]), .C1(r6[14]), .C2(n3277), .Z(n2438) );
  AO222D0BWP12T U749 ( .A1(n3274), .A2(n3055), .B1(write2_in[16]), .B2(n3276), 
        .C1(r6[16]), .C2(n3277), .Z(n2440) );
  AO222D0BWP12T U750 ( .A1(n3274), .A2(n3054), .B1(n3276), .B2(write2_in[17]), 
        .C1(r6[17]), .C2(n3277), .Z(n2441) );
  AO222D0BWP12T U751 ( .A1(n3274), .A2(n3096), .B1(n3276), .B2(write2_in[19]), 
        .C1(r6[19]), .C2(n3277), .Z(n2443) );
  AO222D0BWP12T U752 ( .A1(n3274), .A2(n3095), .B1(n3276), .B2(write2_in[20]), 
        .C1(r6[20]), .C2(n3277), .Z(n2444) );
  AO222D0BWP12T U753 ( .A1(n3274), .A2(n3099), .B1(n3276), .B2(write2_in[22]), 
        .C1(r6[22]), .C2(n3277), .Z(n2446) );
  AO222D0BWP12T U754 ( .A1(n3274), .A2(write1_in[23]), .B1(n3276), .B2(
        write2_in[23]), .C1(r6[23]), .C2(n3277), .Z(n2447) );
  AO222D0BWP12T U755 ( .A1(n3274), .A2(n3097), .B1(n3276), .B2(write2_in[24]), 
        .C1(r6[24]), .C2(n3277), .Z(n2448) );
  AO222D0BWP12T U756 ( .A1(n3274), .A2(n3113), .B1(n3276), .B2(write2_in[25]), 
        .C1(r6[25]), .C2(n3277), .Z(n2449) );
  MOAI22D0BWP12T U757 ( .A1(n3446), .A2(n1297), .B1(pc_out[11]), .B2(n3445), 
        .ZN(n1302) );
  ND4D0BWP12T U758 ( .A1(write2_en), .A2(write2_sel[4]), .A3(n532), .A4(
        write2_sel[3]), .ZN(n120) );
  OR2D0BWP12T U759 ( .A1(write2_sel[0]), .A2(n120), .Z(n369) );
  AO222D0BWP12T U760 ( .A1(n3274), .A2(write1_in[12]), .B1(write2_in[12]), 
        .B2(n3276), .C1(r6[12]), .C2(n3277), .Z(n2436) );
  AO222D0BWP12T U761 ( .A1(n3274), .A2(n177), .B1(n3276), .B2(write2_in[15]), 
        .C1(r6[15]), .C2(n3277), .Z(n2439) );
  AO222D0BWP12T U762 ( .A1(n3274), .A2(n3060), .B1(write2_in[18]), .B2(n3276), 
        .C1(r6[18]), .C2(n3277), .Z(n2442) );
  AO222D0BWP12T U763 ( .A1(n3274), .A2(n3098), .B1(n3276), .B2(write2_in[21]), 
        .C1(r6[21]), .C2(n3277), .Z(n2445) );
  AO222D0BWP12T U764 ( .A1(n3254), .A2(write1_in[14]), .B1(n3255), .B2(
        write2_in[14]), .C1(r5[14]), .C2(n3256), .Z(n2470) );
  AO222D0BWP12T U765 ( .A1(n3254), .A2(n3055), .B1(write2_in[16]), .B2(n3255), 
        .C1(r5[16]), .C2(n3256), .Z(n2472) );
  AO222D0BWP12T U766 ( .A1(n3254), .A2(n3054), .B1(n3255), .B2(write2_in[17]), 
        .C1(r5[17]), .C2(n3256), .Z(n2473) );
  AO222D0BWP12T U767 ( .A1(n3254), .A2(n3096), .B1(n3255), .B2(write2_in[19]), 
        .C1(r5[19]), .C2(n3256), .Z(n2475) );
  AO222D0BWP12T U768 ( .A1(n3254), .A2(n3095), .B1(n3255), .B2(write2_in[20]), 
        .C1(r5[20]), .C2(n3256), .Z(n2476) );
  AO222D0BWP12T U769 ( .A1(n3254), .A2(n3282), .B1(n3255), .B2(write2_in[22]), 
        .C1(r5[22]), .C2(n3256), .Z(n2478) );
  AO222D0BWP12T U770 ( .A1(n3254), .A2(write1_in[23]), .B1(n3255), .B2(
        write2_in[23]), .C1(r5[23]), .C2(n3256), .Z(n2479) );
  AO222D0BWP12T U771 ( .A1(n3254), .A2(n3097), .B1(n3255), .B2(write2_in[24]), 
        .C1(r5[24]), .C2(n3256), .Z(n2480) );
  AO222D0BWP12T U772 ( .A1(n3254), .A2(n3113), .B1(n3255), .B2(write2_in[25]), 
        .C1(r5[25]), .C2(n3256), .Z(n2481) );
  AO222D0BWP12T U773 ( .A1(n3254), .A2(n3108), .B1(n3255), .B2(write2_in[26]), 
        .C1(r5[26]), .C2(n3256), .Z(n2482) );
  AO222D0BWP12T U774 ( .A1(n3518), .A2(write1_in[13]), .B1(write2_in[13]), 
        .B2(n3222), .C1(r4[13]), .C2(n3223), .Z(n2501) );
  IND3D0BWP12T U775 ( .A1(n365), .B1(n360), .B2(write1_sel[3]), .ZN(n544) );
  AO22D1BWP12T U776 ( .A1(n530), .A2(write1_in[2]), .B1(write2_in[2]), .B2(
        n3331), .Z(n2845) );
  AO222D0BWP12T U777 ( .A1(n3254), .A2(write1_in[12]), .B1(write2_in[12]), 
        .B2(n3255), .C1(r5[12]), .C2(n3256), .Z(n2468) );
  AO222D0BWP12T U778 ( .A1(n3254), .A2(n3060), .B1(write2_in[18]), .B2(n3255), 
        .C1(r5[18]), .C2(n3256), .Z(n2474) );
  AO222D0BWP12T U779 ( .A1(n3518), .A2(write1_in[14]), .B1(n3222), .B2(
        write2_in[14]), .C1(r4[14]), .C2(n3223), .Z(n2502) );
  AO222D0BWP12T U780 ( .A1(n3518), .A2(write1_in[15]), .B1(n3222), .B2(
        write2_in[15]), .C1(r4[15]), .C2(n3223), .Z(n2503) );
  AO222D0BWP12T U781 ( .A1(n3518), .A2(n3055), .B1(write2_in[16]), .B2(n3222), 
        .C1(r4[16]), .C2(n3223), .Z(n2504) );
  AO222D0BWP12T U782 ( .A1(n3518), .A2(n3054), .B1(n3222), .B2(write2_in[17]), 
        .C1(r4[17]), .C2(n3223), .Z(n2505) );
  AO222D0BWP12T U783 ( .A1(n3518), .A2(n3096), .B1(n3222), .B2(write2_in[19]), 
        .C1(r4[19]), .C2(n3223), .Z(n2507) );
  AO222D0BWP12T U784 ( .A1(n3518), .A2(n3095), .B1(n3222), .B2(write2_in[20]), 
        .C1(r4[20]), .C2(n3223), .Z(n2508) );
  AO222D0BWP12T U785 ( .A1(n3518), .A2(n3098), .B1(n3222), .B2(write2_in[21]), 
        .C1(r4[21]), .C2(n3223), .Z(n2509) );
  AO222D0BWP12T U786 ( .A1(n3518), .A2(n3099), .B1(n3222), .B2(write2_in[22]), 
        .C1(r4[22]), .C2(n3223), .Z(n2510) );
  AO222D0BWP12T U787 ( .A1(n3518), .A2(write1_in[23]), .B1(n3222), .B2(
        write2_in[23]), .C1(r4[23]), .C2(n3223), .Z(n2511) );
  AO222D0BWP12T U788 ( .A1(n3518), .A2(n3097), .B1(n3222), .B2(write2_in[24]), 
        .C1(r4[24]), .C2(n3223), .Z(n2512) );
  AO222D0BWP12T U789 ( .A1(n3518), .A2(n3113), .B1(n3222), .B2(write2_in[25]), 
        .C1(r4[25]), .C2(n3223), .Z(n2513) );
  AO222D0BWP12T U790 ( .A1(n3518), .A2(n3108), .B1(n3222), .B2(write2_in[26]), 
        .C1(r4[26]), .C2(n3223), .Z(n2514) );
  AO222D0BWP12T U791 ( .A1(n3515), .A2(write1_in[13]), .B1(write2_in[13]), 
        .B2(n3189), .C1(r3[13]), .C2(n3190), .Z(n2533) );
  MOAI22D0BWP12T U792 ( .A1(n3414), .A2(n1485), .B1(n3417), .B2(r1[12]), .ZN(
        n1467) );
  MAOI22D1BWP12T U793 ( .A1(lr[11]), .A2(n1859), .B1(n1787), .B2(n2896), .ZN(
        n1296) );
  AOI21D0BWP12T U794 ( .A1(n531), .A2(n532), .B(n530), .ZN(n602) );
  MOAI22D0BWP12T U795 ( .A1(n3101), .A2(n3102), .B1(n3101), .B2(n3102), .ZN(
        n121) );
  AOI22D0BWP12T U796 ( .A1(n3499), .A2(next_pc_in[11]), .B1(pc_out[11]), .B2(
        n3498), .ZN(n122) );
  OAI21D0BWP12T U797 ( .A1(n3497), .A2(n121), .B(n122), .ZN(n2179) );
  IND2D0BWP12T U798 ( .A1(n3030), .B1(n3031), .ZN(n123) );
  MAOI22D0BWP12T U799 ( .A1(n3032), .A2(n123), .B1(n3032), .B2(n123), .ZN(n124) );
  AO222D0BWP12T U800 ( .A1(n124), .A2(n3505), .B1(pc_out[6]), .B2(n3498), .C1(
        next_pc_in[6]), .C2(n3499), .Z(n2174) );
  AO222D0BWP12T U801 ( .A1(n3518), .A2(write1_in[12]), .B1(write2_in[12]), 
        .B2(n3222), .C1(r4[12]), .C2(n3223), .Z(n2500) );
  AO222D0BWP12T U802 ( .A1(n3518), .A2(n3060), .B1(write2_in[18]), .B2(n3222), 
        .C1(r4[18]), .C2(n3223), .Z(n2506) );
  AO222D0BWP12T U803 ( .A1(n3515), .A2(write1_in[14]), .B1(write2_in[14]), 
        .B2(n3189), .C1(r3[14]), .C2(n3190), .Z(n2534) );
  AO222D0BWP12T U804 ( .A1(n3515), .A2(n177), .B1(write2_in[15]), .B2(n3189), 
        .C1(r3[15]), .C2(n3190), .Z(n2535) );
  AO222D0BWP12T U805 ( .A1(n3515), .A2(n3055), .B1(write2_in[16]), .B2(n3189), 
        .C1(r3[16]), .C2(n3190), .Z(n2536) );
  AO222D0BWP12T U806 ( .A1(n3515), .A2(n3054), .B1(write2_in[17]), .B2(n3189), 
        .C1(r3[17]), .C2(n3190), .Z(n2537) );
  AO222D0BWP12T U807 ( .A1(n3515), .A2(n3096), .B1(write2_in[19]), .B2(n3189), 
        .C1(r3[19]), .C2(n3190), .Z(n2539) );
  AO222D0BWP12T U808 ( .A1(n3515), .A2(n3095), .B1(write2_in[20]), .B2(n3189), 
        .C1(r3[20]), .C2(n3190), .Z(n2540) );
  AO222D0BWP12T U809 ( .A1(n3515), .A2(n3098), .B1(write2_in[21]), .B2(n3189), 
        .C1(r3[21]), .C2(n3190), .Z(n2541) );
  AO222D0BWP12T U810 ( .A1(n3515), .A2(n3099), .B1(write2_in[22]), .B2(n3189), 
        .C1(r3[22]), .C2(n3190), .Z(n2542) );
  AO222D0BWP12T U811 ( .A1(n3515), .A2(write1_in[23]), .B1(write2_in[23]), 
        .B2(n3189), .C1(r3[23]), .C2(n3190), .Z(n2543) );
  AO222D0BWP12T U812 ( .A1(n3515), .A2(n3097), .B1(write2_in[24]), .B2(n3189), 
        .C1(r3[24]), .C2(n3190), .Z(n2544) );
  AO222D0BWP12T U813 ( .A1(n3515), .A2(n3113), .B1(write2_in[25]), .B2(n3189), 
        .C1(r3[25]), .C2(n3190), .Z(n2545) );
  AO222D0BWP12T U814 ( .A1(n3515), .A2(n3108), .B1(write2_in[26]), .B2(n3189), 
        .C1(r3[26]), .C2(n3190), .Z(n2546) );
  AO222D0BWP12T U815 ( .A1(n3516), .A2(write1_in[13]), .B1(write2_in[13]), 
        .B2(n3193), .C1(r2[13]), .C2(n3194), .Z(n2565) );
  INR2D0BWP12T U816 ( .A1(r8[15]), .B1(n1372), .ZN(n1373) );
  MOAI22D0BWP12T U817 ( .A1(n1881), .A2(n2082), .B1(n3445), .B2(pc_out[16]), 
        .ZN(n1206) );
  MOAI22D0BWP12T U818 ( .A1(n3414), .A2(n1547), .B1(n3417), .B2(r1[14]), .ZN(
        n651) );
  IND2D0BWP12T U819 ( .A1(n585), .B1(n419), .ZN(n570) );
  MOAI22D0BWP12T U820 ( .A1(n3547), .A2(n3343), .B1(next_pc_in[30]), .B2(n3499), .ZN(n908) );
  INR2D1BWP12T U821 ( .A1(n369), .B1(n370), .ZN(n1946) );
  OAI22D0BWP12T U822 ( .A1(n3026), .A2(n3068), .B1(n3025), .B2(n3024), .ZN(
        n125) );
  CKND0BWP12T U823 ( .I(pc_out[11]), .ZN(n126) );
  OAI22D0BWP12T U824 ( .A1(n3042), .A2(n3027), .B1(n3028), .B2(n126), .ZN(n127) );
  AOI211D0BWP12T U825 ( .A1(r10[11]), .A2(n3029), .B(n125), .C(n127), .ZN(n128) );
  AOI22D0BWP12T U826 ( .A1(n[3569]), .A2(n3037), .B1(r12[11]), .B2(n3064), 
        .ZN(n129) );
  AOI22D0BWP12T U827 ( .A1(r1[11]), .A2(n3074), .B1(r5[11]), .B2(n3075), .ZN(
        n130) );
  AOI22D0BWP12T U828 ( .A1(r6[11]), .A2(n3077), .B1(r7[11]), .B2(n3076), .ZN(
        n131) );
  AOI22D0BWP12T U829 ( .A1(r2[11]), .A2(n3079), .B1(r3[11]), .B2(n3078), .ZN(
        n132) );
  AOI22D0BWP12T U830 ( .A1(r0[11]), .A2(n3081), .B1(r4[11]), .B2(n3080), .ZN(
        n133) );
  ND4D0BWP12T U831 ( .A1(n130), .A2(n131), .A3(n132), .A4(n133), .ZN(n134) );
  AOI22D0BWP12T U832 ( .A1(r9[11]), .A2(n3063), .B1(n3086), .B2(n134), .ZN(
        n135) );
  ND3D0BWP12T U833 ( .A1(n128), .A2(n129), .A3(n135), .ZN(regD_out[11]) );
  MAOI22D0BWP12T U834 ( .A1(n2950), .A2(n2949), .B1(n2950), .B2(n2949), .ZN(
        n136) );
  AO222D0BWP12T U835 ( .A1(n3505), .A2(n136), .B1(pc_out[3]), .B2(n3498), .C1(
        n3499), .C2(next_pc_in[3]), .Z(n2171) );
  OAI22D0BWP12T U836 ( .A1(write1_in[0]), .A2(n3331), .B1(n530), .B2(
        write2_in[0]), .ZN(n137) );
  AOI22D0BWP12T U837 ( .A1(pc_out[0]), .A2(n3498), .B1(next_pc_in[0]), .B2(
        n3499), .ZN(n138) );
  OAI21D0BWP12T U838 ( .A1(n3497), .A2(n137), .B(n138), .ZN(n2168) );
  IND2D0BWP12T U839 ( .A1(n3056), .B1(n3057), .ZN(n139) );
  CKND2D0BWP12T U840 ( .A1(n3058), .A2(n3059), .ZN(n140) );
  MAOI22D0BWP12T U841 ( .A1(n139), .A2(n140), .B1(n139), .B2(n140), .ZN(n141)
         );
  AOI22D0BWP12T U842 ( .A1(pc_out[9]), .A2(n3498), .B1(next_pc_in[9]), .B2(
        n3499), .ZN(n142) );
  OAI21D0BWP12T U843 ( .A1(n3497), .A2(n141), .B(n142), .ZN(n2177) );
  AO222D0BWP12T U844 ( .A1(n3515), .A2(write1_in[12]), .B1(write2_in[12]), 
        .B2(n3189), .C1(r3[12]), .C2(n3190), .Z(n2532) );
  AO222D0BWP12T U845 ( .A1(n3515), .A2(n3060), .B1(write2_in[18]), .B2(n3189), 
        .C1(r3[18]), .C2(n3190), .Z(n2538) );
  AO222D0BWP12T U846 ( .A1(n3516), .A2(write1_in[14]), .B1(write2_in[14]), 
        .B2(n3193), .C1(r2[14]), .C2(n3194), .Z(n2566) );
  AO222D0BWP12T U847 ( .A1(n3516), .A2(write1_in[15]), .B1(write2_in[15]), 
        .B2(n3193), .C1(r2[15]), .C2(n3194), .Z(n2567) );
  AO222D0BWP12T U848 ( .A1(n3516), .A2(n3055), .B1(write2_in[16]), .B2(n3193), 
        .C1(r2[16]), .C2(n3194), .Z(n2568) );
  AO222D0BWP12T U849 ( .A1(n3516), .A2(n3054), .B1(write2_in[17]), .B2(n3193), 
        .C1(r2[17]), .C2(n3194), .Z(n2569) );
  AO222D0BWP12T U850 ( .A1(n3516), .A2(n3096), .B1(write2_in[19]), .B2(n3193), 
        .C1(r2[19]), .C2(n3194), .Z(n2571) );
  AO222D0BWP12T U851 ( .A1(n3516), .A2(n3095), .B1(write2_in[20]), .B2(n3193), 
        .C1(r2[20]), .C2(n3194), .Z(n2572) );
  AO222D0BWP12T U852 ( .A1(n3516), .A2(n3098), .B1(write2_in[21]), .B2(n3193), 
        .C1(r2[21]), .C2(n3194), .Z(n2573) );
  AO222D0BWP12T U853 ( .A1(n3516), .A2(n3282), .B1(write2_in[22]), .B2(n3193), 
        .C1(r2[22]), .C2(n3194), .Z(n2574) );
  AO222D0BWP12T U854 ( .A1(n3516), .A2(write1_in[23]), .B1(write2_in[23]), 
        .B2(n3193), .C1(r2[23]), .C2(n3194), .Z(n2575) );
  AO222D0BWP12T U855 ( .A1(n3516), .A2(n3097), .B1(write2_in[24]), .B2(n3193), 
        .C1(r2[24]), .C2(n3194), .Z(n2576) );
  AO222D0BWP12T U856 ( .A1(n3516), .A2(n3113), .B1(write2_in[25]), .B2(n3193), 
        .C1(r2[25]), .C2(n3194), .Z(n2577) );
  AO222D0BWP12T U857 ( .A1(n3516), .A2(n3108), .B1(write2_in[26]), .B2(n3193), 
        .C1(r2[26]), .C2(n3194), .Z(n2578) );
  AO222D0BWP12T U858 ( .A1(n3231), .A2(write1_in[13]), .B1(write2_in[13]), 
        .B2(n3232), .C1(r1[13]), .C2(n3233), .Z(n2597) );
  CKND0BWP12T U859 ( .I(tmp1[12]), .ZN(n143) );
  MOAI22D0BWP12T U860 ( .A1(n3378), .A2(n143), .B1(immediate1_in[12]), .B2(
        n1804), .ZN(n1466) );
  IND2D0BWP12T U861 ( .A1(n1837), .B1(r5[15]), .ZN(n1374) );
  MOAI22D1BWP12T U862 ( .A1(n3444), .A2(n1723), .B1(n1859), .B2(lr[7]), .ZN(
        n867) );
  MOAI22D1BWP12T U863 ( .A1(n3436), .A2(n2018), .B1(n1788), .B2(pc_out[5]), 
        .ZN(n698) );
  MOAI22D0BWP12T U864 ( .A1(n1881), .A2(n2900), .B1(n3450), .B2(r4[11]), .ZN(
        n1303) );
  CKND0BWP12T U865 ( .I(n3331), .ZN(n144) );
  OA21D0BWP12T U866 ( .A1(n3318), .A2(n144), .B(n3330), .Z(n3321) );
  IND2D0BWP12T U867 ( .A1(n591), .B1(n419), .ZN(n578) );
  MOAI22D0BWP12T U868 ( .A1(n3533), .A2(n3343), .B1(next_pc_in[29]), .B2(n3499), .ZN(n1603) );
  OAI31D0BWP12T U869 ( .A1(write2_sel[2]), .A2(n546), .A3(n545), .B(n3532), 
        .ZN(n145) );
  NR2D0BWP12T U870 ( .A1(n547), .A2(n145), .ZN(n3201) );
  AO222D0BWP12T U871 ( .A1(n3246), .A2(write1_in[11]), .B1(write2_in[11]), 
        .B2(n1947), .C1(tmp1[11]), .C2(n1946), .Z(n2147) );
  MAOI22D0BWP12T U872 ( .A1(n2845), .A2(n2844), .B1(n2845), .B2(n2844), .ZN(
        n146) );
  AO222D0BWP12T U873 ( .A1(n146), .A2(n3505), .B1(pc_out[2]), .B2(n3498), .C1(
        n3499), .C2(next_pc_in[2]), .Z(n2170) );
  MOAI22D0BWP12T U874 ( .A1(n3093), .A2(n3092), .B1(n3093), .B2(n3092), .ZN(
        n147) );
  AOI22D0BWP12T U875 ( .A1(pc_out[10]), .A2(n3498), .B1(next_pc_in[10]), .B2(
        n3499), .ZN(n148) );
  OAI21D0BWP12T U876 ( .A1(n3497), .A2(n147), .B(n148), .ZN(n2178) );
  MOAI22D0BWP12T U877 ( .A1(n3110), .A2(n3109), .B1(n3110), .B2(n3109), .ZN(
        n149) );
  AOI22D0BWP12T U878 ( .A1(pc_out[13]), .A2(n3498), .B1(n3499), .B2(
        next_pc_in[13]), .ZN(n150) );
  OAI21D0BWP12T U879 ( .A1(n3497), .A2(n149), .B(n150), .ZN(n2181) );
  AO222D0BWP12T U880 ( .A1(n3516), .A2(write1_in[12]), .B1(write2_in[12]), 
        .B2(n3193), .C1(r2[12]), .C2(n3194), .Z(n2564) );
  AO222D0BWP12T U881 ( .A1(n3516), .A2(n3060), .B1(write2_in[18]), .B2(n3193), 
        .C1(r2[18]), .C2(n3194), .Z(n2570) );
  AO222D0BWP12T U882 ( .A1(n3231), .A2(write1_in[14]), .B1(n3232), .B2(
        write2_in[14]), .C1(r1[14]), .C2(n3233), .Z(n2598) );
  AO222D0BWP12T U883 ( .A1(n3231), .A2(n177), .B1(n3232), .B2(write2_in[15]), 
        .C1(r1[15]), .C2(n3233), .Z(n2599) );
  AO222D0BWP12T U884 ( .A1(n3231), .A2(n3055), .B1(write2_in[16]), .B2(n3232), 
        .C1(r1[16]), .C2(n3233), .Z(n2600) );
  AO222D0BWP12T U885 ( .A1(n3231), .A2(n3054), .B1(n3232), .B2(write2_in[17]), 
        .C1(r1[17]), .C2(n3233), .Z(n2601) );
  AO222D0BWP12T U886 ( .A1(n3231), .A2(n3096), .B1(n3232), .B2(write2_in[19]), 
        .C1(r1[19]), .C2(n3233), .Z(n2603) );
  AO222D0BWP12T U887 ( .A1(n3231), .A2(n3095), .B1(n3232), .B2(write2_in[20]), 
        .C1(r1[20]), .C2(n3233), .Z(n2604) );
  AO222D0BWP12T U888 ( .A1(n3231), .A2(n3098), .B1(n3232), .B2(write2_in[21]), 
        .C1(r1[21]), .C2(n3233), .Z(n2605) );
  AO222D0BWP12T U889 ( .A1(n3231), .A2(n3282), .B1(n3232), .B2(write2_in[22]), 
        .C1(r1[22]), .C2(n3233), .Z(n2606) );
  AO222D0BWP12T U890 ( .A1(n3231), .A2(write1_in[23]), .B1(n3232), .B2(
        write2_in[23]), .C1(r1[23]), .C2(n3233), .Z(n2607) );
  AO222D0BWP12T U891 ( .A1(n3231), .A2(n3097), .B1(n3232), .B2(write2_in[24]), 
        .C1(r1[24]), .C2(n3233), .Z(n2608) );
  AO222D0BWP12T U892 ( .A1(n3231), .A2(n3113), .B1(n3232), .B2(write2_in[25]), 
        .C1(r1[25]), .C2(n3233), .Z(n2609) );
  AO222D0BWP12T U893 ( .A1(n3231), .A2(n3108), .B1(n3232), .B2(write2_in[26]), 
        .C1(r1[26]), .C2(n3233), .Z(n2610) );
  MOAI22D0BWP12T U894 ( .A1(n3444), .A2(n1489), .B1(n1788), .B2(pc_out[12]), 
        .ZN(n1479) );
  CKND0BWP12T U895 ( .I(r12[15]), .ZN(n151) );
  MOAI22D0BWP12T U896 ( .A1(n3436), .A2(n151), .B1(immediate1_in[15]), .B2(
        n1804), .ZN(n1388) );
  AO22D0BWP12T U897 ( .A1(r6[17]), .A2(n3412), .B1(r8[17]), .B2(n1473), .Z(
        n612) );
  ND3D0BWP12T U898 ( .A1(n[3573]), .A2(n861), .A3(n1049), .ZN(n863) );
  INR2D0BWP12T U899 ( .A1(r12[14]), .B1(n3436), .ZN(n650) );
  MOAI22D0BWP12T U900 ( .A1(n3404), .A2(n1368), .B1(n3419), .B2(r9[15]), .ZN(
        n1369) );
  MOAI22D0BWP12T U901 ( .A1(n3434), .A2(n2888), .B1(n1380), .B2(tmp1[11]), 
        .ZN(n1305) );
  IND2D0BWP12T U902 ( .A1(n1564), .B1(lr[20]), .ZN(n919) );
  AOI22D0BWP12T U903 ( .A1(pc_out[26]), .A2(n3498), .B1(n3499), .B2(
        next_pc_in[26]), .ZN(n1135) );
  INR2D0BWP12T U904 ( .A1(n359), .B1(write1_sel[2]), .ZN(n419) );
  NR2D0BWP12T U905 ( .A1(n901), .A2(write1_in[29]), .ZN(n902) );
  MOAI22D0BWP12T U906 ( .A1(n3442), .A2(n2864), .B1(n1873), .B2(r5[7]), .ZN(
        n859) );
  MAOI22D0BWP12T U907 ( .A1(n3499), .A2(next_pc_in[21]), .B1(n3343), .B2(n3514), .ZN(n1740) );
  CKND2D0BWP12T U908 ( .A1(n3499), .A2(next_pc_in[31]), .ZN(n3330) );
  AOI22D0BWP12T U909 ( .A1(pc_out[20]), .A2(n3498), .B1(n3499), .B2(
        next_pc_in[20]), .ZN(n3500) );
  INR3D0BWP12T U910 ( .A1(n560), .B1(n545), .B2(n547), .ZN(n3202) );
  MOAI22D0BWP12T U911 ( .A1(n3030), .A2(n3031), .B1(n3030), .B2(n3031), .ZN(
        n152) );
  AO222D0BWP12T U912 ( .A1(n152), .A2(n3505), .B1(n3499), .B2(next_pc_in[5]), 
        .C1(pc_out[5]), .C2(n3498), .Z(n2173) );
  AOI21D0BWP12T U913 ( .A1(n[3569]), .A2(n3186), .B(reset), .ZN(n153) );
  CKND2D0BWP12T U914 ( .A1(n3184), .A2(write1_in[11]), .ZN(n154) );
  OAI211D0BWP12T U915 ( .A1(n2993), .A2(n2902), .B(n153), .C(n154), .ZN(
        spin[11]) );
  AO222D0BWP12T U916 ( .A1(n3231), .A2(write1_in[12]), .B1(write2_in[12]), 
        .B2(n3232), .C1(r1[12]), .C2(n3233), .Z(n2596) );
  AO222D0BWP12T U917 ( .A1(n3517), .A2(write1_in[13]), .B1(write2_in[13]), 
        .B2(n3218), .C1(r0[13]), .C2(n3219), .Z(n2629) );
  AO222D0BWP12T U918 ( .A1(n3517), .A2(write1_in[14]), .B1(n3218), .B2(
        write2_in[14]), .C1(r0[14]), .C2(n3219), .Z(n2630) );
  AO222D0BWP12T U919 ( .A1(n3517), .A2(write1_in[15]), .B1(n3218), .B2(
        write2_in[15]), .C1(r0[15]), .C2(n3219), .Z(n2631) );
  AO222D0BWP12T U920 ( .A1(n3517), .A2(n3055), .B1(write2_in[16]), .B2(n3218), 
        .C1(r0[16]), .C2(n3219), .Z(n2632) );
  AO222D0BWP12T U921 ( .A1(n3517), .A2(n3054), .B1(n3218), .B2(write2_in[17]), 
        .C1(r0[17]), .C2(n3219), .Z(n2633) );
  AO222D0BWP12T U922 ( .A1(n3517), .A2(n3060), .B1(write2_in[18]), .B2(n3218), 
        .C1(r0[18]), .C2(n3219), .Z(n2634) );
  AO222D0BWP12T U923 ( .A1(n3517), .A2(n3096), .B1(n3218), .B2(write2_in[19]), 
        .C1(r0[19]), .C2(n3219), .Z(n2635) );
  AO222D0BWP12T U924 ( .A1(n3517), .A2(n3095), .B1(n3218), .B2(write2_in[20]), 
        .C1(r0[20]), .C2(n3219), .Z(n2636) );
  AO222D0BWP12T U925 ( .A1(n3517), .A2(n3098), .B1(n3218), .B2(write2_in[21]), 
        .C1(r0[21]), .C2(n3219), .Z(n2637) );
  AO222D0BWP12T U926 ( .A1(n3517), .A2(n3282), .B1(n3218), .B2(write2_in[22]), 
        .C1(r0[22]), .C2(n3219), .Z(n2638) );
  AO222D0BWP12T U927 ( .A1(n3517), .A2(write1_in[23]), .B1(n3218), .B2(
        write2_in[23]), .C1(r0[23]), .C2(n3219), .Z(n2639) );
  AO222D0BWP12T U928 ( .A1(n3517), .A2(n3097), .B1(n3218), .B2(write2_in[24]), 
        .C1(r0[24]), .C2(n3219), .Z(n2640) );
  AO222D0BWP12T U929 ( .A1(n3517), .A2(n3113), .B1(n3218), .B2(write2_in[25]), 
        .C1(r0[25]), .C2(n3219), .Z(n2641) );
  AO222D0BWP12T U930 ( .A1(n3517), .A2(n3108), .B1(n3218), .B2(write2_in[26]), 
        .C1(r0[26]), .C2(n3219), .Z(n2642) );
  NR2XD1BWP12T U931 ( .A1(n3285), .A2(n3497), .ZN(n3290) );
  TPNR2D2BWP12T U932 ( .A1(n1359), .A2(n1357), .ZN(n155) );
  TPNR3D2BWP12T U933 ( .A1(n1358), .A2(n1360), .A3(n156), .ZN(n1366) );
  TPOAI22D2BWP12T U934 ( .A1(n3404), .A2(n1356), .B1(n2909), .B2(n3434), .ZN(
        n1359) );
  TPOAI22D1BWP12T U935 ( .A1(n3414), .A2(n2929), .B1(n1810), .B2(n2932), .ZN(
        n1357) );
  TPND2D2BWP12T U936 ( .A1(n1366), .A2(n1365), .ZN(regA_out[8]) );
  AOI21D2BWP12T U937 ( .A1(write1_in[16]), .A2(n530), .B(n496), .ZN(n157) );
  TPAOI21D1BWP12T U938 ( .A1(write1_in[16]), .A2(n530), .B(n496), .ZN(n3138)
         );
  RCIAO21D0BWP12T U939 ( .A1(n455), .A2(n158), .B(n1397), .ZN(n1399) );
  IOA21D2BWP12T U940 ( .A1(write1_in[25]), .A2(n530), .B(n1128), .ZN(n3311) );
  OR2D2BWP12T U941 ( .A1(n1934), .A2(n3100), .Z(n3110) );
  INVD2P3BWP12T U942 ( .I(n3320), .ZN(n899) );
  TPND2D2BWP12T U943 ( .A1(n335), .A2(n334), .ZN(regB_out[21]) );
  ND2D4BWP12T U944 ( .A1(n1049), .A2(n614), .ZN(n1426) );
  TPND2D4BWP12T U945 ( .A1(n1047), .A2(n1049), .ZN(n224) );
  RCOAI21D1BWP12T U946 ( .A1(n1442), .A2(n3497), .B(n1441), .ZN(n2191) );
  INR2D2BWP12T U947 ( .A1(n1699), .B1(n1700), .ZN(n1701) );
  ND2XD0BWP12T U948 ( .A1(n3412), .A2(r6[4]), .ZN(n740) );
  RCAOI21D1BWP12T U949 ( .A1(n3412), .A2(r6[2]), .B(n1281), .ZN(n1283) );
  AOI21D0BWP12T U950 ( .A1(n3412), .A2(r6[0]), .B(n456), .ZN(n460) );
  RCAOI21D1BWP12T U951 ( .A1(n3412), .A2(r6[12]), .B(n1465), .ZN(n1468) );
  NR2XD1BWP12T U952 ( .A1(n1628), .A2(n1627), .ZN(n1632) );
  AN2XD8BWP12T U953 ( .A1(n212), .A2(readA_sel[0]), .Z(n159) );
  CKND2D2BWP12T U954 ( .A1(n3412), .A2(r6[15]), .ZN(n1376) );
  INVD3BWP12T U955 ( .I(n1674), .ZN(n160) );
  INVD6BWP12T U956 ( .I(n1674), .ZN(n161) );
  INVD4BWP12T U957 ( .I(n1674), .ZN(n1889) );
  NR2D4BWP12T U958 ( .A1(n1911), .A2(n1710), .ZN(n1711) );
  ND2D4BWP12T U959 ( .A1(n1109), .A2(n1108), .ZN(regB_out[15]) );
  MOAI22D1BWP12T U960 ( .A1(n2941), .A2(n1881), .B1(n3419), .B2(r9[9]), .ZN(
        n1185) );
  INVD1BWP12T U961 ( .I(r9[9]), .ZN(n2984) );
  DCCKND4BWP12T U962 ( .I(write1_in[24]), .ZN(n162) );
  TPAOI31D2BWP12T U963 ( .A1(write1_in[23]), .A2(write1_in[24]), .A3(n530), 
        .B(n487), .ZN(n488) );
  INVD8BWP12T U964 ( .I(n168), .ZN(n1911) );
  TPNR2D2BWP12T U965 ( .A1(write1_in[26]), .A2(n888), .ZN(n893) );
  TPAOI21D4BWP12T U966 ( .A1(write1_in[17]), .A2(n530), .B(n495), .ZN(n3250)
         );
  NR2XD1BWP12T U967 ( .A1(n3138), .A2(n881), .ZN(n882) );
  CKND2D2BWP12T U968 ( .A1(n1352), .A2(n1351), .ZN(regB_out[19]) );
  INVD3BWP12T U969 ( .I(n276), .ZN(n1697) );
  BUFFD2BWP12T U970 ( .I(n1705), .Z(n1892) );
  INVD3BWP12T U971 ( .I(n1705), .ZN(n1587) );
  CKND2D2BWP12T U972 ( .A1(n1598), .A2(n1597), .ZN(regB_out[24]) );
  RCOAI22D0BWP12T U973 ( .A1(n1652), .A2(n3070), .B1(n2819), .B2(n1896), .ZN(
        n734) );
  INR2D1BWP12T U974 ( .A1(r3[7]), .B1(n1704), .ZN(n1708) );
  INVD1BWP12T U975 ( .I(n1564), .ZN(n164) );
  INVD6BWP12T U976 ( .I(n296), .ZN(n1571) );
  ND2D3BWP12T U977 ( .A1(n252), .A2(n256), .ZN(n165) );
  CKND2D2BWP12T U978 ( .A1(n252), .A2(n256), .ZN(n276) );
  TPNR3D2BWP12T U979 ( .A1(n819), .A2(n818), .A3(n178), .ZN(n826) );
  DCCKND4BWP12T U980 ( .I(readB_sel[2]), .ZN(n250) );
  CKND0BWP12T U981 ( .I(n1909), .ZN(n167) );
  INVD4BWP12T U982 ( .I(n377), .ZN(n1909) );
  ND2D3BWP12T U983 ( .A1(n3103), .A2(n3102), .ZN(n1934) );
  INVD3BWP12T U984 ( .I(n526), .ZN(n527) );
  TPOAI21D1BWP12T U985 ( .A1(n3284), .A2(n3331), .B(n3283), .ZN(n171) );
  AN2D8BWP12T U986 ( .A1(n281), .A2(n283), .Z(n168) );
  ND2D3BWP12T U987 ( .A1(n1527), .A2(r12[13]), .ZN(n169) );
  CKND2D2BWP12T U988 ( .A1(n1918), .A2(r4[13]), .ZN(n170) );
  BUFFXD4BWP12T U989 ( .I(n753), .Z(n1527) );
  TPOAI21D1BWP12T U990 ( .A1(n1887), .A2(n2869), .B(n955), .ZN(n961) );
  NR4D1BWP12T U991 ( .A1(n1350), .A2(n1349), .A3(n1348), .A4(n1347), .ZN(n1351) );
  NR4D2BWP12T U992 ( .A1(n734), .A2(n733), .A3(n732), .A4(n731), .ZN(n735) );
  NR2XD1BWP12T U993 ( .A1(n1891), .A2(n1890), .ZN(n1906) );
  NR4D1BWP12T U994 ( .A1(n3457), .A2(n3456), .A3(n3455), .A4(n3454), .ZN(n3458) );
  TPNR2D3BWP12T U995 ( .A1(n3442), .A2(n1344), .ZN(n664) );
  OR2D2BWP12T U996 ( .A1(n1240), .A2(n1239), .Z(n1241) );
  ND3D1BWP12T U997 ( .A1(n1459), .A2(n184), .A3(n1458), .ZN(n1460) );
  CKBD4BWP12T U998 ( .I(write1_in[31]), .Z(n3275) );
  TPOAI21D1BWP12T U999 ( .A1(n3284), .A2(n3331), .B(n3283), .ZN(n3286) );
  ND3XD3BWP12T U1000 ( .A1(n3503), .A2(n3327), .A3(n1027), .ZN(n1036) );
  ND3XD3BWP12T U1001 ( .A1(n1552), .A2(n1551), .A3(n1550), .ZN(regB_out[14])
         );
  TPOAI21D4BWP12T U1002 ( .A1(n519), .A2(n3331), .B(n880), .ZN(n1942) );
  DCCKND4BWP12T U1003 ( .I(readB_sel[1]), .ZN(n251) );
  INVD12BWP12T U1004 ( .I(n3419), .ZN(n3402) );
  CKND2D4BWP12T U1005 ( .A1(n281), .A2(n286), .ZN(n1704) );
  AN2XD2BWP12T U1006 ( .A1(n1027), .A2(n3327), .Z(n540) );
  ND2D3BWP12T U1007 ( .A1(n878), .A2(n877), .ZN(n886) );
  TPND2D2BWP12T U1008 ( .A1(n3092), .A2(n3093), .ZN(n3100) );
  RCOAI21D1BWP12T U1009 ( .A1(n1945), .A2(n3497), .B(n1944), .ZN(n2186) );
  XNR2D1BWP12T U1010 ( .A1(n1943), .A2(n1942), .ZN(n1945) );
  TPNR2D1BWP12T U1011 ( .A1(write1_in[27]), .A2(n3318), .ZN(n3319) );
  ND3D0BWP12T U1012 ( .A1(n3327), .A2(n1027), .A3(n3503), .ZN(n534) );
  DCCKND4BWP12T U1013 ( .I(n1622), .ZN(n1787) );
  INVD3BWP12T U1014 ( .I(write1_in[28]), .ZN(n3153) );
  ND2XD4BWP12T U1015 ( .A1(n861), .A2(n1049), .ZN(n3446) );
  MOAI22D1BWP12T U1016 ( .A1(n1519), .A2(n1247), .B1(n168), .B2(r1[26]), .ZN(
        n1249) );
  ND3XD3BWP12T U1017 ( .A1(n852), .A2(n851), .A3(n850), .ZN(regB_out[8]) );
  IND3D2BWP12T U1018 ( .A1(n1029), .B1(n3505), .B2(n173), .ZN(n1032) );
  NR2D2BWP12T U1019 ( .A1(n452), .A2(n451), .ZN(n453) );
  TPAOI21D1BWP12T U1020 ( .A1(write1_in[27]), .A2(n530), .B(n3318), .ZN(n173)
         );
  TPAOI21D1BWP12T U1021 ( .A1(write1_in[27]), .A2(n530), .B(n3318), .ZN(n174)
         );
  NR2D1BWP12T U1022 ( .A1(n1605), .A2(n3497), .ZN(n1599) );
  TPAOI21D4BWP12T U1023 ( .A1(write1_in[27]), .A2(n530), .B(n3318), .ZN(n1028)
         );
  TPND2D2BWP12T U1024 ( .A1(n281), .A2(n280), .ZN(n282) );
  INVD1BWP12T U1025 ( .I(n1726), .ZN(n175) );
  MOAI22D1BWP12T U1026 ( .A1(n1519), .A2(n1209), .B1(n168), .B2(r1[16]), .ZN(
        n299) );
  ND2D4BWP12T U1027 ( .A1(n1026), .A2(n1025), .ZN(regB_out[13]) );
  INR3D4BWP12T U1028 ( .A1(n1906), .B1(n1905), .B2(n1904), .ZN(n1931) );
  IND3D1BWP12T U1029 ( .A1(n1535), .B1(n1534), .B2(n1533), .ZN(n1536) );
  MOAI22D0BWP12T U1030 ( .A1(n1887), .A2(n2947), .B1(n1674), .B2(r5[9]), .ZN(
        n1154) );
  INR2D2BWP12T U1031 ( .A1(r11[6]), .B1(n1887), .ZN(n1891) );
  TPND2D3BWP12T U1032 ( .A1(n281), .A2(n277), .ZN(n307) );
  AOI21D1BWP12T U1033 ( .A1(write1_in[4]), .A2(n530), .B(n509), .ZN(n2938) );
  RCIAO22D1BWP12T U1034 ( .B1(n1918), .B2(r4[4]), .A1(n1920), .A2(n176), .ZN(
        n1164) );
  INVD2BWP12T U1035 ( .I(n753), .ZN(n1920) );
  INVD3BWP12T U1036 ( .I(write1_in[18]), .ZN(n519) );
  ND3XD4BWP12T U1037 ( .A1(n1331), .A2(n1330), .A3(n1329), .ZN(regB_out[28])
         );
  TPOAI22D1BWP12T U1038 ( .A1(n1659), .A2(n915), .B1(n1519), .B2(n914), .ZN(
        n917) );
  TPNR2D3BWP12T U1039 ( .A1(n3110), .A2(n1937), .ZN(n3137) );
  INVD2BWP12T U1040 ( .I(n1256), .ZN(n1257) );
  NR2D2BWP12T U1041 ( .A1(n1266), .A2(n1265), .ZN(n1273) );
  TPND3D2BWP12T U1042 ( .A1(n1259), .A2(n1258), .A3(n1257), .ZN(n1266) );
  RCAOI22D1BWP12T U1043 ( .A1(n1526), .A2(tmp1[4]), .B1(n1571), .B2(r8[4]), 
        .ZN(n1163) );
  RCAOI22D1BWP12T U1044 ( .A1(n1921), .A2(tmp1[3]), .B1(n1571), .B2(r8[3]), 
        .ZN(n1263) );
  TPOAI22D1BWP12T U1045 ( .A1(n1887), .A2(n2802), .B1(n161), .B2(n1614), .ZN(
        n1510) );
  TPOAI22D1BWP12T U1046 ( .A1(n1887), .A2(n3360), .B1(n161), .B2(n3353), .ZN(
        n1078) );
  TPOAI22D1BWP12T U1047 ( .A1(n1887), .A2(n1968), .B1(n161), .B2(n1485), .ZN(
        n1488) );
  TPOAI22D1BWP12T U1048 ( .A1(n1887), .A2(n2963), .B1(n161), .B2(n3005), .ZN(
        n996) );
  ND3XD4BWP12T U1049 ( .A1(n982), .A2(n981), .A3(n980), .ZN(regB_out[5]) );
  CKND2D2BWP12T U1050 ( .A1(n1907), .A2(immediate2_in[6]), .ZN(n1908) );
  ND2D1BWP12T U1051 ( .A1(n1907), .A2(immediate2_in[30]), .ZN(n797) );
  ND2D1BWP12T U1052 ( .A1(n1907), .A2(immediate2_in[13]), .ZN(n1002) );
  OAI21D1BWP12T U1053 ( .A1(n1608), .A2(n1605), .B(n891), .ZN(n913) );
  ND2D4BWP12T U1054 ( .A1(n1664), .A2(r12[2]), .ZN(n1665) );
  OA22D2BWP12T U1055 ( .A1(n1911), .A2(n1334), .B1(n1519), .B2(n1333), .Z(
        n1336) );
  INVD6BWP12T U1056 ( .I(n1703), .ZN(n1575) );
  AOI22D1BWP12T U1057 ( .A1(n1575), .A2(pc_out[15]), .B1(n1915), .B2(r6[15]), 
        .ZN(n1095) );
  MOAI22D0BWP12T U1058 ( .A1(n1486), .A2(n1896), .B1(n1690), .B2(n[3568]), 
        .ZN(n1487) );
  MOAI22D0BWP12T U1059 ( .A1(n1238), .A2(n1896), .B1(n1690), .B2(n[3554]), 
        .ZN(n1239) );
  BUFFD2BWP12T U1060 ( .I(n1690), .Z(n1898) );
  DCCKND4BWP12T U1061 ( .I(n1690), .ZN(n1652) );
  TPNR2D4BWP12T U1062 ( .A1(n1127), .A2(n488), .ZN(n3327) );
  IND3D1BWP12T U1063 ( .A1(n3328), .B1(n3327), .B2(n3339), .ZN(n3329) );
  ND3XD4BWP12T U1064 ( .A1(n1570), .A2(n1569), .A3(n1568), .ZN(regB_out[25])
         );
  DCCKND4BWP12T U1065 ( .I(readB_sel[3]), .ZN(n261) );
  MOAI22D1BWP12T U1066 ( .A1(n1670), .A2(n1669), .B1(n1668), .B2(
        immediate2_in[2]), .ZN(n1671) );
  CKND0BWP12T U1067 ( .I(write1_in[31]), .ZN(n3511) );
  BUFFXD6BWP12T U1068 ( .I(n377), .Z(n1714) );
  INVD2BWP12T U1069 ( .I(n3307), .ZN(n3300) );
  OA22D2BWP12T U1070 ( .A1(n1911), .A2(n447), .B1(n1519), .B2(n446), .Z(n449)
         );
  TPNR2D2BWP12T U1071 ( .A1(n1012), .A2(n1011), .ZN(n1026) );
  INVD6BWP12T U1072 ( .I(n282), .ZN(n1674) );
  TPOAI21D4BWP12T U1073 ( .A1(n524), .A2(n3331), .B(n523), .ZN(n3102) );
  TPOAI21D1BWP12T U1074 ( .A1(n522), .A2(n3331), .B(n521), .ZN(n3103) );
  INVD2BWP12T U1075 ( .I(write1_in[12]), .ZN(n522) );
  TPND2D1BWP12T U1076 ( .A1(n900), .A2(n899), .ZN(n903) );
  INVD2BWP12T U1077 ( .I(n1007), .ZN(n1008) );
  OA22D2BWP12T U1078 ( .A1(n1659), .A2(n1613), .B1(n1519), .B2(n1950), .Z(n183) );
  TPAOI21D1BWP12T U1079 ( .A1(n3290), .A2(n3289), .B(n3288), .ZN(n3291) );
  AO222D0BWP12T U1080 ( .A1(n3246), .A2(write1_in[9]), .B1(n1947), .B2(
        write2_in[9]), .C1(n1946), .C2(tmp1[9]), .Z(n2145) );
  TPND2D3BWP12T U1081 ( .A1(n3057), .A2(n498), .ZN(n502) );
  ND2D4BWP12T U1082 ( .A1(write1_in[9]), .A2(n530), .ZN(n3057) );
  BUFFD3BWP12T U1083 ( .I(n174), .Z(n1038) );
  ND2D3BWP12T U1084 ( .A1(n1524), .A2(n1525), .ZN(regB_out[1]) );
  INVD3BWP12T U1085 ( .I(n3504), .ZN(n3503) );
  TPND2D3BWP12T U1086 ( .A1(n517), .A2(n3107), .ZN(n884) );
  NR2D2BWP12T U1087 ( .A1(n515), .A2(n514), .ZN(n517) );
  NR2D1BWP12T U1088 ( .A1(n370), .A2(n369), .ZN(n1947) );
  INVD2BWP12T U1089 ( .I(n3436), .ZN(n621) );
  INVD1BWP12T U1090 ( .I(n3497), .ZN(n3505) );
  OR2XD1BWP12T U1091 ( .A1(n602), .A2(reset), .Z(n3497) );
  INVD1BWP12T U1092 ( .I(n530), .ZN(n3331) );
  INR2XD2BWP12T U1093 ( .A1(n482), .B1(n544), .ZN(n530) );
  NR2D1BWP12T U1094 ( .A1(n406), .A2(n400), .ZN(n3464) );
  AO22D1BWP12T U1095 ( .A1(n1921), .A2(tmp1[23]), .B1(r8[23]), .B2(n1571), .Z(
        n178) );
  INVD1BWP12T U1096 ( .I(n2704), .ZN(n2803) );
  NR2D1BWP12T U1097 ( .A1(n410), .A2(n403), .ZN(n2704) );
  OR2XD1BWP12T U1098 ( .A1(n1669), .A2(n1974), .Z(n179) );
  INVD1BWP12T U1099 ( .I(pc_out[2]), .ZN(n1679) );
  INVD1BWP12T U1100 ( .I(lr[7]), .ZN(n2767) );
  INVD1BWP12T U1101 ( .I(r2[7]), .ZN(n2849) );
  INVD1BWP12T U1102 ( .I(r3[8]), .ZN(n2909) );
  OA22D1BWP12T U1103 ( .A1(n1652), .A2(n1786), .B1(n1771), .B2(n1896), .Z(n180) );
  AO22D1BWP12T U1104 ( .A1(n1664), .A2(r12[26]), .B1(n1918), .B2(r4[26]), .Z(
        n181) );
  INVD1BWP12T U1105 ( .I(r10[8]), .ZN(n2995) );
  OR2D2BWP12T U1106 ( .A1(n1669), .A2(n1094), .Z(n182) );
  CKND2D2BWP12T U1107 ( .A1(readA_sel[1]), .A2(readA_sel[2]), .ZN(n622) );
  OAI22D1BWP12T U1108 ( .A1(n1519), .A2(n1999), .B1(n1659), .B2(n1658), .ZN(
        n1660) );
  INVD1BWP12T U1109 ( .I(r7[5]), .ZN(n957) );
  INVD1BWP12T U1110 ( .I(r8[7]), .ZN(n2860) );
  OA22D1BWP12T U1111 ( .A1(n1911), .A2(n1457), .B1(n1519), .B2(n1456), .Z(n184) );
  OR2XD1BWP12T U1112 ( .A1(n1714), .A2(n1335), .Z(n185) );
  AN2D1BWP12T U1113 ( .A1(n1069), .A2(r10[13]), .Z(n186) );
  OA22D1BWP12T U1114 ( .A1(n1911), .A2(n374), .B1(n1519), .B2(n373), .Z(n187)
         );
  INVD1BWP12T U1115 ( .I(r7[8]), .ZN(n2931) );
  ND2D1BWP12T U1116 ( .A1(n1862), .A2(n[3575]), .ZN(n188) );
  AN2XD2BWP12T U1117 ( .A1(n1900), .A2(r9[6]), .Z(n189) );
  TPOAI22D1BWP12T U1118 ( .A1(n3416), .A2(n2831), .B1(n2802), .B2(n3393), .ZN(
        n1628) );
  INVD8BWP12T U1119 ( .I(readB_sel[0]), .ZN(n260) );
  DCCKND4BWP12T U1120 ( .I(readA_sel[3]), .ZN(n190) );
  TPNR3D4BWP12T U1121 ( .A1(n190), .A2(readA_sel[0]), .A3(readA_sel[4]), .ZN(
        n200) );
  INVD3BWP12T U1122 ( .I(readA_sel[2]), .ZN(n191) );
  INR2D4BWP12T U1123 ( .A1(readA_sel[1]), .B1(n191), .ZN(n614) );
  CKND2D2BWP12T U1124 ( .A1(n200), .A2(n614), .ZN(n1778) );
  INVD3BWP12T U1125 ( .I(n1778), .ZN(n1219) );
  INVD6BWP12T U1126 ( .I(n1219), .ZN(n3416) );
  INVD1BWP12T U1127 ( .I(lr[22]), .ZN(n378) );
  BUFFXD3BWP12T U1128 ( .I(n200), .Z(n193) );
  INVD4BWP12T U1129 ( .I(readA_sel[1]), .ZN(n192) );
  ND2D4BWP12T U1130 ( .A1(n192), .A2(readA_sel[2]), .ZN(n219) );
  INVD4BWP12T U1131 ( .I(n219), .ZN(n861) );
  INVD1BWP12T U1132 ( .I(r12[22]), .ZN(n194) );
  TPNR3D4BWP12T U1133 ( .A1(readA_sel[4]), .A2(readA_sel[0]), .A3(readA_sel[3]), .ZN(n213) );
  INVD3BWP12T U1134 ( .I(n213), .ZN(n195) );
  NR2XD3BWP12T U1135 ( .A1(n195), .A2(n219), .ZN(n3450) );
  INVD4BWP12T U1136 ( .I(n3450), .ZN(n3390) );
  INVD1BWP12T U1137 ( .I(r4[22]), .ZN(n197) );
  INVD1BWP12T U1138 ( .I(r8[22]), .ZN(n196) );
  TPNR2D3BWP12T U1139 ( .A1(readA_sel[1]), .A2(readA_sel[2]), .ZN(n1047) );
  TPND2D2BWP12T U1140 ( .A1(n200), .A2(n1047), .ZN(n1372) );
  OAI22D1BWP12T U1141 ( .A1(n3390), .A2(n197), .B1(n196), .B2(n1372), .ZN(n210) );
  INVD4BWP12T U1142 ( .I(readA_sel[2]), .ZN(n198) );
  ND2D4BWP12T U1143 ( .A1(n198), .A2(readA_sel[1]), .ZN(n199) );
  INVD6BWP12T U1144 ( .I(n199), .ZN(n225) );
  TPND2D2BWP12T U1145 ( .A1(n225), .A2(n200), .ZN(n201) );
  INVD4BWP12T U1146 ( .I(n201), .ZN(n1069) );
  DCCKND8BWP12T U1147 ( .I(n1069), .ZN(n3452) );
  INVD1BWP12T U1148 ( .I(r10[22]), .ZN(n384) );
  DCCKND4BWP12T U1149 ( .I(n225), .ZN(n202) );
  INVD4BWP12T U1150 ( .I(n202), .ZN(n206) );
  ND2D3BWP12T U1151 ( .A1(readA_sel[3]), .A2(readA_sel[0]), .ZN(n205) );
  INVD3BWP12T U1152 ( .I(readA_sel[4]), .ZN(n203) );
  INVD4BWP12T U1153 ( .I(n203), .ZN(n204) );
  TPNR2D8BWP12T U1154 ( .A1(n205), .A2(n204), .ZN(n1049) );
  ND2D8BWP12T U1155 ( .A1(n206), .A2(n1049), .ZN(n3393) );
  INVD1BWP12T U1156 ( .I(r11[22]), .ZN(n2062) );
  ND2D3BWP12T U1157 ( .A1(n614), .A2(n213), .ZN(n455) );
  BUFFD6BWP12T U1158 ( .I(n455), .Z(n3396) );
  INVD1BWP12T U1159 ( .I(r6[22]), .ZN(n207) );
  TPND2D2BWP12T U1160 ( .A1(n213), .A2(n1047), .ZN(n1617) );
  BUFFD12BWP12T U1161 ( .I(n1617), .Z(n3442) );
  INVD1BWP12T U1162 ( .I(r0[22]), .ZN(n387) );
  OAI22D1BWP12T U1163 ( .A1(n3396), .A2(n207), .B1(n3442), .B2(n387), .ZN(n208) );
  NR4D0BWP12T U1164 ( .A1(n211), .A2(n210), .A3(n209), .A4(n208), .ZN(n230) );
  TPNR2D3BWP12T U1165 ( .A1(readA_sel[4]), .A2(readA_sel[3]), .ZN(n212) );
  ND2D3BWP12T U1166 ( .A1(n159), .A2(n1047), .ZN(n618) );
  BUFFXD6BWP12T U1167 ( .I(n618), .Z(n1810) );
  INVD6BWP12T U1168 ( .I(n1810), .ZN(n3384) );
  AN2D8BWP12T U1169 ( .A1(n225), .A2(n213), .Z(n1622) );
  INVD12BWP12T U1170 ( .I(n1622), .ZN(n3432) );
  INVD1BWP12T U1171 ( .I(r2[22]), .ZN(n373) );
  ND2D1BWP12T U1172 ( .A1(readA_sel[4]), .A2(readA_sel[3]), .ZN(n216) );
  INVD2BWP12T U1173 ( .I(readA_sel[0]), .ZN(n214) );
  INVD2BWP12T U1174 ( .I(n214), .ZN(n215) );
  TPNR2D3BWP12T U1175 ( .A1(n216), .A2(n215), .ZN(n3429) );
  INVD1P75BWP12T U1176 ( .I(n622), .ZN(n217) );
  ND2D4BWP12T U1177 ( .A1(n3429), .A2(n217), .ZN(n1621) );
  BUFFXD6BWP12T U1178 ( .I(n1621), .Z(n3378) );
  INVD1BWP12T U1179 ( .I(tmp1[22]), .ZN(n218) );
  OAI22D1BWP12T U1180 ( .A1(n3432), .A2(n373), .B1(n3378), .B2(n218), .ZN(n223) );
  INVD2P3BWP12T U1181 ( .I(n219), .ZN(n220) );
  ND2D4BWP12T U1182 ( .A1(n159), .A2(n220), .ZN(n1837) );
  INVD3BWP12T U1183 ( .I(n1873), .ZN(n3381) );
  INVD1BWP12T U1184 ( .I(r5[22]), .ZN(n390) );
  INVD1BWP12T U1185 ( .I(r7[22]), .ZN(n386) );
  ND2D3BWP12T U1186 ( .A1(n159), .A2(n614), .ZN(n221) );
  INVD6BWP12T U1187 ( .I(n221), .ZN(n1839) );
  INVD12BWP12T U1188 ( .I(n1839), .ZN(n3444) );
  TPOAI22D1BWP12T U1189 ( .A1(n3381), .A2(n390), .B1(n386), .B2(n3444), .ZN(
        n222) );
  AOI211XD1BWP12T U1190 ( .A1(r1[22]), .A2(n3384), .B(n223), .C(n222), .ZN(
        n229) );
  BUFFXD6BWP12T U1191 ( .I(n3446), .Z(n3404) );
  INVD1BWP12T U1192 ( .I(n[3558]), .ZN(n2063) );
  INVD9BWP12T U1193 ( .I(n224), .ZN(n3419) );
  INVD1BWP12T U1194 ( .I(r9[22]), .ZN(n385) );
  OAI22D1BWP12T U1195 ( .A1(n3404), .A2(n2063), .B1(n3402), .B2(n385), .ZN(
        n227) );
  INVD6BWP12T U1196 ( .I(n1426), .ZN(n3445) );
  INVD4BWP12T U1197 ( .I(n3445), .ZN(n3406) );
  INVD1BWP12T U1198 ( .I(r3[22]), .ZN(n391) );
  TPND2D3BWP12T U1199 ( .A1(n159), .A2(n225), .ZN(n1428) );
  INVD6BWP12T U1200 ( .I(n1428), .ZN(n1646) );
  INVD9BWP12T U1201 ( .I(n1646), .ZN(n3434) );
  OAI22D1BWP12T U1202 ( .A1(n3406), .A2(n3535), .B1(n391), .B2(n3434), .ZN(
        n226) );
  NR2D1BWP12T U1203 ( .A1(n227), .A2(n226), .ZN(n228) );
  INVD1BWP12T U1204 ( .I(lr[27]), .ZN(n1453) );
  INVD1BWP12T U1205 ( .I(r12[27]), .ZN(n231) );
  INVD1BWP12T U1206 ( .I(r4[27]), .ZN(n233) );
  INVD1BWP12T U1207 ( .I(r8[27]), .ZN(n232) );
  BUFFD6BWP12T U1208 ( .I(n1372), .Z(n3435) );
  OAI22D1BWP12T U1209 ( .A1(n3390), .A2(n233), .B1(n232), .B2(n3435), .ZN(n237) );
  INVD1BWP12T U1210 ( .I(r10[27]), .ZN(n1447) );
  INVD1BWP12T U1211 ( .I(r11[27]), .ZN(n2722) );
  INVD1BWP12T U1212 ( .I(r6[27]), .ZN(n234) );
  INVD1BWP12T U1213 ( .I(r0[27]), .ZN(n1445) );
  OAI22D1BWP12T U1214 ( .A1(n3396), .A2(n234), .B1(n3442), .B2(n1445), .ZN(
        n235) );
  NR4D0BWP12T U1215 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .ZN(n249) );
  INVD1BWP12T U1216 ( .I(tmp1[27]), .ZN(n239) );
  INVD1BWP12T U1217 ( .I(r2[27]), .ZN(n1456) );
  OAI22D1BWP12T U1218 ( .A1(n3378), .A2(n239), .B1(n1456), .B2(n3432), .ZN(
        n243) );
  INVD1BWP12T U1219 ( .I(r7[27]), .ZN(n1444) );
  INVD1BWP12T U1220 ( .I(r5[27]), .ZN(n1446) );
  TPND2D2BWP12T U1221 ( .A1(n3384), .A2(r1[27]), .ZN(n240) );
  IND2D2BWP12T U1222 ( .A1(n241), .B1(n240), .ZN(n242) );
  INVD1BWP12T U1223 ( .I(n[3553]), .ZN(n244) );
  INVD1BWP12T U1224 ( .I(r9[27]), .ZN(n1448) );
  OAI22D1BWP12T U1225 ( .A1(n3404), .A2(n244), .B1(n3402), .B2(n1448), .ZN(
        n246) );
  INVD1BWP12T U1226 ( .I(r3[27]), .ZN(n1443) );
  OAI22D1BWP12T U1227 ( .A1(n3406), .A2(n3538), .B1(n1443), .B2(n3434), .ZN(
        n245) );
  NR2D1BWP12T U1228 ( .A1(n246), .A2(n245), .ZN(n247) );
  ND3D2BWP12T U1229 ( .A1(n249), .A2(n248), .A3(n247), .ZN(regA_out[27]) );
  NR2D8BWP12T U1230 ( .A1(n251), .A2(n250), .ZN(n277) );
  INVD6BWP12T U1231 ( .I(n277), .ZN(n964) );
  INVD3BWP12T U1232 ( .I(n964), .ZN(n253) );
  TPNR2D2BWP12T U1233 ( .A1(readB_sel[0]), .A2(readB_sel[3]), .ZN(n252) );
  INVD4BWP12T U1234 ( .I(readB_sel[4]), .ZN(n256) );
  CKND3BWP12T U1235 ( .I(n165), .ZN(n965) );
  ND2D8BWP12T U1236 ( .A1(n253), .A2(n965), .ZN(n1654) );
  IND2D1BWP12T U1237 ( .A1(n1654), .B1(r6[11]), .ZN(n255) );
  INR2D4BWP12T U1238 ( .A1(readB_sel[1]), .B1(readB_sel[2]), .ZN(n286) );
  ND2D4BWP12T U1239 ( .A1(n1697), .A2(n286), .ZN(n1519) );
  TPNR3D4BWP12T U1240 ( .A1(n260), .A2(readB_sel[4]), .A3(readB_sel[3]), .ZN(
        n281) );
  TPNR2D3BWP12T U1241 ( .A1(readB_sel[2]), .A2(readB_sel[1]), .ZN(n283) );
  INVD4BWP12T U1242 ( .I(n168), .ZN(n1659) );
  INVD1BWP12T U1243 ( .I(r1[11]), .ZN(n2882) );
  TPOAI22D1BWP12T U1244 ( .A1(n1519), .A2(n2896), .B1(n1659), .B2(n2882), .ZN(
        n254) );
  BUFFD2BWP12T U1245 ( .I(n277), .Z(n258) );
  NR2D4BWP12T U1246 ( .A1(n260), .A2(n261), .ZN(n257) );
  ND2D4BWP12T U1247 ( .A1(n257), .A2(n256), .ZN(n285) );
  INVD4BWP12T U1248 ( .I(n285), .ZN(n278) );
  ND2D8BWP12T U1249 ( .A1(n258), .A2(n278), .ZN(n1703) );
  BUFFXD6BWP12T U1250 ( .I(n1703), .Z(n1917) );
  ND2D2BWP12T U1251 ( .A1(readB_sel[4]), .A2(readB_sel[3]), .ZN(n266) );
  TPNR3D4BWP12T U1252 ( .A1(n964), .A2(n260), .A3(n266), .ZN(n1713) );
  BUFFXD4BWP12T U1253 ( .I(n1713), .Z(n1668) );
  BUFFXD6BWP12T U1254 ( .I(n1668), .Z(n1567) );
  INVD1BWP12T U1255 ( .I(lr[11]), .ZN(n3027) );
  TPNR3D4BWP12T U1256 ( .A1(n261), .A2(readB_sel[4]), .A3(readB_sel[0]), .ZN(
        n287) );
  TPND2D2BWP12T U1257 ( .A1(n287), .A2(n277), .ZN(n377) );
  INVD2BWP12T U1258 ( .I(n1909), .ZN(n1564) );
  INR2D2BWP12T U1259 ( .A1(lr[11]), .B1(n1564), .ZN(n262) );
  TPAOI21D2BWP12T U1260 ( .A1(immediate2_in[11]), .A2(n1567), .B(n262), .ZN(
        n263) );
  ND3D1BWP12T U1261 ( .A1(n265), .A2(n264), .A3(n263), .ZN(n274) );
  TPND2D2BWP12T U1262 ( .A1(n287), .A2(n283), .ZN(n296) );
  BUFFXD3BWP12T U1263 ( .I(n296), .Z(n1922) );
  INR2D2BWP12T U1264 ( .A1(n260), .B1(n266), .ZN(n267) );
  DCCKND4BWP12T U1265 ( .I(n267), .ZN(n268) );
  INR2D4BWP12T U1266 ( .A1(n277), .B1(n268), .ZN(n1692) );
  BUFFXD6BWP12T U1267 ( .I(n1692), .Z(n1526) );
  AOI22D1BWP12T U1268 ( .A1(n1571), .A2(r8[11]), .B1(tmp1[11]), .B2(n1526), 
        .ZN(n272) );
  CKND3BWP12T U1269 ( .I(readB_sel[2]), .ZN(n269) );
  TPNR2D3BWP12T U1270 ( .A1(n269), .A2(readB_sel[1]), .ZN(n280) );
  AN2XD4BWP12T U1271 ( .A1(n287), .A2(n280), .Z(n753) );
  DCCKND4BWP12T U1272 ( .I(n280), .ZN(n275) );
  BUFFXD12BWP12T U1273 ( .I(n270), .Z(n1918) );
  AOI22D1BWP12T U1274 ( .A1(n1527), .A2(r12[11]), .B1(n1918), .B2(r4[11]), 
        .ZN(n271) );
  TPNR2D1BWP12T U1275 ( .A1(n274), .A2(n273), .ZN(n295) );
  BUFFXD12BWP12T U1276 ( .I(n1704), .Z(n1896) );
  TPNR2D2BWP12T U1277 ( .A1(n285), .A2(n275), .ZN(n1690) );
  IOA22D2BWP12T U1278 ( .B1(n2888), .B2(n1896), .A1(n1898), .A2(n[3569]), .ZN(
        n293) );
  INR2D2BWP12T U1279 ( .A1(n283), .B1(n165), .ZN(n1705) );
  INVD1BWP12T U1280 ( .I(r7[11]), .ZN(n2878) );
  BUFFD6BWP12T U1281 ( .I(n307), .Z(n1724) );
  BUFFXD4BWP12T U1282 ( .I(n286), .Z(n279) );
  ND2D8BWP12T U1283 ( .A1(n278), .A2(n279), .ZN(n1675) );
  BUFFXD16BWP12T U1284 ( .I(n1675), .Z(n1887) );
  INVD1BWP12T U1285 ( .I(r11[11]), .ZN(n3026) );
  INVD1BWP12T U1286 ( .I(r5[11]), .ZN(n2884) );
  OAI22D1BWP12T U1287 ( .A1(n1887), .A2(n3026), .B1(n161), .B2(n2884), .ZN(
        n291) );
  INVD2BWP12T U1288 ( .I(n283), .ZN(n284) );
  TPNR2D2BWP12T U1289 ( .A1(n285), .A2(n284), .ZN(n1691) );
  INVD3BWP12T U1290 ( .I(n1691), .ZN(n1590) );
  BUFFD8BWP12T U1291 ( .I(n1590), .Z(n1663) );
  INVD1BWP12T U1292 ( .I(r9[11]), .ZN(n2875) );
  ND2D3BWP12T U1293 ( .A1(n286), .A2(n287), .ZN(n1507) );
  BUFFXD8BWP12T U1294 ( .I(n1507), .Z(n1899) );
  INR2D4BWP12T U1295 ( .A1(r10[11]), .B1(n1899), .ZN(n288) );
  INVD1P75BWP12T U1296 ( .I(n288), .ZN(n289) );
  TPOAI21D1BWP12T U1297 ( .A1(n1663), .A2(n2875), .B(n289), .ZN(n290) );
  NR4D2BWP12T U1298 ( .A1(n293), .A2(n292), .A3(n291), .A4(n290), .ZN(n294) );
  ND2D2BWP12T U1299 ( .A1(n295), .A2(n294), .ZN(regB_out[11]) );
  BUFFD6BWP12T U1300 ( .I(n1692), .Z(n1921) );
  AOI22D1BWP12T U1301 ( .A1(n1921), .A2(tmp1[16]), .B1(r8[16]), .B2(n1571), 
        .ZN(n305) );
  INVD6BWP12T U1302 ( .I(n1909), .ZN(n1669) );
  INVD1BWP12T U1303 ( .I(lr[16]), .ZN(n2081) );
  NR2D1BWP12T U1304 ( .A1(n1669), .A2(n2081), .ZN(n298) );
  AOI22D1BWP12T U1305 ( .A1(n1527), .A2(r12[16]), .B1(n1918), .B2(r4[16]), 
        .ZN(n297) );
  IND2D1BWP12T U1306 ( .A1(n298), .B1(n297), .ZN(n304) );
  INVD15BWP12T U1307 ( .I(n1654), .ZN(n1915) );
  AOI22D1BWP12T U1308 ( .A1(n1575), .A2(pc_out[16]), .B1(r6[16]), .B2(n1915), 
        .ZN(n302) );
  INVD1BWP12T U1309 ( .I(r2[16]), .ZN(n1209) );
  INVD1P75BWP12T U1310 ( .I(n299), .ZN(n301) );
  ND3D2BWP12T U1311 ( .A1(n302), .A2(n301), .A3(n300), .ZN(n303) );
  INR3XD2BWP12T U1312 ( .A1(n305), .B1(n304), .B2(n303), .ZN(n315) );
  INVD1BWP12T U1313 ( .I(n[3564]), .ZN(n1204) );
  INVD1BWP12T U1314 ( .I(r3[16]), .ZN(n1211) );
  OAI22D1BWP12T U1315 ( .A1(n1652), .A2(n1204), .B1(n1211), .B2(n1896), .ZN(
        n313) );
  INVD0BWP12T U1316 ( .I(r9[16]), .ZN(n306) );
  INVD1BWP12T U1317 ( .I(r10[16]), .ZN(n2082) );
  BUFFD6BWP12T U1318 ( .I(n1507), .Z(n1592) );
  OAI22D1BWP12T U1319 ( .A1(n1663), .A2(n306), .B1(n2082), .B2(n1592), .ZN(
        n312) );
  INVD1BWP12T U1320 ( .I(r0[16]), .ZN(n1223) );
  INVD1BWP12T U1321 ( .I(r7[16]), .ZN(n1222) );
  BUFFD6BWP12T U1322 ( .I(n307), .Z(n1895) );
  INVD1BWP12T U1323 ( .I(r11[16]), .ZN(n309) );
  CKND1BWP12T U1324 ( .I(r5[16]), .ZN(n308) );
  TPOAI22D1BWP12T U1325 ( .A1(n1887), .A2(n309), .B1(n160), .B2(n308), .ZN(
        n310) );
  NR4D1BWP12T U1326 ( .A1(n313), .A2(n312), .A3(n311), .A4(n310), .ZN(n314) );
  ND2D3BWP12T U1327 ( .A1(n315), .A2(n314), .ZN(regB_out[16]) );
  AOI22D1BWP12T U1328 ( .A1(n1921), .A2(tmp1[21]), .B1(r8[21]), .B2(n1571), 
        .ZN(n326) );
  INVD1BWP12T U1329 ( .I(lr[21]), .ZN(n1777) );
  NR2D1BWP12T U1330 ( .A1(n167), .A2(n1777), .ZN(n317) );
  BUFFD6BWP12T U1331 ( .I(n753), .Z(n1664) );
  AOI22D1BWP12T U1332 ( .A1(n1664), .A2(r12[21]), .B1(n1918), .B2(r4[21]), 
        .ZN(n316) );
  AOI22D1BWP12T U1333 ( .A1(n1575), .A2(pc_out[21]), .B1(n1915), .B2(r6[21]), 
        .ZN(n323) );
  CKND1BWP12T U1334 ( .I(r2[21]), .ZN(n319) );
  CKND1BWP12T U1335 ( .I(r1[21]), .ZN(n318) );
  TPOAI22D1BWP12T U1336 ( .A1(n1519), .A2(n319), .B1(n1911), .B2(n318), .ZN(
        n320) );
  INVD1BWP12T U1337 ( .I(n320), .ZN(n322) );
  BUFFD6BWP12T U1338 ( .I(n1713), .Z(n1907) );
  INR3XD2BWP12T U1339 ( .A1(n326), .B1(n325), .B2(n324), .ZN(n335) );
  INVD0BWP12T U1340 ( .I(r11[21]), .ZN(n327) );
  INVD1BWP12T U1341 ( .I(r5[21]), .ZN(n1795) );
  TPOAI22D1BWP12T U1342 ( .A1(n1887), .A2(n327), .B1(n1889), .B2(n1795), .ZN(
        n331) );
  BUFFD6BWP12T U1343 ( .I(n1590), .Z(n1553) );
  CKND1BWP12T U1344 ( .I(r10[21]), .ZN(n3463) );
  TPNR2D1BWP12T U1345 ( .A1(n329), .A2(n328), .ZN(n330) );
  INVD1BWP12T U1346 ( .I(n[3559]), .ZN(n1786) );
  INVD1BWP12T U1347 ( .I(r3[21]), .ZN(n1771) );
  IND3D2BWP12T U1348 ( .A1(n331), .B1(n330), .B2(n180), .ZN(n333) );
  INVD1BWP12T U1349 ( .I(r0[21]), .ZN(n1796) );
  INVD1BWP12T U1350 ( .I(r7[21]), .ZN(n1794) );
  TPOAI22D2BWP12T U1351 ( .A1(n1587), .A2(n1796), .B1(n1794), .B2(n1895), .ZN(
        n332) );
  NR2XD2BWP12T U1352 ( .A1(n333), .A2(n332), .ZN(n334) );
  INVD1BWP12T U1353 ( .I(tmp1[26]), .ZN(n336) );
  INVD1BWP12T U1354 ( .I(r2[26]), .ZN(n1247) );
  OAI22D1BWP12T U1355 ( .A1(n3378), .A2(n336), .B1(n1247), .B2(n3432), .ZN(
        n338) );
  BUFFXD8BWP12T U1356 ( .I(n1837), .Z(n3414) );
  INVD1BWP12T U1357 ( .I(r5[26]), .ZN(n1236) );
  INVD1BWP12T U1358 ( .I(r7[26]), .ZN(n1232) );
  OAI22D1BWP12T U1359 ( .A1(n3414), .A2(n1236), .B1(n1232), .B2(n3444), .ZN(
        n337) );
  AOI211D1BWP12T U1360 ( .A1(r1[26]), .A2(n3384), .B(n338), .C(n337), .ZN(n352) );
  INVD1BWP12T U1361 ( .I(lr[26]), .ZN(n1243) );
  INVD1BWP12T U1362 ( .I(r12[26]), .ZN(n339) );
  INVD1BWP12T U1363 ( .I(r4[26]), .ZN(n341) );
  INVD1BWP12T U1364 ( .I(r8[26]), .ZN(n340) );
  OAI22D1BWP12T U1365 ( .A1(n3390), .A2(n341), .B1(n340), .B2(n3435), .ZN(n345) );
  INVD1BWP12T U1366 ( .I(r11[26]), .ZN(n1237) );
  INVD1BWP12T U1367 ( .I(r10[26]), .ZN(n1230) );
  OAI22D1BWP12T U1368 ( .A1(n3393), .A2(n1237), .B1(n1230), .B2(n3452), .ZN(
        n344) );
  INVD1BWP12T U1369 ( .I(r6[26]), .ZN(n342) );
  INVD1BWP12T U1370 ( .I(r0[26]), .ZN(n1233) );
  OAI22D1BWP12T U1371 ( .A1(n3396), .A2(n342), .B1(n3442), .B2(n1233), .ZN(
        n343) );
  NR4D0BWP12T U1372 ( .A1(n346), .A2(n345), .A3(n344), .A4(n343), .ZN(n351) );
  INVD1BWP12T U1373 ( .I(n[3554]), .ZN(n347) );
  INVD1BWP12T U1374 ( .I(r9[26]), .ZN(n1231) );
  OAI22D1BWP12T U1375 ( .A1(n3404), .A2(n347), .B1(n3402), .B2(n1231), .ZN(
        n349) );
  INVD1BWP12T U1376 ( .I(r3[26]), .ZN(n1238) );
  OAI22D1BWP12T U1377 ( .A1(n3406), .A2(n3537), .B1(n1238), .B2(n3434), .ZN(
        n348) );
  NR2D1BWP12T U1378 ( .A1(n349), .A2(n348), .ZN(n350) );
  INVD4BWP12T U1379 ( .I(reset), .ZN(n3532) );
  AOI211D4BWP12T U1380 ( .A1(n579), .A2(n554), .B(n3231), .C(reset), .ZN(n3233) );
  AOI22D0BWP12T U1381 ( .A1(n3233), .A2(r1[31]), .B1(write2_in[31]), .B2(n3232), .ZN(n353) );
  CKND2D1BWP12T U1382 ( .A1(n354), .A2(n353), .ZN(n2615) );
  INR2D1BWP12T U1383 ( .A1(write1_sel[2]), .B1(write1_sel[1]), .ZN(n584) );
  INVD1BWP12T U1384 ( .I(write1_sel[0]), .ZN(n365) );
  INVD4BWP12T U1385 ( .I(n2872), .ZN(n3184) );
  AOI22D0BWP12T U1386 ( .A1(n3186), .A2(n[3549]), .B1(write2_in[31]), .B2(
        n3185), .ZN(n356) );
  CKND2D1BWP12T U1387 ( .A1(n357), .A2(n356), .ZN(spin[31]) );
  TPNR2D3BWP12T U1388 ( .A1(n585), .A2(n420), .ZN(n3516) );
  NR2D3BWP12T U1389 ( .A1(n420), .A2(n544), .ZN(n3522) );
  INVD1BWP12T U1390 ( .I(r6[1]), .ZN(n1514) );
  OAI222D1BWP12T U1391 ( .A1(n1514), .A2(n3008), .B1(n1953), .B2(n3007), .C1(
        n1954), .C2(n3006), .ZN(n2425) );
  INVD1BWP12T U1392 ( .I(lr[1]), .ZN(n2831) );
  OAI222D1BWP12T U1393 ( .A1(n2831), .A2(n3022), .B1(n1953), .B2(n3020), .C1(
        n1954), .C2(n3018), .ZN(n2201) );
  OAI222D1BWP12T U1394 ( .A1(n1614), .A2(n3004), .B1(n1953), .B2(n3003), .C1(
        n1954), .C2(n3002), .ZN(n2457) );
  INVD1BWP12T U1395 ( .I(r7[1]), .ZN(n1612) );
  OAI222D1BWP12T U1396 ( .A1(n1612), .A2(n3000), .B1(n1953), .B2(n2999), .C1(
        n1954), .C2(n2998), .ZN(n2393) );
  ND4D1BWP12T U1397 ( .A1(write1_sel[3]), .A2(write1_sel[4]), .A3(write1_en), 
        .A4(n365), .ZN(n367) );
  NR2D3BWP12T U1398 ( .A1(n366), .A2(n367), .ZN(n3246) );
  CKND0BWP12T U1399 ( .I(n482), .ZN(n368) );
  OAI21D1BWP12T U1400 ( .A1(n368), .A2(n367), .B(n3532), .ZN(n370) );
  AO222D1BWP12T U1401 ( .A1(n3246), .A2(write1_in[5]), .B1(n1947), .B2(
        write2_in[5]), .C1(n1946), .C2(tmp1[5]), .Z(n2141) );
  AO222D1BWP12T U1402 ( .A1(n3246), .A2(n166), .B1(n1947), .B2(write2_in[8]), 
        .C1(n1946), .C2(tmp1[8]), .Z(n2144) );
  OAI222D1BWP12T U1403 ( .A1(n1672), .A2(n3000), .B1(n2003), .B2(n2999), .C1(
        n2004), .C2(n2998), .ZN(n2394) );
  INVD1BWP12T U1404 ( .I(r6[2]), .ZN(n1653) );
  OAI222D1BWP12T U1405 ( .A1(n1653), .A2(n3008), .B1(n2003), .B2(n3007), .C1(
        n2004), .C2(n3006), .ZN(n2426) );
  INVD1BWP12T U1406 ( .I(r5[2]), .ZN(n1278) );
  OAI222D1BWP12T U1407 ( .A1(n1278), .A2(n3004), .B1(n2003), .B2(n3003), .C1(
        n2004), .C2(n3002), .ZN(n2458) );
  AO222D1BWP12T U1408 ( .A1(n3246), .A2(write1_in[4]), .B1(n1947), .B2(
        write2_in[4]), .C1(n1946), .C2(tmp1[4]), .Z(n2140) );
  AOI21D0BWP12T U1409 ( .A1(n3185), .A2(write2_in[2]), .B(reset), .ZN(n372) );
  TPND2D0BWP12T U1410 ( .A1(n3186), .A2(n[3578]), .ZN(n371) );
  OAI211D1BWP12T U1411 ( .A1(n2872), .A2(n2003), .B(n372), .C(n371), .ZN(
        spin[2]) );
  INVD1BWP12T U1412 ( .I(lr[2]), .ZN(n1670) );
  OAI222D1BWP12T U1413 ( .A1(n1670), .A2(n3022), .B1(n2003), .B2(n3020), .C1(
        n2004), .C2(n3018), .ZN(n2202) );
  AOI22D1BWP12T U1414 ( .A1(n1921), .A2(tmp1[22]), .B1(r8[22]), .B2(n1571), 
        .ZN(n376) );
  CKND1BWP12T U1415 ( .I(r1[22]), .ZN(n374) );
  AOI22D1BWP12T U1416 ( .A1(n1664), .A2(r12[22]), .B1(n1918), .B2(r4[22]), 
        .ZN(n375) );
  ND3D1BWP12T U1417 ( .A1(n376), .A2(n187), .A3(n375), .ZN(n383) );
  AOI22D1BWP12T U1418 ( .A1(n1575), .A2(pc_out[22]), .B1(r6[22]), .B2(n1915), 
        .ZN(n381) );
  TPNR2D2BWP12T U1419 ( .A1(n383), .A2(n382), .ZN(n397) );
  OAI22D1BWP12T U1420 ( .A1(n1553), .A2(n385), .B1(n384), .B2(n1592), .ZN(n389) );
  OAI22D1BWP12T U1421 ( .A1(n1587), .A2(n387), .B1(n386), .B2(n1895), .ZN(n388) );
  OR2XD2BWP12T U1422 ( .A1(n389), .A2(n388), .Z(n395) );
  OAI22D1BWP12T U1423 ( .A1(n1652), .A2(n2063), .B1(n391), .B2(n1896), .ZN(
        n392) );
  OR2XD2BWP12T U1424 ( .A1(n393), .A2(n392), .Z(n394) );
  NR2D2BWP12T U1425 ( .A1(n395), .A2(n394), .ZN(n396) );
  ND2D2BWP12T U1426 ( .A1(n397), .A2(n396), .ZN(regB_out[22]) );
  ND2D1BWP12T U1427 ( .A1(readC_sel[1]), .A2(readC_sel[0]), .ZN(n410) );
  ND3D1BWP12T U1428 ( .A1(readC_sel[2]), .A2(readC_sel[3]), .A3(n3492), .ZN(
        n400) );
  OR2XD1BWP12T U1429 ( .A1(n410), .A2(n400), .Z(n2806) );
  INVD1BWP12T U1430 ( .I(readC_sel[1]), .ZN(n399) );
  INVD1BWP12T U1431 ( .I(readC_sel[0]), .ZN(n398) );
  ND2D1BWP12T U1432 ( .A1(n399), .A2(n398), .ZN(n408) );
  OR2XD1BWP12T U1433 ( .A1(n408), .A2(n400), .Z(n2744) );
  AOI22D0BWP12T U1434 ( .A1(pc_out[4]), .A2(n3480), .B1(n3479), .B2(r12[4]), 
        .ZN(n418) );
  ND2D1BWP12T U1435 ( .A1(readC_sel[1]), .A2(n398), .ZN(n407) );
  INVD1BWP12T U1436 ( .I(readC_sel[3]), .ZN(n405) );
  OR2XD1BWP12T U1437 ( .A1(n407), .A2(n403), .Z(n3478) );
  INVD1BWP12T U1438 ( .I(n3473), .ZN(n2779) );
  INVD1BWP12T U1439 ( .I(lr[4]), .ZN(n2843) );
  INVD1BWP12T U1440 ( .I(r11[4]), .ZN(n2011) );
  OAI22D0BWP12T U1441 ( .A1(n2779), .A2(n2843), .B1(n2011), .B2(n2803), .ZN(
        n402) );
  INVD1BWP12T U1442 ( .I(n[3576]), .ZN(n1178) );
  ND2D1BWP12T U1443 ( .A1(readC_sel[0]), .A2(n399), .ZN(n406) );
  INVD1BWP12T U1444 ( .I(n3464), .ZN(n3474) );
  INVD1BWP12T U1445 ( .I(n3475), .ZN(n2805) );
  INVD1BWP12T U1446 ( .I(r9[4]), .ZN(n2842) );
  OAI22D0BWP12T U1447 ( .A1(n1178), .A2(n3474), .B1(n2805), .B2(n2842), .ZN(
        n401) );
  AOI211D0BWP12T U1448 ( .A1(n2810), .A2(r10[4]), .B(n402), .C(n401), .ZN(n417) );
  OR2XD1BWP12T U1449 ( .A1(n408), .A2(n403), .Z(n2800) );
  ND2D1BWP12T U1450 ( .A1(readC_sel[2]), .A2(n405), .ZN(n404) );
  NR2D1BWP12T U1451 ( .A1(n407), .A2(n404), .ZN(n2770) );
  AOI22D0BWP12T U1452 ( .A1(r5[4]), .A2(n3481), .B1(n2770), .B2(r6[4]), .ZN(
        n414) );
  NR2D1BWP12T U1453 ( .A1(n408), .A2(n404), .ZN(n2757) );
  AOI22D0BWP12T U1454 ( .A1(r7[4]), .A2(n3482), .B1(n2757), .B2(r4[4]), .ZN(
        n413) );
  IND2D1BWP12T U1455 ( .A1(readC_sel[2]), .B1(n405), .ZN(n409) );
  AOI22D0BWP12T U1456 ( .A1(r1[4]), .A2(n3484), .B1(n3483), .B2(r2[4]), .ZN(
        n412) );
  AOI22D0BWP12T U1457 ( .A1(r0[4]), .A2(n3486), .B1(n3485), .B2(r3[4]), .ZN(
        n411) );
  ND4D1BWP12T U1458 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(n415) );
  AOI22D0BWP12T U1459 ( .A1(n3493), .A2(r8[4]), .B1(n3492), .B2(n415), .ZN(
        n416) );
  ND3D1BWP12T U1460 ( .A1(n418), .A2(n417), .A3(n416), .ZN(regC_out[4]) );
  INVD1P75BWP12T U1461 ( .I(r1[7]), .ZN(n1710) );
  OAI222D1BWP12T U1462 ( .A1(n1710), .A2(n3012), .B1(n2866), .B2(n3011), .C1(
        n2867), .C2(n3010), .ZN(n2591) );
  INVD1BWP12T U1463 ( .I(r5[7]), .ZN(n1693) );
  OAI222D1BWP12T U1464 ( .A1(n1693), .A2(n3004), .B1(n2866), .B2(n3003), .C1(
        n2867), .C2(n3002), .ZN(n2463) );
  OAI222D1BWP12T U1465 ( .A1(n1723), .A2(n3000), .B1(n2866), .B2(n2999), .C1(
        n2867), .C2(n2998), .ZN(n2399) );
  CKND0BWP12T U1466 ( .I(r9[7]), .ZN(n423) );
  OAI222D1BWP12T U1467 ( .A1(n423), .A2(n3016), .B1(n2866), .B2(n3015), .C1(
        n2867), .C2(n3014), .ZN(n2335) );
  INVD1BWP12T U1468 ( .I(r6[7]), .ZN(n1698) );
  OAI222D1BWP12T U1469 ( .A1(n1698), .A2(n3008), .B1(n2866), .B2(n3007), .C1(
        n2867), .C2(n3006), .ZN(n2431) );
  OAI222D1BWP12T U1470 ( .A1(n2767), .A2(n3022), .B1(n2866), .B2(n3020), .C1(
        n2867), .C2(n3018), .ZN(n2207) );
  INVD0BWP12T U1471 ( .I(r5[5]), .ZN(n424) );
  OAI222D1BWP12T U1472 ( .A1(n424), .A2(n3004), .B1(n2022), .B2(n3003), .C1(
        n2023), .C2(n3002), .ZN(n2461) );
  INVD0BWP12T U1473 ( .I(r9[5]), .ZN(n2733) );
  OAI222D1BWP12T U1474 ( .A1(n2733), .A2(n3016), .B1(n2022), .B2(n3015), .C1(
        n2023), .C2(n3014), .ZN(n2333) );
  TPAOI21D0BWP12T U1475 ( .A1(n3185), .A2(write2_in[3]), .B(reset), .ZN(n426)
         );
  TPND2D0BWP12T U1476 ( .A1(n3186), .A2(n[3577]), .ZN(n425) );
  OAI211D1BWP12T U1477 ( .A1(n2872), .A2(n1961), .B(n426), .C(n425), .ZN(
        spin[3]) );
  INVD1BWP12T U1478 ( .I(r6[5]), .ZN(n966) );
  OAI222D1BWP12T U1479 ( .A1(n966), .A2(n3008), .B1(n2022), .B2(n3007), .C1(
        n2023), .C2(n3006), .ZN(n2429) );
  INVD1BWP12T U1480 ( .I(r7[6]), .ZN(n1894) );
  OAI222D1BWP12T U1481 ( .A1(n1894), .A2(n3000), .B1(n2031), .B2(n2999), .C1(
        n2032), .C2(n2998), .ZN(n2398) );
  INVD1BWP12T U1482 ( .I(r5[3]), .ZN(n1811) );
  OAI222D1BWP12T U1483 ( .A1(n1811), .A2(n3004), .B1(n1961), .B2(n3003), .C1(
        n1962), .C2(n3002), .ZN(n2459) );
  OAI222D1BWP12T U1484 ( .A1(n1816), .A2(n3016), .B1(n1961), .B2(n3015), .C1(
        n1962), .C2(n3014), .ZN(n2331) );
  INVD1BWP12T U1485 ( .I(r7[3]), .ZN(n1807) );
  OAI222D1BWP12T U1486 ( .A1(n1807), .A2(n3000), .B1(n1961), .B2(n2999), .C1(
        n1962), .C2(n2998), .ZN(n2395) );
  OAI222D1BWP12T U1487 ( .A1(n957), .A2(n3000), .B1(n2022), .B2(n2999), .C1(
        n2023), .C2(n2998), .ZN(n2397) );
  INVD1BWP12T U1488 ( .I(r9[1]), .ZN(n2804) );
  OAI222D1BWP12T U1489 ( .A1(n2804), .A2(n3016), .B1(n1953), .B2(n3015), .C1(
        n1954), .C2(n3014), .ZN(n2329) );
  INVD1BWP12T U1490 ( .I(r1[1]), .ZN(n1613) );
  OAI222D1BWP12T U1491 ( .A1(n1613), .A2(n3012), .B1(n1953), .B2(n3011), .C1(
        n1954), .C2(n3010), .ZN(n2585) );
  OAI222D1BWP12T U1492 ( .A1(n1413), .A2(n3022), .B1(n2031), .B2(n3020), .C1(
        n2032), .C2(n3018), .ZN(n2206) );
  INVD1BWP12T U1493 ( .I(lr[5]), .ZN(n975) );
  OAI222D1BWP12T U1494 ( .A1(n975), .A2(n3022), .B1(n2022), .B2(n3020), .C1(
        n2023), .C2(n3018), .ZN(n2205) );
  INVD1BWP12T U1495 ( .I(lr[3]), .ZN(n2851) );
  OAI222D1BWP12T U1496 ( .A1(n2851), .A2(n3022), .B1(n1961), .B2(n3020), .C1(
        n1962), .C2(n3018), .ZN(n2203) );
  TPAOI21D0BWP12T U1497 ( .A1(n3185), .A2(write2_in[5]), .B(reset), .ZN(n428)
         );
  TPND2D0BWP12T U1498 ( .A1(n3186), .A2(n[3575]), .ZN(n427) );
  OAI211D1BWP12T U1499 ( .A1(n2872), .A2(n2022), .B(n428), .C(n427), .ZN(
        spin[5]) );
  INVD0BWP12T U1500 ( .I(r9[6]), .ZN(n2873) );
  OAI222D1BWP12T U1501 ( .A1(n2873), .A2(n3016), .B1(n2031), .B2(n3015), .C1(
        n2032), .C2(n3014), .ZN(n2334) );
  CKND0BWP12T U1502 ( .I(r6[3]), .ZN(n429) );
  OAI222D1BWP12T U1503 ( .A1(n429), .A2(n3008), .B1(n1961), .B2(n3007), .C1(
        n1962), .C2(n3006), .ZN(n2427) );
  CKND0BWP12T U1504 ( .I(r6[6]), .ZN(n430) );
  OAI222D1BWP12T U1505 ( .A1(n430), .A2(n3008), .B1(n2031), .B2(n3007), .C1(
        n2032), .C2(n3006), .ZN(n2430) );
  INVD1BWP12T U1506 ( .I(r1[5]), .ZN(n976) );
  OAI222D1BWP12T U1507 ( .A1(n976), .A2(n3012), .B1(n2022), .B2(n3011), .C1(
        n2023), .C2(n3010), .ZN(n2589) );
  OAI222D1BWP12T U1508 ( .A1(n1809), .A2(n3012), .B1(n1961), .B2(n3011), .C1(
        n1962), .C2(n3010), .ZN(n2587) );
  INVD1BWP12T U1509 ( .I(r1[6]), .ZN(n1910) );
  OAI222D1BWP12T U1510 ( .A1(n1910), .A2(n3012), .B1(n2031), .B2(n3011), .C1(
        n2032), .C2(n3010), .ZN(n2590) );
  INVD1BWP12T U1511 ( .I(r5[6]), .ZN(n1888) );
  OAI222D1BWP12T U1512 ( .A1(n1888), .A2(n3004), .B1(n2031), .B2(n3003), .C1(
        n2032), .C2(n3002), .ZN(n2462) );
  OAI222D1BWP12T U1513 ( .A1(n2843), .A2(n3022), .B1(n2014), .B2(n3020), .C1(
        n2015), .C2(n3018), .ZN(n2204) );
  INVD0BWP12T U1514 ( .I(r6[4]), .ZN(n431) );
  OAI222D1BWP12T U1515 ( .A1(n431), .A2(n3008), .B1(n2014), .B2(n3007), .C1(
        n2015), .C2(n3006), .ZN(n2428) );
  INVD1BWP12T U1516 ( .I(r1[4]), .ZN(n1174) );
  OAI222D1BWP12T U1517 ( .A1(n1174), .A2(n3012), .B1(n2014), .B2(n3011), .C1(
        n2015), .C2(n3010), .ZN(n2588) );
  AO222D0BWP12T U1518 ( .A1(n3246), .A2(write1_in[6]), .B1(n1947), .B2(
        write2_in[6]), .C1(n1946), .C2(tmp1[6]), .Z(n2142) );
  TPAOI21D0BWP12T U1519 ( .A1(n3185), .A2(write2_in[4]), .B(reset), .ZN(n433)
         );
  TPND2D0BWP12T U1520 ( .A1(n3186), .A2(n[3576]), .ZN(n432) );
  OAI211D1BWP12T U1521 ( .A1(n2872), .A2(n2014), .B(n433), .C(n432), .ZN(
        spin[4]) );
  OAI222D1BWP12T U1522 ( .A1(n2842), .A2(n3016), .B1(n2014), .B2(n3015), .C1(
        n2015), .C2(n3014), .ZN(n2332) );
  INVD1BWP12T U1523 ( .I(r5[4]), .ZN(n741) );
  OAI222D1BWP12T U1524 ( .A1(n741), .A2(n3004), .B1(n2014), .B2(n3003), .C1(
        n2015), .C2(n3002), .ZN(n2460) );
  INVD1BWP12T U1525 ( .I(r7[4]), .ZN(n1177) );
  OAI222D1BWP12T U1526 ( .A1(n1177), .A2(n3000), .B1(n2014), .B2(n2999), .C1(
        n2015), .C2(n2998), .ZN(n2396) );
  OAI222D1BWP12T U1527 ( .A1(n730), .A2(n3004), .B1(n2825), .B2(n3003), .C1(
        n2826), .C2(n3002), .ZN(n2456) );
  INVD1BWP12T U1528 ( .I(r1[0]), .ZN(n716) );
  OAI222D1BWP12T U1529 ( .A1(n716), .A2(n3012), .B1(n2825), .B2(n3011), .C1(
        n2826), .C2(n3010), .ZN(n2584) );
  INVD1BWP12T U1530 ( .I(lr[0]), .ZN(n715) );
  OAI222D1BWP12T U1531 ( .A1(n715), .A2(n3022), .B1(n2825), .B2(n3020), .C1(
        n2826), .C2(n3018), .ZN(n2200) );
  INVD1BWP12T U1532 ( .I(r7[0]), .ZN(n729) );
  OAI222D1BWP12T U1533 ( .A1(n729), .A2(n3000), .B1(n2825), .B2(n2999), .C1(
        n2826), .C2(n2998), .ZN(n2392) );
  CKND0BWP12T U1534 ( .I(r6[0]), .ZN(n434) );
  OAI222D1BWP12T U1535 ( .A1(n434), .A2(n3008), .B1(n2825), .B2(n3007), .C1(
        n2826), .C2(n3006), .ZN(n2424) );
  INVD1BWP12T U1536 ( .I(r1[2]), .ZN(n1658) );
  OAI222D1BWP12T U1537 ( .A1(n1658), .A2(n3012), .B1(n2003), .B2(n3011), .C1(
        n2004), .C2(n3010), .ZN(n2586) );
  OAI222D1BWP12T U1538 ( .A1(n2855), .A2(n3016), .B1(n2003), .B2(n3015), .C1(
        n2004), .C2(n3014), .ZN(n2330) );
  OAI222D1BWP12T U1539 ( .A1(n2711), .A2(n3016), .B1(n2825), .B2(n3015), .C1(
        n2826), .C2(n3014), .ZN(n2328) );
  CKND0BWP12T U1540 ( .I(r9[17]), .ZN(n2038) );
  INVD1BWP12T U1541 ( .I(r10[17]), .ZN(n603) );
  OAI22D1BWP12T U1542 ( .A1(n1663), .A2(n2038), .B1(n603), .B2(n1592), .ZN(
        n439) );
  CKND1BWP12T U1543 ( .I(n[3563]), .ZN(n2039) );
  CKND0BWP12T U1544 ( .I(r3[17]), .ZN(n435) );
  OAI22D1BWP12T U1545 ( .A1(n1652), .A2(n2039), .B1(n435), .B2(n1896), .ZN(
        n437) );
  INVD1BWP12T U1546 ( .I(r11[17]), .ZN(n604) );
  INVD1BWP12T U1547 ( .I(r5[17]), .ZN(n606) );
  INVD1BWP12T U1548 ( .I(r0[17]), .ZN(n440) );
  INVD1BWP12T U1549 ( .I(r7[17]), .ZN(n609) );
  OAI22D1BWP12T U1550 ( .A1(n1587), .A2(n440), .B1(n609), .B2(n1895), .ZN(n441) );
  TPNR2D2BWP12T U1551 ( .A1(n442), .A2(n441), .ZN(n454) );
  AOI22D1BWP12T U1552 ( .A1(n1575), .A2(pc_out[17]), .B1(r6[17]), .B2(n1915), 
        .ZN(n445) );
  AOI22D1BWP12T U1553 ( .A1(n1527), .A2(r12[17]), .B1(n1918), .B2(r4[17]), 
        .ZN(n444) );
  INVD1BWP12T U1554 ( .I(lr[17]), .ZN(n610) );
  AOI22D1BWP12T U1555 ( .A1(n1526), .A2(tmp1[17]), .B1(r8[17]), .B2(n1571), 
        .ZN(n450) );
  CKND1BWP12T U1556 ( .I(r1[17]), .ZN(n447) );
  CKND1BWP12T U1557 ( .I(r2[17]), .ZN(n446) );
  ND3D2BWP12T U1558 ( .A1(n450), .A2(n449), .A3(n448), .ZN(n451) );
  TPND2D2BWP12T U1559 ( .A1(n454), .A2(n453), .ZN(regB_out[17]) );
  INVD4BWP12T U1560 ( .I(n455), .ZN(n3412) );
  INVD1P75BWP12T U1561 ( .I(r2[0]), .ZN(n2824) );
  INVD4BWP12T U1562 ( .I(n1621), .ZN(n1876) );
  ND3D1BWP12T U1563 ( .A1(readA_sel[1]), .A2(readA_sel[0]), .A3(readA_sel[3]), 
        .ZN(n458) );
  ND2D1BWP12T U1564 ( .A1(readA_sel[2]), .A2(readA_sel[4]), .ZN(n457) );
  TPNR2D3BWP12T U1565 ( .A1(n458), .A2(n457), .ZN(n1804) );
  AOI22D1BWP12T U1566 ( .A1(n1876), .A2(tmp1[0]), .B1(n1804), .B2(
        immediate1_in[0]), .ZN(n459) );
  ND2D1BWP12T U1567 ( .A1(n460), .A2(n459), .ZN(n464) );
  INVD1BWP12T U1568 ( .I(n[3580]), .ZN(n3070) );
  INVD1BWP12T U1569 ( .I(r3[0]), .ZN(n2819) );
  OAI22D1BWP12T U1570 ( .A1(n3404), .A2(n3070), .B1(n2819), .B2(n3434), .ZN(
        n463) );
  INVD1BWP12T U1571 ( .I(pc_out[0]), .ZN(n721) );
  OAI22D1BWP12T U1572 ( .A1(n3406), .A2(n721), .B1(n729), .B2(n3444), .ZN(n462) );
  OAI22D1BWP12T U1573 ( .A1(n3414), .A2(n730), .B1(n1810), .B2(n716), .ZN(n461) );
  NR4D0BWP12T U1574 ( .A1(n464), .A2(n463), .A3(n462), .A4(n461), .ZN(n470) );
  OAI22D1BWP12T U1575 ( .A1(n3416), .A2(n715), .B1(n3393), .B2(n3067), .ZN(
        n468) );
  INVD1BWP12T U1576 ( .I(r4[0]), .ZN(n2822) );
  INVD1BWP12T U1577 ( .I(r0[0]), .ZN(n2821) );
  OAI22D1BWP12T U1578 ( .A1(n3390), .A2(n2822), .B1(n2821), .B2(n3442), .ZN(
        n467) );
  INVD1BWP12T U1579 ( .I(r8[0]), .ZN(n2823) );
  INVD4BWP12T U1580 ( .I(n1372), .ZN(n1473) );
  INVD4BWP12T U1581 ( .I(n1473), .ZN(n3387) );
  INVD1BWP12T U1582 ( .I(r12[0]), .ZN(n2820) );
  OAI22D0BWP12T U1583 ( .A1(n2823), .A2(n3387), .B1(n3436), .B2(n2820), .ZN(
        n466) );
  INVD1BWP12T U1584 ( .I(r10[0]), .ZN(n3065) );
  OAI22D1BWP12T U1585 ( .A1(n3402), .A2(n2711), .B1(n3065), .B2(n1881), .ZN(
        n465) );
  NR4D0BWP12T U1586 ( .A1(n468), .A2(n467), .A3(n466), .A4(n465), .ZN(n469) );
  CKND2D1BWP12T U1587 ( .A1(n470), .A2(n469), .ZN(regA_out[0]) );
  AOI22D0BWP12T U1588 ( .A1(n[3554]), .A2(n3464), .B1(n3479), .B2(r12[26]), 
        .ZN(n481) );
  AOI22D0BWP12T U1589 ( .A1(lr[26]), .A2(n3473), .B1(r11[26]), .B2(n2704), 
        .ZN(n472) );
  CKND2D0BWP12T U1590 ( .A1(r9[26]), .A2(n3475), .ZN(n471) );
  OAI211D0BWP12T U1591 ( .A1(n2806), .A2(n3537), .B(n472), .C(n471), .ZN(n473)
         );
  AOI21D0BWP12T U1592 ( .A1(r10[26]), .A2(n2810), .B(n473), .ZN(n480) );
  AOI22D0BWP12T U1593 ( .A1(r5[26]), .A2(n3481), .B1(n2770), .B2(r6[26]), .ZN(
        n477) );
  AOI22D0BWP12T U1594 ( .A1(r7[26]), .A2(n3482), .B1(n2757), .B2(r4[26]), .ZN(
        n476) );
  AOI22D0BWP12T U1595 ( .A1(r1[26]), .A2(n3484), .B1(n3483), .B2(r2[26]), .ZN(
        n475) );
  AOI22D0BWP12T U1596 ( .A1(r0[26]), .A2(n3486), .B1(n3485), .B2(r3[26]), .ZN(
        n474) );
  ND4D1BWP12T U1597 ( .A1(n477), .A2(n476), .A3(n475), .A4(n474), .ZN(n478) );
  AOI22D0BWP12T U1598 ( .A1(n3493), .A2(r8[26]), .B1(n3492), .B2(n478), .ZN(
        n479) );
  ND3D1BWP12T U1599 ( .A1(n481), .A2(n480), .A3(n479), .ZN(regC_out[26]) );
  ND3XD4BWP12T U1600 ( .A1(write1_in[19]), .A2(write1_in[20]), .A3(n530), .ZN(
        n483) );
  CKND3BWP12T U1601 ( .I(n483), .ZN(n486) );
  ND4D0BWP12T U1602 ( .A1(write2_in[22]), .A2(write2_in[21]), .A3(
        write2_in[19]), .A4(write2_in[20]), .ZN(n484) );
  NR2D1BWP12T U1603 ( .A1(n530), .A2(n484), .ZN(n485) );
  TPAOI31D2BWP12T U1604 ( .A1(n486), .A2(write1_in[22]), .A3(write1_in[21]), 
        .B(n485), .ZN(n1127) );
  AN3D2BWP12T U1605 ( .A1(n3331), .A2(write2_in[23]), .A3(write2_in[24]), .Z(
        n487) );
  INVD3BWP12T U1606 ( .I(write1_in[25]), .ZN(n489) );
  INR2D2BWP12T U1607 ( .A1(n530), .B1(n489), .ZN(n490) );
  TPND2D2BWP12T U1608 ( .A1(n490), .A2(write1_in[26]), .ZN(n493) );
  CKND0BWP12T U1609 ( .I(write2_in[25]), .ZN(n491) );
  INR2D1BWP12T U1610 ( .A1(write2_in[26]), .B1(n491), .ZN(n492) );
  ND2D1BWP12T U1611 ( .A1(n3331), .A2(n492), .ZN(n887) );
  TPND2D2BWP12T U1612 ( .A1(n493), .A2(n887), .ZN(n1027) );
  INVD1BWP12T U1613 ( .I(write2_in[17]), .ZN(n494) );
  NR2D1BWP12T U1614 ( .A1(n530), .A2(n494), .ZN(n495) );
  INR2D1BWP12T U1615 ( .A1(write2_in[16]), .B1(n530), .ZN(n496) );
  NR2XD2BWP12T U1616 ( .A1(n3250), .A2(n157), .ZN(n497) );
  INVD1P75BWP12T U1617 ( .I(n497), .ZN(n518) );
  INR2D0BWP12T U1618 ( .A1(write2_in[9]), .B1(n530), .ZN(n3056) );
  INVD1BWP12T U1619 ( .I(n3056), .ZN(n498) );
  CKND2D1BWP12T U1620 ( .A1(n3331), .A2(write2_in[8]), .ZN(n499) );
  CKND3BWP12T U1621 ( .I(n3058), .ZN(n501) );
  INR2D4BWP12T U1622 ( .A1(n502), .B1(n501), .ZN(n1933) );
  TPND2D1BWP12T U1623 ( .A1(write1_in[10]), .A2(n530), .ZN(n504) );
  CKND2D1BWP12T U1624 ( .A1(n3331), .A2(write2_in[10]), .ZN(n503) );
  CKND2D2BWP12T U1625 ( .A1(n504), .A2(n503), .ZN(n3093) );
  INR2D0BWP12T U1626 ( .A1(write2_in[6]), .B1(n530), .ZN(n505) );
  TPAOI21D1BWP12T U1627 ( .A1(write1_in[6]), .A2(n530), .B(n505), .ZN(n3032)
         );
  INR2D0BWP12T U1628 ( .A1(write2_in[5]), .B1(n530), .ZN(n506) );
  AOI21D1BWP12T U1629 ( .A1(write1_in[5]), .A2(n530), .B(n506), .ZN(n3030) );
  TPNR2D1BWP12T U1630 ( .A1(n3032), .A2(n3030), .ZN(n510) );
  ND2XD0BWP12T U1631 ( .A1(n3331), .A2(write2_in[1]), .ZN(n507) );
  TPND2D2BWP12T U1632 ( .A1(n2845), .A2(n2844), .ZN(n2950) );
  INR2D0BWP12T U1633 ( .A1(write2_in[3]), .B1(n530), .ZN(n508) );
  INR2D1BWP12T U1634 ( .A1(write2_in[4]), .B1(n530), .ZN(n509) );
  TPNR3D2BWP12T U1635 ( .A1(n2950), .A2(n2949), .A3(n2938), .ZN(n3031) );
  TPND2D1BWP12T U1636 ( .A1(n510), .A2(n3031), .ZN(n3051) );
  INR2D0BWP12T U1637 ( .A1(write2_in[7]), .B1(n530), .ZN(n511) );
  TPAOI21D1BWP12T U1638 ( .A1(write1_in[7]), .A2(n530), .B(n511), .ZN(n3052)
         );
  TPNR2D3BWP12T U1639 ( .A1(n3051), .A2(n3052), .ZN(n3059) );
  TPND3D2BWP12T U1640 ( .A1(n1933), .A2(n3093), .A3(n3059), .ZN(n515) );
  CKND0BWP12T U1641 ( .I(write2_in[14]), .ZN(n513) );
  CKND0BWP12T U1642 ( .I(write2_in[15]), .ZN(n512) );
  TPNR3D0BWP12T U1643 ( .A1(n530), .A2(n513), .A3(n512), .ZN(n520) );
  NR2D0BWP12T U1644 ( .A1(n520), .A2(n530), .ZN(n514) );
  CKND2D1BWP12T U1645 ( .A1(n3331), .A2(write2_in[13]), .ZN(n516) );
  IOA21D2BWP12T U1646 ( .A1(write1_in[13]), .A2(n530), .B(n516), .ZN(n3107) );
  TPNR2D2BWP12T U1647 ( .A1(n518), .A2(n884), .ZN(n528) );
  ND2D1BWP12T U1648 ( .A1(n3331), .A2(write2_in[18]), .ZN(n880) );
  TPAOI21D2BWP12T U1649 ( .A1(write1_in[14]), .A2(write1_in[15]), .B(n520), 
        .ZN(n525) );
  CKND2D1BWP12T U1650 ( .A1(n3331), .A2(write2_in[12]), .ZN(n521) );
  INVD1P75BWP12T U1651 ( .I(write1_in[11]), .ZN(n524) );
  CKND2D1BWP12T U1652 ( .A1(n3331), .A2(write2_in[11]), .ZN(n523) );
  NR2XD2BWP12T U1653 ( .A1(n525), .A2(n1934), .ZN(n877) );
  TPND2D2BWP12T U1654 ( .A1(n1942), .A2(n877), .ZN(n526) );
  ND2XD3BWP12T U1655 ( .A1(n528), .A2(n527), .ZN(n3504) );
  INVD1BWP12T U1656 ( .I(write2_in[27]), .ZN(n529) );
  CKND2D1BWP12T U1657 ( .A1(n534), .A2(n533), .ZN(n542) );
  NR2D1BWP12T U1658 ( .A1(n3504), .A2(n3497), .ZN(n539) );
  NR2D3BWP12T U1659 ( .A1(next_pc_en_BAR), .A2(n535), .ZN(n3499) );
  TPNR2D0BWP12T U1660 ( .A1(n3343), .A2(n3538), .ZN(n537) );
  AO21D1BWP12T U1661 ( .A1(next_pc_in[27]), .A2(n3499), .B(n537), .Z(n538) );
  TPAOI31D1BWP12T U1662 ( .A1(n540), .A2(n539), .A3(n1038), .B(n538), .ZN(n541) );
  ND2D1BWP12T U1663 ( .A1(n542), .A2(n541), .ZN(n2195) );
  BUFFXD6BWP12T U1664 ( .I(write1_in[30]), .Z(n3226) );
  ND2D1BWP12T U1665 ( .A1(n3226), .A2(n3522), .ZN(n549) );
  AOI22D0BWP12T U1666 ( .A1(write2_in[30]), .A2(n3202), .B1(n3201), .B2(
        r11[30]), .ZN(n548) );
  ND2D1BWP12T U1667 ( .A1(n3226), .A2(n3520), .ZN(n553) );
  ND2D1BWP12T U1668 ( .A1(n593), .A2(n560), .ZN(n550) );
  NR2D1BWP12T U1669 ( .A1(n561), .A2(n591), .ZN(n551) );
  AOI22D0BWP12T U1670 ( .A1(r10[30]), .A2(n3198), .B1(n3197), .B2(
        write2_in[30]), .ZN(n552) );
  ND2D1BWP12T U1671 ( .A1(n3226), .A2(n3515), .ZN(n559) );
  ND2D1BWP12T U1672 ( .A1(n560), .A2(n554), .ZN(n556) );
  INR3D4BWP12T U1673 ( .A1(n556), .B1(reset), .B2(n557), .ZN(n3190) );
  TPNR2D2BWP12T U1674 ( .A1(n557), .A2(n556), .ZN(n3189) );
  AOI22D0BWP12T U1675 ( .A1(r3[30]), .A2(n3190), .B1(n3189), .B2(write2_in[30]), .ZN(n558) );
  ND2D1BWP12T U1676 ( .A1(n3226), .A2(n3516), .ZN(n565) );
  ND2D1BWP12T U1677 ( .A1(n560), .A2(n586), .ZN(n562) );
  NR2D1BWP12T U1678 ( .A1(n561), .A2(n585), .ZN(n563) );
  AOI22D0BWP12T U1679 ( .A1(r2[30]), .A2(n3194), .B1(n3193), .B2(write2_in[30]), .ZN(n564) );
  AOI22D0BWP12T U1680 ( .A1(n3190), .A2(r3[31]), .B1(n3189), .B2(write2_in[31]), .ZN(n566) );
  AOI22D0BWP12T U1681 ( .A1(n3194), .A2(r2[31]), .B1(n3193), .B2(write2_in[31]), .ZN(n568) );
  INVD1BWP12T U1682 ( .I(n570), .ZN(n571) );
  AOI211D4BWP12T U1683 ( .A1(n579), .A2(n586), .B(n571), .C(reset), .ZN(n3219)
         );
  TPNR3D2BWP12T U1684 ( .A1(n571), .A2(n587), .A3(n580), .ZN(n3218) );
  AOI22D0BWP12T U1685 ( .A1(n3219), .A2(r0[31]), .B1(write2_in[31]), .B2(n3218), .ZN(n572) );
  AOI22D0BWP12T U1686 ( .A1(write2_in[31]), .A2(n3202), .B1(n3201), .B2(
        r11[31]), .ZN(n574) );
  AOI22D0BWP12T U1687 ( .A1(write2_in[31]), .A2(n1947), .B1(n1946), .B2(
        tmp1[31]), .ZN(n576) );
  INVD1BWP12T U1688 ( .I(n578), .ZN(n581) );
  AOI211D4BWP12T U1689 ( .A1(n579), .A2(n593), .B(n581), .C(reset), .ZN(n3215)
         );
  TPNR3D2BWP12T U1690 ( .A1(n581), .A2(n596), .A3(n580), .ZN(n3214) );
  AOI22D0BWP12T U1691 ( .A1(n3215), .A2(r8[31]), .B1(write2_in[31]), .B2(n3214), .ZN(n582) );
  INVD0BWP12T U1692 ( .I(n584), .ZN(n592) );
  NR2D1BWP12T U1693 ( .A1(n592), .A2(n585), .ZN(n588) );
  AOI211D4BWP12T U1694 ( .A1(n594), .A2(n586), .B(n588), .C(reset), .ZN(n3223)
         );
  TPNR3D2BWP12T U1695 ( .A1(n588), .A2(n587), .A3(n595), .ZN(n3222) );
  AOI22D0BWP12T U1696 ( .A1(n3223), .A2(r4[31]), .B1(write2_in[31]), .B2(n3222), .ZN(n589) );
  NR2D1BWP12T U1697 ( .A1(n592), .A2(n591), .ZN(n597) );
  AOI211D4BWP12T U1698 ( .A1(n594), .A2(n593), .B(n597), .C(reset), .ZN(n3228)
         );
  TPNR3D2BWP12T U1699 ( .A1(n597), .A2(n596), .A3(n595), .ZN(n3227) );
  AOI22D0BWP12T U1700 ( .A1(n3228), .A2(r12[31]), .B1(write2_in[31]), .B2(
        n3227), .ZN(n598) );
  INVD3BWP12T U1701 ( .I(write1_in[29]), .ZN(n3513) );
  TPAOI21D0BWP12T U1702 ( .A1(n3499), .A2(next_pc_in[1]), .B(reset), .ZN(n601)
         );
  TPND2D0BWP12T U1703 ( .A1(n3498), .A2(pc_out[1]), .ZN(n600) );
  OAI211D0BWP12T U1704 ( .A1(n602), .A2(n2844), .B(n601), .C(n600), .ZN(n2169)
         );
  AO222D0BWP12T U1705 ( .A1(n3184), .A2(write1_in[1]), .B1(n3185), .B2(
        write2_in[1]), .C1(n[3579]), .C2(n3186), .Z(spin[1]) );
  AO222D0BWP12T U1706 ( .A1(n3246), .A2(write1_in[1]), .B1(n1947), .B2(
        write2_in[1]), .C1(n1946), .C2(tmp1[1]), .Z(n2137) );
  AO222D0BWP12T U1707 ( .A1(n3246), .A2(write1_in[3]), .B1(n1947), .B2(
        write2_in[3]), .C1(n1946), .C2(tmp1[3]), .Z(n2139) );
  AO222D0BWP12T U1708 ( .A1(n3184), .A2(write1_in[0]), .B1(n3185), .B2(
        write2_in[0]), .C1(n3186), .C2(n[3580]), .Z(spin[0]) );
  AO222D0BWP12T U1709 ( .A1(n3246), .A2(write1_in[0]), .B1(n1947), .B2(
        write2_in[0]), .C1(n1946), .C2(tmp1[0]), .Z(n2135) );
  ND2D1BWP12T U1710 ( .A1(n3419), .A2(r9[17]), .ZN(n605) );
  OR2XD2BWP12T U1711 ( .A1(n608), .A2(n607), .Z(n613) );
  OAI22D1BWP12T U1712 ( .A1(n3416), .A2(n610), .B1(n609), .B2(n3444), .ZN(n611) );
  TPNR3D2BWP12T U1713 ( .A1(n613), .A2(n612), .A3(n611), .ZN(n636) );
  INVD4BWP12T U1714 ( .I(n3446), .ZN(n1862) );
  ND2D1BWP12T U1715 ( .A1(n1049), .A2(pc_out[17]), .ZN(n616) );
  INVD1BWP12T U1716 ( .I(n614), .ZN(n615) );
  ND2D1BWP12T U1717 ( .A1(n3417), .A2(r1[17]), .ZN(n619) );
  TPND2D1BWP12T U1718 ( .A1(n620), .A2(n619), .ZN(n627) );
  TPND2D2BWP12T U1719 ( .A1(n621), .A2(r12[17]), .ZN(n625) );
  INVD3BWP12T U1720 ( .I(n3429), .ZN(n623) );
  TPNR2D3BWP12T U1721 ( .A1(n623), .A2(n622), .ZN(n1380) );
  ND2D1BWP12T U1722 ( .A1(n1380), .A2(tmp1[17]), .ZN(n624) );
  CKND2D2BWP12T U1723 ( .A1(n625), .A2(n624), .ZN(n626) );
  NR2D2BWP12T U1724 ( .A1(n627), .A2(n626), .ZN(n634) );
  INR2D1BWP12T U1725 ( .A1(r3[17]), .B1(n3434), .ZN(n628) );
  INVD1BWP12T U1726 ( .I(n628), .ZN(n632) );
  BUFFD4BWP12T U1727 ( .I(n3450), .Z(n1853) );
  ND2D1BWP12T U1728 ( .A1(n1853), .A2(r4[17]), .ZN(n631) );
  AOI22D1BWP12T U1729 ( .A1(n629), .A2(r0[17]), .B1(n1622), .B2(r2[17]), .ZN(
        n630) );
  INVD1BWP12T U1730 ( .I(r3[14]), .ZN(n1539) );
  OR2XD1BWP12T U1731 ( .A1(n1428), .A2(n1539), .Z(n642) );
  INVD0BWP12T U1732 ( .I(tmp1[14]), .ZN(n638) );
  ND2D1BWP12T U1733 ( .A1(n1804), .A2(immediate1_in[14]), .ZN(n637) );
  OAI21D1BWP12T U1734 ( .A1(n3378), .A2(n638), .B(n637), .ZN(n640) );
  AN2D1BWP12T U1735 ( .A1(n1473), .A2(r8[14]), .Z(n639) );
  INVD1BWP12T U1736 ( .I(lr[14]), .ZN(n1992) );
  INVD8BWP12T U1737 ( .I(n3393), .ZN(n3418) );
  OAI21D1BWP12T U1738 ( .A1(n3416), .A2(n1992), .B(n643), .ZN(n647) );
  BUFFXD3BWP12T U1739 ( .I(n3419), .Z(n1645) );
  ND2D1BWP12T U1740 ( .A1(n1645), .A2(r9[14]), .ZN(n645) );
  ND2D1BWP12T U1741 ( .A1(n3412), .A2(r6[14]), .ZN(n644) );
  TPNR3D2BWP12T U1742 ( .A1(n648), .A2(n647), .A3(n646), .ZN(n663) );
  INVD1BWP12T U1743 ( .I(r5[14]), .ZN(n1547) );
  INR2D1BWP12T U1744 ( .A1(r7[14]), .B1(n3444), .ZN(n649) );
  NR3D1BWP12T U1745 ( .A1(n651), .A2(n650), .A3(n649), .ZN(n662) );
  BUFFXD6BWP12T U1746 ( .I(n3445), .Z(n1788) );
  ND2D1BWP12T U1747 ( .A1(n1788), .A2(pc_out[14]), .ZN(n660) );
  INR2D1BWP12T U1748 ( .A1(r0[14]), .B1(n3442), .ZN(n659) );
  INR2D1BWP12T U1749 ( .A1(r2[14]), .B1(n1787), .ZN(n652) );
  INVD1BWP12T U1750 ( .I(n652), .ZN(n657) );
  ND2D1BWP12T U1751 ( .A1(n3450), .A2(r4[14]), .ZN(n653) );
  IOA21D2BWP12T U1752 ( .A1(n1069), .A2(r10[14]), .B(n653), .ZN(n655) );
  INR2D1BWP12T U1753 ( .A1(n[3566]), .B1(n3446), .ZN(n654) );
  INR3D2BWP12T U1754 ( .A1(n660), .B1(n659), .B2(n658), .ZN(n661) );
  ND3XD4BWP12T U1755 ( .A1(n663), .A2(n662), .A3(n661), .ZN(regA_out[14]) );
  INVD1BWP12T U1756 ( .I(r0[19]), .ZN(n1344) );
  TPAOI21D1BWP12T U1757 ( .A1(r6[19]), .A2(n3412), .B(n664), .ZN(n668) );
  INVD1BWP12T U1758 ( .I(n665), .ZN(n667) );
  ND3D2BWP12T U1759 ( .A1(n668), .A2(n667), .A3(n666), .ZN(n674) );
  INVD1BWP12T U1760 ( .I(r12[19]), .ZN(n670) );
  BUFFXD8BWP12T U1761 ( .I(n1219), .Z(n1859) );
  OAI21D1BWP12T U1762 ( .A1(n3436), .A2(n670), .B(n669), .ZN(n673) );
  INVD4BWP12T U1763 ( .I(n1069), .ZN(n1881) );
  INVD1BWP12T U1764 ( .I(r10[19]), .ZN(n2070) );
  TPND2D2BWP12T U1765 ( .A1(n3418), .A2(r11[19]), .ZN(n671) );
  OAI21D1BWP12T U1766 ( .A1(n1881), .A2(n2070), .B(n671), .ZN(n672) );
  TPNR3D2BWP12T U1767 ( .A1(n674), .A2(n673), .A3(n672), .ZN(n686) );
  INVD1BWP12T U1768 ( .I(r3[19]), .ZN(n1341) );
  NR2D0BWP12T U1769 ( .A1(n1428), .A2(n1341), .ZN(n677) );
  INVD1BWP12T U1770 ( .I(n[3561]), .ZN(n2069) );
  ND2D1BWP12T U1771 ( .A1(n3419), .A2(r9[19]), .ZN(n675) );
  OAI21D1BWP12T U1772 ( .A1(n3404), .A2(n2069), .B(n675), .ZN(n676) );
  INR3D2BWP12T U1773 ( .A1(n678), .B1(n677), .B2(n676), .ZN(n685) );
  INVD1BWP12T U1774 ( .I(r2[19]), .ZN(n1333) );
  OAI21D1BWP12T U1775 ( .A1(n3432), .A2(n1333), .B(n679), .ZN(n683) );
  INVD1BWP12T U1776 ( .I(r7[19]), .ZN(n1343) );
  NR2D1BWP12T U1777 ( .A1(n3444), .A2(n1343), .ZN(n682) );
  INVD1BWP12T U1778 ( .I(r5[19]), .ZN(n1345) );
  ND2D2BWP12T U1779 ( .A1(n3417), .A2(r1[19]), .ZN(n680) );
  TPOAI21D1BWP12T U1780 ( .A1(n3414), .A2(n1345), .B(n680), .ZN(n681) );
  NR3D1BWP12T U1781 ( .A1(n683), .A2(n682), .A3(n681), .ZN(n684) );
  ND3D2BWP12T U1782 ( .A1(n686), .A2(n685), .A3(n684), .ZN(regA_out[19]) );
  INVD1BWP12T U1783 ( .I(r2[5]), .ZN(n2021) );
  ND2D1BWP12T U1784 ( .A1(n1473), .A2(r8[5]), .ZN(n687) );
  TPOAI21D1BWP12T U1785 ( .A1(n2021), .A2(n3432), .B(n687), .ZN(n694) );
  ND2D1BWP12T U1786 ( .A1(n1804), .A2(immediate1_in[5]), .ZN(n688) );
  IOA21D1BWP12T U1787 ( .A1(r4[5]), .A2(n3450), .B(n688), .ZN(n689) );
  INVD1BWP12T U1788 ( .I(n689), .ZN(n693) );
  INVD1BWP12T U1789 ( .I(r10[5]), .ZN(n2868) );
  NR2D1BWP12T U1790 ( .A1(n1881), .A2(n2868), .ZN(n691) );
  TPNR2D1BWP12T U1791 ( .A1(n691), .A2(n690), .ZN(n692) );
  IND3D2BWP12T U1792 ( .A1(n694), .B1(n693), .B2(n692), .ZN(n700) );
  INR2D2BWP12T U1793 ( .A1(lr[5]), .B1(n3416), .ZN(n695) );
  INVD1P75BWP12T U1794 ( .I(n695), .ZN(n697) );
  CKND2D2BWP12T U1795 ( .A1(n3418), .A2(r11[5]), .ZN(n696) );
  ND3D2BWP12T U1796 ( .A1(n697), .A2(n696), .A3(n188), .ZN(n699) );
  TPNR3D2BWP12T U1797 ( .A1(n700), .A2(n699), .A3(n698), .ZN(n714) );
  AN2D1BWP12T U1798 ( .A1(n3412), .A2(r6[5]), .Z(n712) );
  ND2D1BWP12T U1799 ( .A1(n3419), .A2(r9[5]), .ZN(n702) );
  INVD1BWP12T U1800 ( .I(r3[5]), .ZN(n2020) );
  ND2D1BWP12T U1801 ( .A1(n1646), .A2(r3[5]), .ZN(n701) );
  ND2D1BWP12T U1802 ( .A1(n702), .A2(n701), .ZN(n711) );
  INR2D2BWP12T U1803 ( .A1(r1[5]), .B1(n1810), .ZN(n703) );
  INVD1P75BWP12T U1804 ( .I(n703), .ZN(n706) );
  INR2D2BWP12T U1805 ( .A1(r0[5]), .B1(n3442), .ZN(n704) );
  INVD1P75BWP12T U1806 ( .I(n704), .ZN(n705) );
  ND2D2BWP12T U1807 ( .A1(n706), .A2(n705), .ZN(n710) );
  ND2D1BWP12T U1808 ( .A1(n1876), .A2(tmp1[5]), .ZN(n708) );
  TPND2D1BWP12T U1809 ( .A1(n708), .A2(n707), .ZN(n709) );
  NR4D2BWP12T U1810 ( .A1(n712), .A2(n711), .A3(n710), .A4(n709), .ZN(n713) );
  TPND2D2BWP12T U1811 ( .A1(n714), .A2(n713), .ZN(regA_out[5]) );
  MOAI22D0BWP12T U1812 ( .A1(n715), .A2(n1714), .B1(n1713), .B2(
        immediate2_in[0]), .ZN(n720) );
  TPOAI22D1BWP12T U1813 ( .A1(n1911), .A2(n716), .B1(n1519), .B2(n2824), .ZN(
        n717) );
  AOI22D1BWP12T U1814 ( .A1(n1664), .A2(r12[0]), .B1(n1918), .B2(r4[0]), .ZN(
        n718) );
  ND2D1BWP12T U1815 ( .A1(n1915), .A2(r6[0]), .ZN(n724) );
  INR2D2BWP12T U1816 ( .A1(pc_out[0]), .B1(n1703), .ZN(n722) );
  INVD1BWP12T U1817 ( .I(n722), .ZN(n723) );
  CKND2D1BWP12T U1818 ( .A1(n724), .A2(n723), .ZN(n726) );
  AOI22D1BWP12T U1819 ( .A1(n1921), .A2(tmp1[0]), .B1(n1571), .B2(r8[0]), .ZN(
        n725) );
  IND2XD2BWP12T U1820 ( .A1(n726), .B1(n725), .ZN(n727) );
  TPNR2D2BWP12T U1821 ( .A1(n728), .A2(n727), .ZN(n736) );
  TPOAI22D1BWP12T U1822 ( .A1(n1663), .A2(n2711), .B1(n3065), .B2(n1592), .ZN(
        n733) );
  TPOAI22D1BWP12T U1823 ( .A1(n1587), .A2(n2821), .B1(n729), .B2(n1895), .ZN(
        n732) );
  TPOAI22D2BWP12T U1824 ( .A1(n1887), .A2(n3067), .B1(n1889), .B2(n730), .ZN(
        n731) );
  TPND2D3BWP12T U1825 ( .A1(n736), .A2(n735), .ZN(regB_out[0]) );
  INVD1BWP12T U1826 ( .I(r3[4]), .ZN(n2013) );
  OAI22D1BWP12T U1827 ( .A1(n3404), .A2(n1178), .B1(n2013), .B2(n3434), .ZN(
        n745) );
  AOI22D1BWP12T U1828 ( .A1(n1876), .A2(tmp1[4]), .B1(n1804), .B2(
        immediate1_in[4]), .ZN(n739) );
  INVD1BWP12T U1829 ( .I(r2[4]), .ZN(n2012) );
  ND3D1BWP12T U1830 ( .A1(n740), .A2(n739), .A3(n738), .ZN(n744) );
  OAI22D1BWP12T U1831 ( .A1(n3414), .A2(n741), .B1(n1810), .B2(n1174), .ZN(
        n743) );
  INVD1BWP12T U1832 ( .I(pc_out[4]), .ZN(n1169) );
  OAI22D1BWP12T U1833 ( .A1(n3406), .A2(n1169), .B1(n1177), .B2(n3444), .ZN(
        n742) );
  NR4D0BWP12T U1834 ( .A1(n745), .A2(n744), .A3(n743), .A4(n742), .ZN(n751) );
  OAI22D1BWP12T U1835 ( .A1(n3416), .A2(n2843), .B1(n3393), .B2(n2011), .ZN(
        n749) );
  INVD1BWP12T U1836 ( .I(r4[4]), .ZN(n2010) );
  INVD1BWP12T U1837 ( .I(r0[4]), .ZN(n2007) );
  OAI22D1BWP12T U1838 ( .A1(n3390), .A2(n2010), .B1(n2007), .B2(n3442), .ZN(
        n748) );
  INVD1BWP12T U1839 ( .I(r8[4]), .ZN(n2008) );
  INVD1BWP12T U1840 ( .I(r12[4]), .ZN(n2009) );
  OAI22D1BWP12T U1841 ( .A1(n2008), .A2(n3387), .B1(n3436), .B2(n2009), .ZN(
        n747) );
  INVD1BWP12T U1842 ( .I(r10[4]), .ZN(n2841) );
  OAI22D1BWP12T U1843 ( .A1(n3402), .A2(n2842), .B1(n2841), .B2(n1881), .ZN(
        n746) );
  NR4D0BWP12T U1844 ( .A1(n749), .A2(n748), .A3(n747), .A4(n746), .ZN(n750) );
  NR2D1BWP12T U1845 ( .A1(n1922), .A2(n3542), .ZN(n752) );
  AOI21D1BWP12T U1846 ( .A1(n1921), .A2(tmp1[29]), .B(n752), .ZN(n756) );
  ND2D1BWP12T U1847 ( .A1(n756), .A2(n755), .ZN(n765) );
  INVD1BWP12T U1848 ( .I(lr[29]), .ZN(n2656) );
  RCAOI21D1BWP12T U1849 ( .A1(immediate2_in[29]), .A2(n1668), .B(n757), .ZN(
        n761) );
  AN2D1BWP12T U1850 ( .A1(n168), .A2(r1[29]), .Z(n758) );
  TPNR2D1BWP12T U1851 ( .A1(n759), .A2(n758), .ZN(n760) );
  CKND2D2BWP12T U1852 ( .A1(n761), .A2(n760), .ZN(n764) );
  ND2D1BWP12T U1853 ( .A1(n1915), .A2(r6[29]), .ZN(n762) );
  OAI21D1BWP12T U1854 ( .A1(n1917), .A2(n3533), .B(n762), .ZN(n763) );
  TPNR3D2BWP12T U1855 ( .A1(n765), .A2(n764), .A3(n763), .ZN(n776) );
  INVD2BWP12T U1856 ( .I(n1675), .ZN(n1726) );
  INVD1BWP12T U1857 ( .I(r5[29]), .ZN(n1637) );
  NR2D2BWP12T U1858 ( .A1(n161), .A2(n1637), .ZN(n766) );
  RCAOI21D1BWP12T U1859 ( .A1(n1726), .A2(r11[29]), .B(n766), .ZN(n769) );
  INVD1BWP12T U1860 ( .I(r7[29]), .ZN(n1636) );
  NR2D1BWP12T U1861 ( .A1(n1724), .A2(n1636), .ZN(n767) );
  AOI21D1BWP12T U1862 ( .A1(n1892), .A2(r0[29]), .B(n767), .ZN(n768) );
  TPND2D1BWP12T U1863 ( .A1(n769), .A2(n768), .ZN(n774) );
  ND2D1BWP12T U1864 ( .A1(n1898), .A2(n[3551]), .ZN(n770) );
  OAI21D1BWP12T U1865 ( .A1(n1896), .A2(n3534), .B(n770), .ZN(n773) );
  BUFFXD3BWP12T U1866 ( .I(n1691), .Z(n1900) );
  CKND2D0BWP12T U1867 ( .A1(n1900), .A2(r9[29]), .ZN(n771) );
  OAI21D1BWP12T U1868 ( .A1(n1592), .A2(n3544), .B(n771), .ZN(n772) );
  TPNR3D2BWP12T U1869 ( .A1(n774), .A2(n773), .A3(n772), .ZN(n775) );
  TPND2D2BWP12T U1870 ( .A1(n776), .A2(n775), .ZN(regB_out[29]) );
  INVD1BWP12T U1871 ( .I(lr[24]), .ZN(n2697) );
  INVD1BWP12T U1872 ( .I(r12[24]), .ZN(n2696) );
  INVD1BWP12T U1873 ( .I(r4[24]), .ZN(n778) );
  INVD1BWP12T U1874 ( .I(r8[24]), .ZN(n777) );
  OAI22D0BWP12T U1875 ( .A1(n3390), .A2(n778), .B1(n777), .B2(n1372), .ZN(n782) );
  INVD1BWP12T U1876 ( .I(r10[24]), .ZN(n1591) );
  INVD1BWP12T U1877 ( .I(r11[24]), .ZN(n1588) );
  INVD1BWP12T U1878 ( .I(r6[24]), .ZN(n779) );
  INVD1BWP12T U1879 ( .I(r0[24]), .ZN(n1586) );
  TPOAI22D1BWP12T U1880 ( .A1(n3396), .A2(n779), .B1(n3442), .B2(n1586), .ZN(
        n780) );
  NR4D0BWP12T U1881 ( .A1(n783), .A2(n782), .A3(n781), .A4(n780), .ZN(n795) );
  INVD1BWP12T U1882 ( .I(r2[24]), .ZN(n1577) );
  INVD1BWP12T U1883 ( .I(tmp1[24]), .ZN(n784) );
  INVD1BWP12T U1884 ( .I(r7[24]), .ZN(n1585) );
  ND2D1BWP12T U1885 ( .A1(n787), .A2(n786), .ZN(n788) );
  AOI211D1BWP12T U1886 ( .A1(r1[24]), .A2(n3384), .B(n789), .C(n788), .ZN(n794) );
  INVD1BWP12T U1887 ( .I(n[3556]), .ZN(n790) );
  INVD1BWP12T U1888 ( .I(r9[24]), .ZN(n1589) );
  OAI22D1BWP12T U1889 ( .A1(n3404), .A2(n790), .B1(n3402), .B2(n1589), .ZN(
        n792) );
  INVD1BWP12T U1890 ( .I(pc_out[24]), .ZN(n3295) );
  INVD1BWP12T U1891 ( .I(r3[24]), .ZN(n1584) );
  OAI22D1BWP12T U1892 ( .A1(n3406), .A2(n3295), .B1(n1584), .B2(n3434), .ZN(
        n791) );
  NR2D1BWP12T U1893 ( .A1(n792), .A2(n791), .ZN(n793) );
  AOI22D0BWP12T U1894 ( .A1(n3215), .A2(r8[29]), .B1(write2_in[29]), .B2(n3214), .ZN(n3527) );
  AOI22D0BWP12T U1895 ( .A1(n3219), .A2(r0[29]), .B1(write2_in[29]), .B2(n3218), .ZN(n3525) );
  AOI22D0BWP12T U1896 ( .A1(write2_in[29]), .A2(n3202), .B1(n3201), .B2(
        r11[29]), .ZN(n3530) );
  AOI22D0BWP12T U1897 ( .A1(n3228), .A2(r12[29]), .B1(write2_in[29]), .B2(
        n3227), .ZN(n3529) );
  AOI22D0BWP12T U1898 ( .A1(n3223), .A2(r4[29]), .B1(write2_in[29]), .B2(n3222), .ZN(n3526) );
  AOI22D0BWP12T U1899 ( .A1(n3198), .A2(r10[29]), .B1(n3197), .B2(
        write2_in[29]), .ZN(n3528) );
  AOI22D0BWP12T U1900 ( .A1(n3194), .A2(r2[29]), .B1(n3193), .B2(write2_in[29]), .ZN(n3524) );
  AOI22D0BWP12T U1901 ( .A1(n3190), .A2(r3[29]), .B1(n3189), .B2(write2_in[29]), .ZN(n3523) );
  AOI22D0BWP12T U1902 ( .A1(n3198), .A2(r10[31]), .B1(n3197), .B2(
        write2_in[31]), .ZN(n3531) );
  AOI22D1BWP12T U1903 ( .A1(n1575), .A2(pc_out[30]), .B1(r6[30]), .B2(n1915), 
        .ZN(n804) );
  INVD1BWP12T U1904 ( .I(r2[30]), .ZN(n3376) );
  INVD1BWP12T U1905 ( .I(r1[30]), .ZN(n796) );
  IND2XD1BWP12T U1906 ( .A1(n798), .B1(n797), .ZN(n803) );
  AOI22D1BWP12T U1907 ( .A1(n1571), .A2(r8[30]), .B1(tmp1[30]), .B2(n1526), 
        .ZN(n801) );
  AOI22D1BWP12T U1908 ( .A1(n1664), .A2(r12[30]), .B1(n1918), .B2(r4[30]), 
        .ZN(n800) );
  INVD1BWP12T U1909 ( .I(lr[30]), .ZN(n3386) );
  OR2XD1BWP12T U1910 ( .A1(n1714), .A2(n3386), .Z(n799) );
  ND3D1BWP12T U1911 ( .A1(n801), .A2(n800), .A3(n799), .ZN(n802) );
  INR3XD1BWP12T U1912 ( .A1(n804), .B1(n803), .B2(n802), .ZN(n812) );
  INVD1BWP12T U1913 ( .I(r9[30]), .ZN(n3401) );
  INVD1BWP12T U1914 ( .I(r10[30]), .ZN(n3391) );
  OAI22D1BWP12T U1915 ( .A1(n1553), .A2(n3401), .B1(n3391), .B2(n1592), .ZN(
        n806) );
  INVD1BWP12T U1916 ( .I(r0[30]), .ZN(n3394) );
  INVD1BWP12T U1917 ( .I(r7[30]), .ZN(n3379) );
  OAI22D1BWP12T U1918 ( .A1(n1587), .A2(n3394), .B1(n3379), .B2(n1895), .ZN(
        n805) );
  OR2XD2BWP12T U1919 ( .A1(n806), .A2(n805), .Z(n810) );
  INVD1BWP12T U1920 ( .I(n[3550]), .ZN(n3403) );
  INVD1BWP12T U1921 ( .I(r3[30]), .ZN(n3405) );
  OAI22D1BWP12T U1922 ( .A1(n1652), .A2(n3403), .B1(n3405), .B2(n1896), .ZN(
        n808) );
  INVD1BWP12T U1923 ( .I(r11[30]), .ZN(n3392) );
  INVD1BWP12T U1924 ( .I(r5[30]), .ZN(n3380) );
  OR2XD2BWP12T U1925 ( .A1(n808), .A2(n807), .Z(n809) );
  TPNR2D2BWP12T U1926 ( .A1(n810), .A2(n809), .ZN(n811) );
  TPND2D2BWP12T U1927 ( .A1(n812), .A2(n811), .ZN(regB_out[30]) );
  AOI22D1BWP12T U1928 ( .A1(n1575), .A2(pc_out[23]), .B1(r6[23]), .B2(n1915), 
        .ZN(n814) );
  INVD1BWP12T U1929 ( .I(lr[23]), .ZN(n1974) );
  INVD0BWP12T U1930 ( .I(r1[23]), .ZN(n815) );
  INVD1BWP12T U1931 ( .I(r2[23]), .ZN(n1757) );
  AOI22D1BWP12T U1932 ( .A1(n1664), .A2(r12[23]), .B1(n1918), .B2(r4[23]), 
        .ZN(n816) );
  INVD1BWP12T U1933 ( .I(r3[23]), .ZN(n1764) );
  IOA22D2BWP12T U1934 ( .B1(n1764), .B2(n1896), .A1(n1898), .A2(n[3557]), .ZN(
        n824) );
  INVD1BWP12T U1935 ( .I(r0[23]), .ZN(n1751) );
  INVD0BWP12T U1936 ( .I(r7[23]), .ZN(n820) );
  OAI22D1BWP12T U1937 ( .A1(n1587), .A2(n1751), .B1(n820), .B2(n1895), .ZN(
        n823) );
  INVD1BWP12T U1938 ( .I(r11[23]), .ZN(n1750) );
  INVD1BWP12T U1939 ( .I(r5[23]), .ZN(n1759) );
  OAI22D1BWP12T U1940 ( .A1(n1887), .A2(n1750), .B1(n161), .B2(n1759), .ZN(
        n822) );
  INVD1BWP12T U1941 ( .I(r9[23]), .ZN(n1762) );
  INVD1BWP12T U1942 ( .I(r10[23]), .ZN(n1975) );
  NR4D2BWP12T U1943 ( .A1(n824), .A2(n823), .A3(n822), .A4(n821), .ZN(n825) );
  ND2XD4BWP12T U1944 ( .A1(n826), .A2(n825), .ZN(regB_out[23]) );
  INR2D1BWP12T U1945 ( .A1(r7[8]), .B1(n1724), .ZN(n827) );
  INVD1BWP12T U1946 ( .I(r11[8]), .ZN(n2907) );
  ND2D1BWP12T U1947 ( .A1(n1674), .A2(r5[8]), .ZN(n828) );
  OAI21D1BWP12T U1948 ( .A1(n175), .A2(n2907), .B(n828), .ZN(n836) );
  INR2D1BWP12T U1949 ( .A1(r10[8]), .B1(n1899), .ZN(n831) );
  AOI21D1BWP12T U1950 ( .A1(n1898), .A2(n[3572]), .B(n832), .ZN(n833) );
  ND2D1BWP12T U1951 ( .A1(n834), .A2(n833), .ZN(n835) );
  INR3XD2BWP12T U1952 ( .A1(n837), .B1(n836), .B2(n835), .ZN(n852) );
  INVD1BWP12T U1953 ( .I(pc_out[8]), .ZN(n2997) );
  ND2D1BWP12T U1954 ( .A1(n1915), .A2(r6[8]), .ZN(n838) );
  OAI21D1BWP12T U1955 ( .A1(n1917), .A2(n2997), .B(n838), .ZN(n844) );
  INVD1BWP12T U1956 ( .I(r12[8]), .ZN(n2906) );
  ND2D1BWP12T U1957 ( .A1(n1918), .A2(r4[8]), .ZN(n839) );
  OAI21D1BWP12T U1958 ( .A1(n1920), .A2(n2906), .B(n839), .ZN(n843) );
  CKND0BWP12T U1959 ( .I(n1571), .ZN(n841) );
  INVD1BWP12T U1960 ( .I(r8[8]), .ZN(n2905) );
  TPNR3D2BWP12T U1961 ( .A1(n844), .A2(n843), .A3(n842), .ZN(n851) );
  INVD1BWP12T U1962 ( .I(n1669), .ZN(n846) );
  INVD1BWP12T U1963 ( .I(lr[8]), .ZN(n2996) );
  INVD1BWP12T U1964 ( .I(r2[8]), .ZN(n2908) );
  NR2D1BWP12T U1965 ( .A1(n1519), .A2(n2908), .ZN(n848) );
  INVD1BWP12T U1966 ( .I(r1[8]), .ZN(n2932) );
  NR2D1BWP12T U1967 ( .A1(n1659), .A2(n2932), .ZN(n847) );
  AOI21D1BWP12T U1968 ( .A1(n1853), .A2(r4[7]), .B(n853), .ZN(n860) );
  INVD1BWP12T U1969 ( .I(r0[7]), .ZN(n2864) );
  NR2D1BWP12T U1970 ( .A1(n3432), .A2(n2849), .ZN(n854) );
  ND2D1BWP12T U1971 ( .A1(n3384), .A2(r1[7]), .ZN(n856) );
  ND2D1BWP12T U1972 ( .A1(n1380), .A2(tmp1[7]), .ZN(n855) );
  ND3D1BWP12T U1973 ( .A1(n857), .A2(n856), .A3(n855), .ZN(n858) );
  INR3D2BWP12T U1974 ( .A1(n860), .B1(n859), .B2(n858), .ZN(n875) );
  ND2D1BWP12T U1975 ( .A1(n3419), .A2(r9[7]), .ZN(n862) );
  ND2D1BWP12T U1976 ( .A1(n863), .A2(n862), .ZN(n866) );
  ND2D1BWP12T U1977 ( .A1(n1804), .A2(immediate1_in[7]), .ZN(n864) );
  OAI21D1BWP12T U1978 ( .A1(n3436), .A2(n2846), .B(n864), .ZN(n865) );
  NR3XD0BWP12T U1979 ( .A1(n867), .A2(n866), .A3(n865), .ZN(n873) );
  INVD6BWP12T U1980 ( .I(n3393), .ZN(n1200) );
  INVD1BWP12T U1981 ( .I(r10[7]), .ZN(n2859) );
  NR2D1BWP12T U1982 ( .A1(n1881), .A2(n2859), .ZN(n870) );
  INVD1BWP12T U1983 ( .I(r3[7]), .ZN(n2848) );
  ND2D1BWP12T U1984 ( .A1(n3445), .A2(pc_out[7]), .ZN(n868) );
  OAI21D1BWP12T U1985 ( .A1(n3434), .A2(n2848), .B(n868), .ZN(n869) );
  AN2XD2BWP12T U1986 ( .A1(n873), .A2(n872), .Z(n874) );
  TPND2D3BWP12T U1987 ( .A1(n875), .A2(n874), .ZN(regA_out[7]) );
  CKND4BWP12T U1988 ( .I(n3250), .ZN(n883) );
  CKND2D0BWP12T U1989 ( .A1(n887), .A2(n3331), .ZN(n879) );
  IOA21D0BWP12T U1990 ( .A1(n880), .A2(n3331), .B(n879), .ZN(n881) );
  TPND2D2BWP12T U1991 ( .A1(n883), .A2(n882), .ZN(n885) );
  NR3XD4BWP12T U1992 ( .A1(n886), .A2(n885), .A3(n884), .ZN(n892) );
  INR2D4BWP12T U1993 ( .A1(n887), .B1(write1_in[25]), .ZN(n3320) );
  TPND2D2BWP12T U1994 ( .A1(n892), .A2(n899), .ZN(n889) );
  INVD1BWP12T U1995 ( .I(n887), .ZN(n888) );
  TPNR3D2BWP12T U1996 ( .A1(n889), .A2(n1028), .A3(n893), .ZN(n890) );
  ND2XD3BWP12T U1997 ( .A1(n890), .A2(n3327), .ZN(n1608) );
  INR2D1BWP12T U1998 ( .A1(write2_in[28]), .B1(n530), .ZN(n1037) );
  INR2D1BWP12T U1999 ( .A1(write2_in[30]), .B1(n530), .ZN(n907) );
  TPAOI21D8BWP12T U2000 ( .A1(write1_in[30]), .A2(n530), .B(n907), .ZN(n3345)
         );
  INR2XD2BWP12T U2001 ( .A1(n3505), .B1(n3345), .ZN(n891) );
  INVD1BWP12T U2002 ( .I(n3327), .ZN(n896) );
  CKND0BWP12T U2003 ( .I(n1037), .ZN(n897) );
  INVD2P3BWP12T U2004 ( .I(n892), .ZN(n894) );
  NR2D2BWP12T U2005 ( .A1(n894), .A2(n893), .ZN(n3323) );
  IOA21D2BWP12T U2006 ( .A1(n3153), .A2(n897), .B(n3323), .ZN(n895) );
  NR2XD1BWP12T U2007 ( .A1(n896), .A2(n895), .ZN(n905) );
  INR2D1BWP12T U2008 ( .A1(write2_in[29]), .B1(n897), .ZN(n901) );
  OAI21D0BWP12T U2009 ( .A1(n530), .A2(n901), .B(n3505), .ZN(n898) );
  TPNR2D1BWP12T U2010 ( .A1(n174), .A2(n898), .ZN(n900) );
  TPNR2D1BWP12T U2011 ( .A1(n903), .A2(n902), .ZN(n904) );
  ND3XD3BWP12T U2012 ( .A1(n905), .A2(n904), .A3(n3345), .ZN(n912) );
  INR2XD0BWP12T U2013 ( .A1(write2_in[29]), .B1(n530), .ZN(n3324) );
  TPAOI21D2BWP12T U2014 ( .A1(write1_in[29]), .A2(n530), .B(n3324), .ZN(n1606)
         );
  INVD0BWP12T U2015 ( .I(n907), .ZN(n906) );
  INR2D2BWP12T U2016 ( .A1(n906), .B1(write1_in[30]), .ZN(n3337) );
  INVD1BWP12T U2017 ( .I(n3337), .ZN(n910) );
  NR2D0BWP12T U2018 ( .A1(n907), .A2(n530), .ZN(n3333) );
  NR2D0BWP12T U2019 ( .A1(n3497), .A2(n3333), .ZN(n909) );
  TPAOI31D1BWP12T U2020 ( .A1(n1606), .A2(n910), .A3(n909), .B(n908), .ZN(n911) );
  ND3D2BWP12T U2021 ( .A1(n913), .A2(n912), .A3(n911), .ZN(n2198) );
  AOI22D1BWP12T U2022 ( .A1(n1571), .A2(r8[20]), .B1(tmp1[20]), .B2(n1921), 
        .ZN(n923) );
  INVD0BWP12T U2023 ( .I(r1[20]), .ZN(n915) );
  CKND0BWP12T U2024 ( .I(r2[20]), .ZN(n914) );
  AOI22D1BWP12T U2025 ( .A1(n1575), .A2(pc_out[20]), .B1(r6[20]), .B2(n1915), 
        .ZN(n916) );
  AOI22D1BWP12T U2026 ( .A1(n1664), .A2(r12[20]), .B1(n1918), .B2(r4[20]), 
        .ZN(n920) );
  ND3D1BWP12T U2027 ( .A1(n920), .A2(n919), .A3(n918), .ZN(n921) );
  INR3XD1BWP12T U2028 ( .A1(n923), .B1(n922), .B2(n921), .ZN(n933) );
  CKND0BWP12T U2029 ( .I(r3[20]), .ZN(n924) );
  MOAI22D0BWP12T U2030 ( .A1(n924), .A2(n1896), .B1(n1690), .B2(n[3560]), .ZN(
        n931) );
  INVD1BWP12T U2031 ( .I(r0[20]), .ZN(n1869) );
  INVD1BWP12T U2032 ( .I(r7[20]), .ZN(n925) );
  OAI22D1BWP12T U2033 ( .A1(n1587), .A2(n1869), .B1(n925), .B2(n1895), .ZN(
        n930) );
  CKND1BWP12T U2034 ( .I(r11[20]), .ZN(n2710) );
  INVD0BWP12T U2035 ( .I(r5[20]), .ZN(n926) );
  OAI22D1BWP12T U2036 ( .A1(n175), .A2(n2710), .B1(n160), .B2(n926), .ZN(n929)
         );
  INVD1BWP12T U2037 ( .I(r9[20]), .ZN(n927) );
  INVD1BWP12T U2038 ( .I(r10[20]), .ZN(n1880) );
  TPOAI22D1BWP12T U2039 ( .A1(n1553), .A2(n927), .B1(n1880), .B2(n1592), .ZN(
        n928) );
  NR4D1BWP12T U2040 ( .A1(n931), .A2(n930), .A3(n929), .A4(n928), .ZN(n932) );
  ND2D2BWP12T U2041 ( .A1(n933), .A2(n932), .ZN(regB_out[20]) );
  INVD1BWP12T U2042 ( .I(r12[28]), .ZN(n934) );
  INVD1BWP12T U2043 ( .I(lr[28]), .ZN(n1320) );
  INVD1BWP12T U2044 ( .I(r4[28]), .ZN(n936) );
  INVD1BWP12T U2045 ( .I(r8[28]), .ZN(n935) );
  OAI22D0BWP12T U2046 ( .A1(n3390), .A2(n936), .B1(n935), .B2(n1372), .ZN(n940) );
  INVD1BWP12T U2047 ( .I(r11[28]), .ZN(n2679) );
  INVD1BWP12T U2048 ( .I(r10[28]), .ZN(n1311) );
  OAI22D1BWP12T U2049 ( .A1(n3393), .A2(n2679), .B1(n1311), .B2(n3452), .ZN(
        n939) );
  INVD1BWP12T U2050 ( .I(r6[28]), .ZN(n937) );
  INVD1BWP12T U2051 ( .I(r0[28]), .ZN(n1314) );
  OAI22D1BWP12T U2052 ( .A1(n3396), .A2(n937), .B1(n3442), .B2(n1314), .ZN(
        n938) );
  NR4D0BWP12T U2053 ( .A1(n941), .A2(n940), .A3(n939), .A4(n938), .ZN(n950) );
  INVD1BWP12T U2054 ( .I(n[3552]), .ZN(n2680) );
  INVD1BWP12T U2055 ( .I(r9[28]), .ZN(n1312) );
  OAI22D1BWP12T U2056 ( .A1(n3404), .A2(n2680), .B1(n3402), .B2(n1312), .ZN(
        n943) );
  INVD1BWP12T U2057 ( .I(r3[28]), .ZN(n1310) );
  OAI22D1BWP12T U2058 ( .A1(n3406), .A2(n3539), .B1(n1310), .B2(n3434), .ZN(
        n942) );
  NR2D1BWP12T U2059 ( .A1(n943), .A2(n942), .ZN(n949) );
  TPND2D2BWP12T U2060 ( .A1(n3384), .A2(r1[28]), .ZN(n947) );
  INVD1BWP12T U2061 ( .I(tmp1[28]), .ZN(n944) );
  INVD1BWP12T U2062 ( .I(r2[28]), .ZN(n1322) );
  OAI22D1BWP12T U2063 ( .A1(n3378), .A2(n944), .B1(n1322), .B2(n3432), .ZN(
        n946) );
  INVD1BWP12T U2064 ( .I(r5[28]), .ZN(n1315) );
  INVD1BWP12T U2065 ( .I(r7[28]), .ZN(n1313) );
  OAI22D1BWP12T U2066 ( .A1(n3381), .A2(n1315), .B1(n1313), .B2(n3444), .ZN(
        n945) );
  INR3D0BWP12T U2067 ( .A1(n947), .B1(n946), .B2(n945), .ZN(n948) );
  ND3D1BWP12T U2068 ( .A1(n950), .A2(n949), .A3(n948), .ZN(regA_out[28]) );
  CKND3BWP12T U2069 ( .I(write1_in[29]), .ZN(n3512) );
  AOI21D1BWP12T U2070 ( .A1(n1900), .A2(r9[5]), .B(n951), .ZN(n954) );
  NR2D1BWP12T U2071 ( .A1(n1896), .A2(n2020), .ZN(n952) );
  AOI21D1BWP12T U2072 ( .A1(n1898), .A2(n[3575]), .B(n952), .ZN(n953) );
  TPND2D1BWP12T U2073 ( .A1(n954), .A2(n953), .ZN(n963) );
  INVD1BWP12T U2074 ( .I(r11[5]), .ZN(n2869) );
  ND2D1BWP12T U2075 ( .A1(n1674), .A2(r5[5]), .ZN(n955) );
  TPND2D2BWP12T U2076 ( .A1(n1892), .A2(r0[5]), .ZN(n956) );
  INVD1P75BWP12T U2077 ( .I(n956), .ZN(n959) );
  TPNR2D2BWP12T U2078 ( .A1(n959), .A2(n958), .ZN(n960) );
  IND2D2BWP12T U2079 ( .A1(n961), .B1(n960), .ZN(n962) );
  TPNR2D2BWP12T U2080 ( .A1(n963), .A2(n962), .ZN(n982) );
  CKND0BWP12T U2081 ( .I(pc_out[5]), .ZN(n968) );
  INVD0BWP12T U2082 ( .I(n964), .ZN(n1696) );
  IND3D1BWP12T U2083 ( .A1(n966), .B1(n1696), .B2(n965), .ZN(n967) );
  OAI21D1BWP12T U2084 ( .A1(n968), .A2(n1703), .B(n967), .ZN(n973) );
  INVD1BWP12T U2085 ( .I(r12[5]), .ZN(n2018) );
  ND2D1BWP12T U2086 ( .A1(n1918), .A2(r4[5]), .ZN(n969) );
  TPOAI21D1BWP12T U2087 ( .A1(n1920), .A2(n2018), .B(n969), .ZN(n972) );
  INVD1BWP12T U2088 ( .I(r8[5]), .ZN(n2019) );
  ND2D1BWP12T U2089 ( .A1(n1526), .A2(tmp1[5]), .ZN(n970) );
  TPNR3D2BWP12T U2090 ( .A1(n973), .A2(n972), .A3(n971), .ZN(n981) );
  NR2D1BWP12T U2091 ( .A1(n1519), .A2(n2021), .ZN(n978) );
  NR2D1BWP12T U2092 ( .A1(n1911), .A2(n976), .ZN(n977) );
  NR3D3BWP12T U2093 ( .A1(n979), .A2(n978), .A3(n977), .ZN(n980) );
  INVD1BWP12T U2094 ( .I(pc_out[10]), .ZN(n1401) );
  INR2D1BWP12T U2095 ( .A1(pc_out[10]), .B1(n1917), .ZN(n983) );
  INVD1BWP12T U2096 ( .I(r1[10]), .ZN(n3013) );
  INVD1BWP12T U2097 ( .I(r2[10]), .ZN(n2971) );
  OAI22D1BWP12T U2098 ( .A1(n1659), .A2(n3013), .B1(n1519), .B2(n2971), .ZN(
        n985) );
  INVD1BWP12T U2099 ( .I(n985), .ZN(n988) );
  INVD1BWP12T U2100 ( .I(lr[10]), .ZN(n3023) );
  AOI22D1BWP12T U2101 ( .A1(n1921), .A2(tmp1[10]), .B1(r8[10]), .B2(n1571), 
        .ZN(n991) );
  AOI22D1BWP12T U2102 ( .A1(n1527), .A2(r12[10]), .B1(n1918), .B2(r4[10]), 
        .ZN(n990) );
  ND2D1BWP12T U2103 ( .A1(n991), .A2(n990), .ZN(n992) );
  TPNR2D1BWP12T U2104 ( .A1(n993), .A2(n992), .ZN(n1001) );
  INVD1BWP12T U2105 ( .I(r0[10]), .ZN(n2979) );
  INVD1BWP12T U2106 ( .I(r7[10]), .ZN(n3001) );
  OAI22D1BWP12T U2107 ( .A1(n1587), .A2(n2979), .B1(n3001), .B2(n1724), .ZN(
        n995) );
  TPOAI22D1BWP12T U2108 ( .A1(n1663), .A2(n3017), .B1(n1899), .B2(n2975), .ZN(
        n994) );
  OR2XD2BWP12T U2109 ( .A1(n995), .A2(n994), .Z(n999) );
  INVD1BWP12T U2110 ( .I(n[3570]), .ZN(n1400) );
  INVD1BWP12T U2111 ( .I(r3[10]), .ZN(n2967) );
  OAI22D1BWP12T U2112 ( .A1(n1652), .A2(n1400), .B1(n2967), .B2(n1896), .ZN(
        n997) );
  INVD1BWP12T U2113 ( .I(r11[10]), .ZN(n2963) );
  INVD1BWP12T U2114 ( .I(r5[10]), .ZN(n3005) );
  OR2XD2BWP12T U2115 ( .A1(n997), .A2(n996), .Z(n998) );
  NR2XD2BWP12T U2116 ( .A1(n999), .A2(n998), .ZN(n1000) );
  TPND2D2BWP12T U2117 ( .A1(n1001), .A2(n1000), .ZN(regB_out[10]) );
  AOI22D1BWP12T U2118 ( .A1(n1575), .A2(pc_out[13]), .B1(r6[13]), .B2(n1915), 
        .ZN(n1004) );
  INVD1BWP12T U2119 ( .I(lr[13]), .ZN(n2050) );
  AOI22D1BWP12T U2120 ( .A1(n1921), .A2(tmp1[13]), .B1(r8[13]), .B2(n1571), 
        .ZN(n1010) );
  CKND1BWP12T U2121 ( .I(r1[13]), .ZN(n1006) );
  CKND1BWP12T U2122 ( .I(r2[13]), .ZN(n1005) );
  TPOAI22D1BWP12T U2123 ( .A1(n1659), .A2(n1006), .B1(n1519), .B2(n1005), .ZN(
        n1007) );
  ND3D2BWP12T U2124 ( .A1(n1010), .A2(n1009), .A3(n1008), .ZN(n1011) );
  INVD1BWP12T U2125 ( .I(r9[13]), .ZN(n1015) );
  INR2D2BWP12T U2126 ( .A1(r10[13]), .B1(n1899), .ZN(n1013) );
  OAI21D1BWP12T U2127 ( .A1(n1663), .A2(n1015), .B(n1014), .ZN(n1018) );
  INVD1BWP12T U2128 ( .I(r0[13]), .ZN(n1046) );
  CKND1BWP12T U2129 ( .I(r7[13]), .ZN(n1016) );
  OR2XD2BWP12T U2130 ( .A1(n1018), .A2(n1017), .Z(n1024) );
  INVD1BWP12T U2131 ( .I(n[3567]), .ZN(n2051) );
  INVD1BWP12T U2132 ( .I(r3[13]), .ZN(n1053) );
  OAI22D1BWP12T U2133 ( .A1(n1652), .A2(n2051), .B1(n1053), .B2(n1896), .ZN(
        n1022) );
  INVD1BWP12T U2134 ( .I(r11[13]), .ZN(n1065) );
  CKND1BWP12T U2135 ( .I(r5[13]), .ZN(n1019) );
  TPOAI22D1BWP12T U2136 ( .A1(n1887), .A2(n1065), .B1(n161), .B2(n1019), .ZN(
        n1020) );
  IND2XD2BWP12T U2137 ( .A1(n1022), .B1(n1021), .ZN(n1023) );
  NR2D0BWP12T U2138 ( .A1(n530), .A2(write2_in[28]), .ZN(n1029) );
  TPNR2D0BWP12T U2139 ( .A1(n3343), .A2(n3539), .ZN(n1030) );
  TPAOI21D0BWP12T U2140 ( .A1(next_pc_in[28]), .A2(n3499), .B(n1030), .ZN(
        n1031) );
  TPOAI21D1BWP12T U2141 ( .A1(n1033), .A2(n1032), .B(n1031), .ZN(n1034) );
  AOI21D1BWP12T U2142 ( .A1(n1035), .A2(n1036), .B(n1034), .ZN(n1044) );
  DCCKND4BWP12T U2143 ( .I(n1036), .ZN(n1042) );
  TPNR3D4BWP12T U2144 ( .A1(n1038), .A2(n1037), .A3(n3497), .ZN(n1041) );
  ND2D1BWP12T U2145 ( .A1(write1_in[28]), .A2(n530), .ZN(n1040) );
  ND3XD3BWP12T U2146 ( .A1(n1042), .A2(n1041), .A3(n1040), .ZN(n1043) );
  ND2D2BWP12T U2147 ( .A1(n1044), .A2(n1043), .ZN(n2196) );
  ND2D1BWP12T U2148 ( .A1(n1380), .A2(tmp1[13]), .ZN(n1045) );
  INR2D2BWP12T U2149 ( .A1(r6[13]), .B1(n3396), .ZN(n1052) );
  INVD1BWP12T U2150 ( .I(n1047), .ZN(n1048) );
  INR2D1BWP12T U2151 ( .A1(r9[13]), .B1(n1048), .ZN(n1050) );
  AN2D1BWP12T U2152 ( .A1(n1050), .A2(n1049), .Z(n1051) );
  RCAOI21D1BWP12T U2153 ( .A1(n1473), .A2(r8[13]), .B(n1054), .ZN(n1056) );
  ND2D1BWP12T U2154 ( .A1(n1862), .A2(n[3567]), .ZN(n1055) );
  TPND3D2BWP12T U2155 ( .A1(n1057), .A2(n1056), .A3(n1055), .ZN(n1058) );
  INR3D4BWP12T U2156 ( .A1(n1060), .B1(n1059), .B2(n1058), .ZN(n1076) );
  ND2D1BWP12T U2157 ( .A1(n3417), .A2(r1[13]), .ZN(n1061) );
  OAI21D1BWP12T U2158 ( .A1(n3416), .A2(n2050), .B(n1061), .ZN(n1068) );
  TPND2D2BWP12T U2159 ( .A1(n1788), .A2(pc_out[13]), .ZN(n1063) );
  ND2D1BWP12T U2160 ( .A1(n1873), .A2(r5[13]), .ZN(n1062) );
  TPND2D2BWP12T U2161 ( .A1(n1063), .A2(n1062), .ZN(n1067) );
  ND2D1BWP12T U2162 ( .A1(n1804), .A2(immediate1_in[13]), .ZN(n1064) );
  OAI21D1BWP12T U2163 ( .A1(n3393), .A2(n1065), .B(n1064), .ZN(n1066) );
  TPNR3D2BWP12T U2164 ( .A1(n1068), .A2(n1067), .A3(n1066), .ZN(n1075) );
  INR2D1BWP12T U2165 ( .A1(r12[13]), .B1(n3436), .ZN(n1070) );
  TPNR2D1BWP12T U2166 ( .A1(n1070), .A2(n186), .ZN(n1073) );
  ND2D1BWP12T U2167 ( .A1(n1839), .A2(r7[13]), .ZN(n1072) );
  ND2D1BWP12T U2168 ( .A1(n1622), .A2(r2[13]), .ZN(n1071) );
  AN3D4BWP12T U2169 ( .A1(n1073), .A2(n1072), .A3(n1071), .Z(n1074) );
  ND3D4BWP12T U2170 ( .A1(n1076), .A2(n1075), .A3(n1074), .ZN(regA_out[13]) );
  INVD1BWP12T U2171 ( .I(r11[31]), .ZN(n3360) );
  INVD1BWP12T U2172 ( .I(r5[31]), .ZN(n3353) );
  INVD1BWP12T U2173 ( .I(r3[31]), .ZN(n3370) );
  MOAI22D0BWP12T U2174 ( .A1(n3370), .A2(n1896), .B1(n1690), .B2(n[3549]), 
        .ZN(n1077) );
  AOI22D0BWP12T U2175 ( .A1(n1571), .A2(r8[31]), .B1(tmp1[31]), .B2(n1526), 
        .ZN(n1079) );
  INVD1BWP12T U2176 ( .I(n1079), .ZN(n1080) );
  INVD1BWP12T U2177 ( .I(r9[31]), .ZN(n3368) );
  TPOAI22D1BWP12T U2178 ( .A1(n1553), .A2(n3368), .B1(n1592), .B2(n3510), .ZN(
        n1083) );
  INVD1BWP12T U2179 ( .I(r0[31]), .ZN(n3361) );
  INVD1BWP12T U2180 ( .I(r7[31]), .ZN(n3352) );
  TPOAI22D1BWP12T U2181 ( .A1(n1587), .A2(n3361), .B1(n3352), .B2(n1724), .ZN(
        n1082) );
  OR2D2BWP12T U2182 ( .A1(n1083), .A2(n1082), .Z(n1087) );
  AOI22D1BWP12T U2183 ( .A1(n1575), .A2(pc_out[31]), .B1(r6[31]), .B2(n1915), 
        .ZN(n1085) );
  AOI22D1BWP12T U2184 ( .A1(n1664), .A2(r12[31]), .B1(n1918), .B2(r4[31]), 
        .ZN(n1084) );
  NR2D2BWP12T U2185 ( .A1(n1087), .A2(n1086), .ZN(n1092) );
  INVD0BWP12T U2186 ( .I(r1[31]), .ZN(n1088) );
  INVD1BWP12T U2187 ( .I(r2[31]), .ZN(n3350) );
  OAI22D1BWP12T U2188 ( .A1(n1911), .A2(n1088), .B1(n1519), .B2(n3350), .ZN(
        n1090) );
  INVD1BWP12T U2189 ( .I(lr[31]), .ZN(n3357) );
  ND3D2BWP12T U2190 ( .A1(n1093), .A2(n1092), .A3(n1091), .ZN(regB_out[31]) );
  AOI22D1BWP12T U2191 ( .A1(n1526), .A2(tmp1[15]), .B1(r8[15]), .B2(n1571), 
        .ZN(n1103) );
  INVD1BWP12T U2192 ( .I(lr[15]), .ZN(n1094) );
  AOI22D1BWP12T U2193 ( .A1(n1527), .A2(r12[15]), .B1(n1918), .B2(r4[15]), 
        .ZN(n1100) );
  CKND2D2BWP12T U2194 ( .A1(n1907), .A2(immediate2_in[15]), .ZN(n1099) );
  INVD1BWP12T U2195 ( .I(r2[15]), .ZN(n1377) );
  INVD1BWP12T U2196 ( .I(r1[15]), .ZN(n1096) );
  TPOAI22D2BWP12T U2197 ( .A1(n1519), .A2(n1377), .B1(n1659), .B2(n1096), .ZN(
        n1097) );
  INVD1P75BWP12T U2198 ( .I(n1097), .ZN(n1098) );
  ND3D2BWP12T U2199 ( .A1(n1100), .A2(n1099), .A3(n1098), .ZN(n1101) );
  INR3XD2BWP12T U2200 ( .A1(n1103), .B1(n1102), .B2(n1101), .ZN(n1109) );
  INVD1BWP12T U2201 ( .I(n[3565]), .ZN(n1368) );
  INVD1BWP12T U2202 ( .I(r3[15]), .ZN(n1387) );
  TPOAI22D1BWP12T U2203 ( .A1(n1652), .A2(n1368), .B1(n1387), .B2(n1896), .ZN(
        n1107) );
  INVD1BWP12T U2204 ( .I(r9[15]), .ZN(n2662) );
  INVD1BWP12T U2205 ( .I(r10[15]), .ZN(n1367) );
  INVD1BWP12T U2206 ( .I(r11[15]), .ZN(n2663) );
  MOAI22D1BWP12T U2207 ( .A1(n1887), .A2(n2663), .B1(n1674), .B2(r5[15]), .ZN(
        n1105) );
  INVD1BWP12T U2208 ( .I(r0[15]), .ZN(n1375) );
  INVD1BWP12T U2209 ( .I(r7[15]), .ZN(n1391) );
  TPOAI22D2BWP12T U2210 ( .A1(n1587), .A2(n1375), .B1(n1391), .B2(n1895), .ZN(
        n1104) );
  NR4D2BWP12T U2211 ( .A1(n1107), .A2(n1106), .A3(n1105), .A4(n1104), .ZN(
        n1108) );
  AOI22D1BWP12T U2212 ( .A1(n1921), .A2(tmp1[18]), .B1(r8[18]), .B2(n1571), 
        .ZN(n1117) );
  INVD1BWP12T U2213 ( .I(r1[18]), .ZN(n3423) );
  INVD1BWP12T U2214 ( .I(r2[18]), .ZN(n3431) );
  TPOAI22D1BWP12T U2215 ( .A1(n1911), .A2(n3423), .B1(n1519), .B2(n3431), .ZN(
        n1111) );
  AOI22D1BWP12T U2216 ( .A1(n1527), .A2(r12[18]), .B1(n1918), .B2(r4[18]), 
        .ZN(n1110) );
  AOI22D1BWP12T U2217 ( .A1(n1575), .A2(pc_out[18]), .B1(r6[18]), .B2(n1915), 
        .ZN(n1114) );
  INVD1BWP12T U2218 ( .I(lr[18]), .ZN(n3415) );
  OR2XD1BWP12T U2219 ( .A1(n1714), .A2(n3415), .Z(n1113) );
  INR3XD1BWP12T U2220 ( .A1(n1117), .B1(n1116), .B2(n1115), .ZN(n1124) );
  INVD1BWP12T U2221 ( .I(n[3562]), .ZN(n2099) );
  INVD1BWP12T U2222 ( .I(r3[18]), .ZN(n3433) );
  OAI22D1BWP12T U2223 ( .A1(n1652), .A2(n2099), .B1(n3433), .B2(n1896), .ZN(
        n1122) );
  INVD0BWP12T U2224 ( .I(r9[18]), .ZN(n1118) );
  INVD1BWP12T U2225 ( .I(r10[18]), .ZN(n3453) );
  OAI22D1BWP12T U2226 ( .A1(n1663), .A2(n1118), .B1(n3453), .B2(n1592), .ZN(
        n1121) );
  INVD1BWP12T U2227 ( .I(r0[18]), .ZN(n3441) );
  INVD1BWP12T U2228 ( .I(r7[18]), .ZN(n3443) );
  OAI22D1BWP12T U2229 ( .A1(n1587), .A2(n3441), .B1(n3443), .B2(n1895), .ZN(
        n1120) );
  INVD1BWP12T U2230 ( .I(r11[18]), .ZN(n2098) );
  INVD1BWP12T U2231 ( .I(r5[18]), .ZN(n3413) );
  NR4D1BWP12T U2232 ( .A1(n1122), .A2(n1121), .A3(n1120), .A4(n1119), .ZN(
        n1123) );
  CKND2D2BWP12T U2233 ( .A1(n1124), .A2(n1123), .ZN(regB_out[18]) );
  AOI22D0BWP12T U2234 ( .A1(n3186), .A2(n[3551]), .B1(write2_in[29]), .B2(
        n3185), .ZN(n1125) );
  ND2D1BWP12T U2235 ( .A1(n1126), .A2(n1125), .ZN(spin[29]) );
  TPNR2D3BWP12T U2236 ( .A1(n1127), .A2(n3504), .ZN(n3301) );
  INVD1BWP12T U2237 ( .I(n3301), .ZN(n1133) );
  ND2D1BWP12T U2238 ( .A1(n3331), .A2(write2_in[25]), .ZN(n1128) );
  ND2D1BWP12T U2239 ( .A1(write1_in[23]), .A2(n530), .ZN(n1130) );
  CKND2D1BWP12T U2240 ( .A1(n3331), .A2(write2_in[23]), .ZN(n1129) );
  CKND2D2BWP12T U2241 ( .A1(n1130), .A2(n1129), .ZN(n3299) );
  CKND2D1BWP12T U2242 ( .A1(n3331), .A2(write2_in[24]), .ZN(n1131) );
  RCOAI21D2BWP12T U2243 ( .A1(n162), .A2(n3331), .B(n1131), .ZN(n3307) );
  ND4D1BWP12T U2244 ( .A1(n3311), .A2(n1135), .A3(n3299), .A4(n3307), .ZN(
        n1132) );
  TPNR2D1BWP12T U2245 ( .A1(n1133), .A2(n1132), .ZN(n1142) );
  CKAN2D0BWP12T U2246 ( .A1(n3331), .A2(write2_in[26]), .Z(n1134) );
  AOI21D1BWP12T U2247 ( .A1(write1_in[26]), .A2(n530), .B(n1134), .ZN(n1138)
         );
  INR2D1BWP12T U2248 ( .A1(n3505), .B1(n1138), .ZN(n1137) );
  INVD1BWP12T U2249 ( .I(n1135), .ZN(n1136) );
  NR2D1BWP12T U2250 ( .A1(n1137), .A2(n1136), .ZN(n1141) );
  ND2D1BWP12T U2251 ( .A1(n3301), .A2(n3299), .ZN(n3315) );
  CKAN2D2BWP12T U2252 ( .A1(n1138), .A2(n3311), .Z(n1139) );
  TPND2D2BWP12T U2253 ( .A1(n1139), .A2(n3298), .ZN(n1140) );
  TPOAI22D1BWP12T U2254 ( .A1(n1142), .A2(n1141), .B1(n3315), .B2(n1140), .ZN(
        n2194) );
  AOI22D1BWP12T U2255 ( .A1(n1921), .A2(tmp1[9]), .B1(r8[9]), .B2(n1571), .ZN(
        n1144) );
  AOI22D1BWP12T U2256 ( .A1(n1527), .A2(r12[9]), .B1(n1918), .B2(r4[9]), .ZN(
        n1143) );
  INVD1BWP12T U2257 ( .I(r1[9]), .ZN(n2983) );
  OAI22D1BWP12T U2258 ( .A1(n1659), .A2(n2983), .B1(n1519), .B2(n2943), .ZN(
        n1150) );
  INVD1BWP12T U2259 ( .I(lr[9]), .ZN(n2990) );
  MOAI22D1BWP12T U2260 ( .A1(n2990), .A2(n1669), .B1(n1668), .B2(
        immediate2_in[9]), .ZN(n1149) );
  ND2D1BWP12T U2261 ( .A1(n1915), .A2(r6[9]), .ZN(n1147) );
  INVD1BWP12T U2262 ( .I(pc_out[9]), .ZN(n1194) );
  INR2D1BWP12T U2263 ( .A1(pc_out[9]), .B1(n1703), .ZN(n1145) );
  INVD1BWP12T U2264 ( .I(n1145), .ZN(n1146) );
  ND2D1BWP12T U2265 ( .A1(n1147), .A2(n1146), .ZN(n1148) );
  NR4D0BWP12T U2266 ( .A1(n1151), .A2(n1150), .A3(n1149), .A4(n1148), .ZN(
        n1159) );
  INVD1BWP12T U2267 ( .I(n[3571]), .ZN(n2887) );
  INVD1BWP12T U2268 ( .I(r3[9]), .ZN(n2946) );
  OAI22D1BWP12T U2269 ( .A1(n1652), .A2(n2887), .B1(n2946), .B2(n1896), .ZN(
        n1157) );
  INR2D2BWP12T U2270 ( .A1(r10[9]), .B1(n1899), .ZN(n1152) );
  OAI21D1BWP12T U2271 ( .A1(n1663), .A2(n2984), .B(n1153), .ZN(n1156) );
  INVD1BWP12T U2272 ( .I(r0[9]), .ZN(n2945) );
  INVD1BWP12T U2273 ( .I(r7[9]), .ZN(n2986) );
  OAI22D1BWP12T U2274 ( .A1(n1587), .A2(n2945), .B1(n2986), .B2(n1724), .ZN(
        n1155) );
  INVD1BWP12T U2275 ( .I(r11[9]), .ZN(n2947) );
  NR4D0BWP12T U2276 ( .A1(n1157), .A2(n1156), .A3(n1155), .A4(n1154), .ZN(
        n1158) );
  TPND2D1BWP12T U2277 ( .A1(n1159), .A2(n1158), .ZN(regB_out[9]) );
  INVD3BWP12T U2278 ( .I(write1_in[19]), .ZN(n3094) );
  ND2D1BWP12T U2279 ( .A1(n3331), .A2(write2_in[19]), .ZN(n1160) );
  XNR2D1BWP12T U2280 ( .A1(n3503), .A2(n3502), .ZN(n1162) );
  AOI22D1BWP12T U2281 ( .A1(next_pc_in[19]), .A2(n3499), .B1(n3498), .B2(
        pc_out[19]), .ZN(n1161) );
  TPOAI21D1BWP12T U2282 ( .A1(n1162), .A2(n3497), .B(n1161), .ZN(n2187) );
  TPND2D1BWP12T U2283 ( .A1(n1164), .A2(n1163), .ZN(n1168) );
  INR2D2BWP12T U2284 ( .A1(r10[4]), .B1(n1899), .ZN(n1165) );
  INVD1P75BWP12T U2285 ( .I(n1165), .ZN(n1166) );
  TPOAI21D1BWP12T U2286 ( .A1(n1663), .A2(n2842), .B(n1166), .ZN(n1167) );
  TPNR2D2BWP12T U2287 ( .A1(n1168), .A2(n1167), .ZN(n1184) );
  MOAI22D0BWP12T U2288 ( .A1(n2843), .A2(n1669), .B1(n1713), .B2(
        immediate2_in[4]), .ZN(n1173) );
  OR2D2BWP12T U2289 ( .A1(n1703), .A2(n1169), .Z(n1171) );
  ND2D3BWP12T U2290 ( .A1(n1915), .A2(r6[4]), .ZN(n1170) );
  TPND2D1BWP12T U2291 ( .A1(n1171), .A2(n1170), .ZN(n1172) );
  TPNR2D2BWP12T U2292 ( .A1(n1173), .A2(n1172), .ZN(n1183) );
  OAI22D1BWP12T U2293 ( .A1(n1911), .A2(n1174), .B1(n1519), .B2(n2012), .ZN(
        n1176) );
  MOAI22D1BWP12T U2294 ( .A1(n1887), .A2(n2011), .B1(n1674), .B2(r5[4]), .ZN(
        n1175) );
  TPNR2D2BWP12T U2295 ( .A1(n1175), .A2(n1176), .ZN(n1182) );
  OAI22D1BWP12T U2296 ( .A1(n1587), .A2(n2007), .B1(n1177), .B2(n1724), .ZN(
        n1180) );
  OAI22D1BWP12T U2297 ( .A1(n1652), .A2(n1178), .B1(n2013), .B2(n1896), .ZN(
        n1179) );
  TPNR2D2BWP12T U2298 ( .A1(n1180), .A2(n1179), .ZN(n1181) );
  ND4D4BWP12T U2299 ( .A1(n1184), .A2(n1183), .A3(n1182), .A4(n1181), .ZN(
        regB_out[4]) );
  INVD1BWP12T U2300 ( .I(r4[9]), .ZN(n2944) );
  INVD1BWP12T U2301 ( .I(r8[9]), .ZN(n2942) );
  INVD1BWP12T U2302 ( .I(r12[9]), .ZN(n2948) );
  OAI22D1BWP12T U2303 ( .A1(n2942), .A2(n3387), .B1(n3436), .B2(n2948), .ZN(
        n1186) );
  INVD1BWP12T U2304 ( .I(r10[9]), .ZN(n2941) );
  NR4D1BWP12T U2305 ( .A1(n1188), .A2(n1187), .A3(n1186), .A4(n1185), .ZN(
        n1199) );
  AOI21D1BWP12T U2306 ( .A1(n3412), .A2(r6[9]), .B(n1189), .ZN(n1191) );
  AOI22D1BWP12T U2307 ( .A1(n1876), .A2(tmp1[9]), .B1(n1804), .B2(
        immediate1_in[9]), .ZN(n1190) );
  TPND2D1BWP12T U2308 ( .A1(n1191), .A2(n1190), .ZN(n1193) );
  OAI22D2BWP12T U2309 ( .A1(n3446), .A2(n2887), .B1(n2946), .B2(n3434), .ZN(
        n1192) );
  TPNR2D2BWP12T U2310 ( .A1(n1193), .A2(n1192), .ZN(n1198) );
  OAI22D1BWP12T U2311 ( .A1(n3406), .A2(n1194), .B1(n2986), .B2(n3444), .ZN(
        n1196) );
  INVD1BWP12T U2312 ( .I(r5[9]), .ZN(n2987) );
  OAI22D1BWP12T U2313 ( .A1(n3414), .A2(n2987), .B1(n1810), .B2(n2983), .ZN(
        n1195) );
  TPNR2D1BWP12T U2314 ( .A1(n1196), .A2(n1195), .ZN(n1197) );
  ND3D2BWP12T U2315 ( .A1(n1199), .A2(n1198), .A3(n1197), .ZN(regA_out[9]) );
  ND2D1BWP12T U2316 ( .A1(n1876), .A2(tmp1[16]), .ZN(n1203) );
  ND2D1BWP12T U2317 ( .A1(n3419), .A2(r9[16]), .ZN(n1202) );
  ND3D1BWP12T U2318 ( .A1(n1203), .A2(n1202), .A3(n1201), .ZN(n1207) );
  NR2D1BWP12T U2319 ( .A1(n1204), .A2(n3404), .ZN(n1205) );
  NR3D1BWP12T U2320 ( .A1(n1207), .A2(n1206), .A3(n1205), .ZN(n1229) );
  ND2D1BWP12T U2321 ( .A1(n3412), .A2(r6[16]), .ZN(n1218) );
  ND2D1BWP12T U2322 ( .A1(n3417), .A2(r1[16]), .ZN(n1208) );
  INVD1BWP12T U2323 ( .I(r8[16]), .ZN(n1210) );
  TPOAI22D1BWP12T U2324 ( .A1(n3435), .A2(n1210), .B1(n3432), .B2(n1209), .ZN(
        n1213) );
  TPNR2D1BWP12T U2325 ( .A1(n3434), .A2(n1211), .ZN(n1212) );
  TPNR2D1BWP12T U2326 ( .A1(n1213), .A2(n1212), .ZN(n1215) );
  ND2D1BWP12T U2327 ( .A1(n1873), .A2(r5[16]), .ZN(n1214) );
  TPND2D1BWP12T U2328 ( .A1(n1215), .A2(n1214), .ZN(n1216) );
  INR3D2BWP12T U2329 ( .A1(n1218), .B1(n1217), .B2(n1216), .ZN(n1228) );
  ND2D1BWP12T U2330 ( .A1(n1219), .A2(lr[16]), .ZN(n1220) );
  ND2D1BWP12T U2331 ( .A1(n1221), .A2(n1220), .ZN(n1226) );
  INR2D1BWP12T U2332 ( .A1(r7[16]), .B1(n3444), .ZN(n1225) );
  ND3D2BWP12T U2333 ( .A1(n1229), .A2(n1228), .A3(n1227), .ZN(regA_out[16]) );
  TPOAI22D1BWP12T U2334 ( .A1(n1553), .A2(n1231), .B1(n1230), .B2(n1592), .ZN(
        n1235) );
  OR2XD2BWP12T U2335 ( .A1(n1235), .A2(n1234), .Z(n1242) );
  OAI22D1BWP12T U2336 ( .A1(n1887), .A2(n1237), .B1(n1889), .B2(n1236), .ZN(
        n1240) );
  NR2D1BWP12T U2337 ( .A1(n1714), .A2(n1243), .ZN(n1245) );
  IND2XD1BWP12T U2338 ( .A1(n1245), .B1(n1244), .ZN(n1246) );
  AO22XD2BWP12T U2339 ( .A1(n1921), .A2(tmp1[26]), .B1(r8[26]), .B2(n1571), 
        .Z(n1250) );
  ND3XD3BWP12T U2340 ( .A1(n1254), .A2(n1253), .A3(n1252), .ZN(regB_out[26])
         );
  INVD1BWP12T U2341 ( .I(n1255), .ZN(n1259) );
  AOI22D2BWP12T U2342 ( .A1(n1527), .A2(r12[3]), .B1(n1918), .B2(r4[3]), .ZN(
        n1258) );
  TPOAI22D1BWP12T U2343 ( .A1(n1519), .A2(n1960), .B1(n1659), .B2(n1809), .ZN(
        n1256) );
  INR2D1BWP12T U2344 ( .A1(pc_out[3]), .B1(n1703), .ZN(n1260) );
  INVD1BWP12T U2345 ( .I(n1260), .ZN(n1262) );
  ND2D1BWP12T U2346 ( .A1(n1915), .A2(r6[3]), .ZN(n1261) );
  TPND2D1BWP12T U2347 ( .A1(n1262), .A2(n1261), .ZN(n1264) );
  IND2XD2BWP12T U2348 ( .A1(n1264), .B1(n1263), .ZN(n1265) );
  INVD1BWP12T U2349 ( .I(n[3577]), .ZN(n2853) );
  INVD1BWP12T U2350 ( .I(r3[3]), .ZN(n1958) );
  OAI22D1BWP12T U2351 ( .A1(n1652), .A2(n2853), .B1(n1958), .B2(n1896), .ZN(
        n1271) );
  TPND2D1BWP12T U2352 ( .A1(n1674), .A2(r5[3]), .ZN(n1267) );
  TPOAI21D1BWP12T U2353 ( .A1(n1887), .A2(n2852), .B(n1267), .ZN(n1268) );
  NR4D1BWP12T U2354 ( .A1(n1271), .A2(n1270), .A3(n1269), .A4(n1268), .ZN(
        n1272) );
  TPND2D2BWP12T U2355 ( .A1(n1273), .A2(n1272), .ZN(regB_out[3]) );
  INVD1BWP12T U2356 ( .I(r11[2]), .ZN(n2755) );
  OAI22D1BWP12T U2357 ( .A1(n3416), .A2(n1670), .B1(n3393), .B2(n2755), .ZN(
        n1277) );
  INVD1BWP12T U2358 ( .I(r4[2]), .ZN(n2001) );
  INVD1BWP12T U2359 ( .I(r0[2]), .ZN(n1998) );
  OAI22D1BWP12T U2360 ( .A1(n3390), .A2(n2001), .B1(n1998), .B2(n3442), .ZN(
        n1276) );
  INVD1BWP12T U2361 ( .I(r12[2]), .ZN(n2000) );
  OAI22D1BWP12T U2362 ( .A1(n1673), .A2(n3387), .B1(n3436), .B2(n2000), .ZN(
        n1275) );
  INVD1BWP12T U2363 ( .I(r10[2]), .ZN(n2854) );
  OAI22D1BWP12T U2364 ( .A1(n3402), .A2(n2855), .B1(n2854), .B2(n3452), .ZN(
        n1274) );
  NR4D0BWP12T U2365 ( .A1(n1277), .A2(n1276), .A3(n1275), .A4(n1274), .ZN(
        n1288) );
  OAI22D1BWP12T U2366 ( .A1(n3406), .A2(n1679), .B1(n1672), .B2(n3444), .ZN(
        n1280) );
  OAI22D1BWP12T U2367 ( .A1(n3414), .A2(n1278), .B1(n1810), .B2(n1658), .ZN(
        n1279) );
  INVD1BWP12T U2368 ( .I(r2[2]), .ZN(n1999) );
  NR2D2BWP12T U2369 ( .A1(n3432), .A2(n1999), .ZN(n1281) );
  AOI22D1BWP12T U2370 ( .A1(n1876), .A2(tmp1[2]), .B1(n1804), .B2(
        immediate1_in[2]), .ZN(n1282) );
  ND2D1BWP12T U2371 ( .A1(n1283), .A2(n1282), .ZN(n1285) );
  INVD1BWP12T U2372 ( .I(n[3578]), .ZN(n2856) );
  INVD1BWP12T U2373 ( .I(r3[2]), .ZN(n2002) );
  OAI22D1BWP12T U2374 ( .A1(n3404), .A2(n2856), .B1(n2002), .B2(n3434), .ZN(
        n1284) );
  ND3D1BWP12T U2375 ( .A1(n1288), .A2(n1287), .A3(n1286), .ZN(regA_out[2]) );
  ND2D1BWP12T U2376 ( .A1(n3417), .A2(r1[11]), .ZN(n1289) );
  OAI21D1BWP12T U2377 ( .A1(n3444), .A2(n2878), .B(n1289), .ZN(n1295) );
  INVD1BWP12T U2378 ( .I(r6[11]), .ZN(n2880) );
  AOI21D1BWP12T U2379 ( .A1(n1873), .A2(r5[11]), .B(n1290), .ZN(n1293) );
  AOI21D1BWP12T U2380 ( .A1(n3418), .A2(r11[11]), .B(n1291), .ZN(n1292) );
  INR3D2BWP12T U2381 ( .A1(n1296), .B1(n1295), .B2(n1294), .ZN(n1309) );
  INVD1BWP12T U2382 ( .I(r10[11]), .ZN(n2900) );
  INVD1BWP12T U2383 ( .I(n[3569]), .ZN(n1297) );
  INVD1BWP12T U2384 ( .I(r12[11]), .ZN(n2898) );
  ND2D1BWP12T U2385 ( .A1(n1804), .A2(immediate1_in[11]), .ZN(n1299) );
  NR3D1BWP12T U2386 ( .A1(n1303), .A2(n1302), .A3(n1301), .ZN(n1308) );
  INVD1BWP12T U2387 ( .I(r8[11]), .ZN(n3025) );
  INR3D2BWP12T U2388 ( .A1(n1306), .B1(n1305), .B2(n1304), .ZN(n1307) );
  ND3XD3BWP12T U2389 ( .A1(n1309), .A2(n1308), .A3(n1307), .ZN(regA_out[11])
         );
  OAI22D1BWP12T U2390 ( .A1(n1652), .A2(n2680), .B1(n1310), .B2(n1896), .ZN(
        n1319) );
  OAI22D1BWP12T U2391 ( .A1(n1553), .A2(n1312), .B1(n1311), .B2(n1592), .ZN(
        n1318) );
  OAI22D1BWP12T U2392 ( .A1(n1587), .A2(n1314), .B1(n1313), .B2(n1895), .ZN(
        n1317) );
  TPOAI22D1BWP12T U2393 ( .A1(n1887), .A2(n2679), .B1(n160), .B2(n1315), .ZN(
        n1316) );
  NR4D1BWP12T U2394 ( .A1(n1319), .A2(n1318), .A3(n1317), .A4(n1316), .ZN(
        n1331) );
  NR2D1BWP12T U2395 ( .A1(n167), .A2(n1320), .ZN(n1324) );
  INVD0BWP12T U2396 ( .I(r1[28]), .ZN(n1321) );
  OAI22D0BWP12T U2397 ( .A1(n1519), .A2(n1322), .B1(n1911), .B2(n1321), .ZN(
        n1323) );
  INR3D2BWP12T U2398 ( .A1(n1325), .B1(n1324), .B2(n1323), .ZN(n1330) );
  AOI22D1BWP12T U2399 ( .A1(n1575), .A2(pc_out[28]), .B1(r6[28]), .B2(n1915), 
        .ZN(n1328) );
  AOI22D1BWP12T U2400 ( .A1(n1664), .A2(r12[28]), .B1(n1918), .B2(r4[28]), 
        .ZN(n1326) );
  AOI22D1BWP12T U2401 ( .A1(n1921), .A2(tmp1[19]), .B1(r8[19]), .B2(n1571), 
        .ZN(n1340) );
  AOI22D1BWP12T U2402 ( .A1(n1664), .A2(r12[19]), .B1(n1918), .B2(r4[19]), 
        .ZN(n1332) );
  IOA21D1BWP12T U2403 ( .A1(n1907), .A2(immediate2_in[19]), .B(n1332), .ZN(
        n1339) );
  INVD3BWP12T U2404 ( .I(n1703), .ZN(n1532) );
  CKND1BWP12T U2405 ( .I(r1[19]), .ZN(n1334) );
  CKND0BWP12T U2406 ( .I(lr[19]), .ZN(n1335) );
  INR3D2BWP12T U2407 ( .A1(n1340), .B1(n1339), .B2(n1338), .ZN(n1352) );
  OAI22D1BWP12T U2408 ( .A1(n1652), .A2(n2069), .B1(n1341), .B2(n1896), .ZN(
        n1350) );
  CKND0BWP12T U2409 ( .I(r9[19]), .ZN(n1342) );
  OAI22D1BWP12T U2410 ( .A1(n1553), .A2(n1342), .B1(n2070), .B2(n1592), .ZN(
        n1349) );
  OAI22D1BWP12T U2411 ( .A1(n1587), .A2(n1344), .B1(n1343), .B2(n1895), .ZN(
        n1348) );
  CKND0BWP12T U2412 ( .I(r11[19]), .ZN(n1346) );
  OAI22D1BWP12T U2413 ( .A1(n1887), .A2(n1346), .B1(n160), .B2(n1345), .ZN(
        n1347) );
  AOI21D1BWP12T U2414 ( .A1(n3412), .A2(r6[8]), .B(n1353), .ZN(n1355) );
  AOI22D1BWP12T U2415 ( .A1(n1876), .A2(tmp1[8]), .B1(n1804), .B2(
        immediate1_in[8]), .ZN(n1354) );
  INVD1BWP12T U2416 ( .I(n[3572]), .ZN(n1356) );
  INVD1BWP12T U2417 ( .I(r5[8]), .ZN(n2929) );
  OAI22D1BWP12T U2418 ( .A1(n3416), .A2(n2996), .B1(n3393), .B2(n2907), .ZN(
        n1364) );
  INVD1BWP12T U2419 ( .I(r4[8]), .ZN(n2903) );
  INVD1BWP12T U2420 ( .I(r0[8]), .ZN(n2904) );
  INVD1BWP12T U2421 ( .I(r9[8]), .ZN(n2935) );
  OAI22D1BWP12T U2422 ( .A1(n3402), .A2(n2935), .B1(n2995), .B2(n3452), .ZN(
        n1361) );
  NR4D0BWP12T U2423 ( .A1(n1364), .A2(n1363), .A3(n1362), .A4(n1361), .ZN(
        n1365) );
  NR2D1BWP12T U2424 ( .A1(n1881), .A2(n1367), .ZN(n1370) );
  INR3D2BWP12T U2425 ( .A1(n1371), .B1(n1370), .B2(n1369), .ZN(n1396) );
  AOI21D1BWP12T U2426 ( .A1(n1853), .A2(r4[15]), .B(n1373), .ZN(n1386) );
  OAI21D1BWP12T U2427 ( .A1(n3442), .A2(n1375), .B(n1374), .ZN(n1385) );
  INVD1P75BWP12T U2428 ( .I(n1376), .ZN(n1379) );
  INR2D2BWP12T U2429 ( .A1(r2[15]), .B1(n1787), .ZN(n1378) );
  TPNR2D2BWP12T U2430 ( .A1(n1379), .A2(n1378), .ZN(n1383) );
  ND2D1BWP12T U2431 ( .A1(n3417), .A2(r1[15]), .ZN(n1382) );
  ND2D1BWP12T U2432 ( .A1(n1380), .A2(tmp1[15]), .ZN(n1381) );
  INR3D2BWP12T U2433 ( .A1(n1386), .B1(n1385), .B2(n1384), .ZN(n1395) );
  OR2D2BWP12T U2434 ( .A1(n1389), .A2(n1388), .Z(n1393) );
  TPNR2D2BWP12T U2435 ( .A1(n1393), .A2(n1392), .ZN(n1394) );
  ND3D2BWP12T U2436 ( .A1(n1396), .A2(n1395), .A3(n1394), .ZN(regA_out[15]) );
  NR2D2BWP12T U2437 ( .A1(n1787), .A2(n2971), .ZN(n1397) );
  AOI22D1BWP12T U2438 ( .A1(n1876), .A2(tmp1[10]), .B1(immediate1_in[10]), 
        .B2(n1804), .ZN(n1398) );
  OAI22D1BWP12T U2439 ( .A1(n3404), .A2(n1400), .B1(n2967), .B2(n3434), .ZN(
        n1404) );
  OAI22D1BWP12T U2440 ( .A1(n3406), .A2(n1401), .B1(n3001), .B2(n3444), .ZN(
        n1403) );
  OAI22D1BWP12T U2441 ( .A1(n3414), .A2(n3005), .B1(n1810), .B2(n3013), .ZN(
        n1402) );
  NR4D0BWP12T U2442 ( .A1(n1405), .A2(n1404), .A3(n1403), .A4(n1402), .ZN(
        n1411) );
  OAI22D1BWP12T U2443 ( .A1(n3416), .A2(n3023), .B1(n3393), .B2(n2963), .ZN(
        n1409) );
  INVD1BWP12T U2444 ( .I(r4[10]), .ZN(n2951) );
  OAI22D1BWP12T U2445 ( .A1(n3390), .A2(n2951), .B1(n2979), .B2(n3442), .ZN(
        n1408) );
  INVD1BWP12T U2446 ( .I(r8[10]), .ZN(n2959) );
  INVD1BWP12T U2447 ( .I(r12[10]), .ZN(n2955) );
  OAI22D1BWP12T U2448 ( .A1(n2959), .A2(n3387), .B1(n3436), .B2(n2955), .ZN(
        n1407) );
  INVD1BWP12T U2449 ( .I(r10[10]), .ZN(n2975) );
  NR4D0BWP12T U2450 ( .A1(n1409), .A2(n1408), .A3(n1407), .A4(n1406), .ZN(
        n1410) );
  INVD1BWP12T U2451 ( .I(lr[6]), .ZN(n1413) );
  INVD1BWP12T U2452 ( .I(r10[6]), .ZN(n1412) );
  TPOAI22D2BWP12T U2453 ( .A1(n3416), .A2(n1413), .B1(n1881), .B2(n1412), .ZN(
        n1415) );
  INR2D2BWP12T U2454 ( .A1(r0[6]), .B1(n3442), .ZN(n1414) );
  TPNR2D2BWP12T U2455 ( .A1(n1415), .A2(n1414), .ZN(n1421) );
  INR2D2BWP12T U2456 ( .A1(r8[6]), .B1(n3387), .ZN(n1419) );
  INVD1BWP12T U2457 ( .I(n[3574]), .ZN(n1417) );
  ND2D1BWP12T U2458 ( .A1(n1804), .A2(immediate1_in[6]), .ZN(n1416) );
  OAI21D1BWP12T U2459 ( .A1(n3446), .A2(n1417), .B(n1416), .ZN(n1418) );
  TPND2D2BWP12T U2460 ( .A1(n1421), .A2(n1420), .ZN(n1425) );
  INVD1BWP12T U2461 ( .I(r2[6]), .ZN(n2030) );
  NR2D1BWP12T U2462 ( .A1(n3432), .A2(n2030), .ZN(n1422) );
  OR2D2BWP12T U2463 ( .A1(n1423), .A2(n1422), .Z(n1424) );
  INVD1BWP12T U2464 ( .I(pc_out[6]), .ZN(n2874) );
  OR2XD1BWP12T U2465 ( .A1(n1426), .A2(n2874), .Z(n1427) );
  OAI21D1BWP12T U2466 ( .A1(n1810), .A2(n1910), .B(n1427), .ZN(n1432) );
  INVD1BWP12T U2467 ( .I(r3[6]), .ZN(n2029) );
  INVD1BWP12T U2468 ( .I(r11[6]), .ZN(n2027) );
  OAI22D1BWP12T U2469 ( .A1(n1428), .A2(n2029), .B1(n3393), .B2(n2027), .ZN(
        n1431) );
  INR2D1BWP12T U2470 ( .A1(r4[6]), .B1(n3390), .ZN(n1430) );
  INR2D1BWP12T U2471 ( .A1(r5[6]), .B1(n1837), .ZN(n1429) );
  NR4D0BWP12T U2472 ( .A1(n1432), .A2(n1431), .A3(n1430), .A4(n1429), .ZN(
        n1438) );
  ND2D1BWP12T U2473 ( .A1(n1876), .A2(tmp1[6]), .ZN(n1434) );
  ND2D1BWP12T U2474 ( .A1(n3412), .A2(r6[6]), .ZN(n1433) );
  ND2D1BWP12T U2475 ( .A1(n1434), .A2(n1433), .ZN(n1436) );
  INVD1BWP12T U2476 ( .I(r12[6]), .ZN(n2026) );
  OAI22D1BWP12T U2477 ( .A1(n2026), .A2(n3436), .B1(n3444), .B2(n1894), .ZN(
        n1435) );
  NR2D1BWP12T U2478 ( .A1(n1436), .A2(n1435), .ZN(n1437) );
  ND3D2BWP12T U2479 ( .A1(n1439), .A2(n1438), .A3(n1437), .ZN(regA_out[6]) );
  XNR2D1BWP12T U2480 ( .A1(n3301), .A2(n3299), .ZN(n1442) );
  INVD1BWP12T U2481 ( .I(pc_out[23]), .ZN(n1765) );
  TPNR2D0BWP12T U2482 ( .A1(n3343), .A2(n1765), .ZN(n1440) );
  AOI21D1BWP12T U2483 ( .A1(next_pc_in[23]), .A2(n3499), .B(n1440), .ZN(n1441)
         );
  MOAI22D1BWP12T U2484 ( .A1(n1443), .A2(n1896), .B1(n1898), .B2(n[3553]), 
        .ZN(n1452) );
  OAI22D1BWP12T U2485 ( .A1(n1587), .A2(n1445), .B1(n1444), .B2(n1895), .ZN(
        n1451) );
  NR4D0BWP12T U2486 ( .A1(n1452), .A2(n1451), .A3(n1450), .A4(n1449), .ZN(
        n1464) );
  AOI22D2BWP12T U2487 ( .A1(n1571), .A2(r8[27]), .B1(tmp1[27]), .B2(n1921), 
        .ZN(n1462) );
  NR2D1BWP12T U2488 ( .A1(n1564), .A2(n1453), .ZN(n1455) );
  AOI22D1BWP12T U2489 ( .A1(n1664), .A2(r12[27]), .B1(n1918), .B2(r4[27]), 
        .ZN(n1454) );
  AOI22D1BWP12T U2490 ( .A1(n1575), .A2(pc_out[27]), .B1(r6[27]), .B2(n1915), 
        .ZN(n1459) );
  INVD1BWP12T U2491 ( .I(r1[27]), .ZN(n1457) );
  INR3D2BWP12T U2492 ( .A1(n1462), .B1(n1461), .B2(n1460), .ZN(n1463) );
  TPND2D2BWP12T U2493 ( .A1(n1464), .A2(n1463), .ZN(regB_out[27]) );
  INVD1BWP12T U2494 ( .I(r2[12]), .ZN(n1497) );
  NR2D1BWP12T U2495 ( .A1(n1787), .A2(n1497), .ZN(n1465) );
  INVD1BWP12T U2496 ( .I(r5[12]), .ZN(n1485) );
  INVD1BWP12T U2497 ( .I(r0[12]), .ZN(n1490) );
  INVD1BWP12T U2498 ( .I(r10[12]), .ZN(n3038) );
  NR2D1BWP12T U2499 ( .A1(n1881), .A2(n3038), .ZN(n1469) );
  RCIAO21D0BWP12T U2500 ( .A1(n3442), .A2(n1490), .B(n1469), .ZN(n1470) );
  IND2XD2BWP12T U2501 ( .A1(n1471), .B1(n1470), .ZN(n1478) );
  INVD1BWP12T U2502 ( .I(lr[12]), .ZN(n3041) );
  ND2D1BWP12T U2503 ( .A1(n3418), .A2(r11[12]), .ZN(n1472) );
  OAI21D1BWP12T U2504 ( .A1(n3416), .A2(n3041), .B(n1472), .ZN(n1477) );
  AN2D1BWP12T U2505 ( .A1(n3419), .A2(r9[12]), .Z(n1475) );
  AOI22D0BWP12T U2506 ( .A1(n1473), .A2(r8[12]), .B1(r4[12]), .B2(n3450), .ZN(
        n1474) );
  TPNR3D2BWP12T U2507 ( .A1(n1478), .A2(n1477), .A3(n1476), .ZN(n1483) );
  ND2D1BWP12T U2508 ( .A1(n1862), .A2(n[3568]), .ZN(n1481) );
  INVD1BWP12T U2509 ( .I(r3[12]), .ZN(n1486) );
  NR2D1BWP12T U2510 ( .A1(n3434), .A2(n1486), .ZN(n1480) );
  INVD1BWP12T U2511 ( .I(r7[12]), .ZN(n1489) );
  ND3D2BWP12T U2512 ( .A1(n1484), .A2(n1483), .A3(n1482), .ZN(regA_out[12]) );
  INVD1BWP12T U2513 ( .I(r11[12]), .ZN(n1968) );
  OAI22D1BWP12T U2514 ( .A1(n1587), .A2(n1490), .B1(n1489), .B2(n1724), .ZN(
        n1495) );
  INVD1BWP12T U2515 ( .I(r9[12]), .ZN(n1493) );
  INR2D1BWP12T U2516 ( .A1(r10[12]), .B1(n1899), .ZN(n1491) );
  INVD1BWP12T U2517 ( .I(n1491), .ZN(n1492) );
  INVD1BWP12T U2518 ( .I(r1[12]), .ZN(n1498) );
  TPOAI22D1BWP12T U2519 ( .A1(n1659), .A2(n1498), .B1(n1519), .B2(n1497), .ZN(
        n1500) );
  NR2D1BWP12T U2520 ( .A1(n1714), .A2(n3041), .ZN(n1499) );
  RCAOI211D1BWP12T U2521 ( .A1(n1668), .A2(immediate2_in[12]), .B(n1500), .C(
        n1499), .ZN(n1505) );
  AOI22D1BWP12T U2522 ( .A1(n1575), .A2(pc_out[12]), .B1(r6[12]), .B2(n1915), 
        .ZN(n1503) );
  AOI22D0BWP12T U2523 ( .A1(n1571), .A2(r8[12]), .B1(n1526), .B2(tmp1[12]), 
        .ZN(n1502) );
  AOI22D1BWP12T U2524 ( .A1(n1664), .A2(r12[12]), .B1(n1918), .B2(r4[12]), 
        .ZN(n1501) );
  AN3XD2BWP12T U2525 ( .A1(n1503), .A2(n1502), .A3(n1501), .Z(n1504) );
  ND3XD4BWP12T U2526 ( .A1(n1506), .A2(n1505), .A3(n1504), .ZN(regB_out[12])
         );
  INVD1BWP12T U2527 ( .I(n[3579]), .ZN(n2832) );
  INVD1BWP12T U2528 ( .I(r3[1]), .ZN(n1951) );
  OAI22D1BWP12T U2529 ( .A1(n1652), .A2(n2832), .B1(n1951), .B2(n1896), .ZN(
        n1513) );
  INR2D1BWP12T U2530 ( .A1(r10[1]), .B1(n1507), .ZN(n1508) );
  INVD1BWP12T U2531 ( .I(n1508), .ZN(n1509) );
  OAI21D1BWP12T U2532 ( .A1(n1663), .A2(n2804), .B(n1509), .ZN(n1512) );
  MOAI22D0BWP12T U2533 ( .A1(n1612), .A2(n1724), .B1(n1705), .B2(r0[1]), .ZN(
        n1511) );
  NR4D1BWP12T U2534 ( .A1(n1513), .A2(n1512), .A3(n1511), .A4(n1510), .ZN(
        n1525) );
  ND2D1BWP12T U2535 ( .A1(n1915), .A2(r6[1]), .ZN(n1516) );
  ND2D1BWP12T U2536 ( .A1(n1516), .A2(n1515), .ZN(n1518) );
  MOAI22D0BWP12T U2537 ( .A1(n2831), .A2(n1714), .B1(n1713), .B2(
        immediate2_in[1]), .ZN(n1517) );
  OR2D2BWP12T U2538 ( .A1(n1518), .A2(n1517), .Z(n1523) );
  INVD1BWP12T U2539 ( .I(r2[1]), .ZN(n1950) );
  AOI22D2BWP12T U2540 ( .A1(n1664), .A2(r12[1]), .B1(n1918), .B2(r4[1]), .ZN(
        n1520) );
  ND3D2BWP12T U2541 ( .A1(n1521), .A2(n183), .A3(n1520), .ZN(n1522) );
  TPNR2D2BWP12T U2542 ( .A1(n1523), .A2(n1522), .ZN(n1524) );
  AOI22D2BWP12T U2543 ( .A1(n1571), .A2(r8[14]), .B1(tmp1[14]), .B2(n1526), 
        .ZN(n1538) );
  AOI22D2BWP12T U2544 ( .A1(n1527), .A2(r12[14]), .B1(n1918), .B2(r4[14]), 
        .ZN(n1529) );
  ND2D2BWP12T U2545 ( .A1(n1529), .A2(n1528), .ZN(n1537) );
  CKND0BWP12T U2546 ( .I(r2[14]), .ZN(n1530) );
  MOAI22D1BWP12T U2547 ( .A1(n1519), .A2(n1530), .B1(n168), .B2(r1[14]), .ZN(
        n1531) );
  INVD1BWP12T U2548 ( .I(n1531), .ZN(n1534) );
  RCAOI22D2BWP12T U2549 ( .A1(n1532), .A2(pc_out[14]), .B1(r6[14]), .B2(n1915), 
        .ZN(n1533) );
  INR3XD1BWP12T U2550 ( .A1(n1538), .B1(n1537), .B2(n1536), .ZN(n1552) );
  MOAI22D1BWP12T U2551 ( .A1(n1539), .A2(n1896), .B1(n1898), .B2(n[3566]), 
        .ZN(n1544) );
  INVD1BWP12T U2552 ( .I(r9[14]), .ZN(n1542) );
  TPNR2D1BWP12T U2553 ( .A1(n1544), .A2(n1543), .ZN(n1551) );
  INVD0BWP12T U2554 ( .I(r0[14]), .ZN(n1546) );
  INVD0BWP12T U2555 ( .I(r7[14]), .ZN(n1545) );
  OAI22D1BWP12T U2556 ( .A1(n1587), .A2(n1546), .B1(n1545), .B2(n1724), .ZN(
        n1549) );
  INVD1BWP12T U2557 ( .I(r11[14]), .ZN(n1991) );
  OAI22D1BWP12T U2558 ( .A1(n1887), .A2(n1991), .B1(n161), .B2(n1547), .ZN(
        n1548) );
  TPNR2D1BWP12T U2559 ( .A1(n1549), .A2(n1548), .ZN(n1550) );
  INVD1BWP12T U2560 ( .I(r9[25]), .ZN(n1846) );
  INVD1BWP12T U2561 ( .I(r10[25]), .ZN(n1828) );
  OAI22D1BWP12T U2562 ( .A1(n1553), .A2(n1846), .B1(n1828), .B2(n1592), .ZN(
        n1555) );
  INVD1BWP12T U2563 ( .I(r0[25]), .ZN(n1829) );
  INVD1BWP12T U2564 ( .I(r7[25]), .ZN(n1835) );
  OAI22D1BWP12T U2565 ( .A1(n1587), .A2(n1829), .B1(n1835), .B2(n1895), .ZN(
        n1554) );
  OR2XD2BWP12T U2566 ( .A1(n1555), .A2(n1554), .Z(n1559) );
  INVD1BWP12T U2567 ( .I(r11[25]), .ZN(n1827) );
  INVD1BWP12T U2568 ( .I(r5[25]), .ZN(n1836) );
  TPOAI22D1BWP12T U2569 ( .A1(n1887), .A2(n1827), .B1(n160), .B2(n1836), .ZN(
        n1557) );
  INVD1BWP12T U2570 ( .I(n[3555]), .ZN(n2549) );
  INVD1BWP12T U2571 ( .I(r3[25]), .ZN(n1847) );
  AOI22D1BWP12T U2572 ( .A1(n1921), .A2(tmp1[25]), .B1(r8[25]), .B2(n1571), 
        .ZN(n1562) );
  AOI22D1BWP12T U2573 ( .A1(n1664), .A2(r12[25]), .B1(n1918), .B2(r4[25]), 
        .ZN(n1560) );
  AN3XD2BWP12T U2574 ( .A1(n1562), .A2(n1561), .A3(n1560), .Z(n1569) );
  INVD1BWP12T U2575 ( .I(r2[25]), .ZN(n1841) );
  INVD1BWP12T U2576 ( .I(r1[25]), .ZN(n1563) );
  INVD1BWP12T U2577 ( .I(lr[25]), .ZN(n1824) );
  NR2D1BWP12T U2578 ( .A1(n1564), .A2(n1824), .ZN(n1565) );
  RCAOI211D1BWP12T U2579 ( .A1(n1567), .A2(immediate2_in[25]), .B(n1566), .C(
        n1565), .ZN(n1568) );
  AOI22D1BWP12T U2580 ( .A1(n1921), .A2(tmp1[24]), .B1(r8[24]), .B2(n1571), 
        .ZN(n1574) );
  AOI22D1BWP12T U2581 ( .A1(n1664), .A2(r12[24]), .B1(n1918), .B2(r4[24]), 
        .ZN(n1573) );
  OR2XD1BWP12T U2582 ( .A1(n1669), .A2(n2697), .Z(n1572) );
  ND3D1BWP12T U2583 ( .A1(n1574), .A2(n1573), .A3(n1572), .ZN(n1583) );
  CKND1BWP12T U2584 ( .I(r1[24]), .ZN(n1576) );
  TPOAI22D1BWP12T U2585 ( .A1(n1519), .A2(n1577), .B1(n1911), .B2(n1576), .ZN(
        n1578) );
  TPNR2D1BWP12T U2586 ( .A1(n1583), .A2(n1582), .ZN(n1598) );
  MOAI22D0BWP12T U2587 ( .A1(n1584), .A2(n1896), .B1(n1690), .B2(n[3556]), 
        .ZN(n1596) );
  OAI22D1BWP12T U2588 ( .A1(n1587), .A2(n1586), .B1(n1585), .B2(n1895), .ZN(
        n1595) );
  MOAI22D1BWP12T U2589 ( .A1(n1887), .A2(n1588), .B1(n1674), .B2(r5[24]), .ZN(
        n1594) );
  NR4D0BWP12T U2590 ( .A1(n1596), .A2(n1595), .A3(n1594), .A4(n1593), .ZN(
        n1597) );
  DCCKND4BWP12T U2591 ( .I(n1608), .ZN(n3341) );
  ND3XD1BWP12T U2592 ( .A1(n3341), .A2(n1599), .A3(n1606), .ZN(n1611) );
  CKND0BWP12T U2593 ( .I(n3324), .ZN(n1600) );
  AO21D0BWP12T U2594 ( .A1(n3331), .A2(n1600), .B(n3497), .Z(n1601) );
  AOI21D1BWP12T U2595 ( .A1(n1605), .A2(n1604), .B(n1603), .ZN(n1610) );
  NR2XD2BWP12T U2596 ( .A1(n1606), .A2(n3497), .ZN(n1607) );
  ND2XD0BWP12T U2597 ( .A1(n1608), .A2(n1607), .ZN(n1609) );
  ND3D1BWP12T U2598 ( .A1(n1611), .A2(n1610), .A3(n1609), .ZN(n2197) );
  INVD1BWP12T U2599 ( .I(pc_out[1]), .ZN(n2807) );
  INVD1BWP12T U2600 ( .I(r4[1]), .ZN(n1949) );
  INVD1BWP12T U2601 ( .I(r0[1]), .ZN(n1952) );
  OAI22D1BWP12T U2602 ( .A1(n3390), .A2(n1949), .B1(n1952), .B2(n1617), .ZN(
        n1619) );
  INVD1BWP12T U2603 ( .I(tmp1[1]), .ZN(n1620) );
  TPNR2D2BWP12T U2604 ( .A1(n1621), .A2(n1620), .ZN(n1626) );
  ND2D4BWP12T U2605 ( .A1(n3412), .A2(r6[1]), .ZN(n1625) );
  IND4D4BWP12T U2606 ( .A1(n1626), .B1(n1625), .B2(n1624), .B3(n1623), .ZN(
        n1627) );
  INVD1BWP12T U2607 ( .I(r8[1]), .ZN(n2801) );
  INVD1BWP12T U2608 ( .I(r12[1]), .ZN(n1948) );
  INVD1BWP12T U2609 ( .I(r10[1]), .ZN(n2829) );
  ND4D1BWP12T U2610 ( .A1(n1634), .A2(n1633), .A3(n1632), .A4(n1631), .ZN(
        regA_out[1]) );
  INVD1BWP12T U2611 ( .I(tmp1[29]), .ZN(n1635) );
  OAI22D1BWP12T U2612 ( .A1(n3378), .A2(n1635), .B1(n3540), .B2(n3432), .ZN(
        n1639) );
  OAI22D1BWP12T U2613 ( .A1(n3414), .A2(n1637), .B1(n1636), .B2(n3444), .ZN(
        n1638) );
  AOI211D1BWP12T U2614 ( .A1(r1[29]), .A2(n3384), .B(n1639), .C(n1638), .ZN(
        n1651) );
  OAI22D1BWP12T U2615 ( .A1(n3390), .A2(n3543), .B1(n3542), .B2(n3435), .ZN(
        n1643) );
  OAI22D1BWP12T U2616 ( .A1(n3393), .A2(n3545), .B1(n3544), .B2(n3452), .ZN(
        n1642) );
  INVD1BWP12T U2617 ( .I(r6[29]), .ZN(n1640) );
  OAI22D1BWP12T U2618 ( .A1(n3396), .A2(n1640), .B1(n3442), .B2(n3546), .ZN(
        n1641) );
  NR4D0BWP12T U2619 ( .A1(n1644), .A2(n1643), .A3(n1642), .A4(n1641), .ZN(
        n1650) );
  AOI22D1BWP12T U2620 ( .A1(n1862), .A2(n[3551]), .B1(n1645), .B2(r9[29]), 
        .ZN(n1648) );
  AOI22D0BWP12T U2621 ( .A1(n1646), .A2(r3[29]), .B1(pc_out[29]), .B2(n3445), 
        .ZN(n1647) );
  AN2XD2BWP12T U2622 ( .A1(n1648), .A2(n1647), .Z(n1649) );
  ND3D2BWP12T U2623 ( .A1(n1651), .A2(n1650), .A3(n1649), .ZN(regA_out[29]) );
  OAI22D1BWP12T U2624 ( .A1(n1652), .A2(n2856), .B1(n2002), .B2(n1896), .ZN(
        n1657) );
  OR2XD1BWP12T U2625 ( .A1(n1654), .A2(n1653), .Z(n1655) );
  TPNR2D2BWP12T U2626 ( .A1(n1657), .A2(n1656), .ZN(n1689) );
  INR2D4BWP12T U2627 ( .A1(r10[2]), .B1(n1899), .ZN(n1661) );
  DCCKND4BWP12T U2628 ( .I(n1661), .ZN(n1662) );
  TPOAI21D4BWP12T U2629 ( .A1(n1663), .A2(n2855), .B(n1662), .ZN(n1667) );
  IOA21D2BWP12T U2630 ( .A1(n1892), .A2(r0[2]), .B(n1665), .ZN(n1666) );
  NR3XD4BWP12T U2631 ( .A1(n1660), .A2(n1666), .A3(n1667), .ZN(n1688) );
  INVD1BWP12T U2632 ( .I(n1671), .ZN(n1687) );
  INVD1BWP12T U2633 ( .I(r8[2]), .ZN(n1673) );
  TPOAI22D2BWP12T U2634 ( .A1(n1922), .A2(n1673), .B1(n1895), .B2(n1672), .ZN(
        n1685) );
  ND2D1BWP12T U2635 ( .A1(n1674), .A2(r5[2]), .ZN(n1678) );
  INR2D1BWP12T U2636 ( .A1(r11[2]), .B1(n1675), .ZN(n1676) );
  TPND2D2BWP12T U2637 ( .A1(n1678), .A2(n1677), .ZN(n1684) );
  ND2D3BWP12T U2638 ( .A1(n1918), .A2(r4[2]), .ZN(n1682) );
  INR2D4BWP12T U2639 ( .A1(pc_out[2]), .B1(n1703), .ZN(n1680) );
  CKND3BWP12T U2640 ( .I(n1680), .ZN(n1681) );
  ND2XD4BWP12T U2641 ( .A1(n1682), .A2(n1681), .ZN(n1683) );
  NR3XD4BWP12T U2642 ( .A1(n1685), .A2(n1684), .A3(n1683), .ZN(n1686) );
  ND4D4BWP12T U2643 ( .A1(n1689), .A2(n1688), .A3(n1687), .A4(n1686), .ZN(
        regB_out[2]) );
  AOI22D1BWP12T U2644 ( .A1(n1691), .A2(r9[7]), .B1(n1690), .B2(n[3573]), .ZN(
        n1722) );
  ND2D1BWP12T U2645 ( .A1(n1692), .A2(tmp1[7]), .ZN(n1695) );
  INR2D4BWP12T U2646 ( .A1(r5[7]), .B1(n1889), .ZN(n1694) );
  INR2D4BWP12T U2647 ( .A1(n1695), .B1(n1694), .ZN(n1702) );
  IND3D1BWP12T U2648 ( .A1(n1698), .B1(n1697), .B2(n1696), .ZN(n1699) );
  INR2D4BWP12T U2649 ( .A1(r8[7]), .B1(n1922), .ZN(n1700) );
  TPND2D2BWP12T U2650 ( .A1(n1702), .A2(n1701), .ZN(n1721) );
  INR2D2BWP12T U2651 ( .A1(pc_out[7]), .B1(n1703), .ZN(n1709) );
  TPND2D1BWP12T U2652 ( .A1(n1705), .A2(r0[7]), .ZN(n1706) );
  INVD1P75BWP12T U2653 ( .I(n1706), .ZN(n1707) );
  TPNR3D2BWP12T U2654 ( .A1(n1709), .A2(n1708), .A3(n1707), .ZN(n1719) );
  INR2D4BWP12T U2655 ( .A1(r2[7]), .B1(n1519), .ZN(n1712) );
  TPNR2D2BWP12T U2656 ( .A1(n1712), .A2(n1711), .ZN(n1718) );
  INR2D4BWP12T U2657 ( .A1(lr[7]), .B1(n1714), .ZN(n1715) );
  INR2D2BWP12T U2658 ( .A1(n1716), .B1(n1715), .ZN(n1717) );
  ND3D2BWP12T U2659 ( .A1(n1719), .A2(n1718), .A3(n1717), .ZN(n1720) );
  INR3D2BWP12T U2660 ( .A1(n1722), .B1(n1721), .B2(n1720), .ZN(n1734) );
  NR2XD2BWP12T U2661 ( .A1(n1724), .A2(n1723), .ZN(n1725) );
  INVD1P75BWP12T U2662 ( .I(n1725), .ZN(n1732) );
  MOAI22D1BWP12T U2663 ( .A1(n1920), .A2(n2846), .B1(n1726), .B2(r11[7]), .ZN(
        n1731) );
  INVD2BWP12T U2664 ( .I(n1918), .ZN(n1729) );
  INR2D4BWP12T U2665 ( .A1(r10[7]), .B1(n1899), .ZN(n1727) );
  INVD1P75BWP12T U2666 ( .I(n1727), .ZN(n1728) );
  RCOAI21D2BWP12T U2667 ( .A1(n1729), .A2(n2865), .B(n1728), .ZN(n1730) );
  INR3D2BWP12T U2668 ( .A1(n1732), .B1(n1731), .B2(n1730), .ZN(n1733) );
  ND2XD3BWP12T U2669 ( .A1(n1734), .A2(n1733), .ZN(regB_out[7]) );
  TPND2D2BWP12T U2670 ( .A1(n3503), .A2(n3502), .ZN(n1742) );
  INR2D0BWP12T U2671 ( .A1(write2_in[21]), .B1(n530), .ZN(n1735) );
  AOI21D1BWP12T U2672 ( .A1(write1_in[21]), .A2(n530), .B(n1735), .ZN(n3289)
         );
  INVD0BWP12T U2673 ( .I(write2_in[20]), .ZN(n1736) );
  TPNR2D0BWP12T U2674 ( .A1(n530), .A2(n1736), .ZN(n1737) );
  NR2D1BWP12T U2675 ( .A1(n3506), .A2(n3497), .ZN(n1738) );
  CKND2D1BWP12T U2676 ( .A1(n3506), .A2(n3505), .ZN(n1741) );
  OA21D1BWP12T U2677 ( .A1(n3289), .A2(n1741), .B(n1740), .Z(n1745) );
  NR2D1BWP12T U2678 ( .A1(n3289), .A2(n3497), .ZN(n1743) );
  ND2D1BWP12T U2679 ( .A1(n1743), .A2(n1742), .ZN(n1744) );
  INVD1BWP12T U2680 ( .I(r12[23]), .ZN(n1747) );
  INVD1BWP12T U2681 ( .I(r4[23]), .ZN(n1749) );
  INVD1BWP12T U2682 ( .I(r8[23]), .ZN(n1748) );
  OAI22D1BWP12T U2683 ( .A1(n3390), .A2(n1749), .B1(n1748), .B2(n3435), .ZN(
        n1755) );
  INVD1BWP12T U2684 ( .I(r6[23]), .ZN(n1752) );
  NR4D0BWP12T U2685 ( .A1(n1756), .A2(n1755), .A3(n1754), .A4(n1753), .ZN(
        n1770) );
  INVD1BWP12T U2686 ( .I(tmp1[23]), .ZN(n1758) );
  OAI22D2BWP12T U2687 ( .A1(n3378), .A2(n1758), .B1(n1757), .B2(n3432), .ZN(
        n1761) );
  MOAI22D1BWP12T U2688 ( .A1(n3381), .A2(n1759), .B1(r7[23]), .B2(n1839), .ZN(
        n1760) );
  RCAOI211D1BWP12T U2689 ( .A1(r1[23]), .A2(n3384), .B(n1761), .C(n1760), .ZN(
        n1769) );
  INVD1BWP12T U2690 ( .I(n[3557]), .ZN(n1763) );
  OAI22D1BWP12T U2691 ( .A1(n3404), .A2(n1763), .B1(n3402), .B2(n1762), .ZN(
        n1767) );
  OAI22D1BWP12T U2692 ( .A1(n3406), .A2(n1765), .B1(n1764), .B2(n3434), .ZN(
        n1766) );
  NR2D1BWP12T U2693 ( .A1(n1767), .A2(n1766), .ZN(n1768) );
  ND3D2BWP12T U2694 ( .A1(n1770), .A2(n1769), .A3(n1768), .ZN(regA_out[23]) );
  INR2D1BWP12T U2695 ( .A1(r10[21]), .B1(n1881), .ZN(n1773) );
  NR2D1BWP12T U2696 ( .A1(n3434), .A2(n1771), .ZN(n1772) );
  NR2D2BWP12T U2697 ( .A1(n1773), .A2(n1772), .ZN(n1775) );
  ND2D1BWP12T U2698 ( .A1(n1876), .A2(tmp1[21]), .ZN(n1774) );
  TPND2D2BWP12T U2699 ( .A1(n1775), .A2(n1774), .ZN(n1784) );
  INVD1BWP12T U2700 ( .I(n3412), .ZN(n3363) );
  INVD1BWP12T U2701 ( .I(r6[21]), .ZN(n1776) );
  MOAI22D1BWP12T U2702 ( .A1(n3363), .A2(n1776), .B1(n621), .B2(r12[21]), .ZN(
        n1783) );
  ND2D3BWP12T U2703 ( .A1(n3384), .A2(r1[21]), .ZN(n1781) );
  OR2XD1BWP12T U2704 ( .A1(n1778), .A2(n1777), .Z(n1780) );
  ND2D3BWP12T U2705 ( .A1(n3418), .A2(r11[21]), .ZN(n1779) );
  ND3XD3BWP12T U2706 ( .A1(n1781), .A2(n1780), .A3(n1779), .ZN(n1782) );
  TPNR3D2BWP12T U2707 ( .A1(n1784), .A2(n1783), .A3(n1782), .ZN(n1802) );
  ND2D1BWP12T U2708 ( .A1(n3419), .A2(r9[21]), .ZN(n1785) );
  OAI21D1BWP12T U2709 ( .A1(n3404), .A2(n1786), .B(n1785), .ZN(n1793) );
  INR2D2BWP12T U2710 ( .A1(r2[21]), .B1(n1787), .ZN(n1790) );
  TPND2D2BWP12T U2711 ( .A1(n1788), .A2(pc_out[21]), .ZN(n1789) );
  IND2D4BWP12T U2712 ( .A1(n1790), .B1(n1789), .ZN(n1791) );
  OAI22D1BWP12T U2713 ( .A1(n3381), .A2(n1795), .B1(n3444), .B2(n1794), .ZN(
        n1799) );
  INR2D1BWP12T U2714 ( .A1(r8[21]), .B1(n3435), .ZN(n1797) );
  ND3D2BWP12T U2715 ( .A1(n1802), .A2(n1801), .A3(n1800), .ZN(regA_out[21]) );
  TPNR2D3BWP12T U2716 ( .A1(n3432), .A2(n1960), .ZN(n1803) );
  TPAOI21D2BWP12T U2717 ( .A1(n3412), .A2(r6[3]), .B(n1803), .ZN(n1806) );
  AOI22D1BWP12T U2718 ( .A1(n1876), .A2(tmp1[3]), .B1(n1804), .B2(
        immediate1_in[3]), .ZN(n1805) );
  TPND2D2BWP12T U2719 ( .A1(n1806), .A2(n1805), .ZN(n1815) );
  OAI22D1BWP12T U2720 ( .A1(n3446), .A2(n2853), .B1(n1958), .B2(n3434), .ZN(
        n1814) );
  INVD1BWP12T U2721 ( .I(pc_out[3]), .ZN(n1808) );
  OAI22D1BWP12T U2722 ( .A1(n3406), .A2(n1808), .B1(n1807), .B2(n3444), .ZN(
        n1813) );
  OAI22D1BWP12T U2723 ( .A1(n3414), .A2(n1811), .B1(n1810), .B2(n1809), .ZN(
        n1812) );
  NR4D0BWP12T U2724 ( .A1(n1815), .A2(n1814), .A3(n1813), .A4(n1812), .ZN(
        n1822) );
  OAI22D1BWP12T U2725 ( .A1(n3416), .A2(n2851), .B1(n3393), .B2(n2852), .ZN(
        n1820) );
  INVD1BWP12T U2726 ( .I(r4[3]), .ZN(n1957) );
  INVD1BWP12T U2727 ( .I(r8[3]), .ZN(n1955) );
  INVD1BWP12T U2728 ( .I(r12[3]), .ZN(n2850) );
  OAI22D1BWP12T U2729 ( .A1(n1955), .A2(n3387), .B1(n3436), .B2(n2850), .ZN(
        n1818) );
  INVD1BWP12T U2730 ( .I(r10[3]), .ZN(n1959) );
  NR4D0BWP12T U2731 ( .A1(n1820), .A2(n1819), .A3(n1818), .A4(n1817), .ZN(
        n1821) );
  TPND2D1BWP12T U2732 ( .A1(n1822), .A2(n1821), .ZN(regA_out[3]) );
  INVD1BWP12T U2733 ( .I(r12[25]), .ZN(n1823) );
  INVD1BWP12T U2734 ( .I(r4[25]), .ZN(n1826) );
  INVD1BWP12T U2735 ( .I(r8[25]), .ZN(n1825) );
  OAI22D1BWP12T U2736 ( .A1(n3390), .A2(n1826), .B1(n3435), .B2(n1825), .ZN(
        n1833) );
  INVD1BWP12T U2737 ( .I(r6[25]), .ZN(n1830) );
  NR4D0BWP12T U2738 ( .A1(n1834), .A2(n1833), .A3(n1832), .A4(n1831), .ZN(
        n1852) );
  INVD1BWP12T U2739 ( .I(tmp1[25]), .ZN(n1840) );
  OAI22D1BWP12T U2740 ( .A1(n3432), .A2(n1841), .B1(n3378), .B2(n1840), .ZN(
        n1844) );
  INR3XD1BWP12T U2741 ( .A1(n1845), .B1(n1844), .B2(n1843), .ZN(n1851) );
  OAI22D1BWP12T U2742 ( .A1(n3404), .A2(n2549), .B1(n3402), .B2(n1846), .ZN(
        n1849) );
  OAI22D1BWP12T U2743 ( .A1(n3406), .A2(n3536), .B1(n1847), .B2(n3434), .ZN(
        n1848) );
  NR2D1BWP12T U2744 ( .A1(n1849), .A2(n1848), .ZN(n1850) );
  TPND3D1BWP12T U2745 ( .A1(n1852), .A2(n1851), .A3(n1850), .ZN(regA_out[25])
         );
  INR2D1BWP12T U2746 ( .A1(r3[20]), .B1(n3434), .ZN(n1858) );
  ND2D1BWP12T U2747 ( .A1(n1853), .A2(r4[20]), .ZN(n1857) );
  INVD1BWP12T U2748 ( .I(r8[20]), .ZN(n2709) );
  NR2D1BWP12T U2749 ( .A1(n3435), .A2(n2709), .ZN(n1855) );
  IND3D1BWP12T U2750 ( .A1(n1858), .B1(n1857), .B2(n1856), .ZN(n1868) );
  INVD1BWP12T U2751 ( .I(r12[20]), .ZN(n1861) );
  ND2D1BWP12T U2752 ( .A1(n1859), .A2(lr[20]), .ZN(n1860) );
  OAI21D1BWP12T U2753 ( .A1(n3436), .A2(n1861), .B(n1860), .ZN(n1867) );
  ND2D1BWP12T U2754 ( .A1(n3445), .A2(pc_out[20]), .ZN(n1865) );
  ND2D1BWP12T U2755 ( .A1(n3419), .A2(r9[20]), .ZN(n1864) );
  ND2D1BWP12T U2756 ( .A1(n1862), .A2(n[3560]), .ZN(n1863) );
  ND3D1BWP12T U2757 ( .A1(n1865), .A2(n1864), .A3(n1863), .ZN(n1866) );
  TPNR2D1BWP12T U2758 ( .A1(n3442), .A2(n1869), .ZN(n1872) );
  INVD1BWP12T U2759 ( .I(r6[20]), .ZN(n1870) );
  TPNR2D3BWP12T U2760 ( .A1(n3396), .A2(n1870), .ZN(n1871) );
  AOI22D1BWP12T U2761 ( .A1(n3417), .A2(r1[20]), .B1(n1873), .B2(r5[20]), .ZN(
        n1874) );
  ND2D1BWP12T U2762 ( .A1(n1875), .A2(n1874), .ZN(n1884) );
  INR2D1BWP12T U2763 ( .A1(r2[20]), .B1(n3432), .ZN(n1878) );
  ND2D1BWP12T U2764 ( .A1(n1876), .A2(tmp1[20]), .ZN(n1877) );
  IND2XD1BWP12T U2765 ( .A1(n1878), .B1(n1877), .ZN(n1883) );
  OAI21D1BWP12T U2766 ( .A1(n1881), .A2(n1880), .B(n1879), .ZN(n1882) );
  NR3D1BWP12T U2767 ( .A1(n1884), .A2(n1883), .A3(n1882), .ZN(n1885) );
  NR2D2BWP12T U2768 ( .A1(n161), .A2(n1888), .ZN(n1890) );
  ND2D1BWP12T U2769 ( .A1(n1892), .A2(r0[6]), .ZN(n1893) );
  OAI21D1BWP12T U2770 ( .A1(n1895), .A2(n1894), .B(n1893), .ZN(n1905) );
  NR2D1BWP12T U2771 ( .A1(n1896), .A2(n2029), .ZN(n1897) );
  AOI21D2BWP12T U2772 ( .A1(n1898), .A2(n[3574]), .B(n1897), .ZN(n1903) );
  INR2D1BWP12T U2773 ( .A1(r10[6]), .B1(n1899), .ZN(n1901) );
  TPNR2D2BWP12T U2774 ( .A1(n1901), .A2(n189), .ZN(n1902) );
  CKND2D2BWP12T U2775 ( .A1(n1903), .A2(n1902), .ZN(n1904) );
  IOA21D2BWP12T U2776 ( .A1(n164), .A2(lr[6]), .B(n1908), .ZN(n1914) );
  NR2D1BWP12T U2777 ( .A1(n1519), .A2(n2030), .ZN(n1913) );
  TPNR3D2BWP12T U2778 ( .A1(n1914), .A2(n1913), .A3(n1912), .ZN(n1930) );
  ND2D1BWP12T U2779 ( .A1(n1915), .A2(r6[6]), .ZN(n1916) );
  OAI21D1BWP12T U2780 ( .A1(n1920), .A2(n2026), .B(n1919), .ZN(n1927) );
  TPND2D2BWP12T U2781 ( .A1(n1921), .A2(tmp1[6]), .ZN(n1925) );
  INVD1BWP12T U2782 ( .I(r8[6]), .ZN(n2024) );
  INR2D2BWP12T U2783 ( .A1(r8[6]), .B1(n1922), .ZN(n1923) );
  INVD1P75BWP12T U2784 ( .I(n1923), .ZN(n1924) );
  TPND2D1BWP12T U2785 ( .A1(n1925), .A2(n1924), .ZN(n1926) );
  TPNR3D2BWP12T U2786 ( .A1(n1928), .A2(n1927), .A3(n1926), .ZN(n1929) );
  ND3XD3BWP12T U2787 ( .A1(n1931), .A2(n1930), .A3(n1929), .ZN(regB_out[6]) );
  CKND3BWP12T U2788 ( .I(n3059), .ZN(n1932) );
  INR2D4BWP12T U2789 ( .A1(n1933), .B1(n1932), .ZN(n3092) );
  CKND2D1BWP12T U2790 ( .A1(write1_in[14]), .A2(n530), .ZN(n1936) );
  CKND2D0BWP12T U2791 ( .A1(n3331), .A2(write2_in[14]), .ZN(n1935) );
  CKND2D2BWP12T U2792 ( .A1(n3111), .A2(n3107), .ZN(n1937) );
  ND2D1BWP12T U2793 ( .A1(write1_in[15]), .A2(n530), .ZN(n1939) );
  CKND2D0BWP12T U2794 ( .A1(n3331), .A2(write2_in[15]), .ZN(n1938) );
  ND2D1BWP12T U2795 ( .A1(n1939), .A2(n1938), .ZN(n3136) );
  INVD1BWP12T U2796 ( .I(n157), .ZN(n1940) );
  AN2XD2BWP12T U2797 ( .A1(n3136), .A2(n1940), .Z(n1941) );
  TPND2D2BWP12T U2798 ( .A1(n3137), .A2(n1941), .ZN(n3251) );
  TPNR2D2BWP12T U2799 ( .A1(n3251), .A2(n163), .ZN(n1943) );
  AOI22D1BWP12T U2800 ( .A1(next_pc_in[18]), .A2(n3499), .B1(n3498), .B2(
        pc_out[18]), .ZN(n1944) );
  AO222D0BWP12T U2801 ( .A1(n3246), .A2(write1_in[7]), .B1(n1947), .B2(
        write2_in[7]), .C1(n1946), .C2(tmp1[7]), .Z(n2143) );
  AO222D0BWP12T U2802 ( .A1(n3246), .A2(write1_in[2]), .B1(n1947), .B2(
        write2_in[2]), .C1(n1946), .C2(tmp1[2]), .Z(n2138) );
  AN2XD2BWP12T U2803 ( .A1(next_cpsr_in[2]), .A2(n3532), .Z(cpsrin[2]) );
  OAI222D1BWP12T U2804 ( .A1(n1954), .A2(n2958), .B1(n1953), .B2(n2957), .C1(
        n2956), .C2(n1948), .ZN(n2233) );
  OAI222D1BWP12T U2805 ( .A1(n1954), .A2(n2954), .B1(n1953), .B2(n2953), .C1(
        n2952), .C2(n1949), .ZN(n2489) );
  OAI222D1BWP12T U2806 ( .A1(n1954), .A2(n2962), .B1(n1953), .B2(n2961), .C1(
        n2960), .C2(n2801), .ZN(n2361) );
  OAI222D1BWP12T U2807 ( .A1(n1954), .A2(n2966), .B1(n1953), .B2(n2965), .C1(
        n2964), .C2(n2802), .ZN(n2265) );
  OAI222D1BWP12T U2808 ( .A1(n1954), .A2(n2978), .B1(n1953), .B2(n2977), .C1(
        n2976), .C2(n2829), .ZN(n2297) );
  OAI222D1BWP12T U2809 ( .A1(n1954), .A2(n2974), .B1(n1953), .B2(n2973), .C1(
        n2972), .C2(n1950), .ZN(n2553) );
  OAI222D1BWP12T U2810 ( .A1(n1954), .A2(n2970), .B1(n1953), .B2(n2969), .C1(
        n2968), .C2(n1951), .ZN(n2521) );
  OAI222D1BWP12T U2811 ( .A1(n1954), .A2(n2982), .B1(n1953), .B2(n2981), .C1(
        n2980), .C2(n1952), .ZN(n2617) );
  OAI222D1BWP12T U2812 ( .A1(n1962), .A2(n2962), .B1(n1961), .B2(n2961), .C1(
        n2960), .C2(n1955), .ZN(n2363) );
  OAI222D1BWP12T U2813 ( .A1(n1962), .A2(n2982), .B1(n1961), .B2(n2981), .C1(
        n2980), .C2(n1956), .ZN(n2619) );
  OAI222D1BWP12T U2814 ( .A1(n1962), .A2(n2966), .B1(n1961), .B2(n2965), .C1(
        n2964), .C2(n2852), .ZN(n2267) );
  OAI222D1BWP12T U2815 ( .A1(n1962), .A2(n2958), .B1(n1961), .B2(n2957), .C1(
        n2956), .C2(n2850), .ZN(n2235) );
  OAI222D1BWP12T U2816 ( .A1(n1962), .A2(n2954), .B1(n1961), .B2(n2953), .C1(
        n2952), .C2(n1957), .ZN(n2491) );
  OAI222D1BWP12T U2817 ( .A1(n1962), .A2(n2970), .B1(n1961), .B2(n2969), .C1(
        n2968), .C2(n1958), .ZN(n2523) );
  OAI222D1BWP12T U2818 ( .A1(n1962), .A2(n2978), .B1(n1961), .B2(n2977), .C1(
        n2976), .C2(n1959), .ZN(n2299) );
  OAI222D1BWP12T U2819 ( .A1(n1962), .A2(n2974), .B1(n1961), .B2(n2973), .C1(
        n2972), .C2(n1960), .ZN(n2555) );
  AOI22D0BWP12T U2820 ( .A1(n[3568]), .A2(n3464), .B1(n3480), .B2(pc_out[12]), 
        .ZN(n1973) );
  AOI22D0BWP12T U2821 ( .A1(n3479), .A2(r12[12]), .B1(r9[12]), .B2(n3475), 
        .ZN(n1972) );
  AOI22D0BWP12T U2822 ( .A1(r5[12]), .A2(n3481), .B1(n2770), .B2(r6[12]), .ZN(
        n1966) );
  AOI22D0BWP12T U2823 ( .A1(r7[12]), .A2(n3482), .B1(n2757), .B2(r4[12]), .ZN(
        n1965) );
  AOI22D0BWP12T U2824 ( .A1(r1[12]), .A2(n3484), .B1(n3483), .B2(r2[12]), .ZN(
        n1964) );
  AOI22D0BWP12T U2825 ( .A1(r0[12]), .A2(n3486), .B1(n3485), .B2(r3[12]), .ZN(
        n1963) );
  ND4D1BWP12T U2826 ( .A1(n1966), .A2(n1965), .A3(n1964), .A4(n1963), .ZN(
        n1967) );
  AOI22D0BWP12T U2827 ( .A1(r8[12]), .A2(n3493), .B1(n1967), .B2(n3492), .ZN(
        n1971) );
  OAI22D0BWP12T U2828 ( .A1(n2779), .A2(n3041), .B1(n1968), .B2(n2803), .ZN(
        n1969) );
  AOI21D0BWP12T U2829 ( .A1(r10[12]), .A2(n2810), .B(n1969), .ZN(n1970) );
  ND4D1BWP12T U2830 ( .A1(n1973), .A2(n1972), .A3(n1971), .A4(n1970), .ZN(
        regC_out[12]) );
  OAI22D0BWP12T U2831 ( .A1(n3478), .A2(n1975), .B1(n2779), .B2(n1974), .ZN(
        n1976) );
  AOI21D0BWP12T U2832 ( .A1(n[3557]), .A2(n3464), .B(n1976), .ZN(n1985) );
  AOI22D0BWP12T U2833 ( .A1(r5[23]), .A2(n3481), .B1(n2770), .B2(r6[23]), .ZN(
        n1980) );
  AOI22D0BWP12T U2834 ( .A1(r7[23]), .A2(n3482), .B1(n2757), .B2(r4[23]), .ZN(
        n1979) );
  AOI22D0BWP12T U2835 ( .A1(r1[23]), .A2(n3484), .B1(n3483), .B2(r2[23]), .ZN(
        n1978) );
  AOI22D0BWP12T U2836 ( .A1(r0[23]), .A2(n3486), .B1(n3485), .B2(r3[23]), .ZN(
        n1977) );
  ND4D1BWP12T U2837 ( .A1(n1980), .A2(n1979), .A3(n1978), .A4(n1977), .ZN(
        n1981) );
  AOI22D0BWP12T U2838 ( .A1(r8[23]), .A2(n3493), .B1(n1981), .B2(n3492), .ZN(
        n1984) );
  AOI22D0BWP12T U2839 ( .A1(r11[23]), .A2(n2704), .B1(n3475), .B2(r9[23]), 
        .ZN(n1983) );
  AOI22D0BWP12T U2840 ( .A1(pc_out[23]), .A2(n3480), .B1(n3479), .B2(r12[23]), 
        .ZN(n1982) );
  ND4D1BWP12T U2841 ( .A1(n1985), .A2(n1984), .A3(n1983), .A4(n1982), .ZN(
        regC_out[23]) );
  AOI22D0BWP12T U2842 ( .A1(n[3566]), .A2(n3464), .B1(n3480), .B2(pc_out[14]), 
        .ZN(n1997) );
  AOI22D0BWP12T U2843 ( .A1(n3479), .A2(r12[14]), .B1(r9[14]), .B2(n3475), 
        .ZN(n1996) );
  AOI22D0BWP12T U2844 ( .A1(r5[14]), .A2(n3481), .B1(n2770), .B2(r6[14]), .ZN(
        n1989) );
  AOI22D0BWP12T U2845 ( .A1(r7[14]), .A2(n3482), .B1(n2757), .B2(r4[14]), .ZN(
        n1988) );
  AOI22D0BWP12T U2846 ( .A1(r1[14]), .A2(n3484), .B1(n3483), .B2(r2[14]), .ZN(
        n1987) );
  AOI22D0BWP12T U2847 ( .A1(r0[14]), .A2(n3486), .B1(n3485), .B2(r3[14]), .ZN(
        n1986) );
  ND4D1BWP12T U2848 ( .A1(n1989), .A2(n1988), .A3(n1987), .A4(n1986), .ZN(
        n1990) );
  AOI22D0BWP12T U2849 ( .A1(r8[14]), .A2(n3493), .B1(n1990), .B2(n3492), .ZN(
        n1995) );
  OAI22D0BWP12T U2850 ( .A1(n2779), .A2(n1992), .B1(n1991), .B2(n2803), .ZN(
        n1993) );
  AOI21D0BWP12T U2851 ( .A1(r10[14]), .A2(n2810), .B(n1993), .ZN(n1994) );
  ND4D1BWP12T U2852 ( .A1(n1997), .A2(n1996), .A3(n1995), .A4(n1994), .ZN(
        regC_out[14]) );
  OAI222D1BWP12T U2853 ( .A1(n2004), .A2(n2982), .B1(n2003), .B2(n2981), .C1(
        n2980), .C2(n1998), .ZN(n2618) );
  OAI222D1BWP12T U2854 ( .A1(n2004), .A2(n2966), .B1(n2003), .B2(n2965), .C1(
        n2964), .C2(n2755), .ZN(n2266) );
  OAI222D1BWP12T U2855 ( .A1(n2004), .A2(n2974), .B1(n2003), .B2(n2973), .C1(
        n2972), .C2(n1999), .ZN(n2554) );
  OAI222D1BWP12T U2856 ( .A1(n2004), .A2(n2958), .B1(n2003), .B2(n2957), .C1(
        n2956), .C2(n2000), .ZN(n2234) );
  OAI222D1BWP12T U2857 ( .A1(n2004), .A2(n2978), .B1(n2003), .B2(n2977), .C1(
        n2976), .C2(n2854), .ZN(n2298) );
  OAI222D1BWP12T U2858 ( .A1(n2004), .A2(n2954), .B1(n2003), .B2(n2953), .C1(
        n2952), .C2(n2001), .ZN(n2490) );
  OAI222D1BWP12T U2859 ( .A1(n2004), .A2(n2962), .B1(n2003), .B2(n2961), .C1(
        n2960), .C2(n1673), .ZN(n2362) );
  OAI222D1BWP12T U2860 ( .A1(n2004), .A2(n2970), .B1(n2003), .B2(n2969), .C1(
        n2968), .C2(n2002), .ZN(n2522) );
  TPAOI21D0BWP12T U2861 ( .A1(n3185), .A2(write2_in[6]), .B(reset), .ZN(n2006)
         );
  TPND2D0BWP12T U2862 ( .A1(n3186), .A2(n[3574]), .ZN(n2005) );
  OAI211D1BWP12T U2863 ( .A1(n2872), .A2(n2031), .B(n2006), .C(n2005), .ZN(
        spin[6]) );
  OAI222D1BWP12T U2864 ( .A1(n2015), .A2(n2982), .B1(n2014), .B2(n2981), .C1(
        n2980), .C2(n2007), .ZN(n2620) );
  OAI222D1BWP12T U2865 ( .A1(n2015), .A2(n2962), .B1(n2014), .B2(n2961), .C1(
        n2960), .C2(n2008), .ZN(n2364) );
  OAI222D1BWP12T U2866 ( .A1(n2015), .A2(n2958), .B1(n2014), .B2(n2957), .C1(
        n2956), .C2(n2009), .ZN(n2236) );
  OAI222D1BWP12T U2867 ( .A1(n2015), .A2(n2954), .B1(n2014), .B2(n2953), .C1(
        n2952), .C2(n2010), .ZN(n2492) );
  OAI222D1BWP12T U2868 ( .A1(n2015), .A2(n2966), .B1(n2014), .B2(n2965), .C1(
        n2964), .C2(n2011), .ZN(n2268) );
  OAI222D1BWP12T U2869 ( .A1(n2015), .A2(n2974), .B1(n2014), .B2(n2973), .C1(
        n2972), .C2(n2012), .ZN(n2556) );
  OAI222D1BWP12T U2870 ( .A1(n2015), .A2(n2970), .B1(n2014), .B2(n2969), .C1(
        n2968), .C2(n2013), .ZN(n2524) );
  OAI222D1BWP12T U2871 ( .A1(n2015), .A2(n2978), .B1(n2014), .B2(n2977), .C1(
        n2976), .C2(n2841), .ZN(n2300) );
  CKND0BWP12T U2872 ( .I(r0[5]), .ZN(n2016) );
  OAI222D1BWP12T U2873 ( .A1(n2023), .A2(n2982), .B1(n2022), .B2(n2981), .C1(
        n2980), .C2(n2016), .ZN(n2621) );
  INVD0BWP12T U2874 ( .I(r4[5]), .ZN(n2017) );
  OAI222D1BWP12T U2875 ( .A1(n2023), .A2(n2954), .B1(n2022), .B2(n2953), .C1(
        n2952), .C2(n2017), .ZN(n2493) );
  OAI222D1BWP12T U2876 ( .A1(n2023), .A2(n2958), .B1(n2022), .B2(n2957), .C1(
        n2956), .C2(n2018), .ZN(n2237) );
  OAI222D1BWP12T U2877 ( .A1(n2023), .A2(n2962), .B1(n2022), .B2(n2961), .C1(
        n2960), .C2(n2019), .ZN(n2365) );
  OAI222D1BWP12T U2878 ( .A1(n2023), .A2(n2966), .B1(n2022), .B2(n2965), .C1(
        n2964), .C2(n2869), .ZN(n2269) );
  OAI222D1BWP12T U2879 ( .A1(n2023), .A2(n2978), .B1(n2022), .B2(n2977), .C1(
        n2976), .C2(n2868), .ZN(n2301) );
  OAI222D1BWP12T U2880 ( .A1(n2023), .A2(n2970), .B1(n2022), .B2(n2969), .C1(
        n2968), .C2(n2020), .ZN(n2525) );
  OAI222D1BWP12T U2881 ( .A1(n2023), .A2(n2974), .B1(n2022), .B2(n2973), .C1(
        n2972), .C2(n2021), .ZN(n2557) );
  OAI222D1BWP12T U2882 ( .A1(n2032), .A2(n2962), .B1(n2031), .B2(n2961), .C1(
        n2960), .C2(n2024), .ZN(n2366) );
  INVD0BWP12T U2883 ( .I(r0[6]), .ZN(n2025) );
  OAI222D1BWP12T U2884 ( .A1(n2032), .A2(n2982), .B1(n2031), .B2(n2981), .C1(
        n2980), .C2(n2025), .ZN(n2622) );
  OAI222D1BWP12T U2885 ( .A1(n2032), .A2(n2958), .B1(n2031), .B2(n2957), .C1(
        n2956), .C2(n2026), .ZN(n2238) );
  OAI222D1BWP12T U2886 ( .A1(n2032), .A2(n2966), .B1(n2031), .B2(n2965), .C1(
        n2964), .C2(n2027), .ZN(n2270) );
  CKND0BWP12T U2887 ( .I(r4[6]), .ZN(n2028) );
  OAI222D1BWP12T U2888 ( .A1(n2032), .A2(n2954), .B1(n2031), .B2(n2953), .C1(
        n2952), .C2(n2028), .ZN(n2494) );
  OAI222D1BWP12T U2889 ( .A1(n2032), .A2(n2978), .B1(n2031), .B2(n2977), .C1(
        n2976), .C2(n1412), .ZN(n2302) );
  OAI222D1BWP12T U2890 ( .A1(n2032), .A2(n2970), .B1(n2031), .B2(n2969), .C1(
        n2968), .C2(n2029), .ZN(n2526) );
  OAI222D1BWP12T U2891 ( .A1(n2032), .A2(n2974), .B1(n2031), .B2(n2973), .C1(
        n2972), .C2(n2030), .ZN(n2558) );
  AOI22D0BWP12T U2892 ( .A1(lr[17]), .A2(n3473), .B1(n3480), .B2(pc_out[17]), 
        .ZN(n2044) );
  AOI22D0BWP12T U2893 ( .A1(n3479), .A2(r12[17]), .B1(r11[17]), .B2(n2704), 
        .ZN(n2043) );
  AOI22D0BWP12T U2894 ( .A1(r5[17]), .A2(n3481), .B1(n2770), .B2(r6[17]), .ZN(
        n2036) );
  AOI22D0BWP12T U2895 ( .A1(r7[17]), .A2(n3482), .B1(n2757), .B2(r4[17]), .ZN(
        n2035) );
  AOI22D0BWP12T U2896 ( .A1(r1[17]), .A2(n3484), .B1(n3483), .B2(r2[17]), .ZN(
        n2034) );
  AOI22D0BWP12T U2897 ( .A1(r0[17]), .A2(n3486), .B1(n3485), .B2(r3[17]), .ZN(
        n2033) );
  ND4D1BWP12T U2898 ( .A1(n2036), .A2(n2035), .A3(n2034), .A4(n2033), .ZN(
        n2037) );
  AOI22D0BWP12T U2899 ( .A1(r8[17]), .A2(n3493), .B1(n2037), .B2(n3492), .ZN(
        n2042) );
  OAI22D0BWP12T U2900 ( .A1(n2039), .A2(n3474), .B1(n2805), .B2(n2038), .ZN(
        n2040) );
  AOI21D0BWP12T U2901 ( .A1(r10[17]), .A2(n2810), .B(n2040), .ZN(n2041) );
  ND4D1BWP12T U2902 ( .A1(n2044), .A2(n2043), .A3(n2042), .A4(n2041), .ZN(
        regC_out[17]) );
  AOI22D0BWP12T U2903 ( .A1(pc_out[13]), .A2(n3480), .B1(n3479), .B2(r12[13]), 
        .ZN(n2056) );
  AOI22D0BWP12T U2904 ( .A1(r5[13]), .A2(n3481), .B1(n2770), .B2(r6[13]), .ZN(
        n2048) );
  AOI22D0BWP12T U2905 ( .A1(r7[13]), .A2(n3482), .B1(n2757), .B2(r4[13]), .ZN(
        n2047) );
  AOI22D0BWP12T U2906 ( .A1(r1[13]), .A2(n3484), .B1(n3483), .B2(r2[13]), .ZN(
        n2046) );
  AOI22D0BWP12T U2907 ( .A1(r0[13]), .A2(n3486), .B1(n3485), .B2(r3[13]), .ZN(
        n2045) );
  ND4D1BWP12T U2908 ( .A1(n2048), .A2(n2047), .A3(n2046), .A4(n2045), .ZN(
        n2049) );
  AOI22D0BWP12T U2909 ( .A1(r8[13]), .A2(n3493), .B1(n2049), .B2(n3492), .ZN(
        n2055) );
  AOI22D0BWP12T U2910 ( .A1(r11[13]), .A2(n2704), .B1(n3475), .B2(r9[13]), 
        .ZN(n2054) );
  OAI22D0BWP12T U2911 ( .A1(n2051), .A2(n3474), .B1(n2779), .B2(n2050), .ZN(
        n2052) );
  AOI21D0BWP12T U2912 ( .A1(r10[13]), .A2(n2810), .B(n2052), .ZN(n2053) );
  ND4D1BWP12T U2913 ( .A1(n2056), .A2(n2055), .A3(n2054), .A4(n2053), .ZN(
        regC_out[13]) );
  AOI22D0BWP12T U2914 ( .A1(lr[22]), .A2(n3473), .B1(n3480), .B2(pc_out[22]), 
        .ZN(n2068) );
  AOI22D0BWP12T U2915 ( .A1(n3479), .A2(r12[22]), .B1(r9[22]), .B2(n3475), 
        .ZN(n2067) );
  AOI22D0BWP12T U2916 ( .A1(r5[22]), .A2(n3481), .B1(n2770), .B2(r6[22]), .ZN(
        n2060) );
  AOI22D0BWP12T U2917 ( .A1(r7[22]), .A2(n3482), .B1(n2757), .B2(r4[22]), .ZN(
        n2059) );
  AOI22D0BWP12T U2918 ( .A1(r1[22]), .A2(n3484), .B1(n3483), .B2(r2[22]), .ZN(
        n2058) );
  AOI22D0BWP12T U2919 ( .A1(r0[22]), .A2(n3486), .B1(n3485), .B2(r3[22]), .ZN(
        n2057) );
  ND4D1BWP12T U2920 ( .A1(n2060), .A2(n2059), .A3(n2058), .A4(n2057), .ZN(
        n2061) );
  AOI22D0BWP12T U2921 ( .A1(r8[22]), .A2(n3493), .B1(n2061), .B2(n3492), .ZN(
        n2066) );
  OAI22D0BWP12T U2922 ( .A1(n2063), .A2(n3474), .B1(n2803), .B2(n2062), .ZN(
        n2064) );
  AOI21D0BWP12T U2923 ( .A1(r10[22]), .A2(n2810), .B(n2064), .ZN(n2065) );
  ND4D1BWP12T U2924 ( .A1(n2068), .A2(n2067), .A3(n2066), .A4(n2065), .ZN(
        regC_out[22]) );
  OAI22D0BWP12T U2925 ( .A1(n3478), .A2(n2070), .B1(n3474), .B2(n2069), .ZN(
        n2071) );
  AOI21D0BWP12T U2926 ( .A1(lr[19]), .A2(n3473), .B(n2071), .ZN(n2080) );
  AOI22D0BWP12T U2927 ( .A1(r5[19]), .A2(n3481), .B1(n2770), .B2(r6[19]), .ZN(
        n2075) );
  AOI22D0BWP12T U2928 ( .A1(r7[19]), .A2(n3482), .B1(n2757), .B2(r4[19]), .ZN(
        n2074) );
  AOI22D0BWP12T U2929 ( .A1(r1[19]), .A2(n3484), .B1(n3483), .B2(r2[19]), .ZN(
        n2073) );
  AOI22D0BWP12T U2930 ( .A1(r0[19]), .A2(n3486), .B1(n3485), .B2(r3[19]), .ZN(
        n2072) );
  ND4D1BWP12T U2931 ( .A1(n2075), .A2(n2074), .A3(n2073), .A4(n2072), .ZN(
        n2076) );
  AOI22D0BWP12T U2932 ( .A1(r8[19]), .A2(n3493), .B1(n2076), .B2(n3492), .ZN(
        n2079) );
  AOI22D0BWP12T U2933 ( .A1(r11[19]), .A2(n2704), .B1(n3475), .B2(r9[19]), 
        .ZN(n2078) );
  AOI22D0BWP12T U2934 ( .A1(pc_out[19]), .A2(n3480), .B1(n3479), .B2(r12[19]), 
        .ZN(n2077) );
  ND4D1BWP12T U2935 ( .A1(n2080), .A2(n2079), .A3(n2078), .A4(n2077), .ZN(
        regC_out[19]) );
  OAI22D0BWP12T U2936 ( .A1(n3478), .A2(n2082), .B1(n2779), .B2(n2081), .ZN(
        n2083) );
  AOI21D0BWP12T U2937 ( .A1(n[3564]), .A2(n3464), .B(n2083), .ZN(n2092) );
  AOI22D0BWP12T U2938 ( .A1(r5[16]), .A2(n3481), .B1(n2770), .B2(r6[16]), .ZN(
        n2087) );
  AOI22D0BWP12T U2939 ( .A1(r7[16]), .A2(n3482), .B1(n2757), .B2(r4[16]), .ZN(
        n2086) );
  AOI22D0BWP12T U2940 ( .A1(r1[16]), .A2(n3484), .B1(n3483), .B2(r2[16]), .ZN(
        n2085) );
  AOI22D0BWP12T U2941 ( .A1(r0[16]), .A2(n3486), .B1(n3485), .B2(r3[16]), .ZN(
        n2084) );
  ND4D1BWP12T U2942 ( .A1(n2087), .A2(n2086), .A3(n2085), .A4(n2084), .ZN(
        n2088) );
  AOI22D0BWP12T U2943 ( .A1(r8[16]), .A2(n3493), .B1(n2088), .B2(n3492), .ZN(
        n2091) );
  AOI22D0BWP12T U2944 ( .A1(r11[16]), .A2(n2704), .B1(n3475), .B2(r9[16]), 
        .ZN(n2090) );
  AOI22D0BWP12T U2945 ( .A1(pc_out[16]), .A2(n3480), .B1(n3479), .B2(r12[16]), 
        .ZN(n2089) );
  ND4D1BWP12T U2946 ( .A1(n2092), .A2(n2091), .A3(n2090), .A4(n2089), .ZN(
        regC_out[16]) );
  AOI22D0BWP12T U2947 ( .A1(lr[18]), .A2(n3473), .B1(n3480), .B2(pc_out[18]), 
        .ZN(n2104) );
  AOI22D0BWP12T U2948 ( .A1(n3479), .A2(r12[18]), .B1(r9[18]), .B2(n3475), 
        .ZN(n2103) );
  AOI22D0BWP12T U2949 ( .A1(r5[18]), .A2(n3481), .B1(n2770), .B2(r6[18]), .ZN(
        n2096) );
  AOI22D0BWP12T U2950 ( .A1(r7[18]), .A2(n3482), .B1(n2757), .B2(r4[18]), .ZN(
        n2095) );
  AOI22D0BWP12T U2951 ( .A1(r1[18]), .A2(n3484), .B1(n3483), .B2(r2[18]), .ZN(
        n2094) );
  AOI22D0BWP12T U2952 ( .A1(r0[18]), .A2(n3486), .B1(n3485), .B2(r3[18]), .ZN(
        n2093) );
  ND4D1BWP12T U2953 ( .A1(n2096), .A2(n2095), .A3(n2094), .A4(n2093), .ZN(
        n2097) );
  AOI22D0BWP12T U2954 ( .A1(r8[18]), .A2(n3493), .B1(n2097), .B2(n3492), .ZN(
        n2102) );
  OAI22D0BWP12T U2955 ( .A1(n2099), .A2(n3474), .B1(n2803), .B2(n2098), .ZN(
        n2100) );
  AOI21D0BWP12T U2956 ( .A1(r10[18]), .A2(n2810), .B(n2100), .ZN(n2101) );
  ND4D1BWP12T U2957 ( .A1(n2104), .A2(n2103), .A3(n2102), .A4(n2101), .ZN(
        regC_out[18]) );
  AOI21D0BWP12T U2958 ( .A1(n3185), .A2(write2_in[7]), .B(reset), .ZN(n2106)
         );
  ND2XD0BWP12T U2959 ( .A1(n3186), .A2(n[3573]), .ZN(n2105) );
  OAI211D1BWP12T U2960 ( .A1(n2872), .A2(n2866), .B(n2106), .C(n2105), .ZN(
        spin[7]) );
  AOI22D0BWP12T U2961 ( .A1(n[3574]), .A2(n3464), .B1(n3479), .B2(r12[6]), 
        .ZN(n2116) );
  AOI22D0BWP12T U2962 ( .A1(r5[6]), .A2(n3481), .B1(n2770), .B2(r6[6]), .ZN(
        n2110) );
  AOI22D0BWP12T U2963 ( .A1(r7[6]), .A2(n3482), .B1(n2757), .B2(r4[6]), .ZN(
        n2109) );
  AOI22D0BWP12T U2964 ( .A1(r1[6]), .A2(n3484), .B1(n3483), .B2(r2[6]), .ZN(
        n2108) );
  AOI22D0BWP12T U2965 ( .A1(r0[6]), .A2(n3486), .B1(n3485), .B2(r3[6]), .ZN(
        n2107) );
  ND4D1BWP12T U2966 ( .A1(n2110), .A2(n2109), .A3(n2108), .A4(n2107), .ZN(
        n2111) );
  AOI22D0BWP12T U2967 ( .A1(r8[6]), .A2(n3493), .B1(n2111), .B2(n3492), .ZN(
        n2115) );
  AOI22D0BWP12T U2968 ( .A1(r11[6]), .A2(n2704), .B1(n3475), .B2(r9[6]), .ZN(
        n2114) );
  OAI22D0BWP12T U2969 ( .A1(n2874), .A2(n2806), .B1(n2779), .B2(n1413), .ZN(
        n2112) );
  AOI21D0BWP12T U2970 ( .A1(r10[6]), .A2(n2810), .B(n2112), .ZN(n2113) );
  ND4D1BWP12T U2971 ( .A1(n2116), .A2(n2115), .A3(n2114), .A4(n2113), .ZN(
        regC_out[6]) );
  AOI22D0BWP12T U2972 ( .A1(pc_out[9]), .A2(n3480), .B1(n3479), .B2(r12[9]), 
        .ZN(n2126) );
  AOI22D0BWP12T U2973 ( .A1(r5[9]), .A2(n3481), .B1(n2770), .B2(r6[9]), .ZN(
        n2120) );
  AOI22D0BWP12T U2974 ( .A1(r7[9]), .A2(n3482), .B1(n2757), .B2(r4[9]), .ZN(
        n2119) );
  AOI22D0BWP12T U2975 ( .A1(r1[9]), .A2(n3484), .B1(n3483), .B2(r2[9]), .ZN(
        n2118) );
  AOI22D0BWP12T U2976 ( .A1(r0[9]), .A2(n3486), .B1(n3485), .B2(r3[9]), .ZN(
        n2117) );
  ND4D1BWP12T U2977 ( .A1(n2120), .A2(n2119), .A3(n2118), .A4(n2117), .ZN(
        n2121) );
  AOI22D0BWP12T U2978 ( .A1(r8[9]), .A2(n3493), .B1(n2121), .B2(n3492), .ZN(
        n2125) );
  AOI22D0BWP12T U2979 ( .A1(r11[9]), .A2(n2704), .B1(n3475), .B2(r9[9]), .ZN(
        n2124) );
  OAI22D0BWP12T U2980 ( .A1(n2887), .A2(n3474), .B1(n2779), .B2(n2990), .ZN(
        n2122) );
  AOI21D0BWP12T U2981 ( .A1(r10[9]), .A2(n2810), .B(n2122), .ZN(n2123) );
  ND4D1BWP12T U2982 ( .A1(n2126), .A2(n2125), .A3(n2124), .A4(n2123), .ZN(
        regC_out[9]) );
  AOI22D0BWP12T U2983 ( .A1(pc_out[30]), .A2(n3480), .B1(n3479), .B2(r12[30]), 
        .ZN(n2261) );
  AOI22D0BWP12T U2984 ( .A1(r5[30]), .A2(n3481), .B1(n2770), .B2(r6[30]), .ZN(
        n2130) );
  AOI22D0BWP12T U2985 ( .A1(r7[30]), .A2(n3482), .B1(n2757), .B2(r4[30]), .ZN(
        n2129) );
  AOI22D0BWP12T U2986 ( .A1(r1[30]), .A2(n3484), .B1(n3483), .B2(r2[30]), .ZN(
        n2128) );
  AOI22D0BWP12T U2987 ( .A1(r0[30]), .A2(n3486), .B1(n3485), .B2(r3[30]), .ZN(
        n2127) );
  ND4D1BWP12T U2988 ( .A1(n2130), .A2(n2129), .A3(n2128), .A4(n2127), .ZN(
        n2131) );
  AOI22D0BWP12T U2989 ( .A1(r8[30]), .A2(n3493), .B1(n2131), .B2(n3492), .ZN(
        n2136) );
  AOI22D0BWP12T U2990 ( .A1(r11[30]), .A2(n2704), .B1(n3475), .B2(r9[30]), 
        .ZN(n2134) );
  OAI22D0BWP12T U2991 ( .A1(n3403), .A2(n3474), .B1(n2779), .B2(n3386), .ZN(
        n2132) );
  AOI21D0BWP12T U2992 ( .A1(r10[30]), .A2(n2810), .B(n2132), .ZN(n2133) );
  ND4D1BWP12T U2993 ( .A1(n2261), .A2(n2136), .A3(n2134), .A4(n2133), .ZN(
        regC_out[30]) );
  AOI22D0BWP12T U2994 ( .A1(lr[25]), .A2(n3473), .B1(n3479), .B2(r12[25]), 
        .ZN(n2650) );
  AOI22D0BWP12T U2995 ( .A1(r5[25]), .A2(n3481), .B1(n2770), .B2(r6[25]), .ZN(
        n2389) );
  AOI22D0BWP12T U2996 ( .A1(r7[25]), .A2(n3482), .B1(n2757), .B2(r4[25]), .ZN(
        n2327) );
  AOI22D0BWP12T U2997 ( .A1(r1[25]), .A2(n3484), .B1(n3483), .B2(r2[25]), .ZN(
        n2325) );
  AOI22D0BWP12T U2998 ( .A1(r0[25]), .A2(n3486), .B1(n3485), .B2(r3[25]), .ZN(
        n2293) );
  ND4D1BWP12T U2999 ( .A1(n2389), .A2(n2327), .A3(n2325), .A4(n2293), .ZN(
        n2517) );
  AOI22D0BWP12T U3000 ( .A1(r8[25]), .A2(n3493), .B1(n2517), .B2(n3492), .ZN(
        n2649) );
  AOI22D0BWP12T U3001 ( .A1(r11[25]), .A2(n2704), .B1(n3475), .B2(r9[25]), 
        .ZN(n2648) );
  OAI22D0BWP12T U3002 ( .A1(n3536), .A2(n2806), .B1(n2549), .B2(n3474), .ZN(
        n2581) );
  AOI21D0BWP12T U3003 ( .A1(r10[25]), .A2(n2810), .B(n2581), .ZN(n2645) );
  ND4D1BWP12T U3004 ( .A1(n2650), .A2(n2649), .A3(n2648), .A4(n2645), .ZN(
        regC_out[25]) );
  AOI22D0BWP12T U3005 ( .A1(n[3551]), .A2(n3464), .B1(n3479), .B2(r12[29]), 
        .ZN(n2661) );
  AOI22D0BWP12T U3006 ( .A1(r5[29]), .A2(n3481), .B1(n2770), .B2(r6[29]), .ZN(
        n2654) );
  AOI22D0BWP12T U3007 ( .A1(r7[29]), .A2(n3482), .B1(n2757), .B2(r4[29]), .ZN(
        n2653) );
  AOI22D0BWP12T U3008 ( .A1(r1[29]), .A2(n3484), .B1(n3483), .B2(r2[29]), .ZN(
        n2652) );
  AOI22D0BWP12T U3009 ( .A1(r0[29]), .A2(n3486), .B1(n3485), .B2(r3[29]), .ZN(
        n2651) );
  ND4D1BWP12T U3010 ( .A1(n2654), .A2(n2653), .A3(n2652), .A4(n2651), .ZN(
        n2655) );
  AOI22D0BWP12T U3011 ( .A1(r8[29]), .A2(n3493), .B1(n2655), .B2(n3492), .ZN(
        n2660) );
  AOI22D0BWP12T U3012 ( .A1(r11[29]), .A2(n2704), .B1(n3475), .B2(r9[29]), 
        .ZN(n2659) );
  OAI22D0BWP12T U3013 ( .A1(n3533), .A2(n2806), .B1(n2779), .B2(n2656), .ZN(
        n2657) );
  AOI21D0BWP12T U3014 ( .A1(r10[29]), .A2(n2810), .B(n2657), .ZN(n2658) );
  ND4D1BWP12T U3015 ( .A1(n2661), .A2(n2660), .A3(n2659), .A4(n2658), .ZN(
        regC_out[29]) );
  AOI22D0BWP12T U3016 ( .A1(lr[15]), .A2(n3473), .B1(n3464), .B2(n[3565]), 
        .ZN(n2673) );
  AOI22D0BWP12T U3017 ( .A1(pc_out[15]), .A2(n3480), .B1(n3479), .B2(r12[15]), 
        .ZN(n2672) );
  OAI22D0BWP12T U3018 ( .A1(n2803), .A2(n2663), .B1(n2662), .B2(n2805), .ZN(
        n2664) );
  AOI21D0BWP12T U3019 ( .A1(r10[15]), .A2(n2810), .B(n2664), .ZN(n2671) );
  AOI22D0BWP12T U3020 ( .A1(r5[15]), .A2(n3481), .B1(n2770), .B2(r6[15]), .ZN(
        n2668) );
  AOI22D0BWP12T U3021 ( .A1(r7[15]), .A2(n3482), .B1(n2757), .B2(r4[15]), .ZN(
        n2667) );
  AOI22D0BWP12T U3022 ( .A1(r1[15]), .A2(n3484), .B1(n3483), .B2(r2[15]), .ZN(
        n2666) );
  AOI22D0BWP12T U3023 ( .A1(r0[15]), .A2(n3486), .B1(n3485), .B2(r3[15]), .ZN(
        n2665) );
  ND4D1BWP12T U3024 ( .A1(n2668), .A2(n2667), .A3(n2666), .A4(n2665), .ZN(
        n2669) );
  AOI22D0BWP12T U3025 ( .A1(r8[15]), .A2(n3493), .B1(n2669), .B2(n3492), .ZN(
        n2670) );
  ND4D1BWP12T U3026 ( .A1(n2673), .A2(n2672), .A3(n2671), .A4(n2670), .ZN(
        regC_out[15]) );
  AOI22D0BWP12T U3027 ( .A1(lr[28]), .A2(n3473), .B1(n3480), .B2(pc_out[28]), 
        .ZN(n2685) );
  AOI22D0BWP12T U3028 ( .A1(n3479), .A2(r12[28]), .B1(r9[28]), .B2(n3475), 
        .ZN(n2684) );
  AOI22D0BWP12T U3029 ( .A1(r5[28]), .A2(n3481), .B1(n2770), .B2(r6[28]), .ZN(
        n2677) );
  AOI22D0BWP12T U3030 ( .A1(r7[28]), .A2(n3482), .B1(n2757), .B2(r4[28]), .ZN(
        n2676) );
  AOI22D0BWP12T U3031 ( .A1(r1[28]), .A2(n3484), .B1(n3483), .B2(r2[28]), .ZN(
        n2675) );
  AOI22D0BWP12T U3032 ( .A1(r0[28]), .A2(n3486), .B1(n3485), .B2(r3[28]), .ZN(
        n2674) );
  ND4D1BWP12T U3033 ( .A1(n2677), .A2(n2676), .A3(n2675), .A4(n2674), .ZN(
        n2678) );
  AOI22D0BWP12T U3034 ( .A1(r8[28]), .A2(n3493), .B1(n2678), .B2(n3492), .ZN(
        n2683) );
  OAI22D0BWP12T U3035 ( .A1(n2680), .A2(n3474), .B1(n2803), .B2(n2679), .ZN(
        n2681) );
  AOI21D0BWP12T U3036 ( .A1(r10[28]), .A2(n2810), .B(n2681), .ZN(n2682) );
  ND4D1BWP12T U3037 ( .A1(n2685), .A2(n2684), .A3(n2683), .A4(n2682), .ZN(
        regC_out[28]) );
  AOI22D0BWP12T U3038 ( .A1(n[3570]), .A2(n3464), .B1(n3480), .B2(pc_out[10]), 
        .ZN(n2695) );
  AOI22D0BWP12T U3039 ( .A1(n3479), .A2(r12[10]), .B1(r9[10]), .B2(n3475), 
        .ZN(n2694) );
  AOI22D0BWP12T U3040 ( .A1(r5[10]), .A2(n3481), .B1(n2770), .B2(r6[10]), .ZN(
        n2689) );
  AOI22D0BWP12T U3041 ( .A1(r7[10]), .A2(n3482), .B1(n2757), .B2(r4[10]), .ZN(
        n2688) );
  AOI22D0BWP12T U3042 ( .A1(r1[10]), .A2(n3484), .B1(n3483), .B2(r2[10]), .ZN(
        n2687) );
  AOI22D0BWP12T U3043 ( .A1(r0[10]), .A2(n3486), .B1(n3485), .B2(r3[10]), .ZN(
        n2686) );
  ND4D1BWP12T U3044 ( .A1(n2689), .A2(n2688), .A3(n2687), .A4(n2686), .ZN(
        n2690) );
  AOI22D0BWP12T U3045 ( .A1(r8[10]), .A2(n3493), .B1(n2690), .B2(n3492), .ZN(
        n2693) );
  OAI22D0BWP12T U3046 ( .A1(n2779), .A2(n3023), .B1(n2963), .B2(n2803), .ZN(
        n2691) );
  AOI21D0BWP12T U3047 ( .A1(r10[10]), .A2(n2810), .B(n2691), .ZN(n2692) );
  ND4D1BWP12T U3048 ( .A1(n2695), .A2(n2694), .A3(n2693), .A4(n2692), .ZN(
        regC_out[10]) );
  AOI22D0BWP12T U3049 ( .A1(n[3556]), .A2(n3464), .B1(n3480), .B2(pc_out[24]), 
        .ZN(n2708) );
  OAI22D0BWP12T U3050 ( .A1(n2779), .A2(n2697), .B1(n2696), .B2(n2744), .ZN(
        n2698) );
  AOI21D0BWP12T U3051 ( .A1(r10[24]), .A2(n2810), .B(n2698), .ZN(n2707) );
  AOI22D0BWP12T U3052 ( .A1(r5[24]), .A2(n3481), .B1(n2770), .B2(r6[24]), .ZN(
        n2702) );
  AOI22D0BWP12T U3053 ( .A1(r7[24]), .A2(n3482), .B1(n2757), .B2(r4[24]), .ZN(
        n2701) );
  AOI22D0BWP12T U3054 ( .A1(r1[24]), .A2(n3484), .B1(n3483), .B2(r2[24]), .ZN(
        n2700) );
  AOI22D0BWP12T U3055 ( .A1(r0[24]), .A2(n3486), .B1(n3485), .B2(r3[24]), .ZN(
        n2699) );
  ND4D1BWP12T U3056 ( .A1(n2702), .A2(n2701), .A3(n2700), .A4(n2699), .ZN(
        n2703) );
  AOI22D0BWP12T U3057 ( .A1(r8[24]), .A2(n3493), .B1(n2703), .B2(n3492), .ZN(
        n2706) );
  AOI22D0BWP12T U3058 ( .A1(r11[24]), .A2(n2704), .B1(n3475), .B2(r9[24]), 
        .ZN(n2705) );
  ND4D1BWP12T U3059 ( .A1(n2708), .A2(n2707), .A3(n2706), .A4(n2705), .ZN(
        regC_out[24]) );
  AOI22D0BWP12T U3060 ( .A1(lr[0]), .A2(n3473), .B1(n3464), .B2(n[3580]), .ZN(
        n2721) );
  AOI22D0BWP12T U3061 ( .A1(pc_out[0]), .A2(n3480), .B1(n3479), .B2(r12[0]), 
        .ZN(n2720) );
  OAI22D0BWP12T U3062 ( .A1(n2803), .A2(n3067), .B1(n2711), .B2(n2805), .ZN(
        n2712) );
  AOI21D0BWP12T U3063 ( .A1(r10[0]), .A2(n2810), .B(n2712), .ZN(n2719) );
  AOI22D0BWP12T U3064 ( .A1(r5[0]), .A2(n3481), .B1(n2770), .B2(r6[0]), .ZN(
        n2716) );
  AOI22D0BWP12T U3065 ( .A1(r7[0]), .A2(n3482), .B1(n2757), .B2(r4[0]), .ZN(
        n2715) );
  AOI22D0BWP12T U3066 ( .A1(r1[0]), .A2(n3484), .B1(n3483), .B2(r2[0]), .ZN(
        n2714) );
  AOI22D0BWP12T U3067 ( .A1(r0[0]), .A2(n3486), .B1(n3485), .B2(r3[0]), .ZN(
        n2713) );
  ND4D1BWP12T U3068 ( .A1(n2716), .A2(n2715), .A3(n2714), .A4(n2713), .ZN(
        n2717) );
  AOI22D0BWP12T U3069 ( .A1(r8[0]), .A2(n3493), .B1(n2717), .B2(n3492), .ZN(
        n2718) );
  ND4D1BWP12T U3070 ( .A1(n2721), .A2(n2720), .A3(n2719), .A4(n2718), .ZN(
        regC_out[0]) );
  AOI22D0BWP12T U3071 ( .A1(lr[27]), .A2(n3473), .B1(n3464), .B2(n[3553]), 
        .ZN(n2732) );
  OAI22D0BWP12T U3072 ( .A1(n3538), .A2(n2806), .B1(n2803), .B2(n2722), .ZN(
        n2723) );
  AOI21D0BWP12T U3073 ( .A1(r10[27]), .A2(n2810), .B(n2723), .ZN(n2731) );
  AOI22D0BWP12T U3074 ( .A1(n3479), .A2(r12[27]), .B1(r9[27]), .B2(n3475), 
        .ZN(n2730) );
  AOI22D0BWP12T U3075 ( .A1(r5[27]), .A2(n3481), .B1(n2770), .B2(r6[27]), .ZN(
        n2727) );
  AOI22D0BWP12T U3076 ( .A1(r7[27]), .A2(n3482), .B1(n2757), .B2(r4[27]), .ZN(
        n2726) );
  AOI22D0BWP12T U3077 ( .A1(r1[27]), .A2(n3484), .B1(n3483), .B2(r2[27]), .ZN(
        n2725) );
  AOI22D0BWP12T U3078 ( .A1(r0[27]), .A2(n3486), .B1(n3485), .B2(r3[27]), .ZN(
        n2724) );
  ND4D1BWP12T U3079 ( .A1(n2727), .A2(n2726), .A3(n2725), .A4(n2724), .ZN(
        n2728) );
  AOI22D0BWP12T U3080 ( .A1(r8[27]), .A2(n3493), .B1(n2728), .B2(n3492), .ZN(
        n2729) );
  ND4D1BWP12T U3081 ( .A1(n2732), .A2(n2731), .A3(n2730), .A4(n2729), .ZN(
        regC_out[27]) );
  AOI22D0BWP12T U3082 ( .A1(lr[5]), .A2(n3473), .B1(n3464), .B2(n[3575]), .ZN(
        n2743) );
  AOI22D0BWP12T U3083 ( .A1(pc_out[5]), .A2(n3480), .B1(n3479), .B2(r12[5]), 
        .ZN(n2742) );
  OAI22D0BWP12T U3084 ( .A1(n2803), .A2(n2869), .B1(n2733), .B2(n2805), .ZN(
        n2734) );
  AOI21D0BWP12T U3085 ( .A1(r10[5]), .A2(n2810), .B(n2734), .ZN(n2741) );
  AOI22D0BWP12T U3086 ( .A1(r5[5]), .A2(n3481), .B1(n2770), .B2(r6[5]), .ZN(
        n2738) );
  AOI22D0BWP12T U3087 ( .A1(r7[5]), .A2(n3482), .B1(n2757), .B2(r4[5]), .ZN(
        n2737) );
  AOI22D0BWP12T U3088 ( .A1(r1[5]), .A2(n3484), .B1(n3483), .B2(r2[5]), .ZN(
        n2736) );
  AOI22D0BWP12T U3089 ( .A1(r0[5]), .A2(n3486), .B1(n3485), .B2(r3[5]), .ZN(
        n2735) );
  ND4D1BWP12T U3090 ( .A1(n2738), .A2(n2737), .A3(n2736), .A4(n2735), .ZN(
        n2739) );
  AOI22D0BWP12T U3091 ( .A1(r8[5]), .A2(n3493), .B1(n2739), .B2(n3492), .ZN(
        n2740) );
  ND4D1BWP12T U3092 ( .A1(n2743), .A2(n2742), .A3(n2741), .A4(n2740), .ZN(
        regC_out[5]) );
  AOI22D0BWP12T U3093 ( .A1(lr[3]), .A2(n3473), .B1(n3464), .B2(n[3577]), .ZN(
        n2754) );
  AOI22D0BWP12T U3094 ( .A1(n3480), .A2(pc_out[3]), .B1(r9[3]), .B2(n3475), 
        .ZN(n2753) );
  OAI22D0BWP12T U3095 ( .A1(n2803), .A2(n2852), .B1(n2850), .B2(n2744), .ZN(
        n2745) );
  AOI21D0BWP12T U3096 ( .A1(r10[3]), .A2(n2810), .B(n2745), .ZN(n2752) );
  AOI22D0BWP12T U3097 ( .A1(r5[3]), .A2(n3481), .B1(n2770), .B2(r6[3]), .ZN(
        n2749) );
  AOI22D0BWP12T U3098 ( .A1(r7[3]), .A2(n3482), .B1(n2757), .B2(r4[3]), .ZN(
        n2748) );
  AOI22D0BWP12T U3099 ( .A1(r1[3]), .A2(n3484), .B1(n3483), .B2(r2[3]), .ZN(
        n2747) );
  AOI22D0BWP12T U3100 ( .A1(r0[3]), .A2(n3486), .B1(n3485), .B2(r3[3]), .ZN(
        n2746) );
  ND4D1BWP12T U3101 ( .A1(n2749), .A2(n2748), .A3(n2747), .A4(n2746), .ZN(
        n2750) );
  AOI22D0BWP12T U3102 ( .A1(r8[3]), .A2(n3493), .B1(n2750), .B2(n3492), .ZN(
        n2751) );
  ND4D1BWP12T U3103 ( .A1(n2754), .A2(n2753), .A3(n2752), .A4(n2751), .ZN(
        regC_out[3]) );
  AOI22D0BWP12T U3104 ( .A1(lr[2]), .A2(n3473), .B1(n3464), .B2(n[3578]), .ZN(
        n2766) );
  AOI22D0BWP12T U3105 ( .A1(pc_out[2]), .A2(n3480), .B1(n3479), .B2(r12[2]), 
        .ZN(n2765) );
  OAI22D0BWP12T U3106 ( .A1(n2803), .A2(n2755), .B1(n2854), .B2(n3478), .ZN(
        n2756) );
  AOI21D0BWP12T U3107 ( .A1(r8[2]), .A2(n3493), .B(n2756), .ZN(n2764) );
  AOI22D0BWP12T U3108 ( .A1(r5[2]), .A2(n3481), .B1(n2770), .B2(r6[2]), .ZN(
        n2761) );
  AOI22D0BWP12T U3109 ( .A1(r7[2]), .A2(n3482), .B1(n2757), .B2(r4[2]), .ZN(
        n2760) );
  AOI22D0BWP12T U3110 ( .A1(r1[2]), .A2(n3484), .B1(n3483), .B2(r2[2]), .ZN(
        n2759) );
  AOI22D0BWP12T U3111 ( .A1(r0[2]), .A2(n3486), .B1(n3485), .B2(r3[2]), .ZN(
        n2758) );
  ND4D1BWP12T U3112 ( .A1(n2761), .A2(n2760), .A3(n2759), .A4(n2758), .ZN(
        n2762) );
  AOI22D0BWP12T U3113 ( .A1(r9[2]), .A2(n3475), .B1(n2762), .B2(n3492), .ZN(
        n2763) );
  ND4D1BWP12T U3114 ( .A1(n2766), .A2(n2765), .A3(n2764), .A4(n2763), .ZN(
        regC_out[2]) );
  AOI22D0BWP12T U3115 ( .A1(pc_out[7]), .A2(n3480), .B1(n3479), .B2(r12[7]), 
        .ZN(n2778) );
  OAI22D0BWP12T U3116 ( .A1(n2779), .A2(n2767), .B1(n2860), .B2(n2800), .ZN(
        n2769) );
  CKND0BWP12T U3117 ( .I(n[3573]), .ZN(n2861) );
  CKND0BWP12T U3118 ( .I(r11[7]), .ZN(n2847) );
  OAI22D0BWP12T U3119 ( .A1(n2861), .A2(n3474), .B1(n2803), .B2(n2847), .ZN(
        n2768) );
  AOI211D0BWP12T U3120 ( .A1(n2810), .A2(r10[7]), .B(n2769), .C(n2768), .ZN(
        n2777) );
  AOI22D0BWP12T U3121 ( .A1(r5[7]), .A2(n3481), .B1(n2770), .B2(r6[7]), .ZN(
        n2774) );
  AOI22D0BWP12T U3122 ( .A1(r7[7]), .A2(n3482), .B1(n2757), .B2(r4[7]), .ZN(
        n2773) );
  AOI22D0BWP12T U3123 ( .A1(r1[7]), .A2(n3484), .B1(n3483), .B2(r2[7]), .ZN(
        n2772) );
  AOI22D0BWP12T U3124 ( .A1(r0[7]), .A2(n3486), .B1(n3485), .B2(r3[7]), .ZN(
        n2771) );
  ND4D1BWP12T U3125 ( .A1(n2774), .A2(n2773), .A3(n2772), .A4(n2771), .ZN(
        n2775) );
  AOI22D0BWP12T U3126 ( .A1(n3475), .A2(r9[7]), .B1(n3492), .B2(n2775), .ZN(
        n2776) );
  ND3D1BWP12T U3127 ( .A1(n2778), .A2(n2777), .A3(n2776), .ZN(regC_out[7]) );
  AOI22D0BWP12T U3128 ( .A1(n[3569]), .A2(n3464), .B1(n3480), .B2(pc_out[11]), 
        .ZN(n2789) );
  OAI22D0BWP12T U3129 ( .A1(n2779), .A2(n3027), .B1(n3025), .B2(n2800), .ZN(
        n2781) );
  OAI22D0BWP12T U3130 ( .A1(n2803), .A2(n3026), .B1(n2875), .B2(n2805), .ZN(
        n2780) );
  AOI211D0BWP12T U3131 ( .A1(n2810), .A2(r10[11]), .B(n2781), .C(n2780), .ZN(
        n2788) );
  AOI22D0BWP12T U3132 ( .A1(r5[11]), .A2(n3481), .B1(n2770), .B2(r6[11]), .ZN(
        n2785) );
  AOI22D0BWP12T U3133 ( .A1(r7[11]), .A2(n3482), .B1(n2757), .B2(r4[11]), .ZN(
        n2784) );
  AOI22D0BWP12T U3134 ( .A1(r1[11]), .A2(n3484), .B1(n3483), .B2(r2[11]), .ZN(
        n2783) );
  AOI22D0BWP12T U3135 ( .A1(r0[11]), .A2(n3486), .B1(n3485), .B2(r3[11]), .ZN(
        n2782) );
  ND4D1BWP12T U3136 ( .A1(n2785), .A2(n2784), .A3(n2783), .A4(n2782), .ZN(
        n2786) );
  AOI22D0BWP12T U3137 ( .A1(n3479), .A2(r12[11]), .B1(n3492), .B2(n2786), .ZN(
        n2787) );
  ND3D1BWP12T U3138 ( .A1(n2789), .A2(n2788), .A3(n2787), .ZN(regC_out[11]) );
  AOI22D0BWP12T U3139 ( .A1(lr[8]), .A2(n3473), .B1(n3464), .B2(n[3572]), .ZN(
        n2799) );
  OAI22D0BWP12T U3140 ( .A1(n2803), .A2(n2907), .B1(n2995), .B2(n3478), .ZN(
        n2791) );
  OAI22D0BWP12T U3141 ( .A1(n2997), .A2(n2806), .B1(n2805), .B2(n2935), .ZN(
        n2790) );
  AOI211D0BWP12T U3142 ( .A1(n3493), .A2(r8[8]), .B(n2791), .C(n2790), .ZN(
        n2798) );
  AOI22D0BWP12T U3143 ( .A1(r5[8]), .A2(n3481), .B1(n2770), .B2(r6[8]), .ZN(
        n2795) );
  AOI22D0BWP12T U3144 ( .A1(r7[8]), .A2(n3482), .B1(n2757), .B2(r4[8]), .ZN(
        n2794) );
  AOI22D0BWP12T U3145 ( .A1(r1[8]), .A2(n3484), .B1(n3483), .B2(r2[8]), .ZN(
        n2793) );
  AOI22D0BWP12T U3146 ( .A1(r0[8]), .A2(n3486), .B1(n3485), .B2(r3[8]), .ZN(
        n2792) );
  ND4D1BWP12T U3147 ( .A1(n2795), .A2(n2794), .A3(n2793), .A4(n2792), .ZN(
        n2796) );
  AOI22D0BWP12T U3148 ( .A1(n3479), .A2(r12[8]), .B1(n3492), .B2(n2796), .ZN(
        n2797) );
  ND3D1BWP12T U3149 ( .A1(n2799), .A2(n2798), .A3(n2797), .ZN(regC_out[8]) );
  AOI22D0BWP12T U3150 ( .A1(lr[1]), .A2(n3473), .B1(n3464), .B2(n[3579]), .ZN(
        n2818) );
  OAI22D0BWP12T U3151 ( .A1(n2803), .A2(n2802), .B1(n2801), .B2(n2800), .ZN(
        n2809) );
  OAI22D0BWP12T U3152 ( .A1(n2807), .A2(n2806), .B1(n2805), .B2(n2804), .ZN(
        n2808) );
  AOI211D0BWP12T U3153 ( .A1(n2810), .A2(r10[1]), .B(n2809), .C(n2808), .ZN(
        n2817) );
  AOI22D0BWP12T U3154 ( .A1(r5[1]), .A2(n3481), .B1(n2770), .B2(r6[1]), .ZN(
        n2814) );
  AOI22D0BWP12T U3155 ( .A1(r7[1]), .A2(n3482), .B1(n2757), .B2(r4[1]), .ZN(
        n2813) );
  AOI22D0BWP12T U3156 ( .A1(r1[1]), .A2(n3484), .B1(n3483), .B2(r2[1]), .ZN(
        n2812) );
  AOI22D0BWP12T U3157 ( .A1(r0[1]), .A2(n3486), .B1(n3485), .B2(r3[1]), .ZN(
        n2811) );
  ND4D1BWP12T U3158 ( .A1(n2814), .A2(n2813), .A3(n2812), .A4(n2811), .ZN(
        n2815) );
  AOI22D0BWP12T U3159 ( .A1(n3479), .A2(r12[1]), .B1(n3492), .B2(n2815), .ZN(
        n2816) );
  ND3D1BWP12T U3160 ( .A1(n2818), .A2(n2817), .A3(n2816), .ZN(regC_out[1]) );
  OAI222D1BWP12T U3161 ( .A1(n2826), .A2(n2970), .B1(n2825), .B2(n2969), .C1(
        n2968), .C2(n2819), .ZN(n2520) );
  OAI222D1BWP12T U3162 ( .A1(n2826), .A2(n2958), .B1(n2825), .B2(n2957), .C1(
        n2956), .C2(n2820), .ZN(n2232) );
  OAI222D1BWP12T U3163 ( .A1(n2826), .A2(n2978), .B1(n2825), .B2(n2977), .C1(
        n2976), .C2(n3065), .ZN(n2296) );
  OAI222D1BWP12T U3164 ( .A1(n2826), .A2(n2982), .B1(n2825), .B2(n2981), .C1(
        n2980), .C2(n2821), .ZN(n2616) );
  OAI222D1BWP12T U3165 ( .A1(n2826), .A2(n2954), .B1(n2825), .B2(n2953), .C1(
        n2952), .C2(n2822), .ZN(n2488) );
  OAI222D1BWP12T U3166 ( .A1(n2826), .A2(n2962), .B1(n2825), .B2(n2961), .C1(
        n2960), .C2(n2823), .ZN(n2360) );
  OAI222D1BWP12T U3167 ( .A1(n2826), .A2(n2966), .B1(n2825), .B2(n2965), .C1(
        n2964), .C2(n3067), .ZN(n2264) );
  OAI222D1BWP12T U3168 ( .A1(n2826), .A2(n2974), .B1(n2825), .B2(n2973), .C1(
        n2972), .C2(n2824), .ZN(n2552) );
  ND2D1BWP12T U3169 ( .A1(readD_sel[0]), .A2(readD_sel[1]), .ZN(n2837) );
  INVD1BWP12T U3170 ( .I(readD_sel[4]), .ZN(n3086) );
  ND3D1BWP12T U3171 ( .A1(readD_sel[3]), .A2(readD_sel[2]), .A3(n3086), .ZN(
        n2830) );
  NR2D1BWP12T U3172 ( .A1(n2837), .A2(n2830), .ZN(n3061) );
  INVD1BWP12T U3173 ( .I(readD_sel[2]), .ZN(n2833) );
  ND3D1BWP12T U3174 ( .A1(readD_sel[3]), .A2(n3086), .A3(n2833), .ZN(n2828) );
  NR2D1BWP12T U3175 ( .A1(n2837), .A2(n2828), .ZN(n2994) );
  OR2XD1BWP12T U3176 ( .A1(readD_sel[1]), .A2(readD_sel[0]), .Z(n2839) );
  NR2D1BWP12T U3177 ( .A1(n2839), .A2(n2830), .ZN(n3064) );
  INVD1BWP12T U3178 ( .I(readD_sel[0]), .ZN(n2827) );
  OR2XD1BWP12T U3179 ( .A1(readD_sel[1]), .A2(n2827), .Z(n2835) );
  NR2D1BWP12T U3180 ( .A1(n2835), .A2(n2828), .ZN(n3063) );
  NR2D1BWP12T U3181 ( .A1(n2839), .A2(n2828), .ZN(n3073) );
  ND2D1BWP12T U3182 ( .A1(readD_sel[1]), .A2(n2827), .ZN(n2836) );
  NR2D1BWP12T U3183 ( .A1(n2836), .A2(n2828), .ZN(n3029) );
  INVD1BWP12T U3184 ( .I(n3029), .ZN(n3066) );
  NR2D1BWP12T U3185 ( .A1(n2835), .A2(n2830), .ZN(n3037) );
  INVD1BWP12T U3186 ( .I(n3037), .ZN(n3069) );
  NR2D1BWP12T U3187 ( .A1(n2836), .A2(n2830), .ZN(n3062) );
  INVD1BWP12T U3188 ( .I(n3062), .ZN(n3042) );
  INVD1BWP12T U3189 ( .I(readD_sel[3]), .ZN(n2834) );
  ND2D1BWP12T U3190 ( .A1(readD_sel[2]), .A2(n2834), .ZN(n2840) );
  NR2D1BWP12T U3191 ( .A1(n2840), .A2(n2835), .ZN(n3075) );
  ND2D1BWP12T U3192 ( .A1(n2834), .A2(n2833), .ZN(n2838) );
  NR2D1BWP12T U3193 ( .A1(n2838), .A2(n2835), .ZN(n3074) );
  NR2D1BWP12T U3194 ( .A1(n2836), .A2(n2840), .ZN(n3077) );
  NR2D1BWP12T U3195 ( .A1(n2837), .A2(n2840), .ZN(n3076) );
  NR2D1BWP12T U3196 ( .A1(n2838), .A2(n2836), .ZN(n3079) );
  NR2D1BWP12T U3197 ( .A1(n2837), .A2(n2838), .ZN(n3078) );
  NR2D1BWP12T U3198 ( .A1(n2838), .A2(n2839), .ZN(n3081) );
  NR2D1BWP12T U3199 ( .A1(n2840), .A2(n2839), .ZN(n3080) );
  INVD0BWP12T U3200 ( .I(n3063), .ZN(n2886) );
  OAI222D1BWP12T U3201 ( .A1(n2867), .A2(n2962), .B1(n2866), .B2(n2961), .C1(
        n2960), .C2(n2860), .ZN(n2367) );
  OAI222D1BWP12T U3202 ( .A1(n2867), .A2(n2958), .B1(n2866), .B2(n2957), .C1(
        n2956), .C2(n2846), .ZN(n2239) );
  OAI222D1BWP12T U3203 ( .A1(n2867), .A2(n2966), .B1(n2866), .B2(n2965), .C1(
        n2964), .C2(n2847), .ZN(n2271) );
  OAI222D1BWP12T U3204 ( .A1(n2867), .A2(n2970), .B1(n2866), .B2(n2969), .C1(
        n2968), .C2(n2848), .ZN(n2527) );
  OAI222D1BWP12T U3205 ( .A1(n2867), .A2(n2974), .B1(n2866), .B2(n2973), .C1(
        n2972), .C2(n2849), .ZN(n2559) );
  OAI222D1BWP12T U3206 ( .A1(n2867), .A2(n2978), .B1(n2866), .B2(n2977), .C1(
        n2976), .C2(n2859), .ZN(n2303) );
  CKND0BWP12T U3207 ( .I(n3064), .ZN(n2920) );
  INVD1BWP12T U3208 ( .I(n2994), .ZN(n3068) );
  TPAOI21D0BWP12T U3209 ( .A1(n3185), .A2(write2_in[8]), .B(reset), .ZN(n2858)
         );
  TPND2D0BWP12T U3210 ( .A1(n3186), .A2(n[3572]), .ZN(n2857) );
  OAI211D1BWP12T U3211 ( .A1(n2872), .A2(n2934), .B(n2858), .C(n2857), .ZN(
        spin[8]) );
  CKND0BWP12T U3212 ( .I(n3073), .ZN(n3024) );
  TPAOI21D0BWP12T U3213 ( .A1(n3185), .A2(write2_in[9]), .B(reset), .ZN(n2863)
         );
  TPND2D0BWP12T U3214 ( .A1(n3186), .A2(n[3571]), .ZN(n2862) );
  OAI211D1BWP12T U3215 ( .A1(n2872), .A2(n2989), .B(n2863), .C(n2862), .ZN(
        spin[9]) );
  OAI222D1BWP12T U3216 ( .A1(n2867), .A2(n2982), .B1(n2866), .B2(n2981), .C1(
        n2980), .C2(n2864), .ZN(n2623) );
  OAI222D1BWP12T U3217 ( .A1(n2867), .A2(n2954), .B1(n2866), .B2(n2953), .C1(
        n2952), .C2(n2865), .ZN(n2495) );
  TPAOI21D0BWP12T U3218 ( .A1(n3185), .A2(write2_in[10]), .B(reset), .ZN(n2871) );
  TPND2D0BWP12T U3219 ( .A1(n3186), .A2(n[3570]), .ZN(n2870) );
  OAI211D1BWP12T U3220 ( .A1(n2872), .A2(n3021), .B(n2871), .C(n2870), .ZN(
        spin[10]) );
  CKND0BWP12T U3221 ( .I(n3061), .ZN(n3028) );
  OAI22D1BWP12T U3222 ( .A1(n3016), .A2(n2875), .B1(n3014), .B2(n2902), .ZN(
        n2876) );
  AO21D1BWP12T U3223 ( .A1(write1_in[11]), .A2(n3269), .B(n2876), .Z(n2339) );
  OAI22D1BWP12T U3224 ( .A1(n3022), .A2(n3027), .B1(n3018), .B2(n2902), .ZN(
        n2877) );
  AO21D1BWP12T U3225 ( .A1(write1_in[11]), .A2(n3259), .B(n2877), .Z(n2211) );
  OAI22D1BWP12T U3226 ( .A1(n3000), .A2(n2878), .B1(n2998), .B2(n2902), .ZN(
        n2879) );
  AO21D1BWP12T U3227 ( .A1(write1_in[11]), .A2(n3264), .B(n2879), .Z(n2403) );
  OAI22D1BWP12T U3228 ( .A1(n3008), .A2(n2880), .B1(n3006), .B2(n2902), .ZN(
        n2881) );
  AO21D1BWP12T U3229 ( .A1(write1_in[11]), .A2(n3274), .B(n2881), .Z(n2435) );
  OAI22D1BWP12T U3230 ( .A1(n3012), .A2(n2882), .B1(n3010), .B2(n2902), .ZN(
        n2883) );
  AO21D1BWP12T U3231 ( .A1(write1_in[11]), .A2(n3231), .B(n2883), .Z(n2595) );
  OAI22D1BWP12T U3232 ( .A1(n3004), .A2(n2884), .B1(n3002), .B2(n2902), .ZN(
        n2885) );
  AO21D1BWP12T U3233 ( .A1(write1_in[11]), .A2(n3254), .B(n2885), .Z(n2467) );
  OAI22D1BWP12T U3234 ( .A1(n2968), .A2(n2888), .B1(n2970), .B2(n2902), .ZN(
        n2889) );
  AO21D1BWP12T U3235 ( .A1(write1_in[11]), .A2(n3515), .B(n2889), .Z(n2531) );
  CKND0BWP12T U3236 ( .I(r4[11]), .ZN(n2890) );
  OAI22D1BWP12T U3237 ( .A1(n2952), .A2(n2890), .B1(n2954), .B2(n2902), .ZN(
        n2891) );
  AO21D1BWP12T U3238 ( .A1(write1_in[11]), .A2(n3518), .B(n2891), .Z(n2499) );
  OAI22D1BWP12T U3239 ( .A1(n2966), .A2(n2902), .B1(n2964), .B2(n3026), .ZN(
        n2892) );
  AO21D1BWP12T U3240 ( .A1(write1_in[11]), .A2(n3522), .B(n2892), .Z(n2275) );
  OAI22D1BWP12T U3241 ( .A1(n2980), .A2(n2893), .B1(n2982), .B2(n2902), .ZN(
        n2894) );
  AO21D1BWP12T U3242 ( .A1(write1_in[11]), .A2(n3517), .B(n2894), .Z(n2627) );
  OAI22D1BWP12T U3243 ( .A1(n2960), .A2(n3025), .B1(n2962), .B2(n2902), .ZN(
        n2895) );
  AO21D1BWP12T U3244 ( .A1(write1_in[11]), .A2(n3519), .B(n2895), .Z(n2371) );
  OAI22D1BWP12T U3245 ( .A1(n2972), .A2(n2896), .B1(n2974), .B2(n2902), .ZN(
        n2897) );
  AO21D1BWP12T U3246 ( .A1(write1_in[11]), .A2(n3516), .B(n2897), .Z(n2563) );
  OAI22D1BWP12T U3247 ( .A1(n2956), .A2(n2898), .B1(n2958), .B2(n2902), .ZN(
        n2899) );
  AO21D1BWP12T U3248 ( .A1(write1_in[11]), .A2(n3521), .B(n2899), .Z(n2243) );
  OAI22D1BWP12T U3249 ( .A1(n2976), .A2(n2900), .B1(n2978), .B2(n2902), .ZN(
        n2901) );
  AO21D1BWP12T U3250 ( .A1(write1_in[11]), .A2(n3520), .B(n2901), .Z(n2307) );
  INVD0BWP12T U3251 ( .I(n3185), .ZN(n2993) );
  AO222D1BWP12T U3252 ( .A1(n3246), .A2(write1_in[10]), .B1(n1947), .B2(
        write2_in[10]), .C1(n1946), .C2(tmp1[10]), .Z(n2146) );
  OAI222D1BWP12T U3253 ( .A1(n2933), .A2(n2954), .B1(n2934), .B2(n2953), .C1(
        n2952), .C2(n2903), .ZN(n2496) );
  OAI222D1BWP12T U3254 ( .A1(n2933), .A2(n2982), .B1(n2934), .B2(n2981), .C1(
        n2980), .C2(n2904), .ZN(n2624) );
  OAI222D1BWP12T U3255 ( .A1(n2933), .A2(n2962), .B1(n2934), .B2(n2961), .C1(
        n2960), .C2(n2905), .ZN(n2368) );
  OAI222D1BWP12T U3256 ( .A1(n2933), .A2(n2958), .B1(n2934), .B2(n2957), .C1(
        n2956), .C2(n2906), .ZN(n2240) );
  OAI222D1BWP12T U3257 ( .A1(n2933), .A2(n2966), .B1(n2934), .B2(n2965), .C1(
        n2964), .C2(n2907), .ZN(n2272) );
  OAI222D1BWP12T U3258 ( .A1(n2933), .A2(n2978), .B1(n2934), .B2(n2977), .C1(
        n2976), .C2(n2995), .ZN(n2304) );
  OAI222D1BWP12T U3259 ( .A1(n2933), .A2(n2974), .B1(n2934), .B2(n2973), .C1(
        n2972), .C2(n2908), .ZN(n2560) );
  OAI222D1BWP12T U3260 ( .A1(n2933), .A2(n2970), .B1(n2934), .B2(n2969), .C1(
        n2968), .C2(n2909), .ZN(n2528) );
  TPND2D0BWP12T U3261 ( .A1(write1_in[13]), .A2(n3274), .ZN(n2911) );
  AOI22D0BWP12T U3262 ( .A1(n3277), .A2(r6[13]), .B1(n3276), .B2(write2_in[13]), .ZN(n2910) );
  ND2D1BWP12T U3263 ( .A1(n2911), .A2(n2910), .ZN(n2437) );
  TPND2D0BWP12T U3264 ( .A1(write1_in[13]), .A2(n3259), .ZN(n2913) );
  AOI22D0BWP12T U3265 ( .A1(n3261), .A2(lr[13]), .B1(n3260), .B2(write2_in[13]), .ZN(n2912) );
  ND2D1BWP12T U3266 ( .A1(n2913), .A2(n2912), .ZN(n2213) );
  TPND2D0BWP12T U3267 ( .A1(write1_in[13]), .A2(n3264), .ZN(n2915) );
  AOI22D0BWP12T U3268 ( .A1(n3266), .A2(r7[13]), .B1(n3265), .B2(write2_in[13]), .ZN(n2914) );
  ND2D1BWP12T U3269 ( .A1(n2915), .A2(n2914), .ZN(n2405) );
  TPND2D0BWP12T U3270 ( .A1(write1_in[13]), .A2(n3254), .ZN(n2917) );
  AOI22D0BWP12T U3271 ( .A1(n3256), .A2(r5[13]), .B1(n3255), .B2(write2_in[13]), .ZN(n2916) );
  ND2D1BWP12T U3272 ( .A1(n2917), .A2(n2916), .ZN(n2469) );
  TPND2D0BWP12T U3273 ( .A1(write1_in[13]), .A2(n3269), .ZN(n2919) );
  AOI22D0BWP12T U3274 ( .A1(n3271), .A2(r9[13]), .B1(n3270), .B2(write2_in[13]), .ZN(n2918) );
  ND2D1BWP12T U3275 ( .A1(n2919), .A2(n2918), .ZN(n2341) );
  TPND2D0BWP12T U3276 ( .A1(write1_in[13]), .A2(n3519), .ZN(n2922) );
  AOI22D0BWP12T U3277 ( .A1(n3215), .A2(r8[13]), .B1(n3214), .B2(write2_in[13]), .ZN(n2921) );
  ND2D1BWP12T U3278 ( .A1(n2922), .A2(n2921), .ZN(n2373) );
  TPND2D0BWP12T U3279 ( .A1(write1_in[13]), .A2(n3521), .ZN(n2924) );
  AOI22D0BWP12T U3280 ( .A1(n3228), .A2(r12[13]), .B1(n3227), .B2(
        write2_in[13]), .ZN(n2923) );
  ND2D1BWP12T U3281 ( .A1(n2924), .A2(n2923), .ZN(n2245) );
  TPND2D0BWP12T U3282 ( .A1(write1_in[13]), .A2(n3522), .ZN(n2926) );
  AOI22D0BWP12T U3283 ( .A1(n3202), .A2(write2_in[13]), .B1(n3201), .B2(
        r11[13]), .ZN(n2925) );
  ND2D1BWP12T U3284 ( .A1(n2926), .A2(n2925), .ZN(n2277) );
  TPND2D0BWP12T U3285 ( .A1(write1_in[13]), .A2(n3184), .ZN(n2928) );
  AOI22D0BWP12T U3286 ( .A1(n3186), .A2(n[3567]), .B1(n3185), .B2(
        write2_in[13]), .ZN(n2927) );
  ND2D1BWP12T U3287 ( .A1(n2928), .A2(n2927), .ZN(spin[13]) );
  OAI222D1BWP12T U3288 ( .A1(n2929), .A2(n3004), .B1(n2934), .B2(n3003), .C1(
        n2933), .C2(n3002), .ZN(n2464) );
  INVD0BWP12T U3289 ( .I(r6[8]), .ZN(n2930) );
  OAI222D1BWP12T U3290 ( .A1(n2930), .A2(n3008), .B1(n2934), .B2(n3007), .C1(
        n2933), .C2(n3006), .ZN(n2432) );
  OAI222D1BWP12T U3291 ( .A1(n2931), .A2(n3000), .B1(n2934), .B2(n2999), .C1(
        n2933), .C2(n2998), .ZN(n2400) );
  OAI222D1BWP12T U3292 ( .A1(n2932), .A2(n3012), .B1(n2934), .B2(n3011), .C1(
        n2933), .C2(n3010), .ZN(n2592) );
  OAI222D1BWP12T U3293 ( .A1(n2996), .A2(n3022), .B1(n2934), .B2(n3020), .C1(
        n2933), .C2(n3018), .ZN(n2208) );
  OAI222D1BWP12T U3294 ( .A1(n2935), .A2(n3016), .B1(n2934), .B2(n3015), .C1(
        n2933), .C2(n3014), .ZN(n2336) );
  TPND2D0BWP12T U3295 ( .A1(write1_in[13]), .A2(n3246), .ZN(n2937) );
  AOI22D0BWP12T U3296 ( .A1(n1946), .A2(tmp1[13]), .B1(n1947), .B2(
        write2_in[13]), .ZN(n2936) );
  ND2D1BWP12T U3297 ( .A1(n2937), .A2(n2936), .ZN(n2149) );
  NR2D1BWP12T U3298 ( .A1(n2950), .A2(n2949), .ZN(n2939) );
  XNR2D1BWP12T U3299 ( .A1(n2939), .A2(n2938), .ZN(n2940) );
  AO222D1BWP12T U3300 ( .A1(n2940), .A2(n3505), .B1(n3498), .B2(pc_out[4]), 
        .C1(n3499), .C2(next_pc_in[4]), .Z(n2172) );
  OAI222D1BWP12T U3301 ( .A1(n2988), .A2(n2978), .B1(n2989), .B2(n2977), .C1(
        n2976), .C2(n2941), .ZN(n2305) );
  OAI222D1BWP12T U3302 ( .A1(n2988), .A2(n2962), .B1(n2989), .B2(n2961), .C1(
        n2960), .C2(n2942), .ZN(n2369) );
  OAI222D1BWP12T U3303 ( .A1(n2988), .A2(n2974), .B1(n2989), .B2(n2973), .C1(
        n2972), .C2(n2943), .ZN(n2561) );
  OAI222D1BWP12T U3304 ( .A1(n2988), .A2(n2954), .B1(n2989), .B2(n2953), .C1(
        n2952), .C2(n2944), .ZN(n2497) );
  OAI222D1BWP12T U3305 ( .A1(n2988), .A2(n2982), .B1(n2989), .B2(n2981), .C1(
        n2980), .C2(n2945), .ZN(n2625) );
  OAI222D1BWP12T U3306 ( .A1(n2988), .A2(n2970), .B1(n2989), .B2(n2969), .C1(
        n2968), .C2(n2946), .ZN(n2529) );
  OAI222D1BWP12T U3307 ( .A1(n2988), .A2(n2966), .B1(n2989), .B2(n2965), .C1(
        n2964), .C2(n2947), .ZN(n2273) );
  OAI222D1BWP12T U3308 ( .A1(n2988), .A2(n2958), .B1(n2989), .B2(n2957), .C1(
        n2956), .C2(n2948), .ZN(n2241) );
  OAI222D1BWP12T U3309 ( .A1(n3019), .A2(n2954), .B1(n3021), .B2(n2953), .C1(
        n2952), .C2(n2951), .ZN(n2498) );
  OAI222D1BWP12T U3310 ( .A1(n3019), .A2(n2958), .B1(n3021), .B2(n2957), .C1(
        n2956), .C2(n2955), .ZN(n2242) );
  OAI222D1BWP12T U3311 ( .A1(n3019), .A2(n2962), .B1(n3021), .B2(n2961), .C1(
        n2960), .C2(n2959), .ZN(n2370) );
  OAI222D1BWP12T U3312 ( .A1(n3019), .A2(n2966), .B1(n3021), .B2(n2965), .C1(
        n2964), .C2(n2963), .ZN(n2274) );
  OAI222D1BWP12T U3313 ( .A1(n3019), .A2(n2970), .B1(n3021), .B2(n2969), .C1(
        n2968), .C2(n2967), .ZN(n2530) );
  OAI222D1BWP12T U3314 ( .A1(n3019), .A2(n2974), .B1(n3021), .B2(n2973), .C1(
        n2972), .C2(n2971), .ZN(n2562) );
  OAI222D1BWP12T U3315 ( .A1(n3019), .A2(n2978), .B1(n3021), .B2(n2977), .C1(
        n2976), .C2(n2975), .ZN(n2306) );
  OAI222D1BWP12T U3316 ( .A1(n3019), .A2(n2982), .B1(n3021), .B2(n2981), .C1(
        n2980), .C2(n2979), .ZN(n2626) );
  OAI222D1BWP12T U3317 ( .A1(n2983), .A2(n3012), .B1(n2989), .B2(n3011), .C1(
        n2988), .C2(n3010), .ZN(n2593) );
  OAI222D1BWP12T U3318 ( .A1(n2984), .A2(n3016), .B1(n2989), .B2(n3015), .C1(
        n2988), .C2(n3014), .ZN(n2337) );
  INVD0BWP12T U3319 ( .I(r6[9]), .ZN(n2985) );
  OAI222D1BWP12T U3320 ( .A1(n2985), .A2(n3008), .B1(n2989), .B2(n3007), .C1(
        n2988), .C2(n3006), .ZN(n2433) );
  OAI222D1BWP12T U3321 ( .A1(n2986), .A2(n3000), .B1(n2989), .B2(n2999), .C1(
        n2988), .C2(n2998), .ZN(n2401) );
  OAI222D1BWP12T U3322 ( .A1(n2987), .A2(n3004), .B1(n2989), .B2(n3003), .C1(
        n2988), .C2(n3002), .ZN(n2465) );
  OAI222D1BWP12T U3323 ( .A1(n2990), .A2(n3022), .B1(n2989), .B2(n3020), .C1(
        n2988), .C2(n3018), .ZN(n2209) );
  TPND2D0BWP12T U3324 ( .A1(write1_in[13]), .A2(n3520), .ZN(n2992) );
  AOI22D0BWP12T U3325 ( .A1(n3198), .A2(r10[13]), .B1(n3197), .B2(
        write2_in[13]), .ZN(n2991) );
  ND2D1BWP12T U3326 ( .A1(n2992), .A2(n2991), .ZN(n2309) );
  OAI222D1BWP12T U3327 ( .A1(n3001), .A2(n3000), .B1(n3021), .B2(n2999), .C1(
        n3019), .C2(n2998), .ZN(n2402) );
  OAI222D1BWP12T U3328 ( .A1(n3005), .A2(n3004), .B1(n3021), .B2(n3003), .C1(
        n3019), .C2(n3002), .ZN(n2466) );
  INVD1BWP12T U3329 ( .I(r6[10]), .ZN(n3009) );
  OAI222D1BWP12T U3330 ( .A1(n3009), .A2(n3008), .B1(n3021), .B2(n3007), .C1(
        n3019), .C2(n3006), .ZN(n2434) );
  OAI222D1BWP12T U3331 ( .A1(n3013), .A2(n3012), .B1(n3021), .B2(n3011), .C1(
        n3019), .C2(n3010), .ZN(n2594) );
  OAI222D1BWP12T U3332 ( .A1(n3017), .A2(n3016), .B1(n3021), .B2(n3015), .C1(
        n3019), .C2(n3014), .ZN(n2338) );
  OAI222D1BWP12T U3333 ( .A1(n3023), .A2(n3022), .B1(n3021), .B2(n3020), .C1(
        n3019), .C2(n3018), .ZN(n2210) );
  AOI22D0BWP12T U3334 ( .A1(r5[12]), .A2(n3075), .B1(n3074), .B2(r1[12]), .ZN(
        n3036) );
  AOI22D0BWP12T U3335 ( .A1(r0[12]), .A2(n3081), .B1(n3080), .B2(r4[12]), .ZN(
        n3035) );
  AOI22D0BWP12T U3336 ( .A1(r6[12]), .A2(n3077), .B1(n3076), .B2(r7[12]), .ZN(
        n3034) );
  AOI22D0BWP12T U3337 ( .A1(r2[12]), .A2(n3079), .B1(n3078), .B2(r3[12]), .ZN(
        n3033) );
  AN4XD1BWP12T U3338 ( .A1(n3036), .A2(n3035), .A3(n3034), .A4(n3033), .Z(
        n3047) );
  AOI22D0BWP12T U3339 ( .A1(n[3568]), .A2(n3037), .B1(n3064), .B2(r12[12]), 
        .ZN(n3046) );
  NR2D0BWP12T U3340 ( .A1(n3066), .A2(n3038), .ZN(n3044) );
  CKND2D0BWP12T U3341 ( .A1(pc_out[12]), .A2(n3061), .ZN(n3040) );
  AOI22D0BWP12T U3342 ( .A1(r9[12]), .A2(n3063), .B1(r11[12]), .B2(n2994), 
        .ZN(n3039) );
  OAI211D0BWP12T U3343 ( .A1(n3042), .A2(n3041), .B(n3040), .C(n3039), .ZN(
        n3043) );
  AOI211D0BWP12T U3344 ( .A1(n3073), .A2(r8[12]), .B(n3044), .C(n3043), .ZN(
        n3045) );
  OAI211D1BWP12T U3345 ( .A1(n3047), .A2(readD_sel[4]), .B(n3046), .C(n3045), 
        .ZN(regD_out[12]) );
  XNR2XD0BWP12T U3346 ( .A1(n3058), .A2(n3059), .ZN(n3049) );
  AOI22D1BWP12T U3347 ( .A1(next_pc_in[8]), .A2(n3499), .B1(n3498), .B2(
        pc_out[8]), .ZN(n3048) );
  OAI21D1BWP12T U3348 ( .A1(n3049), .A2(n3497), .B(n3048), .ZN(n2176) );
  INVD1BWP12T U3349 ( .I(write1_in[16]), .ZN(n3050) );
  CKXOR2D1BWP12T U3350 ( .A1(n3052), .A2(n3051), .Z(n3053) );
  AO222D1BWP12T U3351 ( .A1(n3053), .A2(n3505), .B1(n3498), .B2(pc_out[7]), 
        .C1(n3499), .C2(next_pc_in[7]), .Z(n2175) );
  AOI22D0BWP12T U3352 ( .A1(lr[0]), .A2(n3062), .B1(n3061), .B2(pc_out[0]), 
        .ZN(n3091) );
  AOI22D0BWP12T U3353 ( .A1(r12[0]), .A2(n3064), .B1(n3063), .B2(r9[0]), .ZN(
        n3090) );
  NR2D0BWP12T U3354 ( .A1(n3066), .A2(n3065), .ZN(n3072) );
  OAI22D0BWP12T U3355 ( .A1(n3070), .A2(n3069), .B1(n3068), .B2(n3067), .ZN(
        n3071) );
  RCAOI211D0BWP12T U3356 ( .A1(n3073), .A2(r8[0]), .B(n3072), .C(n3071), .ZN(
        n3089) );
  AOI22D0BWP12T U3357 ( .A1(r5[0]), .A2(n3075), .B1(n3074), .B2(r1[0]), .ZN(
        n3085) );
  AOI22D0BWP12T U3358 ( .A1(r6[0]), .A2(n3077), .B1(n3076), .B2(r7[0]), .ZN(
        n3084) );
  AOI22D0BWP12T U3359 ( .A1(r2[0]), .A2(n3079), .B1(n3078), .B2(r3[0]), .ZN(
        n3083) );
  AOI22D0BWP12T U3360 ( .A1(r0[0]), .A2(n3081), .B1(n3080), .B2(r4[0]), .ZN(
        n3082) );
  ND4D1BWP12T U3361 ( .A1(n3085), .A2(n3084), .A3(n3083), .A4(n3082), .ZN(
        n3087) );
  CKND2D1BWP12T U3362 ( .A1(n3087), .A2(n3086), .ZN(n3088) );
  ND4D1BWP12T U3363 ( .A1(n3091), .A2(n3090), .A3(n3089), .A4(n3088), .ZN(
        regD_out[0]) );
  CKBD1BWP12T U3364 ( .I(write1_in[20]), .Z(n3095) );
  BUFFD2BWP12T U3365 ( .I(write1_in[24]), .Z(n3097) );
  BUFFXD4BWP12T U3366 ( .I(write1_in[22]), .Z(n3282) );
  BUFFD2BWP12T U3367 ( .I(n3282), .Z(n3099) );
  BUFFXD12BWP12T U3368 ( .I(write1_in[26]), .Z(n3108) );
  INVD1BWP12T U3369 ( .I(n3100), .ZN(n3101) );
  ND2D1BWP12T U3370 ( .A1(n3102), .A2(n3101), .ZN(n3104) );
  XOR2XD1BWP12T U3371 ( .A1(n3104), .A2(n3103), .Z(n3106) );
  AOI22D1BWP12T U3372 ( .A1(next_pc_in[12]), .A2(n3499), .B1(n3498), .B2(
        pc_out[12]), .ZN(n3105) );
  OAI21D1BWP12T U3373 ( .A1(n3106), .A2(n3497), .B(n3105), .ZN(n2180) );
  INVD1BWP12T U3374 ( .I(n3107), .ZN(n3109) );
  NR2D1BWP12T U3375 ( .A1(n3110), .A2(n3109), .ZN(n3112) );
  BUFFXD4BWP12T U3376 ( .I(write1_in[25]), .Z(n3113) );
  CKND2D1BWP12T U3377 ( .A1(n3150), .A2(n3231), .ZN(n3115) );
  AOI22D0BWP12T U3378 ( .A1(n3233), .A2(r1[27]), .B1(write2_in[27]), .B2(n3232), .ZN(n3114) );
  ND2D1BWP12T U3379 ( .A1(n3115), .A2(n3114), .ZN(n2611) );
  CKND2D1BWP12T U3380 ( .A1(n3150), .A2(n3264), .ZN(n3117) );
  AOI22D0BWP12T U3381 ( .A1(n3266), .A2(r7[27]), .B1(write2_in[27]), .B2(n3265), .ZN(n3116) );
  ND2D1BWP12T U3382 ( .A1(n3117), .A2(n3116), .ZN(n2419) );
  CKND2D1BWP12T U3383 ( .A1(n3150), .A2(n3259), .ZN(n3119) );
  AOI22D0BWP12T U3384 ( .A1(n3261), .A2(lr[27]), .B1(write2_in[27]), .B2(n3260), .ZN(n3118) );
  ND2D1BWP12T U3385 ( .A1(n3119), .A2(n3118), .ZN(n2227) );
  CKND2D1BWP12T U3386 ( .A1(n3150), .A2(n3274), .ZN(n3121) );
  AOI22D0BWP12T U3387 ( .A1(n3277), .A2(r6[27]), .B1(write2_in[27]), .B2(n3276), .ZN(n3120) );
  ND2D1BWP12T U3388 ( .A1(n3121), .A2(n3120), .ZN(n2451) );
  CKND2D1BWP12T U3389 ( .A1(n3150), .A2(n3254), .ZN(n3123) );
  AOI22D0BWP12T U3390 ( .A1(n3256), .A2(r5[27]), .B1(write2_in[27]), .B2(n3255), .ZN(n3122) );
  ND2D1BWP12T U3391 ( .A1(n3123), .A2(n3122), .ZN(n2483) );
  CKND2D1BWP12T U3392 ( .A1(n3150), .A2(n3269), .ZN(n3125) );
  AOI22D0BWP12T U3393 ( .A1(n3271), .A2(r9[27]), .B1(write2_in[27]), .B2(n3270), .ZN(n3124) );
  ND2D1BWP12T U3394 ( .A1(n3125), .A2(n3124), .ZN(n2355) );
  CKND2D1BWP12T U3395 ( .A1(n3150), .A2(n3246), .ZN(n3127) );
  AOI22D0BWP12T U3396 ( .A1(write2_in[27]), .A2(n1947), .B1(n1946), .B2(
        tmp1[27]), .ZN(n3126) );
  ND2D1BWP12T U3397 ( .A1(n3127), .A2(n3126), .ZN(n2163) );
  CKND2D1BWP12T U3398 ( .A1(n3150), .A2(n3184), .ZN(n3129) );
  AOI22D0BWP12T U3399 ( .A1(n3186), .A2(n[3553]), .B1(write2_in[27]), .B2(
        n3185), .ZN(n3128) );
  ND2D1BWP12T U3400 ( .A1(n3129), .A2(n3128), .ZN(spin[27]) );
  CKND2D1BWP12T U3401 ( .A1(n3150), .A2(n3515), .ZN(n3131) );
  AOI22D0BWP12T U3402 ( .A1(n3190), .A2(r3[27]), .B1(n3189), .B2(write2_in[27]), .ZN(n3130) );
  ND2D1BWP12T U3403 ( .A1(n3131), .A2(n3130), .ZN(n2547) );
  CKND2D1BWP12T U3404 ( .A1(n3150), .A2(n3516), .ZN(n3133) );
  AOI22D0BWP12T U3405 ( .A1(n3194), .A2(r2[27]), .B1(n3193), .B2(write2_in[27]), .ZN(n3132) );
  ND2D1BWP12T U3406 ( .A1(n3133), .A2(n3132), .ZN(n2579) );
  CKND2D1BWP12T U3407 ( .A1(n3150), .A2(n3520), .ZN(n3135) );
  AOI22D0BWP12T U3408 ( .A1(n3198), .A2(r10[27]), .B1(n3197), .B2(
        write2_in[27]), .ZN(n3134) );
  ND2D1BWP12T U3409 ( .A1(n3135), .A2(n3134), .ZN(n2323) );
  ND2D1BWP12T U3410 ( .A1(n3137), .A2(n3136), .ZN(n3139) );
  XNR2D1BWP12T U3411 ( .A1(n3139), .A2(n157), .ZN(n3141) );
  AOI22D1BWP12T U3412 ( .A1(next_pc_in[16]), .A2(n3499), .B1(n3498), .B2(
        pc_out[16]), .ZN(n3140) );
  OAI21D1BWP12T U3413 ( .A1(n3141), .A2(n3497), .B(n3140), .ZN(n2184) );
  CKND2D1BWP12T U3414 ( .A1(n3150), .A2(n3522), .ZN(n3143) );
  AOI22D0BWP12T U3415 ( .A1(write2_in[27]), .A2(n3202), .B1(n3201), .B2(
        r11[27]), .ZN(n3142) );
  ND2D1BWP12T U3416 ( .A1(n3143), .A2(n3142), .ZN(n2291) );
  CKND2D1BWP12T U3417 ( .A1(n3150), .A2(n3519), .ZN(n3145) );
  AOI22D0BWP12T U3418 ( .A1(n3215), .A2(r8[27]), .B1(write2_in[27]), .B2(n3214), .ZN(n3144) );
  ND2D1BWP12T U3419 ( .A1(n3145), .A2(n3144), .ZN(n2387) );
  CKND2D1BWP12T U3420 ( .A1(n3150), .A2(n3517), .ZN(n3147) );
  AOI22D0BWP12T U3421 ( .A1(n3219), .A2(r0[27]), .B1(write2_in[27]), .B2(n3218), .ZN(n3146) );
  ND2D1BWP12T U3422 ( .A1(n3147), .A2(n3146), .ZN(n2643) );
  CKND2D1BWP12T U3423 ( .A1(n3150), .A2(n3518), .ZN(n3149) );
  AOI22D0BWP12T U3424 ( .A1(n3223), .A2(r4[27]), .B1(write2_in[27]), .B2(n3222), .ZN(n3148) );
  ND2D1BWP12T U3425 ( .A1(n3149), .A2(n3148), .ZN(n2515) );
  CKND2D1BWP12T U3426 ( .A1(n3150), .A2(n3521), .ZN(n3152) );
  AOI22D0BWP12T U3427 ( .A1(n3228), .A2(r12[27]), .B1(write2_in[27]), .B2(
        n3227), .ZN(n3151) );
  ND2D1BWP12T U3428 ( .A1(n3152), .A2(n3151), .ZN(n2259) );
  CKND2D1BWP12T U3429 ( .A1(n3211), .A2(n3231), .ZN(n3155) );
  AOI22D0BWP12T U3430 ( .A1(n3233), .A2(r1[28]), .B1(write2_in[28]), .B2(n3232), .ZN(n3154) );
  ND2D1BWP12T U3431 ( .A1(n3155), .A2(n3154), .ZN(n2612) );
  CKND2D1BWP12T U3432 ( .A1(n3211), .A2(n3254), .ZN(n3157) );
  AOI22D0BWP12T U3433 ( .A1(n3256), .A2(r5[28]), .B1(write2_in[28]), .B2(n3255), .ZN(n3156) );
  ND2D1BWP12T U3434 ( .A1(n3157), .A2(n3156), .ZN(n2484) );
  CKND2D1BWP12T U3435 ( .A1(n3211), .A2(n3264), .ZN(n3159) );
  AOI22D0BWP12T U3436 ( .A1(n3266), .A2(r7[28]), .B1(write2_in[28]), .B2(n3265), .ZN(n3158) );
  ND2D1BWP12T U3437 ( .A1(n3159), .A2(n3158), .ZN(n2420) );
  CKND2D1BWP12T U3438 ( .A1(n3211), .A2(n3274), .ZN(n3161) );
  AOI22D0BWP12T U3439 ( .A1(n3277), .A2(r6[28]), .B1(write2_in[28]), .B2(n3276), .ZN(n3160) );
  ND2D1BWP12T U3440 ( .A1(n3161), .A2(n3160), .ZN(n2452) );
  CKND2D1BWP12T U3441 ( .A1(n3211), .A2(n3259), .ZN(n3163) );
  AOI22D0BWP12T U3442 ( .A1(n3261), .A2(lr[28]), .B1(write2_in[28]), .B2(n3260), .ZN(n3162) );
  ND2D1BWP12T U3443 ( .A1(n3163), .A2(n3162), .ZN(n2228) );
  CKND2D1BWP12T U3444 ( .A1(n3211), .A2(n3269), .ZN(n3165) );
  AOI22D0BWP12T U3445 ( .A1(n3271), .A2(r9[28]), .B1(write2_in[28]), .B2(n3270), .ZN(n3164) );
  ND2D1BWP12T U3446 ( .A1(n3165), .A2(n3164), .ZN(n2356) );
  ND2D1BWP12T U3447 ( .A1(n3226), .A2(n3231), .ZN(n3167) );
  AOI22D0BWP12T U3448 ( .A1(n3233), .A2(r1[30]), .B1(write2_in[30]), .B2(n3232), .ZN(n3166) );
  ND2D1BWP12T U3449 ( .A1(n3167), .A2(n3166), .ZN(n2614) );
  ND2D1BWP12T U3450 ( .A1(n3226), .A2(n3264), .ZN(n3169) );
  AOI22D0BWP12T U3451 ( .A1(n3266), .A2(r7[30]), .B1(write2_in[30]), .B2(n3265), .ZN(n3168) );
  ND2D1BWP12T U3452 ( .A1(n3169), .A2(n3168), .ZN(n2422) );
  ND2D1BWP12T U3453 ( .A1(n3226), .A2(n3254), .ZN(n3171) );
  AOI22D0BWP12T U3454 ( .A1(n3256), .A2(r5[30]), .B1(write2_in[30]), .B2(n3255), .ZN(n3170) );
  ND2D1BWP12T U3455 ( .A1(n3171), .A2(n3170), .ZN(n2486) );
  ND2D1BWP12T U3456 ( .A1(n3226), .A2(n3274), .ZN(n3173) );
  AOI22D0BWP12T U3457 ( .A1(n3277), .A2(r6[30]), .B1(write2_in[30]), .B2(n3276), .ZN(n3172) );
  ND2D1BWP12T U3458 ( .A1(n3173), .A2(n3172), .ZN(n2454) );
  ND2D1BWP12T U3459 ( .A1(n3226), .A2(n3259), .ZN(n3175) );
  AOI22D0BWP12T U3460 ( .A1(n3261), .A2(lr[30]), .B1(write2_in[30]), .B2(n3260), .ZN(n3174) );
  ND2D1BWP12T U3461 ( .A1(n3175), .A2(n3174), .ZN(n2230) );
  ND2D1BWP12T U3462 ( .A1(n3226), .A2(n3269), .ZN(n3177) );
  AOI22D0BWP12T U3463 ( .A1(n3271), .A2(r9[30]), .B1(write2_in[30]), .B2(n3270), .ZN(n3176) );
  ND2D1BWP12T U3464 ( .A1(n3177), .A2(n3176), .ZN(n2358) );
  CKND2D1BWP12T U3465 ( .A1(n3211), .A2(n3246), .ZN(n3179) );
  AOI22D0BWP12T U3466 ( .A1(write2_in[28]), .A2(n1947), .B1(n1946), .B2(
        tmp1[28]), .ZN(n3178) );
  ND2D1BWP12T U3467 ( .A1(n3179), .A2(n3178), .ZN(n2164) );
  ND2D1BWP12T U3468 ( .A1(n3226), .A2(n3246), .ZN(n3181) );
  AOI22D0BWP12T U3469 ( .A1(write2_in[30]), .A2(n1947), .B1(n1946), .B2(
        tmp1[30]), .ZN(n3180) );
  ND2D1BWP12T U3470 ( .A1(n3181), .A2(n3180), .ZN(n2166) );
  CKND2D1BWP12T U3471 ( .A1(n3211), .A2(n3184), .ZN(n3183) );
  AOI22D0BWP12T U3472 ( .A1(n3186), .A2(n[3552]), .B1(write2_in[28]), .B2(
        n3185), .ZN(n3182) );
  ND2D1BWP12T U3473 ( .A1(n3183), .A2(n3182), .ZN(spin[28]) );
  ND2D1BWP12T U3474 ( .A1(n3226), .A2(n3184), .ZN(n3188) );
  AOI22D0BWP12T U3475 ( .A1(n3186), .A2(n[3550]), .B1(write2_in[30]), .B2(
        n3185), .ZN(n3187) );
  ND2D1BWP12T U3476 ( .A1(n3188), .A2(n3187), .ZN(spin[30]) );
  CKND2D1BWP12T U3477 ( .A1(n3211), .A2(n3515), .ZN(n3192) );
  AOI22D0BWP12T U3478 ( .A1(n3190), .A2(r3[28]), .B1(n3189), .B2(write2_in[28]), .ZN(n3191) );
  ND2D1BWP12T U3479 ( .A1(n3192), .A2(n3191), .ZN(n2548) );
  CKND2D1BWP12T U3480 ( .A1(n3211), .A2(n3516), .ZN(n3196) );
  AOI22D0BWP12T U3481 ( .A1(n3194), .A2(r2[28]), .B1(n3193), .B2(write2_in[28]), .ZN(n3195) );
  ND2D1BWP12T U3482 ( .A1(n3196), .A2(n3195), .ZN(n2580) );
  CKND2D1BWP12T U3483 ( .A1(n3211), .A2(n3520), .ZN(n3200) );
  AOI22D0BWP12T U3484 ( .A1(n3198), .A2(r10[28]), .B1(n3197), .B2(
        write2_in[28]), .ZN(n3199) );
  ND2D1BWP12T U3485 ( .A1(n3200), .A2(n3199), .ZN(n2324) );
  CKND2D1BWP12T U3486 ( .A1(n3211), .A2(n3522), .ZN(n3204) );
  AOI22D0BWP12T U3487 ( .A1(write2_in[28]), .A2(n3202), .B1(n3201), .B2(
        r11[28]), .ZN(n3203) );
  ND2D1BWP12T U3488 ( .A1(n3204), .A2(n3203), .ZN(n2292) );
  CKND2D1BWP12T U3489 ( .A1(n3211), .A2(n3517), .ZN(n3206) );
  AOI22D0BWP12T U3490 ( .A1(n3219), .A2(r0[28]), .B1(write2_in[28]), .B2(n3218), .ZN(n3205) );
  ND2D1BWP12T U3491 ( .A1(n3206), .A2(n3205), .ZN(n2644) );
  CKND2D1BWP12T U3492 ( .A1(n3211), .A2(n3519), .ZN(n3208) );
  AOI22D0BWP12T U3493 ( .A1(n3215), .A2(r8[28]), .B1(write2_in[28]), .B2(n3214), .ZN(n3207) );
  ND2D1BWP12T U3494 ( .A1(n3208), .A2(n3207), .ZN(n2388) );
  CKND2D1BWP12T U3495 ( .A1(n3211), .A2(n3518), .ZN(n3210) );
  AOI22D0BWP12T U3496 ( .A1(n3223), .A2(r4[28]), .B1(write2_in[28]), .B2(n3222), .ZN(n3209) );
  ND2D1BWP12T U3497 ( .A1(n3210), .A2(n3209), .ZN(n2516) );
  CKND2D1BWP12T U3498 ( .A1(n3211), .A2(n3521), .ZN(n3213) );
  AOI22D0BWP12T U3499 ( .A1(n3228), .A2(r12[28]), .B1(write2_in[28]), .B2(
        n3227), .ZN(n3212) );
  ND2D1BWP12T U3500 ( .A1(n3213), .A2(n3212), .ZN(n2260) );
  ND2D1BWP12T U3501 ( .A1(n3226), .A2(n3519), .ZN(n3217) );
  AOI22D0BWP12T U3502 ( .A1(n3215), .A2(r8[30]), .B1(write2_in[30]), .B2(n3214), .ZN(n3216) );
  ND2D1BWP12T U3503 ( .A1(n3217), .A2(n3216), .ZN(n2390) );
  ND2D1BWP12T U3504 ( .A1(n3226), .A2(n3517), .ZN(n3221) );
  AOI22D0BWP12T U3505 ( .A1(n3219), .A2(r0[30]), .B1(write2_in[30]), .B2(n3218), .ZN(n3220) );
  ND2D1BWP12T U3506 ( .A1(n3221), .A2(n3220), .ZN(n2646) );
  AOI22D0BWP12T U3507 ( .A1(n3223), .A2(r4[30]), .B1(write2_in[30]), .B2(n3222), .ZN(n3224) );
  ND2D1BWP12T U3508 ( .A1(n3225), .A2(n3224), .ZN(n2518) );
  ND2D1BWP12T U3509 ( .A1(n3226), .A2(n3521), .ZN(n3230) );
  AOI22D0BWP12T U3510 ( .A1(n3228), .A2(r12[30]), .B1(write2_in[30]), .B2(
        n3227), .ZN(n3229) );
  ND2D1BWP12T U3511 ( .A1(n3230), .A2(n3229), .ZN(n2262) );
  AOI22D0BWP12T U3512 ( .A1(n3233), .A2(r1[29]), .B1(write2_in[29]), .B2(n3232), .ZN(n3234) );
  ND2D1BWP12T U3513 ( .A1(n3235), .A2(n3234), .ZN(n2613) );
  ND2D1BWP12T U3514 ( .A1(n3247), .A2(n3259), .ZN(n3237) );
  AOI22D0BWP12T U3515 ( .A1(n3261), .A2(lr[29]), .B1(write2_in[29]), .B2(n3260), .ZN(n3236) );
  ND2D1BWP12T U3516 ( .A1(n3237), .A2(n3236), .ZN(n2229) );
  ND2D1BWP12T U3517 ( .A1(n3247), .A2(n3254), .ZN(n3239) );
  AOI22D0BWP12T U3518 ( .A1(n3256), .A2(r5[29]), .B1(write2_in[29]), .B2(n3255), .ZN(n3238) );
  ND2D1BWP12T U3519 ( .A1(n3239), .A2(n3238), .ZN(n2485) );
  ND2D1BWP12T U3520 ( .A1(n3247), .A2(n3264), .ZN(n3241) );
  AOI22D0BWP12T U3521 ( .A1(n3266), .A2(r7[29]), .B1(write2_in[29]), .B2(n3265), .ZN(n3240) );
  ND2D1BWP12T U3522 ( .A1(n3241), .A2(n3240), .ZN(n2421) );
  CKND2D1BWP12T U3523 ( .A1(n3247), .A2(n3274), .ZN(n3243) );
  AOI22D0BWP12T U3524 ( .A1(n3277), .A2(r6[29]), .B1(write2_in[29]), .B2(n3276), .ZN(n3242) );
  ND2D1BWP12T U3525 ( .A1(n3243), .A2(n3242), .ZN(n2453) );
  ND2D1BWP12T U3526 ( .A1(n3247), .A2(n3269), .ZN(n3245) );
  AOI22D0BWP12T U3527 ( .A1(n3271), .A2(r9[29]), .B1(write2_in[29]), .B2(n3270), .ZN(n3244) );
  ND2D1BWP12T U3528 ( .A1(n3245), .A2(n3244), .ZN(n2357) );
  CKND2D1BWP12T U3529 ( .A1(n3247), .A2(n3246), .ZN(n3249) );
  AOI22D0BWP12T U3530 ( .A1(write2_in[29]), .A2(n1947), .B1(n1946), .B2(
        tmp1[29]), .ZN(n3248) );
  ND2D1BWP12T U3531 ( .A1(n3249), .A2(n3248), .ZN(n2165) );
  XNR2D1BWP12T U3532 ( .A1(n3251), .A2(n163), .ZN(n3253) );
  AOI22D1BWP12T U3533 ( .A1(next_pc_in[17]), .A2(n3499), .B1(n3498), .B2(
        pc_out[17]), .ZN(n3252) );
  OAI21D1BWP12T U3534 ( .A1(n3253), .A2(n3497), .B(n3252), .ZN(n2185) );
  AOI22D0BWP12T U3535 ( .A1(n3256), .A2(r5[31]), .B1(write2_in[31]), .B2(n3255), .ZN(n3257) );
  ND2D1BWP12T U3536 ( .A1(n3258), .A2(n3257), .ZN(n2487) );
  AOI22D0BWP12T U3537 ( .A1(n3261), .A2(lr[31]), .B1(write2_in[31]), .B2(n3260), .ZN(n3262) );
  ND2D1BWP12T U3538 ( .A1(n3263), .A2(n3262), .ZN(n2231) );
  AOI22D0BWP12T U3539 ( .A1(n3266), .A2(r7[31]), .B1(write2_in[31]), .B2(n3265), .ZN(n3267) );
  ND2D1BWP12T U3540 ( .A1(n3268), .A2(n3267), .ZN(n2423) );
  AOI22D0BWP12T U3541 ( .A1(n3271), .A2(r9[31]), .B1(write2_in[31]), .B2(n3270), .ZN(n3272) );
  ND2D1BWP12T U3542 ( .A1(n3273), .A2(n3272), .ZN(n2359) );
  AOI22D0BWP12T U3543 ( .A1(n3277), .A2(r6[31]), .B1(write2_in[31]), .B2(n3276), .ZN(n3278) );
  ND2D1BWP12T U3544 ( .A1(n3279), .A2(n3278), .ZN(n2455) );
  INVD1BWP12T U3545 ( .I(n3506), .ZN(n3280) );
  TPND2D1BWP12T U3546 ( .A1(n3502), .A2(n3280), .ZN(n3281) );
  NR2D1BWP12T U3547 ( .A1(n3281), .A2(n3504), .ZN(n3294) );
  CKND2BWP12T U3548 ( .I(n3282), .ZN(n3284) );
  CKND2D1BWP12T U3549 ( .A1(n3331), .A2(write2_in[22]), .ZN(n3283) );
  INVD1P75BWP12T U3550 ( .I(n3286), .ZN(n3285) );
  INVD1BWP12T U3551 ( .I(n3290), .ZN(n3293) );
  TPNR3D1BWP12T U3552 ( .A1(n171), .A2(n3289), .A3(n3497), .ZN(n3287) );
  TPND2D1BWP12T U3553 ( .A1(n3287), .A2(n3294), .ZN(n3292) );
  MOAI22D0BWP12T U3554 ( .A1(n3343), .A2(n3535), .B1(next_pc_in[22]), .B2(
        n3499), .ZN(n3288) );
  OAI211D1BWP12T U3555 ( .A1(n3294), .A2(n3293), .B(n3291), .C(n3292), .ZN(
        n2190) );
  CKND1BWP12T U3556 ( .I(n3299), .ZN(n3297) );
  MOAI22D0BWP12T U3557 ( .A1(n3343), .A2(n3295), .B1(next_pc_in[24]), .B2(
        n3499), .ZN(n3296) );
  AOI31D1BWP12T U3558 ( .A1(n3297), .A2(n3505), .A3(n3307), .B(n3296), .ZN(
        n3304) );
  IND2D1BWP12T U3559 ( .A1(n3301), .B1(n3298), .ZN(n3303) );
  ND4D1BWP12T U3560 ( .A1(n3301), .A2(n3300), .A3(n3505), .A4(n3299), .ZN(
        n3302) );
  ND3D1BWP12T U3561 ( .A1(n3304), .A2(n3303), .A3(n3302), .ZN(n2192) );
  INR3D0BWP12T U3562 ( .A1(n3307), .B1(n3497), .B2(n3311), .ZN(n3305) );
  INVD1BWP12T U3563 ( .I(n3305), .ZN(n3314) );
  INR2D1BWP12T U3564 ( .A1(n3311), .B1(n3497), .ZN(n3306) );
  TPND2D1BWP12T U3565 ( .A1(n3315), .A2(n3306), .ZN(n3313) );
  NR2D1BWP12T U3566 ( .A1(n3307), .A2(n3497), .ZN(n3310) );
  CKND2D0BWP12T U3567 ( .A1(next_pc_in[25]), .A2(n3499), .ZN(n3308) );
  OAI21D0BWP12T U3568 ( .A1(n3536), .A2(n3343), .B(n3308), .ZN(n3309) );
  AOI21D1BWP12T U3569 ( .A1(n3311), .A2(n3310), .B(n3309), .ZN(n3312) );
  OAI211D1BWP12T U3570 ( .A1(n3315), .A2(n3314), .B(n3313), .C(n3312), .ZN(
        n2193) );
  CKND0BWP12T U3571 ( .I(write2_in[31]), .ZN(n3316) );
  AOI21D0BWP12T U3572 ( .A1(n3331), .A2(n3316), .B(n3497), .ZN(n3317) );
  TPOAI21D1BWP12T U3573 ( .A1(write1_in[31]), .A2(n3331), .B(n3317), .ZN(n3342) );
  INR3D2BWP12T U3574 ( .A1(n3321), .B1(n3320), .B2(n3319), .ZN(n3322) );
  CKND2D2BWP12T U3575 ( .A1(n3323), .A2(n3322), .ZN(n3328) );
  TPND2D3BWP12T U3576 ( .A1(write1_in[28]), .A2(n530), .ZN(n3326) );
  CKND2D0BWP12T U3577 ( .A1(n3324), .A2(write2_in[28]), .ZN(n3325) );
  TPOAI21D1BWP12T U3578 ( .A1(n3513), .A2(n3326), .B(n3325), .ZN(n3339) );
  IOA21D2BWP12T U3579 ( .A1(n3342), .A2(n3330), .B(n3329), .ZN(n3349) );
  ND2D2BWP12T U3580 ( .A1(write1_in[31]), .A2(n530), .ZN(n3336) );
  CKND2D0BWP12T U3581 ( .A1(n3331), .A2(write2_in[31]), .ZN(n3332) );
  IND3D0BWP12T U3582 ( .A1(n3333), .B1(n3332), .B2(n3505), .ZN(n3334) );
  INVD1BWP12T U3583 ( .I(n3334), .ZN(n3335) );
  TPND2D2BWP12T U3584 ( .A1(n3336), .A2(n3335), .ZN(n3338) );
  NR2XD1BWP12T U3585 ( .A1(n3338), .A2(n3337), .ZN(n3340) );
  ND3XD1BWP12T U3586 ( .A1(n3341), .A2(n3340), .A3(n3339), .ZN(n3348) );
  INVD1BWP12T U3587 ( .I(n3342), .ZN(n3346) );
  TPNR2D0BWP12T U3588 ( .A1(n3343), .A2(n3548), .ZN(n3344) );
  AOI21D1BWP12T U3589 ( .A1(n3346), .A2(n3345), .B(n3344), .ZN(n3347) );
  ND3D1BWP12T U3590 ( .A1(n3349), .A2(n3348), .A3(n3347), .ZN(n2199) );
  INVD1BWP12T U3591 ( .I(tmp1[31]), .ZN(n3351) );
  OAI22D1BWP12T U3592 ( .A1(n3378), .A2(n3351), .B1(n3350), .B2(n3432), .ZN(
        n3355) );
  OAI22D1BWP12T U3593 ( .A1(n3414), .A2(n3353), .B1(n3352), .B2(n3444), .ZN(
        n3354) );
  AOI211D1BWP12T U3594 ( .A1(r1[31]), .A2(n3384), .B(n3355), .C(n3354), .ZN(
        n3375) );
  INVD1BWP12T U3595 ( .I(r12[31]), .ZN(n3356) );
  OAI22D1BWP12T U3596 ( .A1(n3416), .A2(n3357), .B1(n3356), .B2(n3436), .ZN(
        n3367) );
  INVD1BWP12T U3597 ( .I(r4[31]), .ZN(n3359) );
  INVD1BWP12T U3598 ( .I(r8[31]), .ZN(n3358) );
  OAI22D1BWP12T U3599 ( .A1(n3390), .A2(n3359), .B1(n3358), .B2(n3387), .ZN(
        n3366) );
  OAI22D1BWP12T U3600 ( .A1(n3393), .A2(n3360), .B1(n3510), .B2(n1881), .ZN(
        n3365) );
  INVD1BWP12T U3601 ( .I(r6[31]), .ZN(n3362) );
  OAI22D1BWP12T U3602 ( .A1(n3363), .A2(n3362), .B1(n3442), .B2(n3361), .ZN(
        n3364) );
  NR4D0BWP12T U3603 ( .A1(n3367), .A2(n3366), .A3(n3365), .A4(n3364), .ZN(
        n3374) );
  INVD1BWP12T U3604 ( .I(n[3549]), .ZN(n3369) );
  OAI22D1BWP12T U3605 ( .A1(n3404), .A2(n3369), .B1(n3402), .B2(n3368), .ZN(
        n3372) );
  OAI22D1BWP12T U3606 ( .A1(n3406), .A2(n3548), .B1(n3370), .B2(n3434), .ZN(
        n3371) );
  NR2D1BWP12T U3607 ( .A1(n3372), .A2(n3371), .ZN(n3373) );
  ND3D1BWP12T U3608 ( .A1(n3375), .A2(n3374), .A3(n3373), .ZN(regA_out[31]) );
  INVD1BWP12T U3609 ( .I(tmp1[30]), .ZN(n3377) );
  OAI22D1BWP12T U3610 ( .A1(n3378), .A2(n3377), .B1(n3376), .B2(n3432), .ZN(
        n3383) );
  OAI22D1BWP12T U3611 ( .A1(n3381), .A2(n3380), .B1(n3379), .B2(n3444), .ZN(
        n3382) );
  AOI211D1BWP12T U3612 ( .A1(r1[30]), .A2(n3384), .B(n3383), .C(n3382), .ZN(
        n3411) );
  INVD1BWP12T U3613 ( .I(r12[30]), .ZN(n3385) );
  OAI22D1BWP12T U3614 ( .A1(n3416), .A2(n3386), .B1(n3385), .B2(n3436), .ZN(
        n3400) );
  INVD1BWP12T U3615 ( .I(r4[30]), .ZN(n3389) );
  INVD1BWP12T U3616 ( .I(r8[30]), .ZN(n3388) );
  OAI22D0BWP12T U3617 ( .A1(n3390), .A2(n3389), .B1(n3388), .B2(n3387), .ZN(
        n3399) );
  OAI22D1BWP12T U3618 ( .A1(n3393), .A2(n3392), .B1(n3391), .B2(n1881), .ZN(
        n3398) );
  INVD1BWP12T U3619 ( .I(r6[30]), .ZN(n3395) );
  OAI22D1BWP12T U3620 ( .A1(n3396), .A2(n3395), .B1(n3442), .B2(n3394), .ZN(
        n3397) );
  NR4D0BWP12T U3621 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(
        n3410) );
  OAI22D1BWP12T U3622 ( .A1(n3404), .A2(n3403), .B1(n3402), .B2(n3401), .ZN(
        n3408) );
  OAI22D0BWP12T U3623 ( .A1(n3406), .A2(n3547), .B1(n3405), .B2(n3434), .ZN(
        n3407) );
  NR2D1BWP12T U3624 ( .A1(n3408), .A2(n3407), .ZN(n3409) );
  ND3D1BWP12T U3625 ( .A1(n3411), .A2(n3410), .A3(n3409), .ZN(regA_out[30]) );
  ND2D1BWP12T U3626 ( .A1(n3412), .A2(r6[18]), .ZN(n3426) );
  OAI22D1BWP12T U3627 ( .A1(n3416), .A2(n3415), .B1(n3414), .B2(n3413), .ZN(
        n3425) );
  INVD1BWP12T U3628 ( .I(n3417), .ZN(n3422) );
  TPND2D2BWP12T U3629 ( .A1(n3418), .A2(r11[18]), .ZN(n3421) );
  ND2D1BWP12T U3630 ( .A1(n3419), .A2(r9[18]), .ZN(n3420) );
  OAI211D1BWP12T U3631 ( .A1(n3423), .A2(n3422), .B(n3421), .C(n3420), .ZN(
        n3424) );
  INR3D0BWP12T U3632 ( .A1(n3426), .B1(n3425), .B2(n3424), .ZN(n3460) );
  INVD1BWP12T U3633 ( .I(tmp1[18]), .ZN(n3427) );
  NR2D1BWP12T U3634 ( .A1(n622), .A2(n3427), .ZN(n3428) );
  CKND2D0BWP12T U3635 ( .A1(n3429), .A2(n3428), .ZN(n3430) );
  OAI21D1BWP12T U3636 ( .A1(n3432), .A2(n3431), .B(n3430), .ZN(n3440) );
  NR2D1BWP12T U3637 ( .A1(n3434), .A2(n3433), .ZN(n3439) );
  INR2D1BWP12T U3638 ( .A1(r8[18]), .B1(n3435), .ZN(n3438) );
  INR2D1BWP12T U3639 ( .A1(r12[18]), .B1(n3436), .ZN(n3437) );
  NR4D0BWP12T U3640 ( .A1(n3440), .A2(n3439), .A3(n3438), .A4(n3437), .ZN(
        n3459) );
  NR2D1BWP12T U3641 ( .A1(n3444), .A2(n3443), .ZN(n3456) );
  ND2D1BWP12T U3642 ( .A1(n3445), .A2(pc_out[18]), .ZN(n3449) );
  INR2D1BWP12T U3643 ( .A1(n[3562]), .B1(n3446), .ZN(n3447) );
  INVD1BWP12T U3644 ( .I(n3447), .ZN(n3448) );
  ND2D1BWP12T U3645 ( .A1(n3449), .A2(n3448), .ZN(n3455) );
  ND2D1BWP12T U3646 ( .A1(n3450), .A2(r4[18]), .ZN(n3451) );
  OAI21D1BWP12T U3647 ( .A1(n3453), .A2(n1881), .B(n3451), .ZN(n3454) );
  ND3D1BWP12T U3648 ( .A1(n3460), .A2(n3459), .A3(n3458), .ZN(regA_out[18]) );
  AOI22D0BWP12T U3649 ( .A1(lr[21]), .A2(n3473), .B1(r8[21]), .B2(n3493), .ZN(
        n3462) );
  AOI22D0BWP12T U3650 ( .A1(r9[21]), .A2(n3475), .B1(r11[21]), .B2(n2704), 
        .ZN(n3461) );
  OAI211D0BWP12T U3651 ( .A1(n3463), .A2(n3478), .B(n3462), .C(n3461), .ZN(
        n3472) );
  AOI22D0BWP12T U3652 ( .A1(n[3559]), .A2(n3464), .B1(n3480), .B2(pc_out[21]), 
        .ZN(n3471) );
  AOI22D0BWP12T U3653 ( .A1(r5[21]), .A2(n3481), .B1(n2770), .B2(r6[21]), .ZN(
        n3468) );
  AOI22D0BWP12T U3654 ( .A1(r7[21]), .A2(n3482), .B1(n2757), .B2(r4[21]), .ZN(
        n3467) );
  AOI22D0BWP12T U3655 ( .A1(r1[21]), .A2(n3484), .B1(n3483), .B2(r2[21]), .ZN(
        n3466) );
  AOI22D0BWP12T U3656 ( .A1(r0[21]), .A2(n3486), .B1(n3485), .B2(r3[21]), .ZN(
        n3465) );
  ND4D1BWP12T U3657 ( .A1(n3468), .A2(n3467), .A3(n3466), .A4(n3465), .ZN(
        n3469) );
  AOI22D0BWP12T U3658 ( .A1(n3479), .A2(r12[21]), .B1(n3492), .B2(n3469), .ZN(
        n3470) );
  IND3D1BWP12T U3659 ( .A1(n3472), .B1(n3471), .B2(n3470), .ZN(regC_out[21])
         );
  AOI22D0BWP12T U3660 ( .A1(lr[31]), .A2(n3473), .B1(r11[31]), .B2(n2704), 
        .ZN(n3477) );
  AOI22D0BWP12T U3661 ( .A1(n[3549]), .A2(n3464), .B1(r9[31]), .B2(n3475), 
        .ZN(n3476) );
  OAI211D0BWP12T U3662 ( .A1(n3510), .A2(n3478), .B(n3477), .C(n3476), .ZN(
        n3496) );
  AOI22D0BWP12T U3663 ( .A1(pc_out[31]), .A2(n3480), .B1(n3479), .B2(r12[31]), 
        .ZN(n3495) );
  AOI22D0BWP12T U3664 ( .A1(r5[31]), .A2(n3481), .B1(n2770), .B2(r6[31]), .ZN(
        n3490) );
  AOI22D0BWP12T U3665 ( .A1(r7[31]), .A2(n3482), .B1(n2757), .B2(r4[31]), .ZN(
        n3489) );
  AOI22D0BWP12T U3666 ( .A1(r1[31]), .A2(n3484), .B1(n3483), .B2(r2[31]), .ZN(
        n3488) );
  AOI22D0BWP12T U3667 ( .A1(r0[31]), .A2(n3486), .B1(n3485), .B2(r3[31]), .ZN(
        n3487) );
  ND4D1BWP12T U3668 ( .A1(n3490), .A2(n3489), .A3(n3488), .A4(n3487), .ZN(
        n3491) );
  AOI22D0BWP12T U3669 ( .A1(n3493), .A2(r8[31]), .B1(n3492), .B2(n3491), .ZN(
        n3494) );
  IND3D1BWP12T U3670 ( .A1(n3496), .B1(n3495), .B2(n3494), .ZN(regC_out[31])
         );
  OAI21D1BWP12T U3671 ( .A1(n3502), .A2(n3501), .B(n3500), .ZN(n3509) );
  ND4D1BWP12T U3672 ( .A1(n3503), .A2(n3505), .A3(n3506), .A4(n3502), .ZN(
        n3508) );
  IND3D1BWP12T U3673 ( .A1(n3506), .B1(n3505), .B2(n3504), .ZN(n3507) );
  IND3D1BWP12T U3674 ( .A1(n3509), .B1(n3508), .B2(n3507), .ZN(n2188) );
endmodule


module ALU_VARIABLE ( a, b, op, c_in, result, c_out, z, n, v );
  input [31:0] a;
  input [31:0] b;
  input [3:0] op;
  output [31:0] result;
  input c_in;
  output c_out, z, n, v;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n272, n273, n274, n275, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103;

  OAI22D1BWP12T U3 ( .A1(n2548), .A2(n2629), .B1(n2627), .B2(n3455), .ZN(n2708) );
  OAI21D1BWP12T U4 ( .A1(n1614), .A2(n1613), .B(n1612), .ZN(n2817) );
  INVD1BWP12T U5 ( .I(n4933), .ZN(n4636) );
  OAI21D1BWP12T U6 ( .A1(n1596), .A2(n1595), .B(n1594), .ZN(n3788) );
  INVD1BWP12T U7 ( .I(n4846), .ZN(n3843) );
  INVD1BWP12T U8 ( .I(n2817), .ZN(n4985) );
  CKBD1BWP12T U9 ( .I(a[1]), .Z(n4911) );
  INVD1BWP12T U10 ( .I(n5102), .ZN(n4209) );
  INR2D1BWP12T U11 ( .A1(op[2]), .B1(op[3]), .ZN(n933) );
  INVD1BWP12T U12 ( .I(n3872), .ZN(n3933) );
  INVD1BWP12T U13 ( .I(n3873), .ZN(n3930) );
  ND2D1BWP12T U14 ( .A1(n932), .A2(n931), .ZN(n5042) );
  XNR2D1BWP12T U15 ( .A1(n3382), .A2(n3381), .ZN(n4267) );
  INR2D1BWP12T U16 ( .A1(op[2]), .B1(op[1]), .ZN(n765) );
  XNR2D1BWP12T U17 ( .A1(n3234), .A2(n3847), .ZN(n2677) );
  XNR2D1BWP12T U18 ( .A1(n4762), .A2(n2666), .ZN(n2670) );
  XOR2D1BWP12T U19 ( .A1(n2694), .A2(n2693), .Z(n2695) );
  OAI22D1BWP12T U20 ( .A1(n2687), .A2(n2686), .B1(n2685), .B2(n2684), .ZN(
        n2694) );
  XNR2D1BWP12T U21 ( .A1(n4761), .A2(n2688), .ZN(n2692) );
  XNR2D1BWP12T U22 ( .A1(n4843), .A2(n4909), .ZN(n2687) );
  OAI22D1BWP12T U23 ( .A1(n2649), .A2(n2647), .B1(n2579), .B2(n2648), .ZN(
        n2673) );
  XNR2D1BWP12T U24 ( .A1(n2591), .A2(n4906), .ZN(n2703) );
  XNR2D1BWP12T U25 ( .A1(n2623), .A2(n4924), .ZN(n2577) );
  XNR2D1BWP12T U26 ( .A1(n2172), .A2(n4699), .ZN(n2550) );
  XNR2D1BWP12T U27 ( .A1(n2167), .A2(n4916), .ZN(n2549) );
  ND2D1BWP12T U28 ( .A1(n2629), .A2(n2547), .ZN(n2627) );
  XNR2D1BWP12T U29 ( .A1(n2167), .A2(n2746), .ZN(n637) );
  XNR2D1BWP12T U30 ( .A1(n2071), .A2(n2742), .ZN(n435) );
  XNR2D1BWP12T U31 ( .A1(n4214), .A2(n341), .ZN(n417) );
  OAI22D1BWP12T U32 ( .A1(n2028), .A2(n2747), .B1(n2748), .B2(n1910), .ZN(
        n2029) );
  XNR2D1BWP12T U33 ( .A1(b[29]), .A2(n2593), .ZN(n2040) );
  XNR2D1BWP12T U34 ( .A1(n2098), .A2(n2742), .ZN(n570) );
  CKND2D2BWP12T U35 ( .A1(n534), .A2(n355), .ZN(n540) );
  ND2D1BWP12T U36 ( .A1(n610), .A2(n356), .ZN(n534) );
  XNR2D1BWP12T U37 ( .A1(n2072), .A2(n2701), .ZN(n531) );
  OAI22D1BWP12T U38 ( .A1(n558), .A2(n2702), .B1(n609), .B2(n2319), .ZN(n664)
         );
  ND2D1BWP12T U39 ( .A1(n645), .A2(n644), .ZN(n647) );
  INVD1BWP12T U40 ( .I(n649), .ZN(n645) );
  INVD1BWP12T U41 ( .I(n1084), .ZN(n1080) );
  OAI22D1BWP12T U42 ( .A1(n2064), .A2(n2647), .B1(n2227), .B2(n2648), .ZN(
        n2147) );
  BUFFD2BWP12T U43 ( .I(n2263), .Z(n2740) );
  ND2D1BWP12T U44 ( .A1(n2009), .A2(n2008), .ZN(n2122) );
  ND2D1BWP12T U45 ( .A1(n1908), .A2(n1907), .ZN(n1946) );
  OAI21D1BWP12T U46 ( .A1(n2007), .A2(n2006), .B(n2005), .ZN(n1907) );
  CKBD1BWP12T U47 ( .I(n2140), .Z(n2136) );
  CKBD1BWP12T U48 ( .I(n2141), .Z(n2135) );
  INR2D1BWP12T U49 ( .A1(n4316), .B1(n2647), .ZN(n440) );
  INVD1BWP12T U50 ( .I(n491), .ZN(n485) );
  OAI21D1BWP12T U51 ( .A1(n2727), .A2(n2726), .B(n2725), .ZN(n2729) );
  ND2D1BWP12T U52 ( .A1(n2727), .A2(n2726), .ZN(n2728) );
  ND2D1BWP12T U53 ( .A1(n1920), .A2(n1919), .ZN(n2533) );
  IND2D1BWP12T U54 ( .A1(n1918), .B1(n1917), .ZN(n1919) );
  INVD1BWP12T U55 ( .I(n2186), .ZN(n2114) );
  INR2D2BWP12T U56 ( .A1(n2082), .B1(n2081), .ZN(n2142) );
  INR2D1BWP12T U57 ( .A1(n2304), .B1(n2080), .ZN(n2081) );
  OAI22D1BWP12T U58 ( .A1(n504), .A2(n2702), .B1(n531), .B2(n2319), .ZN(n548)
         );
  ND2D1BWP12T U59 ( .A1(n541), .A2(n540), .ZN(n618) );
  ND2D1BWP12T U60 ( .A1(n3651), .A2(n771), .ZN(n773) );
  IOA21D1BWP12T U61 ( .A1(n1047), .A2(n1129), .B(n1046), .ZN(n1275) );
  INVD1BWP12T U62 ( .I(n1275), .ZN(n1271) );
  OR2XD1BWP12T U63 ( .A1(n4694), .A2(n4908), .Z(n3935) );
  IND2D1BWP12T U64 ( .A1(n3132), .B1(n3131), .ZN(n3844) );
  INVD1BWP12T U65 ( .I(n4761), .ZN(n4716) );
  HA1D1BWP12T U66 ( .A(n2156), .B(n2155), .CO(n2289), .S(n2230) );
  OR2XD1BWP12T U67 ( .A1(n4695), .A2(n4922), .Z(n3681) );
  NR2D1BWP12T U68 ( .A1(n3754), .A2(n2854), .ZN(n4797) );
  INVD1BWP12T U69 ( .I(n4730), .ZN(n4693) );
  ND2D1BWP12T U70 ( .A1(n4742), .A2(n373), .ZN(n4109) );
  OA21D1BWP12T U71 ( .A1(n4095), .A2(n384), .B(n4096), .Z(n1755) );
  INVD1BWP12T U72 ( .I(n4098), .ZN(n384) );
  OR2XD1BWP12T U73 ( .A1(n4843), .A2(n4921), .Z(n3352) );
  INVD1BWP12T U74 ( .I(n953), .ZN(n3961) );
  ND2D1BWP12T U75 ( .A1(n3294), .A2(n3293), .ZN(n4580) );
  ND2D1BWP12T U76 ( .A1(n3291), .A2(n3902), .ZN(n3294) );
  ND2D1BWP12T U77 ( .A1(n4743), .A2(n4843), .ZN(n3969) );
  INVD1BWP12T U78 ( .I(n4566), .ZN(n4039) );
  ND2D1BWP12T U79 ( .A1(n4889), .A2(n5099), .ZN(n3777) );
  ND2D1BWP12T U80 ( .A1(n4743), .A2(n848), .ZN(n3509) );
  OAI21D1BWP12T U81 ( .A1(n4476), .A2(n2796), .B(n2801), .ZN(n3830) );
  CKBD1BWP12T U82 ( .I(n2442), .Z(n3868) );
  NR2D1BWP12T U83 ( .A1(n2941), .A2(n2828), .ZN(n3802) );
  NR2D1BWP12T U84 ( .A1(n4698), .A2(n2818), .ZN(n3723) );
  AOI21D1BWP12T U85 ( .A1(n2817), .A2(n2816), .B(n2815), .ZN(n3991) );
  NR2D1BWP12T U86 ( .A1(n981), .A2(n980), .ZN(n4035) );
  INVD1BWP12T U87 ( .I(n3777), .ZN(n3903) );
  TPNR2D1BWP12T U88 ( .A1(n1283), .A2(n2624), .ZN(n1373) );
  INVD1BWP12T U89 ( .I(n4316), .ZN(n1283) );
  INR2D1BWP12T U90 ( .A1(n4209), .B1(n4890), .ZN(n3849) );
  INVD2BWP12T U91 ( .I(n3818), .ZN(n4801) );
  FA1D0BWP12T U92 ( .A(n4711), .B(n4933), .CI(n3431), .CO(n2876), .S(n4363) );
  NR2D1BWP12T U93 ( .A1(n1816), .A2(n3818), .ZN(n4833) );
  INVD1BWP12T U94 ( .I(n3213), .ZN(n3534) );
  ND2D1BWP12T U95 ( .A1(n876), .A2(n875), .ZN(n4779) );
  AOI211D1BWP12T U96 ( .A1(n3937), .A2(n3115), .B(n874), .C(n873), .ZN(n875)
         );
  AN2D1BWP12T U97 ( .A1(n3940), .A2(n3126), .Z(n874) );
  INR2D1BWP12T U98 ( .A1(n3114), .B1(n3812), .ZN(n873) );
  NR2D1BWP12T U99 ( .A1(n4806), .A2(n5024), .ZN(n3304) );
  FA1D0BWP12T U100 ( .A(n2853), .B(n3455), .CI(n2852), .CO(n2808), .S(n4516)
         );
  INVD1BWP12T U101 ( .I(n3899), .ZN(n5038) );
  NR2D1BWP12T U102 ( .A1(n4175), .A2(n4174), .ZN(n4860) );
  INR2D1BWP12T U103 ( .A1(n4742), .B1(n4743), .ZN(n4556) );
  AN2D1BWP12T U104 ( .A1(n953), .A2(n5082), .Z(n4562) );
  INR2D1BWP12T U105 ( .A1(n5075), .B1(n3957), .ZN(n4559) );
  INVD1BWP12T U106 ( .I(n4206), .ZN(n4569) );
  NR2D1BWP12T U107 ( .A1(n4843), .A2(n5040), .ZN(n3645) );
  INVD1BWP12T U108 ( .I(n3199), .ZN(n4493) );
  INVD1BWP12T U109 ( .I(n911), .ZN(n904) );
  INVD1BWP12T U110 ( .I(n5042), .ZN(n4167) );
  AOI211D1BWP12T U111 ( .A1(n5099), .A2(n3843), .B(n3013), .C(n3012), .ZN(
        n3014) );
  XNR2D1BWP12T U112 ( .A1(n2963), .A2(n2962), .ZN(n4978) );
  XNR2D1BWP12T U113 ( .A1(n2950), .A2(n2962), .ZN(n4313) );
  TPOAI22D1BWP12T U114 ( .A1(n1551), .A2(n2646), .B1(n2323), .B2(n4257), .ZN(
        n2326) );
  NR2D1BWP12T U115 ( .A1(n3849), .A2(n3645), .ZN(n3899) );
  AN3XD1BWP12T U116 ( .A1(n4830), .A2(n4829), .A3(n5094), .Z(n1008) );
  AN2D1BWP12T U117 ( .A1(n4833), .A2(n5094), .Z(n1006) );
  NR2D1BWP12T U118 ( .A1(n979), .A2(n978), .ZN(n1020) );
  INVD1BWP12T U119 ( .I(n5088), .ZN(n4396) );
  AOI22D1BWP12T U120 ( .A1(n5090), .A2(n5011), .B1(n5010), .B2(n5093), .ZN(
        n5034) );
  IND2D1BWP12T U121 ( .A1(n3202), .B1(n3201), .ZN(n3211) );
  ND4D1BWP12T U122 ( .A1(n3484), .A2(n3483), .A3(n3482), .A4(n3481), .ZN(n3485) );
  ND2D1BWP12T U123 ( .A1(n4994), .A2(n5093), .ZN(n3484) );
  TPOAI22D1BWP12T U124 ( .A1(n1239), .A2(n2747), .B1(n1150), .B2(n2748), .ZN(
        n1229) );
  TPNR2D1BWP12T U125 ( .A1(n1153), .A2(n1152), .ZN(n1228) );
  NR2D1BWP12T U126 ( .A1(n2648), .A2(n1151), .ZN(n1152) );
  NR2D1BWP12T U127 ( .A1(n1159), .A2(n2647), .ZN(n1153) );
  AO21D1BWP12T U128 ( .A1(n4267), .A2(n5085), .B(n3418), .Z(result[8]) );
  INVD1BWP12T U129 ( .I(n3040), .ZN(n323) );
  ND2D1BWP12T U130 ( .A1(n1052), .A2(n1049), .ZN(n1051) );
  INVD1BWP12T U131 ( .I(n1052), .ZN(n1053) );
  OAI22D1BWP12T U132 ( .A1(n2178), .A2(n2625), .B1(n2177), .B2(n2624), .ZN(
        n1985) );
  INVD2BWP12T U133 ( .I(n2643), .ZN(n1870) );
  INVD1BWP12T U134 ( .I(n1863), .ZN(n1881) );
  XNR2D1BWP12T U135 ( .A1(n4726), .A2(n5014), .ZN(n2741) );
  XNR2D1BWP12T U136 ( .A1(n4754), .A2(n4914), .ZN(n2576) );
  XNR2D1BWP12T U137 ( .A1(n4751), .A2(n2593), .ZN(n2645) );
  INVD1BWP12T U138 ( .I(n4465), .ZN(n272) );
  XNR2D1BWP12T U139 ( .A1(n2551), .A2(n2688), .ZN(n2690) );
  INVD1BWP12T U140 ( .I(n554), .ZN(n555) );
  XNR2D1BWP12T U141 ( .A1(n341), .A2(n288), .ZN(n629) );
  INVD2BWP12T U142 ( .I(n1442), .ZN(n631) );
  XOR2D1BWP12T U143 ( .A1(b[3]), .A2(n866), .Z(n643) );
  ND2D1BWP12T U144 ( .A1(n1106), .A2(n1105), .ZN(n1195) );
  INVD1BWP12T U145 ( .I(n1083), .ZN(n1081) );
  TPOAI22D1BWP12T U146 ( .A1(n2090), .A2(n2680), .B1(n2682), .B2(n1953), .ZN(
        n2088) );
  TPOAI22D1BWP12T U147 ( .A1(n1983), .A2(n2643), .B1(n2073), .B2(n1982), .ZN(
        n2179) );
  XOR3D2BWP12T U148 ( .A1(n2007), .A2(n2006), .A3(n2005), .Z(n2128) );
  INVD1BWP12T U149 ( .I(n1998), .ZN(n1875) );
  TPOAI22D1BWP12T U150 ( .A1(n1993), .A2(n2648), .B1(n1906), .B2(n2647), .ZN(
        n2007) );
  XOR3D2BWP12T U151 ( .A1(n2700), .A2(n2699), .A3(n2698), .Z(n2721) );
  XNR2D1BWP12T U152 ( .A1(n2672), .A2(n2671), .ZN(n2700) );
  XNR3D1BWP12T U153 ( .A1(n2697), .A2(n2696), .A3(n2695), .ZN(n2698) );
  OAI22D1BWP12T U154 ( .A1(n2670), .A2(n2669), .B1(n2668), .B2(n2667), .ZN(
        n2671) );
  XNR2D1BWP12T U155 ( .A1(n4740), .A2(n2701), .ZN(n2705) );
  OAI21D1BWP12T U156 ( .A1(n2709), .A2(n2708), .B(n2706), .ZN(n2707) );
  XNR2D1BWP12T U157 ( .A1(n2551), .A2(n2666), .ZN(n1924) );
  XNR2D1BWP12T U158 ( .A1(n4726), .A2(n2701), .ZN(n1921) );
  XNR2D1BWP12T U159 ( .A1(b[22]), .A2(n4906), .ZN(n2592) );
  CKBD1BWP12T U160 ( .I(n2022), .Z(n284) );
  OAI22D1BWP12T U161 ( .A1(n2595), .A2(n2747), .B1(n2748), .B2(n2028), .ZN(
        n2580) );
  TPOAI22D1BWP12T U162 ( .A1(n2577), .A2(n2620), .B1(n2026), .B2(n2218), .ZN(
        n2582) );
  OAI22D1BWP12T U163 ( .A1(n2556), .A2(n2686), .B1(n2685), .B2(n2038), .ZN(
        n2559) );
  TPOAI22D1BWP12T U164 ( .A1(n1931), .A2(n305), .B1(n1930), .B2(n2624), .ZN(
        n1961) );
  INVD1BWP12T U165 ( .I(n631), .ZN(n483) );
  TPOAI22D1BWP12T U166 ( .A1(n1032), .A2(n2647), .B1(n716), .B2(n1442), .ZN(
        n1050) );
  OAI22D1BWP12T U167 ( .A1(n2667), .A2(n741), .B1(n339), .B2(n2669), .ZN(n1035) );
  XNR2D1BWP12T U168 ( .A1(n4738), .A2(n2666), .ZN(n339) );
  OAI22D1BWP12T U169 ( .A1(n1048), .A2(n4257), .B1(n2646), .B2(n742), .ZN(
        n1036) );
  TPOAI22D1BWP12T U170 ( .A1(n568), .A2(n2263), .B1(n2739), .B2(n611), .ZN(
        n616) );
  INVD1BWP12T U171 ( .I(n614), .ZN(n615) );
  TPOAI22D1BWP12T U172 ( .A1(n606), .A2(n2680), .B1(n654), .B2(n2682), .ZN(
        n648) );
  TPNR2D1BWP12T U173 ( .A1(n639), .A2(n638), .ZN(n661) );
  OAI22D1BWP12T U174 ( .A1(n2263), .A2(n643), .B1(n2739), .B2(n743), .ZN(n736)
         );
  INVD1BWP12T U175 ( .I(n1124), .ZN(n1120) );
  INVD1BWP12T U176 ( .I(n1125), .ZN(n1121) );
  ND2D1BWP12T U177 ( .A1(n1207), .A2(n1206), .ZN(n1262) );
  OR2XD2BWP12T U178 ( .A1(n1256), .A2(n1255), .Z(n1254) );
  ND2D1BWP12T U179 ( .A1(n1045), .A2(n1044), .ZN(n1128) );
  XOR3D2BWP12T U180 ( .A1(n1084), .A2(n1083), .A3(n1079), .Z(n1131) );
  INVD1BWP12T U181 ( .I(n1133), .ZN(n1076) );
  CKBD1BWP12T U182 ( .I(n4914), .Z(n1631) );
  CKBD1BWP12T U183 ( .I(n4916), .Z(n1639) );
  INVD1BWP12T U184 ( .I(n2291), .ZN(n2074) );
  OAI22D1BWP12T U185 ( .A1(n2070), .A2(n2748), .B1(n1994), .B2(n2747), .ZN(
        n2078) );
  TPOAI22D1BWP12T U186 ( .A1(n1935), .A2(n2620), .B1(n2095), .B2(n2218), .ZN(
        n2102) );
  OAI22D2BWP12T U187 ( .A1(n2691), .A2(n2000), .B1(n2099), .B2(n2689), .ZN(
        n2107) );
  INVD1BWP12T U188 ( .I(n2145), .ZN(n2146) );
  INVD1BWP12T U189 ( .I(n2403), .ZN(n2276) );
  INVD1BWP12T U190 ( .I(n1249), .ZN(n1250) );
  INVD1BWP12T U191 ( .I(n4733), .ZN(n4694) );
  INVD1BWP12T U192 ( .I(n4257), .ZN(n420) );
  TPOAI22D1BWP12T U193 ( .A1(n437), .A2(n2748), .B1(n2747), .B2(n436), .ZN(
        n443) );
  INVD1BWP12T U194 ( .I(n446), .ZN(n425) );
  OAI22D1BWP12T U195 ( .A1(n415), .A2(n2647), .B1(n1442), .B2(n431), .ZN(n447)
         );
  XNR2D1BWP12T U196 ( .A1(n2167), .A2(n2593), .ZN(n472) );
  IOA21D1BWP12T U197 ( .A1(n2031), .A2(n2030), .B(n2029), .ZN(n2032) );
  INVD1BWP12T U198 ( .I(n2034), .ZN(n2030) );
  OAI22D1BWP12T U199 ( .A1(n2546), .A2(n2669), .B1(n2667), .B2(n1924), .ZN(
        n2598) );
  OA22D1BWP12T U200 ( .A1(n1940), .A2(n2646), .B1(n2040), .B2(n4257), .Z(n2050) );
  INVD1BWP12T U201 ( .I(n2051), .ZN(n2055) );
  NR2D1BWP12T U202 ( .A1(n2053), .A2(n2052), .ZN(n2056) );
  TPOAI22D1BWP12T U203 ( .A1(n561), .A2(n2646), .B1(n560), .B2(n4257), .ZN(
        n583) );
  XNR2D1BWP12T U204 ( .A1(n4316), .A2(n2701), .ZN(n481) );
  ND2D1BWP12T U205 ( .A1(n551), .A2(n550), .ZN(n574) );
  ND2D1BWP12T U206 ( .A1(n549), .A2(n548), .ZN(n550) );
  INVD1BWP12T U207 ( .I(n664), .ZN(n559) );
  ND2D1BWP12T U208 ( .A1(n725), .A2(n724), .ZN(n727) );
  OAI21D1BWP12T U209 ( .A1(n723), .A2(n722), .B(n721), .ZN(n1070) );
  NR2D1BWP12T U210 ( .A1(n720), .A2(n719), .ZN(n723) );
  XOR3D2BWP12T U211 ( .A1(n1043), .A2(n1042), .A3(n1040), .Z(n1124) );
  INVD1BWP12T U212 ( .I(n4759), .ZN(n4687) );
  INVD1BWP12T U213 ( .I(n1264), .ZN(n1269) );
  INVD1BWP12T U214 ( .I(n4762), .ZN(n4714) );
  INVD1BWP12T U215 ( .I(n336), .ZN(n4715) );
  IOA21D1BWP12T U216 ( .A1(n1413), .A2(n1412), .B(n1411), .ZN(n1490) );
  CKBD1BWP12T U217 ( .I(n4914), .Z(n1634) );
  CKBD1BWP12T U218 ( .I(n4914), .Z(n1598) );
  INVD1BWP12T U219 ( .I(n4726), .ZN(n4712) );
  INVD1BWP12T U220 ( .I(n5053), .ZN(n4713) );
  INVD1BWP12T U221 ( .I(n280), .ZN(n4717) );
  INVD1BWP12T U222 ( .I(n4740), .ZN(n4697) );
  XNR2D1BWP12T U223 ( .A1(n2096), .A2(n4699), .ZN(n2153) );
  XNR2D1BWP12T U224 ( .A1(n4628), .A2(n4914), .ZN(n2178) );
  BUFFD2BWP12T U225 ( .I(b[25]), .Z(n2578) );
  ND2D1BWP12T U226 ( .A1(n2068), .A2(n2067), .ZN(n2303) );
  OAI21D1BWP12T U227 ( .A1(n2364), .A2(n2229), .B(n2228), .ZN(n2362) );
  INVD1BWP12T U228 ( .I(b[26]), .ZN(n4695) );
  INVD1BWP12T U229 ( .I(n4749), .ZN(n4705) );
  OR2XD1BWP12T U230 ( .A1(n4739), .A2(n2818), .Z(n3832) );
  NR2D1BWP12T U231 ( .A1(n2136), .A2(n2135), .ZN(n2138) );
  ND2D1BWP12T U232 ( .A1(n2136), .A2(n2135), .ZN(n2137) );
  INVD1BWP12T U233 ( .I(n2201), .ZN(n2204) );
  ND2D1BWP12T U234 ( .A1(n442), .A2(n441), .ZN(n453) );
  NR2D1BWP12T U235 ( .A1(n4749), .A2(n4905), .ZN(n891) );
  ND2D1BWP12T U236 ( .A1(n2729), .A2(n2728), .ZN(n2768) );
  OAI22D1BWP12T U237 ( .A1(n2142), .A2(n2116), .B1(n2115), .B2(n2144), .ZN(
        n2198) );
  NR2D1BWP12T U238 ( .A1(n2143), .A2(n2111), .ZN(n2116) );
  AN2D1BWP12T U239 ( .A1(n2120), .A2(n2119), .Z(n294) );
  OAI22D1BWP12T U240 ( .A1(n4233), .A2(n4954), .B1(n4489), .B2(n4232), .ZN(
        n4234) );
  INVD1BWP12T U241 ( .I(n4955), .ZN(n4233) );
  XOR3D2BWP12T U242 ( .A1(n622), .A2(n623), .A3(n539), .Z(n690) );
  XOR3D2BWP12T U243 ( .A1(n676), .A2(n675), .A3(n674), .Z(n696) );
  ND2D1BWP12T U244 ( .A1(n947), .A2(n946), .ZN(n4040) );
  INVD1BWP12T U245 ( .I(n4753), .ZN(n4673) );
  XOR3D2BWP12T U246 ( .A1(n1072), .A2(n1073), .A3(n1070), .Z(n1139) );
  NR2D1BWP12T U247 ( .A1(n803), .A2(n4932), .ZN(n807) );
  INVD1BWP12T U248 ( .I(n4752), .ZN(n803) );
  OR2XD1BWP12T U249 ( .A1(n4673), .A2(n783), .Z(n3176) );
  TPNR2D1BWP12T U250 ( .A1(n776), .A2(n775), .ZN(n1614) );
  OR2XD1BWP12T U251 ( .A1(n4687), .A2(n2666), .Z(n1607) );
  INVD1BWP12T U252 ( .I(n4927), .ZN(n4638) );
  ND2D1BWP12T U253 ( .A1(n3102), .A2(n3101), .ZN(n3499) );
  IOA21D1BWP12T U254 ( .A1(n1275), .A2(n1274), .B(n1273), .ZN(n1276) );
  OAI21D1BWP12T U255 ( .A1(n4493), .A2(n1807), .B(n1806), .ZN(n3161) );
  INVD1BWP12T U256 ( .I(n4651), .ZN(n4915) );
  TPNR2D2BWP12T U257 ( .A1(n1279), .A2(n1278), .ZN(n3733) );
  INR2D1BWP12T U258 ( .A1(n3509), .B1(n3982), .ZN(n4846) );
  INVD1BWP12T U259 ( .I(n4729), .ZN(n4683) );
  INVD1BWP12T U260 ( .I(n4739), .ZN(n4698) );
  INVD1BWP12T U261 ( .I(n4214), .ZN(n901) );
  XNR2D1BWP12T U262 ( .A1(n2072), .A2(n4916), .ZN(n2235) );
  XNR2D1BWP12T U263 ( .A1(n2167), .A2(n2688), .ZN(n2234) );
  NR2D1BWP12T U264 ( .A1(n1518), .A2(n2263), .ZN(n1519) );
  NR2D1BWP12T U265 ( .A1(n1558), .A2(n2265), .ZN(n1520) );
  XNR2D1BWP12T U266 ( .A1(n4753), .A2(n2679), .ZN(n2164) );
  XNR2D1BWP12T U267 ( .A1(n2578), .A2(n2593), .ZN(n2166) );
  XOR3D1BWP12T U268 ( .A1(n2304), .A2(n2303), .A3(n2302), .Z(n2315) );
  IOA21D1BWP12T U269 ( .A1(n2285), .A2(n2284), .B(n2283), .ZN(n2301) );
  INVD1BWP12T U270 ( .I(n4728), .ZN(n4651) );
  NR2D1BWP12T U271 ( .A1(n2974), .A2(n2973), .ZN(n4154) );
  OAI22D1BWP12T U272 ( .A1(n3459), .A2(n3957), .B1(n3470), .B2(n3961), .ZN(
        n2973) );
  INVD1BWP12T U273 ( .I(n4727), .ZN(n4711) );
  OAI22D1BWP12T U274 ( .A1(n1914), .A2(n1913), .B1(n1912), .B2(n1911), .ZN(
        n2573) );
  CKBD1BWP12T U275 ( .I(n4304), .Z(n4306) );
  ND2D1BWP12T U276 ( .A1(n4046), .A2(n3566), .ZN(n4874) );
  OAI21D1BWP12T U277 ( .A1(n3936), .A2(n2805), .B(n3998), .ZN(n3591) );
  ND2D1BWP12T U278 ( .A1(n4733), .A2(n4908), .ZN(n3998) );
  INVD1BWP12T U279 ( .I(n4559), .ZN(n3462) );
  NR2D1BWP12T U280 ( .A1(n381), .A2(n380), .ZN(n996) );
  OAI21D1BWP12T U281 ( .A1(n961), .A2(n4394), .B(n4221), .ZN(n4115) );
  MUX2D1BWP12T U282 ( .I0(n373), .I1(n4644), .S(n5075), .Z(n2972) );
  ND2D1BWP12T U283 ( .A1(n4743), .A2(n4125), .ZN(n4100) );
  AOI21D1BWP12T U284 ( .A1(n5075), .A2(n3618), .B(n3621), .ZN(n1768) );
  NR2D1BWP12T U285 ( .A1(n3652), .A2(n1771), .ZN(n1773) );
  INVD1BWP12T U286 ( .I(n5077), .ZN(n5045) );
  INVD1BWP12T U287 ( .I(n1774), .ZN(n4102) );
  NR2D1BWP12T U288 ( .A1(n4891), .A2(n3332), .ZN(n3337) );
  INVD1BWP12T U289 ( .I(n4040), .ZN(n3637) );
  BUFFD2BWP12T U290 ( .I(n2172), .Z(n4748) );
  INVD1BWP12T U291 ( .I(n392), .ZN(n370) );
  XOR3D2BWP12T U292 ( .A1(n457), .A2(n458), .A3(n456), .Z(n406) );
  AOI21D1BWP12T U293 ( .A1(n1774), .A2(n822), .B(n821), .ZN(n3213) );
  ND2D1BWP12T U294 ( .A1(n460), .A2(n459), .ZN(n461) );
  ND2D1BWP12T U295 ( .A1(n456), .A2(n455), .ZN(n460) );
  IND2D1BWP12T U296 ( .A1(n458), .B1(n454), .ZN(n455) );
  INVD1BWP12T U297 ( .I(n3358), .ZN(n3652) );
  NR2D1BWP12T U298 ( .A1(n4748), .A2(n4931), .ZN(n3231) );
  CKBD1BWP12T U299 ( .I(n3234), .Z(n4750) );
  INVD1BWP12T U300 ( .I(n3061), .ZN(n3126) );
  NR3D1BWP12T U301 ( .A1(n3506), .A2(n3505), .A3(n3504), .ZN(n3518) );
  AN2D1BWP12T U302 ( .A1(n499), .A2(n498), .Z(n501) );
  AOI21D1BWP12T U303 ( .A1(n1787), .A2(n802), .B(n801), .ZN(n1596) );
  CKND2D2BWP12T U304 ( .A1(n2517), .A2(n2516), .ZN(n3925) );
  ND2D1BWP12T U305 ( .A1(n2530), .A2(n2529), .ZN(n2770) );
  INVD1BWP12T U306 ( .I(n1944), .ZN(n2607) );
  ND3D1BWP12T U307 ( .A1(n921), .A2(n922), .A3(n925), .ZN(n851) );
  ND2D1BWP12T U308 ( .A1(n856), .A2(n855), .ZN(n927) );
  NR2D1BWP12T U309 ( .A1(n4731), .A2(b[26]), .ZN(n855) );
  NR2D1BWP12T U310 ( .A1(n4730), .A2(n4733), .ZN(n856) );
  INVD1BWP12T U311 ( .I(n288), .ZN(n4679) );
  INVD1BWP12T U312 ( .I(n4931), .ZN(n4631) );
  INVD1BWP12T U313 ( .I(n4925), .ZN(n4652) );
  INVD2BWP12T U314 ( .I(n3217), .ZN(n3321) );
  INVD1BWP12T U315 ( .I(n4904), .ZN(n4654) );
  NR2D1BWP12T U316 ( .A1(n3044), .A2(n3043), .ZN(n3046) );
  INVD1BWP12T U317 ( .I(n4743), .ZN(n3902) );
  NR2D1BWP12T U318 ( .A1(n4205), .A2(n4204), .ZN(n4818) );
  AOI31D1BWP12T U319 ( .A1(n4203), .A2(n4202), .A3(n4201), .B(n4743), .ZN(
        n4204) );
  OAI21D1BWP12T U320 ( .A1(n586), .A2(n585), .B(n584), .ZN(n600) );
  ND2D1BWP12T U321 ( .A1(n587), .A2(n588), .ZN(n584) );
  NR2D1BWP12T U322 ( .A1(n587), .A2(n588), .ZN(n585) );
  ND2D1BWP12T U323 ( .A1(n595), .A2(n594), .ZN(n598) );
  ND2D1BWP12T U324 ( .A1(n3523), .A2(n4655), .ZN(n4446) );
  INVD1BWP12T U325 ( .I(n3940), .ZN(n3813) );
  INVD1BWP12T U326 ( .I(n3100), .ZN(n3114) );
  CKND2D2BWP12T U327 ( .A1(n3005), .A2(n863), .ZN(n3812) );
  CKBD1BWP12T U328 ( .I(n4753), .Z(n295) );
  ND2D1BWP12T U329 ( .A1(n759), .A2(n758), .ZN(n760) );
  CKBD1BWP12T U330 ( .I(n1058), .Z(n4930) );
  OR2XD1BWP12T U331 ( .A1(n4752), .A2(n4932), .Z(n4030) );
  OR2XD1BWP12T U332 ( .A1(n803), .A2(n4932), .Z(n4021) );
  XNR2D1BWP12T U333 ( .A1(n4188), .A2(n4187), .ZN(n4506) );
  AOI21D1BWP12T U334 ( .A1(n3844), .A2(n4743), .B(n3139), .ZN(n4861) );
  XNR2D1BWP12T U335 ( .A1(n3095), .A2(n3160), .ZN(n4409) );
  INVD1BWP12T U336 ( .I(n1145), .ZN(n1146) );
  OR2XD2BWP12T U337 ( .A1(n1147), .A2(n1145), .Z(n4146) );
  TPNR2D1BWP12T U338 ( .A1(n1277), .A2(n1276), .ZN(n3731) );
  XNR2D1BWP12T U339 ( .A1(n4478), .A2(n4477), .ZN(n5062) );
  XNR2D1BWP12T U340 ( .A1(n3883), .A2(n3882), .ZN(n4989) );
  XNR2D1BWP12T U341 ( .A1(n3914), .A2(n3913), .ZN(n4372) );
  OAI21D1BWP12T U342 ( .A1(n4367), .A2(n3912), .B(n3911), .ZN(n3914) );
  INVD2BWP12T U343 ( .I(n4916), .ZN(n1856) );
  XNR2D1BWP12T U344 ( .A1(n3686), .A2(n3697), .ZN(n4377) );
  CKBD1BWP12T U345 ( .I(n3669), .Z(n292) );
  INVD1BWP12T U346 ( .I(n273), .ZN(n3673) );
  CKND2D2BWP12T U347 ( .A1(n2511), .A2(n2510), .ZN(n3672) );
  OAI21D1BWP12T U348 ( .A1(n3553), .A2(n3551), .B(n3552), .ZN(n3430) );
  DEL025D1BWP12T U349 ( .I(n1316), .Z(n1311) );
  ND2D1BWP12T U350 ( .A1(n1354), .A2(n1353), .ZN(n1357) );
  INVD1BWP12T U351 ( .I(n1376), .ZN(n1354) );
  INVD1BWP12T U352 ( .I(n1377), .ZN(n1353) );
  INVD1BWP12T U353 ( .I(n1321), .ZN(n1318) );
  OAI22D1BWP12T U354 ( .A1(n1340), .A2(n2682), .B1(n1304), .B2(n2680), .ZN(
        n312) );
  XNR2D1BWP12T U355 ( .A1(n2167), .A2(n2666), .ZN(n1517) );
  XNR2D1BWP12T U356 ( .A1(n2619), .A2(n5014), .ZN(n2266) );
  XNR2D1BWP12T U357 ( .A1(n4753), .A2(n5014), .ZN(n2264) );
  INVD1BWP12T U358 ( .I(n2329), .ZN(n2330) );
  XNR2D1BWP12T U359 ( .A1(n4740), .A2(n2593), .ZN(n2324) );
  INVD1BWP12T U360 ( .I(n1562), .ZN(n1567) );
  NR2D1BWP12T U361 ( .A1(n1543), .A2(n1542), .ZN(n1541) );
  XNR2D1BWP12T U362 ( .A1(n2226), .A2(n2746), .ZN(n1552) );
  IOA21D1BWP12T U363 ( .A1(n1374), .A2(n1373), .B(n1372), .ZN(n1469) );
  TPOAI22D1BWP12T U364 ( .A1(n1368), .A2(n2744), .B1(n1414), .B2(n2743), .ZN(
        n1471) );
  TPOAI22D1BWP12T U365 ( .A1(n1517), .A2(n2667), .B1(n2237), .B2(n2669), .ZN(
        n2258) );
  TPOAI22D1BWP12T U366 ( .A1(n1547), .A2(n2319), .B1(n1464), .B2(n2702), .ZN(
        n1524) );
  TPNR2D1BWP12T U367 ( .A1(n2511), .A2(n2510), .ZN(n273) );
  INVD1BWP12T U368 ( .I(n4889), .ZN(n3566) );
  NR2D2BWP12T U369 ( .A1(n3051), .A2(n4645), .ZN(n3701) );
  OR2XD1BWP12T U370 ( .A1(n4743), .A2(n4843), .Z(n4611) );
  OAI21D1BWP12T U371 ( .A1(n4476), .A2(n2804), .B(n2803), .ZN(n2886) );
  INVD1BWP12T U372 ( .I(n3758), .ZN(n4045) );
  INVD1BWP12T U373 ( .I(n3812), .ZN(n3939) );
  INR2D1BWP12T U374 ( .A1(n790), .B1(n833), .ZN(n932) );
  INVD1BWP12T U375 ( .I(n4731), .ZN(n4696) );
  OAI21D1BWP12T U376 ( .A1(n3991), .A2(n2821), .B(n2820), .ZN(n2929) );
  NR2D1BWP12T U377 ( .A1(n834), .A2(n4910), .ZN(n4244) );
  INVD1BWP12T U378 ( .I(n5075), .ZN(n834) );
  ND2D1BWP12T U379 ( .A1(n4306), .A2(n4305), .ZN(n4307) );
  CKBD1BWP12T U380 ( .I(n3549), .Z(n300) );
  CKBD1BWP12T U381 ( .I(n982), .Z(n4664) );
  FA1D0BWP12T U382 ( .A(n4693), .B(n4909), .CI(n3554), .CO(n3431), .S(n4362)
         );
  OAI21D1BWP12T U383 ( .A1(n4353), .A2(n2837), .B(n2836), .ZN(n3554) );
  AN2D1BWP12T U384 ( .A1(n3274), .A2(n4569), .Z(n949) );
  NR2D1BWP12T U385 ( .A1(n3637), .A2(n4554), .ZN(n948) );
  NR2D1BWP12T U386 ( .A1(n974), .A2(n973), .ZN(n977) );
  INR2D1BWP12T U387 ( .A1(n1754), .B1(n1753), .ZN(n1756) );
  INVD1BWP12T U388 ( .I(n4921), .ZN(n1765) );
  AN2D1BWP12T U389 ( .A1(n4321), .A2(n5090), .Z(n3349) );
  INVD1BWP12T U390 ( .I(n5100), .ZN(n4046) );
  INVD1BWP12T U391 ( .I(n4249), .ZN(n3604) );
  CKBD1BWP12T U392 ( .I(n4316), .Z(n4258) );
  ND2D1BWP12T U393 ( .A1(n4861), .A2(n4843), .ZN(n4865) );
  ND2D1BWP12T U394 ( .A1(n4788), .A2(n4843), .ZN(n4548) );
  INVD1BWP12T U395 ( .I(n4272), .ZN(n1685) );
  AN2XD2BWP12T U396 ( .A1(n599), .A2(n598), .Z(n4272) );
  NR2D1BWP12T U397 ( .A1(n4093), .A2(n4032), .ZN(n2917) );
  ND2D1BWP12T U398 ( .A1(op[3]), .A2(op[0]), .ZN(n911) );
  INVD1BWP12T U399 ( .I(n4032), .ZN(n3754) );
  ND2D1BWP12T U400 ( .A1(n4760), .A2(n4925), .ZN(n3207) );
  INVD1BWP12T U401 ( .I(n4005), .ZN(n4007) );
  NR2D1BWP12T U402 ( .A1(n4592), .A2(n5042), .ZN(n935) );
  XNR2D1BWP12T U403 ( .A1(n832), .A2(n831), .ZN(n4508) );
  INVD1BWP12T U404 ( .I(n4180), .ZN(n4197) );
  NR2D1BWP12T U405 ( .A1(n4178), .A2(n4177), .ZN(n4179) );
  NR2D1BWP12T U406 ( .A1(n4176), .A2(n4860), .ZN(n4177) );
  XNR2D1BWP12T U407 ( .A1(n3092), .A2(n3158), .ZN(n4947) );
  XNR2D1BWP12T U408 ( .A1(n1801), .A2(n1845), .ZN(n4980) );
  MAOI22D0BWP12T U409 ( .A1(n5065), .A2(n5093), .B1(n5064), .B2(n5063), .ZN(
        n5066) );
  XNR2D1BWP12T U410 ( .A1(n4356), .A2(n4986), .ZN(n5071) );
  XOR2D1BWP12T U411 ( .A1(n4293), .A2(n4292), .Z(n5073) );
  OAI21D1BWP12T U412 ( .A1(n1496), .A2(n3867), .B(n3868), .ZN(n1497) );
  NR2D1BWP12T U413 ( .A1(n1489), .A2(n3867), .ZN(n1498) );
  AOI21D1BWP12T U414 ( .A1(n5093), .A2(n4948), .B(n3860), .ZN(n3861) );
  XNR2D1BWP12T U415 ( .A1(n3807), .A2(n3808), .ZN(n4312) );
  XNR2D1BWP12T U416 ( .A1(n3725), .A2(n3724), .ZN(n4993) );
  OAI21D1BWP12T U417 ( .A1(n3991), .A2(n3723), .B(n3805), .ZN(n3725) );
  ND2D1BWP12T U418 ( .A1(n932), .A2(op[3]), .ZN(n4318) );
  AOI211D1BWP12T U419 ( .A1(n4515), .A2(n4103), .B(n3479), .C(n3478), .ZN(
        n3482) );
  MOAI22D0BWP12T U420 ( .A1(n4035), .A2(n3984), .B1(n3449), .B2(n5094), .ZN(
        n3479) );
  ND2D1BWP12T U421 ( .A1(n4363), .A2(n5090), .ZN(n3483) );
  ND2D1BWP12T U422 ( .A1(n4374), .A2(n5088), .ZN(n3481) );
  INVD2BWP12T U423 ( .I(n4924), .ZN(n1342) );
  XNR2D1BWP12T U424 ( .A1(n4753), .A2(n288), .ZN(n1352) );
  XNR2D1BWP12T U425 ( .A1(n2072), .A2(n2688), .ZN(n1242) );
  XNR2D1BWP12T U426 ( .A1(n2167), .A2(n5014), .ZN(n1180) );
  XNR2D1BWP12T U427 ( .A1(n4761), .A2(n2742), .ZN(n1186) );
  XNR2D1BWP12T U428 ( .A1(n4316), .A2(n4924), .ZN(n1240) );
  NR2D1BWP12T U429 ( .A1(n1296), .A2(n1295), .ZN(n1384) );
  TPOAI22D1BWP12T U430 ( .A1(n1360), .A2(n2647), .B1(n1352), .B2(n1442), .ZN(
        n1377) );
  OAI22D2BWP12T U431 ( .A1(n1464), .A2(n2704), .B1(n1350), .B2(n2702), .ZN(
        n1459) );
  INVD1BWP12T U432 ( .I(n1434), .ZN(n1430) );
  OAI22D1BWP12T U433 ( .A1(n1557), .A2(n2682), .B1(n1439), .B2(n2680), .ZN(
        n1540) );
  AOI21D1BWP12T U434 ( .A1(n2343), .A2(n2342), .B(n2341), .ZN(n2468) );
  BUFFD2BWP12T U435 ( .I(b[27]), .Z(n4731) );
  INVD1BWP12T U436 ( .I(n4165), .ZN(n3763) );
  ND2D1BWP12T U437 ( .A1(n4285), .A2(n4284), .ZN(n4286) );
  NR2D1BWP12T U438 ( .A1(n4283), .A2(n4282), .ZN(n4285) );
  AOI21D1BWP12T U439 ( .A1(n4140), .A2(n4139), .B(n5100), .ZN(n4880) );
  IND2D1BWP12T U440 ( .A1(n4136), .B1(n4135), .ZN(n4137) );
  INR2D1BWP12T U441 ( .A1(n5099), .B1(n4852), .ZN(n3338) );
  ND2D1BWP12T U442 ( .A1(n4265), .A2(n5085), .ZN(n3373) );
  OR3XD1BWP12T U443 ( .A1(n5063), .A2(n4853), .A3(n4854), .Z(n3657) );
  XNR2D1BWP12T U444 ( .A1(n3268), .A2(n3267), .ZN(n4276) );
  ND2D1BWP12T U445 ( .A1(n3266), .A2(n3265), .ZN(n3268) );
  AOI211D1BWP12T U446 ( .A1(n4387), .A2(n5088), .B(n3281), .C(n3280), .ZN(
        n3306) );
  AOI211D1BWP12T U447 ( .A1(n4497), .A2(n4103), .B(n3304), .C(n3303), .ZN(
        n3305) );
  ND2D1BWP12T U448 ( .A1(n4516), .A2(n4103), .ZN(n2874) );
  AN2D1BWP12T U449 ( .A1(n4364), .A2(n5090), .Z(n2877) );
  NR2D1BWP12T U450 ( .A1(n4860), .A2(n4707), .ZN(n5095) );
  MAOI22D0BWP12T U451 ( .A1(n4557), .A2(n4556), .B1(n4555), .B2(n4554), .ZN(
        n4572) );
  NR2D1BWP12T U452 ( .A1(n4623), .A2(n4633), .ZN(n5077) );
  XNR2D1BWP12T U453 ( .A1(n4316), .A2(n5079), .ZN(n5091) );
  INVD1BWP12T U454 ( .I(n4633), .ZN(n5083) );
  INVD1BWP12T U455 ( .I(n5048), .ZN(n5080) );
  INVD1BWP12T U456 ( .I(n3645), .ZN(n5098) );
  IOA21D1BWP12T U457 ( .A1(n4988), .A2(n5093), .B(n1680), .ZN(n1681) );
  XNR2D1BWP12T U458 ( .A1(n1604), .A2(n1603), .ZN(n4357) );
  IOA21D1BWP12T U459 ( .A1(n5090), .A2(n4313), .B(n3018), .ZN(n3019) );
  INVD2BWP12T U460 ( .I(a[7]), .ZN(n414) );
  XNR2D1BWP12T U461 ( .A1(n2071), .A2(n2679), .ZN(n1118) );
  TPOAI22D1BWP12T U462 ( .A1(n1186), .A2(n2744), .B1(n1282), .B2(n2743), .ZN(
        n1293) );
  TPOAI22D1BWP12T U463 ( .A1(n1188), .A2(n4257), .B1(n1187), .B2(n2646), .ZN(
        n1247) );
  ND2D1BWP12T U464 ( .A1(n1193), .A2(n1192), .ZN(n1243) );
  INVD1BWP12T U465 ( .I(n1213), .ZN(n1215) );
  ND2D1BWP12T U466 ( .A1(n1238), .A2(n1237), .ZN(n1322) );
  IND2D1BWP12T U467 ( .A1(n1236), .B1(n1235), .ZN(n1237) );
  IOA21D1BWP12T U468 ( .A1(n1236), .A2(n1234), .B(n1233), .ZN(n1238) );
  INVD1BWP12T U469 ( .I(n1232), .ZN(n1233) );
  TPND2D1BWP12T U470 ( .A1(n2413), .A2(n2412), .ZN(n2490) );
  INVD1BWP12T U471 ( .I(n2483), .ZN(n2482) );
  ND4D1BWP12T U472 ( .A1(n1020), .A2(n1019), .A3(n1018), .A4(n1017), .ZN(
        result[2]) );
  AOI211D1BWP12T U473 ( .A1(n4886), .A2(n1008), .B(n1007), .C(n1006), .ZN(
        n1019) );
  ND2D1BWP12T U474 ( .A1(n1794), .A2(n1793), .ZN(result[4]) );
  INR4D0BWP12T U475 ( .A1(n1792), .B1(n1791), .B2(n1790), .B3(n1789), .ZN(
        n1793) );
  NR2D1BWP12T U476 ( .A1(n1761), .A2(n1760), .ZN(n1794) );
  ND2D1BWP12T U477 ( .A1(n3666), .A2(n3665), .ZN(result[6]) );
  ND2D1BWP12T U478 ( .A1(n4266), .A2(n5085), .ZN(n3665) );
  INR2D1BWP12T U479 ( .A1(n3660), .B1(n3659), .ZN(n3666) );
  ND2D1BWP12T U480 ( .A1(n3264), .A2(n3263), .ZN(result[7]) );
  INR3D0BWP12T U481 ( .A1(n3247), .B1(n3246), .B2(n3245), .ZN(n3264) );
  AOI21D1BWP12T U482 ( .A1(n4269), .A2(n5085), .B(n3262), .ZN(n3263) );
  OAI21D2BWP12T U483 ( .A1(n3544), .A2(n4260), .B(n3543), .ZN(result[9]) );
  INVD1BWP12T U484 ( .I(n4268), .ZN(n3544) );
  AN4XD1BWP12T U485 ( .A1(n3542), .A2(n3541), .A3(n3540), .A4(n3539), .Z(n3543) );
  ND4D1BWP12T U486 ( .A1(n5034), .A2(n5033), .A3(n5032), .A4(n5031), .ZN(n5035) );
  TPNR2D1BWP12T U487 ( .A1(n3211), .A2(n3210), .ZN(n3212) );
  MOAI22D0BWP12T U488 ( .A1(n4826), .A2(n5040), .B1(n4393), .B2(n5088), .ZN(
        n3210) );
  TPOAI22D1BWP12T U489 ( .A1(n1118), .A2(n2682), .B1(n2680), .B2(n1060), .ZN(
        n1085) );
  INVD2BWP12T U490 ( .I(n2679), .ZN(n653) );
  XNR2D1BWP12T U491 ( .A1(n2072), .A2(n2666), .ZN(n1119) );
  XNR2D1BWP12T U492 ( .A1(n2619), .A2(n2742), .ZN(n1113) );
  AN2D1BWP12T U493 ( .A1(n1059), .A2(n4316), .Z(n1086) );
  XNR2D1BWP12T U494 ( .A1(n4316), .A2(n2688), .ZN(n1112) );
  ND2D1BWP12T U495 ( .A1(n1163), .A2(n1162), .ZN(n1379) );
  OAI21D1BWP12T U496 ( .A1(n1225), .A2(n1226), .B(n1224), .ZN(n1162) );
  ND2D1BWP12T U497 ( .A1(n1158), .A2(n1157), .ZN(n1324) );
  IOA21D1BWP12T U498 ( .A1(n1156), .A2(n1228), .B(n1227), .ZN(n1158) );
  XOR3D2BWP12T U499 ( .A1(n1248), .A2(n1247), .A3(n1243), .Z(n1211) );
  ND2D1BWP12T U500 ( .A1(n1174), .A2(n1173), .ZN(n1214) );
  ND2D1BWP12T U501 ( .A1(n1172), .A2(n1171), .ZN(n1173) );
  INVD1BWP12T U502 ( .I(n1392), .ZN(n1393) );
  OAI21D1BWP12T U503 ( .A1(n1087), .A2(n1086), .B(n1085), .ZN(n1088) );
  ND2D1BWP12T U504 ( .A1(n2098), .A2(n288), .ZN(n309) );
  INVD1BWP12T U505 ( .I(n288), .ZN(n308) );
  XNR2D1BWP12T U506 ( .A1(n2094), .A2(n2701), .ZN(n1033) );
  XNR2D1BWP12T U507 ( .A1(n4754), .A2(n5014), .ZN(n1348) );
  XNR2D1BWP12T U508 ( .A1(n4753), .A2(n2742), .ZN(n1067) );
  XNR2D1BWP12T U509 ( .A1(n4738), .A2(n2666), .ZN(n1031) );
  INVD1BWP12T U510 ( .I(n2680), .ZN(n748) );
  XOR3D2BWP12T U511 ( .A1(n1214), .A2(n1213), .A3(n1211), .Z(n1260) );
  NR2D1BWP12T U512 ( .A1(n1097), .A2(n1098), .ZN(n1101) );
  NR2D1BWP12T U513 ( .A1(n1196), .A2(n1195), .ZN(n1198) );
  INVD1BWP12T U514 ( .I(n1194), .ZN(n1199) );
  INR3D0BWP12T U515 ( .A1(n4426), .B1(n4923), .B2(n3770), .ZN(n1) );
  MOAI22D0BWP12T U516 ( .A1(n1), .A2(n3771), .B1(n1), .B2(n3771), .ZN(n4427)
         );
  AOI22D0BWP12T U517 ( .A1(n2666), .A2(n4759), .B1(n4760), .B2(n4925), .ZN(n2)
         );
  AOI22D0BWP12T U518 ( .A1(n4924), .A2(n336), .B1(n2688), .B2(n280), .ZN(n3)
         );
  AOI22D0BWP12T U519 ( .A1(n4923), .A2(n4762), .B1(n4761), .B2(n4927), .ZN(n4)
         );
  CKND2D0BWP12T U520 ( .A1(n4765), .A2(n4906), .ZN(n5) );
  ND4D0BWP12T U521 ( .A1(n2), .A2(n3), .A3(n4), .A4(n5), .ZN(n6) );
  AO211D0BWP12T U522 ( .A1(n4910), .A2(n5075), .B(n5076), .C(n6), .Z(n4766) );
  IOA21D0BWP12T U523 ( .A1(n3318), .A2(n848), .B(n4035), .ZN(n3456) );
  CKND2D0BWP12T U524 ( .A1(n4426), .A2(n4425), .ZN(n7) );
  MAOI22D0BWP12T U525 ( .A1(n5051), .A2(n7), .B1(n5051), .B2(n7), .ZN(n5050)
         );
  IND2D0BWP12T U526 ( .A1(n3743), .B1(n3744), .ZN(n3789) );
  IAO21D0BWP12T U527 ( .A1(n4910), .A2(c_in), .B(n961), .ZN(n962) );
  IND2D0BWP12T U528 ( .A1(n4149), .B1(n4150), .ZN(n4187) );
  MAOI22D0BWP12T U529 ( .A1(n3051), .A2(n3128), .B1(n3067), .B2(n4624), .ZN(
        n3190) );
  IND2D0BWP12T U530 ( .A1(n4226), .B1(n4227), .ZN(n4243) );
  AO21D0BWP12T U531 ( .A1(n3988), .A2(n3935), .B(n2829), .Z(n8) );
  AOI31D0BWP12T U532 ( .A1(n2929), .A2(n3935), .A3(n3989), .B(n8), .ZN(n3553)
         );
  CKND2D0BWP12T U533 ( .A1(n4124), .A2(n373), .ZN(n9) );
  MAOI22D0BWP12T U534 ( .A1(n4125), .A2(n9), .B1(n4125), .B2(n9), .ZN(n4419)
         );
  IND2D0BWP12T U535 ( .A1(n4475), .B1(n4474), .ZN(n3785) );
  AN4D0BWP12T U536 ( .A1(n10), .A2(n4109), .A3(n4225), .A4(n1769), .Z(n1771)
         );
  CKND0BWP12T U537 ( .I(n1770), .ZN(n10) );
  MOAI22D0BWP12T U538 ( .A1(n4742), .A2(n3456), .B1(n4742), .B2(n3455), .ZN(
        n3643) );
  IND4D0BWP12T U539 ( .A1(n4838), .B1(n4826), .B2(n4828), .B3(n4827), .ZN(n11)
         );
  OAI21D0BWP12T U540 ( .A1(n4843), .A2(n4836), .B(n4835), .ZN(n12) );
  NR4D0BWP12T U541 ( .A1(n4837), .A2(n4833), .A3(n4834), .A4(n12), .ZN(n13) );
  NR4D0BWP12T U542 ( .A1(n4842), .A2(n4839), .A3(n4841), .A4(n4840), .ZN(n14)
         );
  ND4D0BWP12T U543 ( .A1(n4819), .A2(n4860), .A3(n4853), .A4(n4820), .ZN(n15)
         );
  INR4D0BWP12T U544 ( .A1(n4821), .B1(n4823), .B2(n4822), .B3(n15), .ZN(n16)
         );
  AO31D0BWP12T U545 ( .A1(n4824), .A2(n4825), .A3(n16), .B(n4843), .Z(n17) );
  IND4D0BWP12T U546 ( .A1(n11), .B1(n13), .B2(n14), .B3(n17), .ZN(n4844) );
  IND2D0BWP12T U547 ( .A1(n4189), .B1(n4190), .ZN(n4193) );
  INR2D0BWP12T U548 ( .A1(n963), .B1(n4114), .ZN(n18) );
  OAI21D0BWP12T U549 ( .A1(n961), .A2(n4487), .B(n4229), .ZN(n19) );
  MAOI22D0BWP12T U550 ( .A1(n18), .A2(n19), .B1(n18), .B2(n19), .ZN(n4488) );
  NR2D0BWP12T U551 ( .A1(n3606), .A2(n4921), .ZN(n20) );
  MOAI22D0BWP12T U552 ( .A1(n2746), .A2(n20), .B1(n2746), .B2(n20), .ZN(n4433)
         );
  IOA21D0BWP12T U553 ( .A1(n3999), .A2(n3994), .B(n3998), .ZN(n21) );
  AOI31D1BWP12T U554 ( .A1(n2931), .A2(n3999), .A3(n3995), .B(n21), .ZN(n3555)
         );
  INR2D0BWP12T U555 ( .A1(n4785), .B1(n4546), .ZN(n22) );
  AOI211D0BWP12T U556 ( .A1(n4548), .A2(n4866), .B(n22), .C(n4547), .ZN(n23)
         );
  ND4D0BWP12T U557 ( .A1(n4544), .A2(n4543), .A3(n4821), .A4(n4825), .ZN(n24)
         );
  IND4D0BWP12T U558 ( .A1(n4532), .B1(n4788), .B2(n4860), .B3(n4824), .ZN(n25)
         );
  OAI31D0BWP12T U559 ( .A1(n4784), .A2(n24), .A3(n25), .B(n4605), .ZN(n26) );
  OAI21D0BWP12T U560 ( .A1(n4549), .A2(n4605), .B(n4886), .ZN(n27) );
  ND4D0BWP12T U561 ( .A1(n4550), .A2(n23), .A3(n26), .A4(n27), .ZN(n4776) );
  AOI21D0BWP12T U562 ( .A1(n3829), .A2(n3830), .B(n3828), .ZN(n28) );
  CKND2D0BWP12T U563 ( .A1(n3831), .A2(n3832), .ZN(n29) );
  MAOI22D0BWP12T U564 ( .A1(n28), .A2(n29), .B1(n28), .B2(n29), .ZN(n4509) );
  INR2D0BWP12T U565 ( .A1(n3987), .B1(n3991), .ZN(n30) );
  OAI32D0BWP12T U566 ( .A1(n3988), .A2(n30), .A3(n3990), .B1(n3989), .B2(n3988), .ZN(n31) );
  MAOI22D0BWP12T U567 ( .A1(n31), .A2(n3992), .B1(n31), .B2(n3992), .ZN(n4992)
         );
  IND2D0BWP12T U568 ( .A1(n3602), .B1(n3603), .ZN(n3654) );
  OAI22D0BWP12T U569 ( .A1(n4200), .A2(n4567), .B1(n3812), .B2(n2972), .ZN(n32) );
  AOI21D0BWP12T U570 ( .A1(n3107), .A2(n3471), .B(n32), .ZN(n3946) );
  CKND2D0BWP12T U571 ( .A1(op[2]), .A2(op[1]), .ZN(n33) );
  NR2D0BWP12T U572 ( .A1(n911), .A2(n33), .ZN(n5048) );
  NR2D0BWP12T U573 ( .A1(n4583), .A2(n4582), .ZN(n34) );
  AOI31D0BWP12T U574 ( .A1(n4588), .A2(n4587), .A3(n34), .B(n4890), .ZN(n35)
         );
  NR4D0BWP12T U575 ( .A1(n4591), .A2(n4590), .A3(n4589), .A4(n35), .ZN(n36) );
  INR3D0BWP12T U576 ( .A1(n4581), .B1(n5020), .B2(n5096), .ZN(n37) );
  AOI32D0BWP12T U577 ( .A1(n4580), .A2(n36), .A3(n37), .B1(n4890), .B2(n36), 
        .ZN(n4599) );
  INR2D0BWP12T U578 ( .A1(n4573), .B1(n4545), .ZN(n4866) );
  AN4XD1BWP12T U579 ( .A1(n38), .A2(n4680), .A3(n710), .A4(n1721), .Z(n3142)
         );
  CKND0BWP12T U580 ( .I(n4057), .ZN(n38) );
  CKND2D0BWP12T U581 ( .A1(n2969), .A2(n2968), .ZN(n39) );
  OAI211D0BWP12T U582 ( .A1(n3888), .A2(n2784), .B(n2967), .C(n39), .ZN(n2785)
         );
  AOI21D0BWP12T U583 ( .A1(n3746), .A2(n3696), .B(n3695), .ZN(n40) );
  MAOI22D0BWP12T U584 ( .A1(n40), .A2(n3697), .B1(n40), .B2(n3697), .ZN(n4505)
         );
  NR2D0BWP12T U585 ( .A1(n3606), .A2(n3605), .ZN(n41) );
  MOAI22D0BWP12T U586 ( .A1(n4931), .A2(n41), .B1(n4931), .B2(n41), .ZN(n4432)
         );
  OAI22D1BWP12T U587 ( .A1(n3323), .A2(n4665), .B1(n3322), .B2(n4624), .ZN(n42) );
  OAI22D0BWP12T U588 ( .A1(n3321), .A2(n4636), .B1(n275), .B2(n4664), .ZN(n43)
         );
  NR2D1BWP12T U589 ( .A1(n42), .A2(n43), .ZN(n4173) );
  INR2D0BWP12T U590 ( .A1(n4108), .B1(n975), .ZN(n44) );
  OAI21D0BWP12T U591 ( .A1(n4226), .A2(n4244), .B(n4227), .ZN(n45) );
  MAOI22D0BWP12T U592 ( .A1(n44), .A2(n45), .B1(n44), .B2(n45), .ZN(n4317) );
  CKND0BWP12T U593 ( .I(n4556), .ZN(n46) );
  CKND0BWP12T U594 ( .I(n3902), .ZN(n47) );
  INR2D1BWP12T U595 ( .A1(n4039), .B1(n4555), .ZN(n48) );
  AOI211D1BWP12T U596 ( .A1(n1752), .A2(n47), .B(n48), .C(n4843), .ZN(n49) );
  OAI21D1BWP12T U597 ( .A1(n4172), .A2(n46), .B(n49), .ZN(n1720) );
  AOI222D0BWP12T U598 ( .A1(n3937), .A2(n3953), .B1(n3940), .B2(n3954), .C1(
        n3939), .C2(n3952), .ZN(n50) );
  IOA21D0BWP12T U599 ( .A1(n3941), .A2(n3951), .B(n50), .ZN(n4802) );
  CKND2D0BWP12T U600 ( .A1(n3832), .A2(n3831), .ZN(n51) );
  MAOI22D0BWP12T U601 ( .A1(n3997), .A2(n51), .B1(n3997), .B2(n51), .ZN(n4408)
         );
  IND2D0BWP12T U602 ( .A1(n3029), .B1(n3030), .ZN(n3035) );
  CKND2D0BWP12T U603 ( .A1(n3999), .A2(n3998), .ZN(n52) );
  MAOI22D0BWP12T U604 ( .A1(n3936), .A2(n52), .B1(n3936), .B2(n52), .ZN(n4500)
         );
  IND2D0BWP12T U605 ( .A1(n4446), .B1(n4448), .ZN(n53) );
  MAOI22D0BWP12T U606 ( .A1(n4904), .A2(n53), .B1(n4904), .B2(n53), .ZN(n4443)
         );
  NR4D0BWP12T U607 ( .A1(n4262), .A2(n4265), .A3(n4261), .A4(n4266), .ZN(n54)
         );
  NR3D1BWP12T U608 ( .A1(n4267), .A2(n4268), .A3(n4269), .ZN(n55) );
  IIND4D1BWP12T U609 ( .A1(n4263), .A2(n4264), .B1(n54), .B2(n55), .ZN(n56) );
  NR4D0BWP12T U610 ( .A1(n4275), .A2(n4276), .A3(n5036), .A4(n56), .ZN(n4280)
         );
  NR4D0BWP12T U611 ( .A1(n4964), .A2(n4962), .A3(n4963), .A4(n4961), .ZN(n57)
         );
  NR4D0BWP12T U612 ( .A1(n4953), .A2(n4955), .A3(n4954), .A4(n5092), .ZN(n58)
         );
  IND2D0BWP12T U613 ( .A1(n4957), .B1(n58), .ZN(n59) );
  NR4D0BWP12T U614 ( .A1(n4958), .A2(n4956), .A3(n4960), .A4(n59), .ZN(n60) );
  NR4D0BWP12T U615 ( .A1(n4976), .A2(n5010), .A3(n4977), .A4(n4978), .ZN(n61)
         );
  IND4D0BWP12T U616 ( .A1(n4959), .B1(n57), .B2(n60), .B3(n61), .ZN(n4981) );
  AOI21D1BWP12T U617 ( .A1(n3217), .A2(n848), .B(n3128), .ZN(n3823) );
  OA21D0BWP12T U618 ( .A1(n4486), .A2(n4910), .B(n4487), .Z(n5089) );
  AOI222D0BWP12T U619 ( .A1(n3937), .A2(n3119), .B1(n3940), .B2(n3118), .C1(
        n3811), .C2(n3939), .ZN(n62) );
  IOA21D0BWP12T U620 ( .A1(n3941), .A2(n3810), .B(n62), .ZN(n3559) );
  IND2D0BWP12T U621 ( .A1(n3412), .B1(n3411), .ZN(n3260) );
  MAOI22D0BWP12T U622 ( .A1(n1709), .A2(n1710), .B1(n3323), .B2(n4650), .ZN(
        n63) );
  OA21D0BWP12T U623 ( .A1(n3850), .A2(n275), .B(n63), .Z(n4171) );
  IND2D0BWP12T U624 ( .A1(n4379), .B1(n4492), .ZN(n64) );
  OAI211D1BWP12T U625 ( .A1(n4381), .A2(n895), .B(n4491), .C(n64), .ZN(n1734)
         );
  INR3D0BWP12T U626 ( .A1(n4448), .B1(n4925), .B2(n4058), .ZN(n65) );
  MOAI22D0BWP12T U627 ( .A1(n3187), .A2(n65), .B1(n3187), .B2(n65), .ZN(n4453)
         );
  IOA21D0BWP12T U628 ( .A1(n3161), .A2(n3094), .B(n3093), .ZN(n66) );
  MOAI22D0BWP12T U629 ( .A1(n1844), .A2(n66), .B1(n1844), .B2(n66), .ZN(n4502)
         );
  AO21D0BWP12T U630 ( .A1(n4536), .A2(n4569), .B(n3052), .Z(n4542) );
  CKND0BWP12T U631 ( .I(n3930), .ZN(n67) );
  CKND0BWP12T U632 ( .I(n3989), .ZN(n68) );
  NR3D0BWP12T U633 ( .A1(n3929), .A2(n3928), .A3(n68), .ZN(n69) );
  CKND0BWP12T U634 ( .I(n69), .ZN(n70) );
  OAI32D0BWP12T U635 ( .A1(n68), .A2(n3928), .A3(n3932), .B1(n3931), .B2(n68), 
        .ZN(n71) );
  AOI211D0BWP12T U636 ( .A1(n69), .A2(n3933), .B(n3988), .C(n71), .ZN(n72) );
  OAI31D0BWP12T U637 ( .A1(n4353), .A2(n67), .A3(n70), .B(n72), .ZN(n73) );
  MOAI22D0BWP12T U638 ( .A1(n3992), .A2(n73), .B1(n3992), .B2(n73), .ZN(n4314)
         );
  AOI22D0BWP12T U639 ( .A1(n4751), .A2(n905), .B1(n4633), .B2(n4668), .ZN(n74)
         );
  CKND0BWP12T U640 ( .I(n4751), .ZN(n75) );
  AOI222D0BWP12T U641 ( .A1(n2870), .A2(n4751), .B1(n2870), .B2(op[2]), .C1(
        n4623), .C2(n75), .ZN(n76) );
  MAOI22D0BWP12T U642 ( .A1(n4624), .A2(n5048), .B1(n4624), .B2(n76), .ZN(n77)
         );
  OAI211D0BWP12T U643 ( .A1(n4616), .A2(n5042), .B(n74), .C(n77), .ZN(n2871)
         );
  CKND2D0BWP12T U644 ( .A1(n4394), .A2(n4952), .ZN(n78) );
  MOAI22D0BWP12T U645 ( .A1(n5075), .A2(n78), .B1(n5075), .B2(n78), .ZN(n5087)
         );
  AOI22D0BWP12T U646 ( .A1(n3447), .A2(n3125), .B1(n1822), .B2(n3701), .ZN(n79) );
  CKND2D0BWP12T U647 ( .A1(n953), .A2(n1821), .ZN(n80) );
  OAI211D0BWP12T U648 ( .A1(n3471), .A2(n3959), .B(n79), .C(n80), .ZN(n3291)
         );
  MOAI22D0BWP12T U649 ( .A1(n2916), .A2(n3061), .B1(n3107), .B2(n3115), .ZN(
        n4093) );
  INR3D0BWP12T U650 ( .A1(n4426), .B1(n5051), .B2(n3892), .ZN(n81) );
  MOAI22D0BWP12T U651 ( .A1(n81), .A2(n3053), .B1(n81), .B2(n3053), .ZN(n4430)
         );
  IND2D0BWP12T U652 ( .A1(n3432), .B1(n3433), .ZN(n82) );
  MAOI22D0BWP12T U653 ( .A1(n3434), .A2(n82), .B1(n3434), .B2(n82), .ZN(n4515)
         );
  AOI21D0BWP12T U654 ( .A1(n3788), .A2(n3787), .B(n3786), .ZN(n83) );
  MAOI22D0BWP12T U655 ( .A1(n83), .A2(n3789), .B1(n83), .B2(n3789), .ZN(n4330)
         );
  INR2D0BWP12T U656 ( .A1(n3993), .B1(n3997), .ZN(n84) );
  OAI32D0BWP12T U657 ( .A1(n3994), .A2(n84), .A3(n3996), .B1(n3995), .B2(n3994), .ZN(n85) );
  CKND2D0BWP12T U658 ( .A1(n3999), .A2(n3998), .ZN(n86) );
  MAOI22D0BWP12T U659 ( .A1(n85), .A2(n86), .B1(n85), .B2(n86), .ZN(n4376) );
  CKND0BWP12T U660 ( .I(n4566), .ZN(n87) );
  OAI21D0BWP12T U661 ( .A1(n4521), .A2(n4520), .B(n4707), .ZN(n88) );
  AOI21D0BWP12T U662 ( .A1(n4088), .A2(n87), .B(n88), .ZN(n89) );
  OAI21D0BWP12T U663 ( .A1(n3902), .A2(n3223), .B(n89), .ZN(n4823) );
  CKND0BWP12T U664 ( .I(n848), .ZN(n90) );
  AOI32D0BWP12T U665 ( .A1(n4954), .A2(n90), .A3(n4318), .B1(n848), .B2(n3487), 
        .ZN(n3490) );
  CKND2D0BWP12T U666 ( .A1(n4951), .A2(n4952), .ZN(n91) );
  MOAI22D0BWP12T U667 ( .A1(n5082), .A2(n91), .B1(n5082), .B2(n91), .ZN(n5092)
         );
  IAO21D0BWP12T U668 ( .A1(n4753), .A2(n827), .B(n828), .ZN(n830) );
  CKND0BWP12T U669 ( .I(n4367), .ZN(n92) );
  AOI21D0BWP12T U670 ( .A1(n3781), .A2(n92), .B(n3784), .ZN(n93) );
  MAOI22D0BWP12T U671 ( .A1(n93), .A2(n1844), .B1(n93), .B2(n1844), .ZN(n4411)
         );
  AOI21D0BWP12T U672 ( .A1(n4384), .A2(n3206), .B(n1734), .ZN(n94) );
  MAOI22D0BWP12T U673 ( .A1(n94), .A2(n1735), .B1(n94), .B2(n1735), .ZN(n4392)
         );
  CKND0BWP12T U674 ( .I(n4743), .ZN(n95) );
  OAI221D0BWP12T U675 ( .A1(n4743), .A2(n1655), .B1(n95), .B2(n4585), .C(n4605), .ZN(n4592) );
  IAO21D0BWP12T U676 ( .A1(n3190), .A2(n4685), .B(n3052), .ZN(n4859) );
  NR4D0BWP12T U677 ( .A1(n4467), .A2(n4466), .A3(n4469), .A4(n4468), .ZN(n96)
         );
  NR4D0BWP12T U678 ( .A1(n4444), .A2(n4445), .A3(n4442), .A4(n4443), .ZN(n97)
         );
  ND4D0BWP12T U679 ( .A1(n4454), .A2(n97), .A3(n4455), .A4(n4456), .ZN(n98) );
  NR4D0BWP12T U680 ( .A1(n4433), .A2(n4431), .A3(n4432), .A4(n4430), .ZN(n99)
         );
  NR4D0BWP12T U681 ( .A1(n4429), .A2(n4428), .A3(n4427), .A4(n5050), .ZN(n100)
         );
  NR4D0BWP12T U682 ( .A1(n4422), .A2(n4424), .A3(n4434), .A4(n4423), .ZN(n101)
         );
  ND3D0BWP12T U683 ( .A1(n99), .A2(n100), .A3(n101), .ZN(n102) );
  NR4D0BWP12T U684 ( .A1(n4458), .A2(n4457), .A3(n98), .A4(n102), .ZN(n103) );
  AO31D0BWP12T U685 ( .A1(n4573), .A2(n4470), .A3(n96), .B(n103), .Z(n104) );
  CKND2D0BWP12T U686 ( .A1(n5079), .A2(n104), .ZN(n4471) );
  OAI21D0BWP12T U687 ( .A1(n4353), .A2(n3873), .B(n3872), .ZN(n105) );
  MOAI22D0BWP12T U688 ( .A1(n3882), .A2(n105), .B1(n3882), .B2(n105), .ZN(
        n4358) );
  CKND2D0BWP12T U689 ( .A1(n3589), .A2(n3590), .ZN(n106) );
  MOAI22D0BWP12T U690 ( .A1(n3591), .A2(n106), .B1(n3591), .B2(n106), .ZN(
        n4514) );
  IOA21D0BWP12T U691 ( .A1(n4035), .A2(n3766), .B(n1015), .ZN(n4544) );
  IND2D0BWP12T U692 ( .A1(n4251), .B1(n4801), .ZN(n4787) );
  OR3D0BWP12T U693 ( .A1(n860), .A2(op[3]), .A3(op[2]), .Z(n5102) );
  OAI22D0BWP12T U694 ( .A1(n3812), .A2(n3964), .B1(n3813), .B2(n3951), .ZN(
        n107) );
  AOI21D0BWP12T U695 ( .A1(n3941), .A2(n3688), .B(n107), .ZN(n108) );
  OAI32D0BWP12T U696 ( .A1(n3818), .A2(n3945), .A3(n3960), .B1(n108), .B2(
        n3818), .ZN(n3689) );
  AO222D1BWP12T U697 ( .A1(n3701), .A2(n3126), .B1(n953), .B2(n3115), .C1(
        n3067), .C2(n3114), .Z(n3575) );
  CKND2D0BWP12T U698 ( .A1(n3649), .A2(n3651), .ZN(n109) );
  OAI21D0BWP12T U699 ( .A1(n109), .A2(n4486), .B(n3653), .ZN(n110) );
  MOAI22D0BWP12T U700 ( .A1(n3654), .A2(n110), .B1(n3654), .B2(n110), .ZN(
        n4964) );
  RCIAO21D0BWP12T U701 ( .A1(n4843), .A2(n4921), .B(n3628), .ZN(n3620) );
  INR3D0BWP12T U702 ( .A1(n4426), .B1(n3891), .B2(n3892), .ZN(n111) );
  MOAI22D0BWP12T U703 ( .A1(n111), .A2(n4915), .B1(n111), .B2(n4915), .ZN(
        n4445) );
  CKND0BWP12T U704 ( .I(n3681), .ZN(n112) );
  OA21D0BWP12T U705 ( .A1(n3805), .A2(n112), .B(n3680), .Z(n3931) );
  NR4D0BWP12T U706 ( .A1(n4508), .A2(n4507), .A3(n4506), .A4(n4505), .ZN(n113)
         );
  NR4D0BWP12T U707 ( .A1(n4512), .A2(n4511), .A3(n4510), .A4(n4509), .ZN(n114)
         );
  IND4D0BWP12T U708 ( .A1(n4514), .B1(n113), .B2(n114), .B3(n4513), .ZN(n115)
         );
  NR4D0BWP12T U709 ( .A1(n4485), .A2(n4484), .A3(n4483), .A4(n4482), .ZN(n116)
         );
  NR4D0BWP12T U710 ( .A1(n4481), .A2(n4480), .A3(n4479), .A4(n5062), .ZN(n117)
         );
  NR4D0BWP12T U711 ( .A1(n4497), .A2(n4499), .A3(n4498), .A4(n4500), .ZN(n118)
         );
  ND3D0BWP12T U712 ( .A1(n116), .A2(n117), .A3(n118), .ZN(n119) );
  NR4D0BWP12T U713 ( .A1(n4516), .A2(n4515), .A3(n115), .A4(n119), .ZN(n4944)
         );
  CKND0BWP12T U714 ( .I(n4131), .ZN(n120) );
  OAI21D0BWP12T U715 ( .A1(n4244), .A2(n120), .B(n4132), .ZN(n121) );
  CKND2D0BWP12T U716 ( .A1(n4134), .A2(n4133), .ZN(n122) );
  MOAI22D0BWP12T U717 ( .A1(n121), .A2(n122), .B1(n121), .B2(n122), .ZN(n4323)
         );
  AOI21D0BWP12T U718 ( .A1(n3824), .A2(n4848), .B(n3902), .ZN(n123) );
  INVD1BWP12T U719 ( .I(n3141), .ZN(n124) );
  CKND2D0BWP12T U720 ( .A1(n3766), .A2(n3823), .ZN(n125) );
  OAI31D1BWP12T U721 ( .A1(n3140), .A2(n123), .A3(n124), .B(n125), .ZN(n4788)
         );
  CKND0BWP12T U722 ( .I(n3509), .ZN(n126) );
  OAI32D0BWP12T U723 ( .A1(n4605), .A2(n3567), .A3(n126), .B1(n4573), .B2(
        n4605), .ZN(n127) );
  OAI21D0BWP12T U724 ( .A1(n3191), .A2(n127), .B(n4046), .ZN(n4896) );
  CKND0BWP12T U725 ( .I(n5048), .ZN(n128) );
  MOAI22D0BWP12T U726 ( .A1(n4921), .A2(n128), .B1(n4921), .B2(n1764), .ZN(
        n129) );
  AOI21D0BWP12T U727 ( .A1(n5078), .A2(n4422), .B(n129), .ZN(n130) );
  AOI32D0BWP12T U728 ( .A1(n4633), .A2(n4843), .A3(n1765), .B1(n905), .B2(
        n4843), .ZN(n131) );
  OA211D0BWP12T U729 ( .A1(n4819), .A2(n5098), .B(n130), .C(n131), .Z(n1792)
         );
  IOA21D0BWP12T U730 ( .A1(n5094), .A2(n4842), .B(n3513), .ZN(n132) );
  AOI21D0BWP12T U731 ( .A1(n5090), .A2(n4343), .B(n132), .ZN(n3542) );
  INR2D1BWP12T U732 ( .A1(n3005), .B1(n3436), .ZN(n3097) );
  AO21D1BWP12T U733 ( .A1(n1711), .A2(n4742), .B(n1708), .Z(n1752) );
  OA21D0BWP12T U734 ( .A1(n4035), .A2(n4206), .B(n3644), .Z(n4538) );
  AOI21D0BWP12T U735 ( .A1(n4624), .A2(n4843), .B(n4891), .ZN(n4889) );
  NR4D0BWP12T U736 ( .A1(n4405), .A2(n4404), .A3(n4403), .A4(n4402), .ZN(n133)
         );
  NR2D0BWP12T U737 ( .A1(n4409), .A2(n4408), .ZN(n134) );
  NR4D0BWP12T U738 ( .A1(n4417), .A2(n4416), .A3(n4407), .A4(n4406), .ZN(n135)
         );
  NR4D0BWP12T U739 ( .A1(n4375), .A2(n4374), .A3(n4377), .A4(n4376), .ZN(n136)
         );
  ND4D0BWP12T U740 ( .A1(n133), .A2(n134), .A3(n135), .A4(n136), .ZN(n4473) );
  AOI21D0BWP12T U741 ( .A1(n4333), .A2(n4192), .B(n4191), .ZN(n137) );
  MAOI22D0BWP12T U742 ( .A1(n137), .A2(n4193), .B1(n137), .B2(n4193), .ZN(
        n4341) );
  AO222D1BWP12T U743 ( .A1(n4742), .A2(n4567), .B1(n953), .B2(n2972), .C1(
        n3125), .C2(n3004), .Z(n4607) );
  INR3D0BWP12T U744 ( .A1(n4448), .B1(n4057), .B2(n4058), .ZN(n138) );
  MOAI22D0BWP12T U745 ( .A1(n4932), .A2(n138), .B1(n4932), .B2(n138), .ZN(
        n4440) );
  CKND2D0BWP12T U746 ( .A1(n2930), .A2(n3995), .ZN(n139) );
  MOAI22D0BWP12T U747 ( .A1(n2886), .A2(n139), .B1(n2886), .B2(n139), .ZN(
        n4503) );
  OAI21D0BWP12T U748 ( .A1(n3604), .A2(n4588), .B(n3350), .ZN(n140) );
  AO211D1BWP12T U749 ( .A1(n4094), .A2(n4778), .B(n3349), .C(n140), .Z(n3371)
         );
  NR2D0BWP12T U750 ( .A1(n4704), .A2(n3524), .ZN(n141) );
  AOI211D0BWP12T U751 ( .A1(n5078), .A2(n4444), .B(n141), .C(n3525), .ZN(n142)
         );
  CKND0BWP12T U752 ( .I(n5102), .ZN(n143) );
  AOI22D1BWP12T U753 ( .A1(n4388), .A2(n5088), .B1(n4574), .B2(n143), .ZN(n144) );
  OA211D1BWP12T U754 ( .A1(n4581), .A2(n3526), .B(n142), .C(n144), .Z(n3541)
         );
  CKND0BWP12T U755 ( .I(n4962), .ZN(n145) );
  MOAI22D0BWP12T U756 ( .A1(n4954), .A2(n145), .B1(n4898), .B2(n5099), .ZN(
        n3314) );
  MOAI22D0BWP12T U757 ( .A1(n4914), .A2(n2623), .B1(n4914), .B2(n2623), .ZN(
        n146) );
  OAI22D0BWP12T U758 ( .A1(n2624), .A2(n146), .B1(n306), .B2(n2626), .ZN(n2639) );
  CKND0BWP12T U759 ( .I(n3633), .ZN(n147) );
  OA21D0BWP12T U760 ( .A1(n3627), .A2(n147), .B(n3632), .Z(n819) );
  AOI21D0BWP12T U761 ( .A1(n1769), .A2(n971), .B(n4110), .ZN(n148) );
  CKND2D0BWP12T U762 ( .A1(n4108), .A2(n4109), .ZN(n149) );
  MAOI22D0BWP12T U763 ( .A1(n148), .A2(n149), .B1(n148), .B2(n149), .ZN(n4953)
         );
  AO22D1BWP12T U764 ( .A1(n3051), .A2(n4518), .B1(n4742), .B2(n3767), .Z(n3224) );
  OAI222D0BWP12T U765 ( .A1(n3945), .A2(n1821), .B1(n3812), .B2(n3447), .C1(
        n3813), .C2(n1822), .ZN(n150) );
  AOI21D0BWP12T U766 ( .A1(n3107), .A2(n3458), .B(n150), .ZN(n3938) );
  CKND2D0BWP12T U767 ( .A1(n2970), .A2(n3889), .ZN(n151) );
  NR2D0BWP12T U768 ( .A1(n2965), .A2(n151), .ZN(n152) );
  CKND0BWP12T U769 ( .I(n4367), .ZN(n153) );
  CKND0BWP12T U770 ( .I(n3888), .ZN(n154) );
  AOI21D0BWP12T U771 ( .A1(n2970), .A2(n154), .B(n2969), .ZN(n155) );
  CKND2D0BWP12T U772 ( .A1(n152), .A2(n3910), .ZN(n156) );
  OAI211D0BWP12T U773 ( .A1(n2966), .A2(n151), .B(n155), .C(n156), .ZN(n157)
         );
  AOI31D0BWP12T U774 ( .A1(n152), .A2(n3907), .A3(n153), .B(n157), .ZN(n158)
         );
  MAOI22D0BWP12T U775 ( .A1(n158), .A2(n2971), .B1(n158), .B2(n2971), .ZN(
        n4412) );
  CKND2D0BWP12T U776 ( .A1(n3590), .A2(n3589), .ZN(n159) );
  MAOI22D0BWP12T U777 ( .A1(n3555), .A2(n159), .B1(n3555), .B2(n159), .ZN(
        n4416) );
  CKND2D0BWP12T U778 ( .A1(n3360), .A2(n1784), .ZN(n160) );
  AOI32D0BWP12T U779 ( .A1(n1788), .A2(n4133), .A3(n4132), .B1(n1770), .B2(
        n4133), .ZN(n161) );
  MOAI22D0BWP12T U780 ( .A1(n160), .A2(n161), .B1(n160), .B2(n161), .ZN(n4322)
         );
  CKND0BWP12T U781 ( .I(n4384), .ZN(n162) );
  OAI21D0BWP12T U782 ( .A1(n4378), .A2(n162), .B(n4381), .ZN(n163) );
  MOAI22D0BWP12T U783 ( .A1(n3287), .A2(n163), .B1(n3287), .B2(n163), .ZN(
        n4387) );
  INR3D0BWP12T U784 ( .A1(n4818), .B1(n4817), .B2(n4843), .ZN(n4545) );
  IIND4D0BWP12T U785 ( .A1(n4058), .A2(n4057), .B1(n4680), .B2(n4448), .ZN(
        n164) );
  MAOI22D0BWP12T U786 ( .A1(n2666), .A2(n164), .B1(n2666), .B2(n164), .ZN(
        n4439) );
  IOA21D0BWP12T U787 ( .A1(n4696), .A2(n2885), .B(n3989), .ZN(n165) );
  NR2D0BWP12T U788 ( .A1(n3928), .A2(n3929), .ZN(n166) );
  CKND0BWP12T U789 ( .I(n4353), .ZN(n167) );
  AOI32D0BWP12T U790 ( .A1(n3930), .A2(n166), .A3(n167), .B1(n3933), .B2(n166), 
        .ZN(n168) );
  OAI211D0BWP12T U791 ( .A1(n3928), .A2(n3932), .B(n3931), .C(n168), .ZN(n169)
         );
  MOAI22D0BWP12T U792 ( .A1(n165), .A2(n169), .B1(n165), .B2(n169), .ZN(n4315)
         );
  CKND2D0BWP12T U793 ( .A1(n4492), .A2(n4491), .ZN(n170) );
  MAOI22D0BWP12T U794 ( .A1(n4493), .A2(n170), .B1(n4493), .B2(n170), .ZN(
        n5030) );
  AOI22D0BWP12T U795 ( .A1(n4103), .A2(n5089), .B1(n5087), .B2(n5088), .ZN(
        n171) );
  OAI22D0BWP12T U796 ( .A1(n5082), .A2(n5081), .B1(n5084), .B2(n5083), .ZN(
        n172) );
  MUX2ND0BWP12T U797 ( .I0(n5077), .I1(n5076), .S(n5075), .ZN(n173) );
  NR3D0BWP12T U798 ( .A1(n905), .A2(n5078), .A3(n173), .ZN(n174) );
  MUX2ND0BWP12T U799 ( .I0(n174), .I1(n5080), .S(n5079), .ZN(n175) );
  AOI211D0BWP12T U800 ( .A1(n5085), .A2(n5086), .B(n172), .C(n175), .ZN(n176)
         );
  AOI22D0BWP12T U801 ( .A1(n5090), .A2(n5091), .B1(n5092), .B2(n5093), .ZN(
        n177) );
  CKND0BWP12T U802 ( .I(n5098), .ZN(n178) );
  AOI22D0BWP12T U803 ( .A1(n5074), .A2(n178), .B1(n5097), .B2(n5096), .ZN(n179) );
  ND4D0BWP12T U804 ( .A1(n171), .A2(n176), .A3(n177), .A4(n179), .ZN(n180) );
  AOI21D0BWP12T U805 ( .A1(n5095), .A2(n5094), .B(n180), .ZN(n181) );
  OAI21D0BWP12T U806 ( .A1(n5100), .A2(n5101), .B(n5099), .ZN(n182) );
  OAI211D0BWP12T U807 ( .A1(n5103), .A2(n5102), .B(n181), .C(n182), .ZN(
        result[0]) );
  MOAI22D0BWP12T U808 ( .A1(n288), .A2(b[26]), .B1(n288), .B2(b[26]), .ZN(n183) );
  OAI22D0BWP12T U809 ( .A1(n2647), .A2(n183), .B1(n2648), .B2(n2649), .ZN(
        n2650) );
  MOAI22D0BWP12T U810 ( .A1(n4729), .A2(n5014), .B1(n4729), .B2(n5014), .ZN(
        n184) );
  OAI22D0BWP12T U811 ( .A1(n2739), .A2(n184), .B1(n2740), .B2(n2741), .ZN(
        n2752) );
  CKND2D0BWP12T U812 ( .A1(n3781), .A2(n3783), .ZN(n185) );
  CKND2D0BWP12T U813 ( .A1(n3784), .A2(n3783), .ZN(n186) );
  OAI211D0BWP12T U814 ( .A1(n4367), .A2(n185), .B(n3782), .C(n186), .ZN(n187)
         );
  MOAI22D0BWP12T U815 ( .A1(n3785), .A2(n187), .B1(n3785), .B2(n187), .ZN(
        n4410) );
  CKND0BWP12T U816 ( .I(n4742), .ZN(n188) );
  OAI221D0BWP12T U817 ( .A1(n4742), .A2(n5077), .B1(n188), .B2(n5076), .C(
        n5081), .ZN(n189) );
  MUX2ND0BWP12T U818 ( .I0(n189), .I1(n5048), .S(n373), .ZN(n967) );
  CKND0BWP12T U819 ( .I(n4586), .ZN(n190) );
  OAI22D0BWP12T U820 ( .A1(n4064), .A2(n3902), .B1(n4611), .B2(n3901), .ZN(
        n191) );
  AOI211D0BWP12T U821 ( .A1(n4843), .A2(n190), .B(n4156), .C(n191), .ZN(n4601)
         );
  AOI222D0BWP12T U822 ( .A1(n3937), .A2(n3811), .B1(n3940), .B2(n3119), .C1(
        n3810), .C2(n3939), .ZN(n192) );
  IOA21D0BWP12T U823 ( .A1(n3941), .A2(n2918), .B(n192), .ZN(n2859) );
  AOI21D0BWP12T U824 ( .A1(n3830), .A2(n2970), .B(n2969), .ZN(n193) );
  MAOI22D0BWP12T U825 ( .A1(n193), .A2(n2971), .B1(n193), .B2(n2971), .ZN(
        n4510) );
  MOAI22D0BWP12T U826 ( .A1(n4743), .A2(n3762), .B1(n4743), .B2(n4583), .ZN(
        n5020) );
  IND2D0BWP12T U827 ( .A1(n3551), .B1(n3552), .ZN(n194) );
  MAOI22D0BWP12T U828 ( .A1(n3553), .A2(n194), .B1(n3553), .B2(n194), .ZN(
        n4946) );
  IND2D0BWP12T U829 ( .A1(n3277), .B1(n3972), .ZN(n4829) );
  CKND0BWP12T U830 ( .I(n4628), .ZN(n195) );
  OAI32D0BWP12T U831 ( .A1(n195), .A2(n2746), .A3(n5083), .B1(n5081), .B2(n195), .ZN(n196) );
  CKND0BWP12T U832 ( .I(n4741), .ZN(n197) );
  CKND0BWP12T U833 ( .I(n905), .ZN(n198) );
  OAI221D0BWP12T U834 ( .A1(n4741), .A2(n5077), .B1(n197), .B2(n5076), .C(n198), .ZN(n199) );
  MAOI22D0BWP12T U835 ( .A1(n4627), .A2(n5080), .B1(n4627), .B2(n199), .ZN(
        n200) );
  AOI211D0BWP12T U836 ( .A1(n4433), .A2(n5078), .B(n196), .C(n200), .ZN(n3350)
         );
  IND2D0BWP12T U837 ( .A1(n4542), .B1(n4843), .ZN(n4785) );
  CKND2D0BWP12T U838 ( .A1(n3598), .A2(n3600), .ZN(n201) );
  CKND2D0BWP12T U839 ( .A1(n3601), .A2(n3600), .ZN(n202) );
  OAI211D0BWP12T U840 ( .A1(n4244), .A2(n201), .B(n3599), .C(n202), .ZN(n203)
         );
  MOAI22D0BWP12T U841 ( .A1(n3654), .A2(n203), .B1(n3654), .B2(n203), .ZN(
        n4324) );
  IND3D0BWP12T U842 ( .A1(n3606), .B1(n3233), .B2(n4631), .ZN(n204) );
  MAOI22D0BWP12T U843 ( .A1(n288), .A2(n204), .B1(n288), .B2(n204), .ZN(n4431)
         );
  AOI21D0BWP12T U844 ( .A1(n897), .A2(n4030), .B(n1623), .ZN(n205) );
  IND2D0BWP12T U845 ( .A1(n4049), .B1(n4384), .ZN(n206) );
  CKND2D0BWP12T U846 ( .A1(n893), .A2(n4030), .ZN(n207) );
  AOI32D0BWP12T U847 ( .A1(n4052), .A2(n205), .A3(n206), .B1(n207), .B2(n205), 
        .ZN(n208) );
  CKND2D0BWP12T U848 ( .A1(n4183), .A2(n1642), .ZN(n209) );
  MOAI22D0BWP12T U849 ( .A1(n208), .A2(n209), .B1(n208), .B2(n209), .ZN(n4406)
         );
  NR2D0BWP12T U850 ( .A1(n3488), .A2(n4458), .ZN(n210) );
  AOI211D0BWP12T U851 ( .A1(n3488), .A2(n4458), .B(n4420), .C(n210), .ZN(n3489) );
  OAI21D0BWP12T U852 ( .A1(n4247), .A2(n4817), .B(n4246), .ZN(n211) );
  CKND2D0BWP12T U853 ( .A1(n4582), .A2(n4249), .ZN(n212) );
  ND3D0BWP12T U854 ( .A1(n212), .A2(n211), .A3(n4250), .ZN(n4254) );
  MOAI22D0BWP12T U855 ( .A1(n2746), .A2(n4733), .B1(n2746), .B2(n4733), .ZN(
        n213) );
  OAI22D0BWP12T U856 ( .A1(n2747), .A2(n213), .B1(n2748), .B2(n2749), .ZN(
        n2750) );
  IND2D0BWP12T U857 ( .A1(n3770), .B1(n3142), .ZN(n1829) );
  IND2D0BWP12T U858 ( .A1(n2746), .B1(n1765), .ZN(n3605) );
  XOR3D1BWP12T U859 ( .A1(n2763), .A2(n2762), .A3(n2761), .Z(n321) );
  OAI21D1BWP12T U860 ( .A1(n2774), .A2(n2773), .B(n2772), .ZN(n2775) );
  CKND0BWP12T U861 ( .I(n2593), .ZN(n214) );
  OAI21D0BWP12T U862 ( .A1(n1512), .A2(n214), .B(n2646), .ZN(n4237) );
  CKND0BWP12T U863 ( .I(n4476), .ZN(n215) );
  AO21D0BWP12T U864 ( .A1(n3037), .A2(n215), .B(n3038), .Z(n3887) );
  CKND0BWP12T U865 ( .I(n4739), .ZN(n216) );
  CKND0BWP12T U866 ( .I(n905), .ZN(n217) );
  OAI221D0BWP12T U867 ( .A1(n4739), .A2(n5077), .B1(n216), .B2(n5076), .C(n217), .ZN(n218) );
  MAOI22D0BWP12T U868 ( .A1(n3850), .A2(n5080), .B1(n3850), .B2(n218), .ZN(
        n3851) );
  MAOI22D0BWP12T U869 ( .A1(n3051), .A2(n4036), .B1(n3051), .B2(n4035), .ZN(
        n3694) );
  OAI21D0BWP12T U870 ( .A1(n3029), .A2(n4354), .B(n3030), .ZN(n219) );
  AOI21D0BWP12T U871 ( .A1(n4350), .A2(n1599), .B(n219), .ZN(n3872) );
  CKND0BWP12T U872 ( .I(n3972), .ZN(n220) );
  OAI21D0BWP12T U873 ( .A1(n3464), .A2(n3463), .B(n4158), .ZN(n221) );
  OAI211D1BWP12T U874 ( .A1(n4064), .A2(n220), .B(n4573), .C(n221), .ZN(n222)
         );
  AOI211D1BWP12T U875 ( .A1(n3467), .A2(n3761), .B(n4470), .C(n222), .ZN(n223)
         );
  OA21D1BWP12T U876 ( .A1(n4586), .A2(n3969), .B(n223), .Z(n4600) );
  CKND0BWP12T U877 ( .I(n3997), .ZN(n224) );
  AO21D0BWP12T U878 ( .A1(n3993), .A2(n224), .B(n3996), .Z(n2931) );
  CKND2D0BWP12T U879 ( .A1(n4109), .A2(n4110), .ZN(n225) );
  OAI211D0BWP12T U880 ( .A1(n4486), .A2(n4111), .B(n4108), .C(n225), .ZN(n226)
         );
  CKND2D0BWP12T U881 ( .A1(n4112), .A2(n4134), .ZN(n227) );
  MOAI22D0BWP12T U882 ( .A1(n226), .A2(n227), .B1(n226), .B2(n227), .ZN(n4957)
         );
  OAI21D0BWP12T U883 ( .A1(n4102), .A2(n3626), .B(n3629), .ZN(n228) );
  CKND2D0BWP12T U884 ( .A1(n3627), .A2(n3366), .ZN(n229) );
  MOAI22D0BWP12T U885 ( .A1(n228), .A2(n229), .B1(n228), .B2(n229), .ZN(n4485)
         );
  CKND2D0BWP12T U886 ( .A1(n3529), .A2(n3498), .ZN(n230) );
  MOAI22D0BWP12T U887 ( .A1(n4333), .A2(n230), .B1(n4333), .B2(n230), .ZN(
        n4343) );
  MAOI22D0BWP12T U888 ( .A1(n3902), .A2(n3520), .B1(n3902), .B2(n4248), .ZN(
        n4581) );
  OAI222D0BWP12T U889 ( .A1(n3945), .A2(n3098), .B1(n3812), .B2(n3121), .C1(
        n3813), .C2(n3096), .ZN(n231) );
  AOI21D0BWP12T U890 ( .A1(n3941), .A2(n3104), .B(n231), .ZN(n3203) );
  CKND0BWP12T U891 ( .I(n295), .ZN(n232) );
  CKND0BWP12T U892 ( .I(n905), .ZN(n233) );
  OAI32D0BWP12T U893 ( .A1(n232), .A2(n4926), .A3(n5083), .B1(n233), .B2(n232), 
        .ZN(n234) );
  OAI221D0BWP12T U894 ( .A1(n295), .A2(n5077), .B1(n232), .B2(n5076), .C(n233), 
        .ZN(n235) );
  MAOI22D0BWP12T U895 ( .A1(n4653), .A2(n5080), .B1(n4653), .B2(n235), .ZN(
        n236) );
  AOI211D0BWP12T U896 ( .A1(n5078), .A2(n4453), .B(n234), .C(n236), .ZN(n3188)
         );
  IAO21D0BWP12T U897 ( .A1(n1673), .A2(n3509), .B(n1674), .ZN(n4540) );
  IND2D0BWP12T U898 ( .A1(n3846), .B1(n2901), .ZN(n237) );
  MAOI22D0BWP12T U899 ( .A1(n3040), .A2(n237), .B1(n3040), .B2(n237), .ZN(
        n4438) );
  CKND2D0BWP12T U900 ( .A1(n2928), .A2(n3989), .ZN(n238) );
  MOAI22D0BWP12T U901 ( .A1(n2929), .A2(n238), .B1(n2929), .B2(n238), .ZN(
        n4945) );
  ND3D0BWP12T U902 ( .A1(n4384), .A2(n3206), .A3(n3205), .ZN(n239) );
  OAI211D0BWP12T U903 ( .A1(n3208), .A2(n4052), .B(n3207), .C(n239), .ZN(n240)
         );
  MAOI22D0BWP12T U904 ( .A1(n3209), .A2(n240), .B1(n3209), .B2(n240), .ZN(
        n4393) );
  MOAI22D0BWP12T U905 ( .A1(n4924), .A2(n2619), .B1(n4924), .B2(n2619), .ZN(
        n241) );
  OAI22D0BWP12T U906 ( .A1(n2620), .A2(n241), .B1(n2621), .B2(n2622), .ZN(
        n2640) );
  MOAI22D0BWP12T U907 ( .A1(n4699), .A2(n4749), .B1(n4699), .B2(n4749), .ZN(
        n242) );
  OAI22D0BWP12T U908 ( .A1(n2678), .A2(n242), .B1(n2676), .B2(n2677), .ZN(
        n2697) );
  MOAI22D0BWP12T U909 ( .A1(n2742), .A2(n4727), .B1(n2742), .B2(n4727), .ZN(
        n243) );
  OAI22D0BWP12T U910 ( .A1(n2743), .A2(n243), .B1(n2744), .B2(n2745), .ZN(
        n2751) );
  IND2D0BWP12T U911 ( .A1(n1917), .B1(n1918), .ZN(n1915) );
  OAI21D0BWP12T U912 ( .A1(n2588), .A2(n2587), .B(n2586), .ZN(n2590) );
  INR2D0BWP12T U913 ( .A1(n3128), .B1(n4848), .ZN(n3129) );
  IND2D0BWP12T U914 ( .A1(n2362), .B1(n2361), .ZN(n2249) );
  INR2D0BWP12T U915 ( .A1(n4923), .B1(n1829), .ZN(n1830) );
  MOAI22D0BWP12T U916 ( .A1(n2742), .A2(n4316), .B1(n2742), .B2(n4316), .ZN(
        n244) );
  OAI22D0BWP12T U917 ( .A1(n2744), .A2(n244), .B1(n2743), .B2(n377), .ZN(n382)
         );
  IIND4D0BWP12T U918 ( .A1(n2781), .A2(n3891), .B1(n4651), .B2(n4425), .ZN(
        n3708) );
  CKND2D0BWP12T U919 ( .A1(n3832), .A2(n3828), .ZN(n245) );
  OAI211D0BWP12T U920 ( .A1(n2801), .A2(n2800), .B(n3831), .C(n245), .ZN(n3695) );
  AOI21D0BWP12T U921 ( .A1(n5075), .A2(n962), .B(n4115), .ZN(n246) );
  IND2D0BWP12T U922 ( .A1(n4114), .B1(n963), .ZN(n247) );
  MAOI22D0BWP12T U923 ( .A1(n246), .A2(n247), .B1(n246), .B2(n247), .ZN(n4395)
         );
  AN2D0BWP12T U924 ( .A1(n2608), .A2(n2607), .Z(n2611) );
  OA21D0BWP12T U925 ( .A1(n4238), .A2(n4237), .B(n4239), .Z(n4259) );
  CKND0BWP12T U926 ( .I(n3176), .ZN(n248) );
  OA21D0BWP12T U927 ( .A1(n3172), .A2(n248), .B(n4071), .Z(n4015) );
  CKND0BWP12T U928 ( .I(n2259), .ZN(n249) );
  OAI21D0BWP12T U929 ( .A1(n2261), .A2(n249), .B(n2258), .ZN(n2260) );
  AN2D0BWP12T U930 ( .A1(n4103), .A2(n4495), .Z(n4104) );
  CKND0BWP12T U931 ( .I(n4743), .ZN(n250) );
  OAI21D0BWP12T U932 ( .A1(n3752), .A2(n250), .B(n3769), .ZN(n4824) );
  INR2D0BWP12T U933 ( .A1(n4586), .B1(n3604), .ZN(n3613) );
  CKND0BWP12T U934 ( .I(n3618), .ZN(n251) );
  CKND0BWP12T U935 ( .I(n3231), .ZN(n252) );
  CKND2D0BWP12T U936 ( .A1(n3620), .A2(n252), .ZN(n253) );
  IOA21D0BWP12T U937 ( .A1(n252), .A2(n3619), .B(n3632), .ZN(n254) );
  AOI31D0BWP12T U938 ( .A1(n3621), .A2(n3620), .A3(n252), .B(n254), .ZN(n255)
         );
  OAI31D0BWP12T U939 ( .A1(n5082), .A2(n251), .A3(n253), .B(n255), .ZN(n256)
         );
  MOAI22D0BWP12T U940 ( .A1(n3232), .A2(n256), .B1(n3232), .B2(n256), .ZN(
        n4389) );
  CKND2D0BWP12T U941 ( .A1(n4448), .A2(n4655), .ZN(n257) );
  MAOI22D0BWP12T U942 ( .A1(n4906), .A2(n257), .B1(n4906), .B2(n257), .ZN(
        n4444) );
  CKND0BWP12T U943 ( .I(n3278), .ZN(n258) );
  OAI32D0BWP12T U944 ( .A1(n258), .A2(n4543), .A3(n5040), .B1(n5098), .B2(n258), .ZN(n3281) );
  OAI22D0BWP12T U945 ( .A1(n3945), .A2(n3061), .B1(n3812), .B2(n3099), .ZN(
        n259) );
  AOI21D0BWP12T U946 ( .A1(n3107), .A2(n3114), .B(n259), .ZN(n3557) );
  AOI21D0BWP12T U947 ( .A1(n3199), .A2(n4023), .B(n4026), .ZN(n260) );
  MOAI22D0BWP12T U948 ( .A1(n260), .A2(n3209), .B1(n260), .B2(n3209), .ZN(
        n4480) );
  AO22D0BWP12T U949 ( .A1(n4960), .A2(n5093), .B1(n5090), .B2(n4341), .Z(n4194) );
  CKND2D0BWP12T U950 ( .A1(n3428), .A2(n3429), .ZN(n261) );
  MOAI22D0BWP12T U951 ( .A1(n3430), .A2(n261), .B1(n3430), .B2(n261), .ZN(
        n4994) );
  CKND2D0BWP12T U952 ( .A1(n2930), .A2(n3995), .ZN(n262) );
  MOAI22D0BWP12T U953 ( .A1(n2931), .A2(n262), .B1(n2931), .B2(n262), .ZN(
        n4413) );
  CKND0BWP12T U954 ( .I(n3598), .ZN(n263) );
  CKND0BWP12T U955 ( .I(n3412), .ZN(n264) );
  CKND2D0BWP12T U956 ( .A1(n3409), .A2(n264), .ZN(n265) );
  OAI21D0BWP12T U957 ( .A1(n3412), .A2(n3413), .B(n3411), .ZN(n266) );
  AOI31D0BWP12T U958 ( .A1(n3601), .A2(n3409), .A3(n264), .B(n266), .ZN(n267)
         );
  OAI31D0BWP12T U959 ( .A1(n4244), .A2(n263), .A3(n265), .B(n267), .ZN(n268)
         );
  MOAI22D0BWP12T U960 ( .A1(n3414), .A2(n268), .B1(n3414), .B2(n268), .ZN(
        n4328) );
  OR4D0BWP12T U961 ( .A1(n4311), .A2(n4312), .A3(n4313), .A4(n4315), .Z(n269)
         );
  NR2D0BWP12T U962 ( .A1(n4314), .A2(n269), .ZN(n5005) );
  AN2D0BWP12T U963 ( .A1(n5090), .A2(n4322), .Z(n1789) );
  CKND0BWP12T U964 ( .I(n2808), .ZN(n270) );
  AOI222D0BWP12T U965 ( .A1(n270), .A2(n4103), .B1(n2794), .B2(n5088), .C1(
        n3488), .C2(n5078), .ZN(n2841) );
  IND2D0BWP12T U966 ( .A1(op[2]), .B1(n2870), .ZN(n5076) );
  AO21D0BWP12T U967 ( .A1(n5099), .A2(n4865), .B(n4548), .Z(n4212) );
  AO21D4BWP12T U968 ( .A1(n5009), .A2(n5085), .B(n3485), .Z(result[30]) );
  INVD2BWP12T U969 ( .I(n3420), .ZN(n3545) );
  XOR2XD4BWP12T U970 ( .A1(n2094), .A2(n272), .Z(n2035) );
  TPNR2D2BWP12T U971 ( .A1(n2511), .A2(n2510), .ZN(n3671) );
  OR2XD1BWP12T U972 ( .A1(n2521), .A2(n2520), .Z(n274) );
  TPOAI22D2BWP12T U973 ( .A1(n674), .A2(n673), .B1(n672), .B2(n671), .ZN(n726)
         );
  AO21D2BWP12T U974 ( .A1(n4281), .A2(n5085), .B(n4198), .Z(result[16]) );
  CKND2D2BWP12T U975 ( .A1(n2486), .A2(n2485), .ZN(n2495) );
  IOA21D2BWP12T U976 ( .A1(n2482), .A2(n2481), .B(n2480), .ZN(n2486) );
  INVD1BWP12T U977 ( .I(n2172), .ZN(n347) );
  DCCKND4BWP12T U978 ( .I(n852), .ZN(n2172) );
  XNR2XD4BWP12T U979 ( .A1(n2172), .A2(n5014), .ZN(n1093) );
  XNR2D2BWP12T U980 ( .A1(n2172), .A2(n2742), .ZN(n470) );
  TPND2D2BWP12T U981 ( .A1(n2404), .A2(n2405), .ZN(n2274) );
  NR2D2BWP12T U982 ( .A1(n2404), .A2(n2405), .ZN(n2275) );
  TPOAI22D1BWP12T U983 ( .A1(n2266), .A2(n2265), .B1(n2264), .B2(n2263), .ZN(
        n2372) );
  IOA21D1BWP12T U984 ( .A1(n2262), .A2(n2261), .B(n2260), .ZN(n2347) );
  XNR2XD2BWP12T U985 ( .A1(n2623), .A2(n288), .ZN(n1159) );
  XNR2XD2BWP12T U986 ( .A1(n2623), .A2(n2593), .ZN(n608) );
  NR2D1BWP12T U987 ( .A1(n321), .A2(n2770), .ZN(n2773) );
  INVD1BWP12T U988 ( .I(n1949), .ZN(n1942) );
  OAI21D0BWP12T U989 ( .A1(n2545), .A2(n2544), .B(n2542), .ZN(n2543) );
  ND2D4BWP12T U990 ( .A1(n992), .A2(n5075), .ZN(n275) );
  INVD12BWP12T U991 ( .I(n275), .ZN(n3218) );
  ND2D1BWP12T U992 ( .A1(n3306), .A2(n3305), .ZN(n3315) );
  AO21D4BWP12T U993 ( .A1(n4289), .A2(n5085), .B(n3019), .Z(result[24]) );
  NR4D0BWP12T U994 ( .A1(n4289), .A2(n4288), .A3(n4287), .A4(n4286), .ZN(n4298) );
  AN2D1BWP12T U995 ( .A1(n3673), .A2(n3672), .Z(n3674) );
  OR2XD1BWP12T U996 ( .A1(n1493), .A2(n1492), .Z(n277) );
  TPOAI21D4BWP12T U997 ( .A1(n1406), .A2(n1405), .B(n1404), .ZN(n1492) );
  TPND2D1BWP12T U998 ( .A1(n1570), .A2(n1571), .ZN(n1568) );
  TPOAI22D2BWP12T U999 ( .A1(n429), .A2(n2646), .B1(n4257), .B2(n472), .ZN(
        n476) );
  RCAOI21D4BWP12T U1000 ( .A1(n2205), .A2(n2195), .B(n2194), .ZN(n2203) );
  CKND2D2BWP12T U1001 ( .A1(n1579), .A2(n1578), .ZN(n1580) );
  TPND2D3BWP12T U1002 ( .A1(n1452), .A2(n1451), .ZN(n1579) );
  TPND2D1BWP12T U1003 ( .A1(n2316), .A2(n2317), .ZN(n297) );
  INVD1BWP12T U1004 ( .I(n394), .ZN(n278) );
  TPOAI22D1BWP12T U1005 ( .A1(n2037), .A2(n2624), .B1(n305), .B2(n1930), .ZN(
        n2041) );
  CKND2D2BWP12T U1006 ( .A1(n393), .A2(n392), .ZN(n3340) );
  TPND2D1BWP12T U1007 ( .A1(n1507), .A2(n1506), .ZN(n1511) );
  TPND2D1BWP12T U1008 ( .A1(n1862), .A2(n1879), .ZN(n1865) );
  OAI22D4BWP12T U1009 ( .A1(n642), .A2(n2319), .B1(n609), .B2(n2702), .ZN(n659) );
  BUFFXD4BWP12T U1010 ( .I(b[17]), .Z(n279) );
  BUFFXD3BWP12T U1011 ( .I(b[17]), .Z(n280) );
  BUFFD2BWP12T U1012 ( .I(b[17]), .Z(n4763) );
  ND2D1BWP12T U1013 ( .A1(n1874), .A2(n1873), .ZN(n281) );
  TPND2D3BWP12T U1014 ( .A1(n1874), .A2(n1873), .ZN(n2043) );
  IOA21D2BWP12T U1015 ( .A1(n2197), .A2(n2198), .B(n2124), .ZN(n2606) );
  OAI22D1BWP12T U1016 ( .A1(n1974), .A2(n1903), .B1(n1902), .B2(n1901), .ZN(
        n2574) );
  IND3D4BWP12T U1017 ( .A1(n2631), .B1(n1884), .B2(n2634), .ZN(n1885) );
  OAI21D2BWP12T U1018 ( .A1(n2477), .A2(n2470), .B(n2469), .ZN(n282) );
  OAI21D2BWP12T U1019 ( .A1(n2477), .A2(n2470), .B(n2469), .ZN(n2506) );
  XOR3XD4BWP12T U1020 ( .A1(n1950), .A2(n1949), .A3(n1948), .Z(n283) );
  ND3D2BWP12T U1021 ( .A1(n285), .A2(n286), .A3(n287), .ZN(n1950) );
  TPOAI22D4BWP12T U1022 ( .A1(n2322), .A2(n2743), .B1(n1550), .B2(n2744), .ZN(
        n2327) );
  INVD1BWP12T U1023 ( .I(n1484), .ZN(n1486) );
  XNR2XD2BWP12T U1024 ( .A1(n2167), .A2(n2742), .ZN(n537) );
  XNR2XD4BWP12T U1025 ( .A1(n2167), .A2(n4914), .ZN(n1930) );
  NR2XD2BWP12T U1026 ( .A1(n1939), .A2(n1938), .ZN(n2045) );
  XOR3D2BWP12T U1027 ( .A1(n1961), .A2(n1960), .A3(n1959), .Z(n2126) );
  ND2D1BWP12T U1028 ( .A1(n1961), .A2(n1960), .ZN(n285) );
  ND2D1BWP12T U1029 ( .A1(n1961), .A2(n1959), .ZN(n286) );
  ND2D1BWP12T U1030 ( .A1(n1960), .A2(n1959), .ZN(n287) );
  OAI21D1BWP12T U1031 ( .A1(n2130), .A2(n2131), .B(n2128), .ZN(n2009) );
  TPOAI22D4BWP12T U1032 ( .A1(n1909), .A2(n2689), .B1(n2027), .B2(n2691), .ZN(
        n2034) );
  OAI22D4BWP12T U1033 ( .A1(n1515), .A2(n2643), .B1(n1894), .B2(n1856), .ZN(
        n2261) );
  TPOAI22D2BWP12T U1034 ( .A1(n1983), .A2(n2641), .B1(n1895), .B2(n2643), .ZN(
        n1955) );
  XNR2XD8BWP12T U1035 ( .A1(n4914), .A2(n4728), .ZN(n2643) );
  CKND0BWP12T U1036 ( .I(n2401), .ZN(n2386) );
  TPNR2D3BWP12T U1037 ( .A1(n2519), .A2(n2518), .ZN(n3547) );
  DCCKND4BWP12T U1038 ( .I(n1402), .ZN(n345) );
  BUFFXD8BWP12T U1039 ( .I(a[7]), .Z(n288) );
  XNR2D2BWP12T U1040 ( .A1(n3088), .A2(n3087), .ZN(n4284) );
  INVD3BWP12T U1041 ( .I(n1785), .ZN(n289) );
  INVD2BWP12T U1042 ( .I(n4560), .ZN(n1785) );
  TPND2D3BWP12T U1043 ( .A1(n1390), .A2(n1389), .ZN(n1446) );
  INR2XD2BWP12T U1044 ( .A1(n4316), .B1(n2634), .ZN(n1984) );
  OAI22D4BWP12T U1045 ( .A1(n1933), .A2(n2632), .B1(n2018), .B2(n2634), .ZN(
        n2060) );
  TPND2D1BWP12T U1046 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2XD4BWP12T U1047 ( .A1(n2071), .A2(n1883), .Z(n1929) );
  INVD4BWP12T U1048 ( .I(n4699), .ZN(n1883) );
  ND2D4BWP12T U1049 ( .A1(n2515), .A2(n2514), .ZN(n3921) );
  XNR2XD2BWP12T U1050 ( .A1(n2591), .A2(n2746), .ZN(n1994) );
  OAI22D0BWP12T U1051 ( .A1(n2037), .A2(n2624), .B1(n305), .B2(n1930), .ZN(
        n290) );
  TPNR2D1BWP12T U1052 ( .A1(n3846), .A2(n4907), .ZN(n3848) );
  BUFFXD3BWP12T U1053 ( .I(a[0]), .Z(n4910) );
  TPOAI21D1BWP12T U1054 ( .A1(n4293), .A2(n2447), .B(n2446), .ZN(n291) );
  TPOAI21D1BWP12T U1055 ( .A1(n4293), .A2(n2447), .B(n2446), .ZN(n3796) );
  OAI22D1BWP12T U1056 ( .A1(n1980), .A2(n2702), .B1(n1904), .B2(n2319), .ZN(
        n293) );
  OAI22D1BWP12T U1057 ( .A1(n1980), .A2(n2702), .B1(n1904), .B2(n2319), .ZN(
        n1967) );
  XNR2D1BWP12T U1058 ( .A1(n2243), .A2(n4906), .ZN(n1904) );
  NR2D4BWP12T U1059 ( .A1(n2509), .A2(n2508), .ZN(n3798) );
  XOR3D2BWP12T U1060 ( .A1(n2010), .A2(n294), .A3(n2121), .Z(n2196) );
  INVD2BWP12T U1061 ( .I(n2122), .ZN(n2010) );
  INVD3BWP12T U1062 ( .I(n2464), .ZN(n2336) );
  TPOAI22D2BWP12T U1063 ( .A1(n1561), .A2(n2647), .B1(n1442), .B2(n1441), .ZN(
        n335) );
  TPND2D1BWP12T U1064 ( .A1(n4303), .A2(n4302), .ZN(n4308) );
  TPND2D2BWP12T U1065 ( .A1(n2121), .A2(n2012), .ZN(n2015) );
  INVD2BWP12T U1066 ( .I(n1448), .ZN(n1450) );
  TPNR2D2BWP12T U1067 ( .A1(n283), .A2(n320), .ZN(n1972) );
  TPOAI21D1BWP12T U1068 ( .A1(n2344), .A2(n2346), .B(n2345), .ZN(n2239) );
  TPND2D1BWP12T U1069 ( .A1(n1469), .A2(n1468), .ZN(n1473) );
  XNR2D1BWP12T U1070 ( .A1(n848), .A2(n3748), .ZN(n2630) );
  TPNR2D2BWP12T U1071 ( .A1(n3051), .A2(n4912), .ZN(n975) );
  INVD4BWP12T U1072 ( .I(n610), .ZN(n296) );
  DCCKND8BWP12T U1073 ( .I(n1307), .ZN(n610) );
  OAI21D1BWP12T U1074 ( .A1(n3213), .A2(n826), .B(n825), .ZN(n3199) );
  AOI21D1BWP12T U1075 ( .A1(n2886), .A2(n3995), .B(n3994), .ZN(n3936) );
  TPND2D2BWP12T U1076 ( .A1(n1419), .A2(n1418), .ZN(n1564) );
  XNR2D2BWP12T U1077 ( .A1(n4761), .A2(n2679), .ZN(n1937) );
  XOR3XD4BWP12T U1078 ( .A1(n2316), .A2(n2317), .A3(n2315), .Z(n2434) );
  ND2D1BWP12T U1079 ( .A1(n2316), .A2(n2315), .ZN(n298) );
  ND2D1BWP12T U1080 ( .A1(n2317), .A2(n2315), .ZN(n299) );
  ND3D2BWP12T U1081 ( .A1(n297), .A2(n298), .A3(n299), .ZN(n2311) );
  INVD2BWP12T U1082 ( .I(n2311), .ZN(n2305) );
  TPND2D1BWP12T U1083 ( .A1(n2310), .A2(n2311), .ZN(n2307) );
  TPOAI22D2BWP12T U1084 ( .A1(n1439), .A2(n2682), .B1(n1340), .B2(n2680), .ZN(
        n1415) );
  TPND2D3BWP12T U1085 ( .A1(n2519), .A2(n2518), .ZN(n3549) );
  TPOAI22D2BWP12T U1086 ( .A1(n314), .A2(n4257), .B1(n2646), .B2(n1188), .ZN(
        n1378) );
  INVD2BWP12T U1087 ( .I(n4295), .ZN(n3920) );
  CKND2D2BWP12T U1088 ( .A1(n283), .A2(n320), .ZN(n1971) );
  OAI31D2BWP12T U1089 ( .A1(n5009), .A2(n5008), .A3(n5007), .B(n5006), .ZN(z)
         );
  TPOAI22D2BWP12T U1090 ( .A1(n1896), .A2(n2678), .B1(n2676), .B2(n2097), .ZN(
        n1954) );
  TPOAI22D1BWP12T U1091 ( .A1(n2324), .A2(n2646), .B1(n2166), .B2(n4257), .ZN(
        n2271) );
  DEL025D1BWP12T U1092 ( .I(n2528), .Z(n301) );
  XNR2D2BWP12T U1093 ( .A1(n2071), .A2(n4914), .ZN(n2223) );
  BUFFXD8BWP12T U1094 ( .I(b[4]), .Z(n2071) );
  INR2D2BWP12T U1095 ( .A1(n2504), .B1(n2503), .ZN(n302) );
  INR2D2BWP12T U1096 ( .A1(n2504), .B1(n2503), .ZN(n3794) );
  INVD2BWP12T U1097 ( .I(n3171), .ZN(n4008) );
  XNR2XD4BWP12T U1098 ( .A1(n764), .A2(n763), .ZN(n4282) );
  XNR2D2BWP12T U1099 ( .A1(n2742), .A2(b[20]), .ZN(n1550) );
  XNR2D2BWP12T U1100 ( .A1(b[20]), .A2(n2593), .ZN(n1367) );
  OAI21D1BWP12T U1101 ( .A1(n2313), .A2(n2314), .B(n2312), .ZN(n2294) );
  CKND2D2BWP12T U1102 ( .A1(n1569), .A2(n1568), .ZN(n1575) );
  ND2D3BWP12T U1103 ( .A1(n1495), .A2(n1494), .ZN(n2442) );
  XNR3XD4BWP12T U1104 ( .A1(n1944), .A2(n2605), .A3(n2606), .ZN(n303) );
  TPOAI22D2BWP12T U1105 ( .A1(n2320), .A2(n2319), .B1(n2318), .B2(n2702), .ZN(
        n2369) );
  TPNR2D1BWP12T U1106 ( .A1(n1583), .A2(n1582), .ZN(n304) );
  TPNR2D1BWP12T U1107 ( .A1(n1583), .A2(n1582), .ZN(n2443) );
  CKND2D2BWP12T U1108 ( .A1(n2379), .A2(n2381), .ZN(n2224) );
  TPND2D3BWP12T U1109 ( .A1(n1345), .A2(n1344), .ZN(n305) );
  TPND2D3BWP12T U1110 ( .A1(n1345), .A2(n1344), .ZN(n306) );
  TPND2D3BWP12T U1111 ( .A1(n1343), .A2(n1342), .ZN(n1345) );
  TPND2D2BWP12T U1112 ( .A1(n1345), .A2(n1344), .ZN(n2625) );
  TPND2D2BWP12T U1113 ( .A1(n307), .A2(n308), .ZN(n310) );
  TPND2D2BWP12T U1114 ( .A1(n309), .A2(n310), .ZN(n1032) );
  CKND3BWP12T U1115 ( .I(n2098), .ZN(n307) );
  BUFFXD8BWP12T U1116 ( .I(b[9]), .Z(n2098) );
  CKBD4BWP12T U1117 ( .I(n2098), .Z(n4765) );
  BUFFD2BWP12T U1118 ( .I(n4291), .Z(n311) );
  TPOAI22D1BWP12T U1119 ( .A1(n1340), .A2(n2682), .B1(n1304), .B2(n2680), .ZN(
        n1334) );
  AO21D0BWP12T U1120 ( .A1(n5085), .A2(n4300), .B(n4084), .Z(n) );
  XNR2XD2BWP12T U1121 ( .A1(b[3]), .A2(n4914), .ZN(n2222) );
  OA21XD0BWP12T U1122 ( .A1(n905), .A2(n3056), .B(n4726), .Z(n3057) );
  INVD2BWP12T U1123 ( .I(n1280), .ZN(n313) );
  INVD1BWP12T U1124 ( .I(n313), .ZN(n314) );
  XNR2XD8BWP12T U1125 ( .A1(n4764), .A2(n2593), .ZN(n1280) );
  TPND2D1BWP12T U1126 ( .A1(n1380), .A2(n1378), .ZN(n1381) );
  NR2D2BWP12T U1127 ( .A1(n4686), .A2(n4742), .ZN(n953) );
  TPOAI21D1BWP12T U1128 ( .A1(n4008), .A2(n1024), .B(n1027), .ZN(n764) );
  XOR2D1BWP12T U1129 ( .A1(n3664), .A2(n3663), .Z(n4266) );
  INVD1BWP12T U1130 ( .I(n2481), .ZN(n315) );
  TPND2D3BWP12T U1131 ( .A1(n1477), .A2(n1476), .ZN(n1481) );
  CKND2D2BWP12T U1132 ( .A1(n553), .A2(n552), .ZN(n691) );
  TPOAI22D2BWP12T U1133 ( .A1(n1936), .A2(n2740), .B1(n2058), .B2(n2739), .ZN(
        n2047) );
  OR2D2BWP12T U1134 ( .A1(n335), .A2(n1554), .Z(n316) );
  TPND2D2BWP12T U1135 ( .A1(n3797), .A2(n3795), .ZN(n3667) );
  INVD2BWP12T U1136 ( .I(n699), .ZN(n688) );
  INVD2BWP12T U1137 ( .I(n699), .ZN(n700) );
  XNR2XD2BWP12T U1138 ( .A1(n4738), .A2(n2701), .ZN(n504) );
  INVD12BWP12T U1139 ( .I(n2701), .ZN(n319) );
  ND2D4BWP12T U1140 ( .A1(n1075), .A2(n1074), .ZN(n1132) );
  BUFFXD0BWP12T U1141 ( .I(n853), .Z(n317) );
  INVD6BWP12T U1142 ( .I(b[5]), .ZN(n853) );
  XNR2XD2BWP12T U1143 ( .A1(n4761), .A2(n2593), .ZN(n1109) );
  XOR2XD4BWP12T U1144 ( .A1(n2094), .A2(n1810), .Z(n2233) );
  DCCKND12BWP12T U1145 ( .I(n1810), .ZN(n2688) );
  IOA21D1BWP12T U1146 ( .A1(n2203), .A2(n2204), .B(n2202), .ZN(n2199) );
  INVD1BWP12T U1147 ( .I(n1489), .ZN(n318) );
  NR2D2BWP12T U1148 ( .A1(n3022), .A2(n3020), .ZN(n3865) );
  INVD12BWP12T U1149 ( .I(n861), .ZN(n4926) );
  TPOAI22D4BWP12T U1150 ( .A1(n2173), .A2(n2220), .B1(n2218), .B2(n2221), .ZN(
        n2215) );
  TPOAI22D2BWP12T U1151 ( .A1(n1951), .A2(n2632), .B1(n348), .B2(n2634), .ZN(
        n1960) );
  XNR2XD2BWP12T U1152 ( .A1(n2072), .A2(n3040), .ZN(n348) );
  ND2D3BWP12T U1153 ( .A1(n2614), .A2(n2613), .ZN(n2844) );
  XNR2D2BWP12T U1154 ( .A1(n2578), .A2(n2742), .ZN(n2001) );
  BUFFXD8BWP12T U1155 ( .I(n2578), .Z(n4739) );
  XNR2XD4BWP12T U1156 ( .A1(n2094), .A2(n5014), .ZN(n1181) );
  OAI21D4BWP12T U1157 ( .A1(n1058), .A2(a[14]), .B(n1164), .ZN(n707) );
  XOR2XD4BWP12T U1158 ( .A1(n2071), .A2(n1342), .Z(n1548) );
  INVD12BWP12T U1159 ( .I(n1652), .ZN(n4924) );
  TPOAI22D1BWP12T U1160 ( .A1(n1177), .A2(n2702), .B1(n2319), .B2(n1351), .ZN(
        n1295) );
  XOR2XD4BWP12T U1161 ( .A1(n2094), .A2(n319), .Z(n329) );
  TPND2D2BWP12T U1162 ( .A1(n1970), .A2(n1969), .ZN(n320) );
  TPND2D2BWP12T U1163 ( .A1(n1970), .A2(n1969), .ZN(n2062) );
  TPND2D3BWP12T U1164 ( .A1(n1968), .A2(n2125), .ZN(n1970) );
  ND2XD0BWP12T U1165 ( .A1(n2148), .A2(n2147), .ZN(n2067) );
  ND2XD0BWP12T U1166 ( .A1(n1471), .A2(n1470), .ZN(n1472) );
  HA1D2BWP12T U1167 ( .A(n1356), .B(n1355), .CO(n1375), .S(n1301) );
  OA22D2BWP12T U1168 ( .A1(n2244), .A2(n2748), .B1(n2070), .B2(n2747), .Z(
        n2291) );
  BUFFD8BWP12T U1169 ( .I(n471), .Z(n2743) );
  TPND2D2BWP12T U1170 ( .A1(n1888), .A2(n1887), .ZN(n1978) );
  TPND2D2BWP12T U1171 ( .A1(n1457), .A2(n1456), .ZN(n1535) );
  TPND2D1BWP12T U1172 ( .A1(n4741), .A2(n3040), .ZN(n324) );
  TPND2D2BWP12T U1173 ( .A1(n322), .A2(n323), .ZN(n325) );
  CKND2D2BWP12T U1174 ( .A1(n324), .A2(n325), .ZN(n2633) );
  INVD2BWP12T U1175 ( .I(n4741), .ZN(n322) );
  TPAOI22D0BWP12T U1176 ( .A1(n289), .A2(n4562), .B1(n4561), .B2(n4921), .ZN(
        n4203) );
  TPOAI21D4BWP12T U1177 ( .A1(n1027), .A2(n1026), .B(n1025), .ZN(n1028) );
  TPOAI22D4BWP12T U1178 ( .A1(n670), .A2(n2744), .B1(n733), .B2(n2743), .ZN(
        n720) );
  XNR2XD4BWP12T U1179 ( .A1(n2619), .A2(n288), .ZN(n1360) );
  BUFFD6BWP12T U1180 ( .I(b[14]), .Z(n2619) );
  ND2D3BWP12T U1181 ( .A1(n424), .A2(n445), .ZN(n427) );
  IOA21D0BWP12T U1182 ( .A1(n1942), .A2(n1941), .B(n1948), .ZN(n1943) );
  NR2D2BWP12T U1183 ( .A1(n1024), .A2(n1026), .ZN(n1029) );
  XOR3XD4BWP12T U1184 ( .A1(n1950), .A2(n1949), .A3(n1948), .Z(n326) );
  ND2D3BWP12T U1185 ( .A1(n303), .A2(n2520), .ZN(n3425) );
  XOR3XD4BWP12T U1186 ( .A1(n2434), .A2(n2433), .A3(n2432), .Z(n327) );
  OAI22D1BWP12T U1187 ( .A1(n1936), .A2(n2740), .B1(n2058), .B2(n2739), .ZN(
        n328) );
  NR4D1BWP12T U1188 ( .A1(b[22]), .A2(n2591), .A3(n854), .A4(n2551), .ZN(n919)
         );
  OAI22D4BWP12T U1189 ( .A1(n642), .A2(n2702), .B1(n713), .B2(n2704), .ZN(n737) );
  TPNR2D1BWP12T U1190 ( .A1(n1176), .A2(n2702), .ZN(n1179) );
  TPOAI22D4BWP12T U1191 ( .A1(n608), .A2(n607), .B1(n657), .B2(n4257), .ZN(
        n649) );
  TPND2D2BWP12T U1192 ( .A1(n464), .A2(n463), .ZN(n3379) );
  CKND0BWP12T U1193 ( .I(n486), .ZN(n490) );
  XNR3XD4BWP12T U1194 ( .A1(n1944), .A2(n2605), .A3(n2606), .ZN(n2521) );
  INVD9BWP12T U1195 ( .I(n416), .ZN(n2094) );
  XNR2XD2BWP12T U1196 ( .A1(n2167), .A2(n4924), .ZN(n2095) );
  TPND2D1BWP12T U1197 ( .A1(n1888), .A2(n1887), .ZN(n330) );
  IOA21D1BWP12T U1198 ( .A1(n591), .A2(n590), .B(n589), .ZN(n595) );
  BUFFD12BWP12T U1199 ( .I(b[0]), .Z(n5075) );
  OA211D2BWP12T U1200 ( .A1(n4318), .A2(n3728), .B(n3727), .C(n3726), .Z(n3729) );
  TPNR2D2BWP12T U1201 ( .A1(n1361), .A2(n305), .ZN(n1362) );
  TPOAI21D4BWP12T U1202 ( .A1(n1501), .A2(n332), .B(n1499), .ZN(n1503) );
  TPNR2D2BWP12T U1203 ( .A1(n3424), .A2(n3547), .ZN(n2523) );
  OAI21D4BWP12T U1204 ( .A1(n4921), .A2(n4627), .B(n374), .ZN(n360) );
  NR2D4BWP12T U1205 ( .A1(n715), .A2(n714), .ZN(n1052) );
  TPNR2D2BWP12T U1206 ( .A1(n3733), .A2(n3731), .ZN(n2439) );
  INVD6BWP12T U1207 ( .I(b[1]), .ZN(n605) );
  TPND2D1BWP12T U1208 ( .A1(n1054), .A2(n1053), .ZN(n1055) );
  INVD1BWP12T U1209 ( .I(n1054), .ZN(n1049) );
  INVD4BWP12T U1210 ( .I(n2669), .ZN(n706) );
  FA1D4BWP12T U1211 ( .A(n520), .B(n519), .CI(n518), .CO(n578), .S(n522) );
  INVD12BWP12T U1212 ( .I(n411), .ZN(n412) );
  INVD12BWP12T U1213 ( .I(n411), .ZN(n2647) );
  TPNR2D1BWP12T U1214 ( .A1(n4300), .A2(n4299), .ZN(n4310) );
  BUFFXD4BWP12T U1215 ( .I(b[20]), .Z(n2243) );
  XNR2XD2BWP12T U1216 ( .A1(n4763), .A2(n4906), .ZN(n2242) );
  XNR2XD4BWP12T U1217 ( .A1(n5053), .A2(n5014), .ZN(n2563) );
  XNR2XD2BWP12T U1218 ( .A1(n2167), .A2(n2679), .ZN(n1340) );
  TPND2D2BWP12T U1219 ( .A1(n346), .A2(n1401), .ZN(n1390) );
  ND2D1BWP12T U1220 ( .A1(n2015), .A2(n2014), .ZN(n331) );
  XOR3XD4BWP12T U1221 ( .A1(n1998), .A2(n1997), .A3(n1996), .Z(n2130) );
  TPND2D2BWP12T U1222 ( .A1(n1436), .A2(n1435), .ZN(n332) );
  TPND2D2BWP12T U1223 ( .A1(n1436), .A2(n1435), .ZN(n1500) );
  TPOAI21D2BWP12T U1224 ( .A1(n3733), .A2(n3730), .B(n3734), .ZN(n2438) );
  XOR2D2BWP12T U1225 ( .A1(n901), .A2(b[21]), .Z(n1440) );
  OAI21D1BWP12T U1226 ( .A1(n1539), .A2(n1538), .B(n1537), .ZN(n333) );
  OAI21D0BWP12T U1227 ( .A1(n1539), .A2(n1538), .B(n1537), .ZN(n334) );
  TPND2D1BWP12T U1228 ( .A1(n1536), .A2(n1535), .ZN(n1537) );
  TPOAI21D1BWP12T U1229 ( .A1(n1380), .A2(n1378), .B(n1379), .ZN(n1382) );
  TPND2D2BWP12T U1230 ( .A1(n2021), .A2(n2020), .ZN(n2025) );
  AN2D4BWP12T U1231 ( .A1(n1426), .A2(n337), .Z(n354) );
  INVD1BWP12T U1232 ( .I(n2458), .ZN(n2460) );
  RCAOI22D2BWP12T U1233 ( .A1(n2110), .A2(n2296), .B1(n2295), .B2(n2109), .ZN(
        n2144) );
  XOR3D2BWP12T U1234 ( .A1(n2597), .A2(n2598), .A3(n2596), .Z(n2532) );
  TPOAI22D2BWP12T U1235 ( .A1(n1561), .A2(n2647), .B1(n1442), .B2(n1441), .ZN(
        n1553) );
  BUFFXD6BWP12T U1236 ( .I(n4764), .Z(n336) );
  XNR2XD2BWP12T U1237 ( .A1(b[22]), .A2(n2746), .ZN(n2070) );
  XNR2XD2BWP12T U1238 ( .A1(b[22]), .A2(n288), .ZN(n1906) );
  XNR2D2BWP12T U1239 ( .A1(b[22]), .A2(n4214), .ZN(n1551) );
  INVD1BWP12T U1240 ( .I(n3864), .ZN(n1496) );
  INVD1BWP12T U1241 ( .I(n4270), .ZN(n4274) );
  TPOAI21D1BWP12T U1242 ( .A1(n1023), .A2(n1686), .B(n1685), .ZN(n1690) );
  CKND2D2BWP12T U1243 ( .A1(n422), .A2(n446), .ZN(n424) );
  TPOAI21D1BWP12T U1244 ( .A1(n1338), .A2(n1337), .B(n1336), .ZN(n337) );
  OAI21D1BWP12T U1245 ( .A1(n1338), .A2(n1337), .B(n1336), .ZN(n1425) );
  XOR3XD4BWP12T U1246 ( .A1(n2408), .A2(n2407), .A3(n2406), .Z(n2489) );
  INVD2BWP12T U1247 ( .I(n1880), .ZN(n1859) );
  TPOAI21D2BWP12T U1248 ( .A1(n3669), .A2(n3671), .B(n3672), .ZN(n2512) );
  OAI22D4BWP12T U1249 ( .A1(n1925), .A2(n2667), .B1(n1924), .B2(n2669), .ZN(
        n2023) );
  XOR3D2BWP12T U1250 ( .A1(n2378), .A2(n2377), .A3(n2373), .Z(n338) );
  TPOAI22D2BWP12T U1251 ( .A1(n1546), .A2(n1894), .B1(n2236), .B2(n2643), .ZN(
        n2378) );
  CKND2D2BWP12T U1252 ( .A1(n736), .A2(n735), .ZN(n740) );
  RCAOI21D2BWP12T U1253 ( .A1(n767), .A2(n4110), .B(n766), .ZN(n3358) );
  TPOAI22D4BWP12T U1254 ( .A1(n2069), .A2(n2740), .B1(n1981), .B2(n2739), .ZN(
        n2084) );
  TPND2D2BWP12T U1255 ( .A1(n1493), .A2(n1492), .ZN(n3023) );
  INVD2BWP12T U1256 ( .I(n2107), .ZN(n2002) );
  TPOAI22D4BWP12T U1257 ( .A1(n1280), .A2(n2646), .B1(n1367), .B2(n4257), .ZN(
        n1310) );
  OAI22D4BWP12T U1258 ( .A1(n611), .A2(n2263), .B1(n2265), .B2(n643), .ZN(n658) );
  XNR2XD2BWP12T U1259 ( .A1(n4754), .A2(n2593), .ZN(n561) );
  XNR2XD2BWP12T U1260 ( .A1(n4754), .A2(n2701), .ZN(n1177) );
  XNR2XD2BWP12T U1261 ( .A1(n4754), .A2(n2688), .ZN(n2099) );
  XNR2XD2BWP12T U1262 ( .A1(n4754), .A2(n2666), .ZN(n2238) );
  XNR2XD4BWP12T U1263 ( .A1(n4754), .A2(n288), .ZN(n1108) );
  MUX2NXD16BWP12T U1264 ( .I0(n604), .I1(n603), .S(n1164), .ZN(n2680) );
  ND2XD16BWP12T U1265 ( .A1(n413), .A2(n412), .ZN(n1442) );
  OA22D1BWP12T U1266 ( .A1(n1547), .A2(n2319), .B1(n1464), .B2(n2702), .Z(n340) );
  ND2D3BWP12T U1267 ( .A1(n1447), .A2(n1446), .ZN(n1452) );
  TPND2D1BWP12T U1268 ( .A1(n328), .A2(n2046), .ZN(n2048) );
  XNR2XD4BWP12T U1269 ( .A1(n2072), .A2(n3040), .ZN(n1933) );
  DCCKND4BWP12T U1270 ( .I(b[8]), .ZN(n428) );
  INVD6BWP12T U1271 ( .I(n852), .ZN(n341) );
  TPOAI22D1BWP12T U1272 ( .A1(n2178), .A2(n306), .B1(n2177), .B2(n2624), .ZN(
        n2180) );
  IOA21D1BWP12T U1273 ( .A1(n1330), .A2(n1329), .B(n1394), .ZN(n1331) );
  RCAOI21D4BWP12T U1274 ( .A1(n711), .A2(n2667), .B(n710), .ZN(n1054) );
  INVD1BWP12T U1275 ( .I(n4676), .ZN(n342) );
  INVD1BWP12T U1276 ( .I(n2482), .ZN(n343) );
  TPND2D2BWP12T U1277 ( .A1(n1330), .A2(n1329), .ZN(n1395) );
  TPOAI22D1BWP12T U1278 ( .A1(n558), .A2(n2319), .B1(n531), .B2(n2702), .ZN(
        n564) );
  TPOAI22D1BWP12T U1279 ( .A1(n732), .A2(n2748), .B1(n2747), .B2(n1064), .ZN(
        n1043) );
  TPND2D2BWP12T U1280 ( .A1(n345), .A2(n344), .ZN(n346) );
  DCCKND4BWP12T U1281 ( .I(n1403), .ZN(n344) );
  TPND2D2BWP12T U1282 ( .A1(n1382), .A2(n1381), .ZN(n1402) );
  INVD4BWP12T U1283 ( .I(b[6]), .ZN(n852) );
  CKND2D2BWP12T U1284 ( .A1(n1279), .A2(n1278), .ZN(n3734) );
  BUFFD12BWP12T U1285 ( .I(b[16]), .Z(n4761) );
  TPOAI22D4BWP12T U1286 ( .A1(n1181), .A2(n296), .B1(n1093), .B2(n2263), .ZN(
        n1190) );
  TPOAI21D1BWP12T U1287 ( .A1(n2354), .A2(n2353), .B(n2246), .ZN(n2247) );
  XOR3D2BWP12T U1288 ( .A1(n2232), .A2(n2231), .A3(n2230), .Z(n2354) );
  INVD2BWP12T U1289 ( .I(n2355), .ZN(n2246) );
  TPOAI22D2BWP12T U1290 ( .A1(n482), .A2(n2747), .B1(n436), .B2(n2748), .ZN(
        n487) );
  TPOAI22D2BWP12T U1291 ( .A1(n1108), .A2(n1442), .B1(n1151), .B2(n2647), .ZN(
        n1172) );
  TPNR2D1BWP12T U1292 ( .A1(n1536), .A2(n1535), .ZN(n1539) );
  XNR2XD4BWP12T U1293 ( .A1(n2575), .A2(n5014), .ZN(n1518) );
  INVD1BWP12T U1294 ( .I(n2507), .ZN(n2474) );
  FA1D2BWP12T U1295 ( .A(n2327), .B(n2326), .CI(n2325), .CO(n2465), .S(n2409)
         );
  INR2D2BWP12T U1296 ( .A1(n2045), .B1(n328), .ZN(n2049) );
  INVD1BWP12T U1297 ( .I(n3249), .ZN(n3377) );
  BUFFXD4BWP12T U1298 ( .I(b[31]), .Z(n4751) );
  FA1D2BWP12T U1299 ( .A(n2718), .B(n2717), .CI(n2716), .CO(n2719), .S(n2758)
         );
  XNR2XD4BWP12T U1300 ( .A1(n2575), .A2(n2679), .ZN(n2267) );
  OR2D4BWP12T U1301 ( .A1(n652), .A2(n2647), .Z(n633) );
  XNR2XD4BWP12T U1302 ( .A1(n2094), .A2(n288), .ZN(n652) );
  XOR3XD4BWP12T U1303 ( .A1(n1271), .A2(n1274), .A3(n1270), .Z(n1149) );
  RCOAI21D2BWP12T U1304 ( .A1(n4284), .A2(n4260), .B(n3168), .ZN(result[17])
         );
  BUFFXD8BWP12T U1305 ( .I(b[12]), .Z(n2623) );
  IOA21D2BWP12T U1306 ( .A1(n2087), .A2(n2088), .B(n1958), .ZN(n2127) );
  IOA21D2BWP12T U1307 ( .A1(n1957), .A2(n1956), .B(n2086), .ZN(n1958) );
  XNR2XD2BWP12T U1308 ( .A1(n2555), .A2(n4699), .ZN(n1896) );
  BUFFD16BWP12T U1309 ( .I(b[0]), .Z(n4316) );
  CKND2D2BWP12T U1310 ( .A1(n2170), .A2(n2688), .ZN(n1092) );
  INVD2BWP12T U1311 ( .I(n682), .ZN(n683) );
  TPND2D2BWP12T U1312 ( .A1(n682), .A2(n684), .ZN(n627) );
  RCOAI21D2BWP12T U1313 ( .A1(n682), .A2(n684), .B(n685), .ZN(n628) );
  NR2D0BWP12T U1314 ( .A1(n3844), .A2(n4707), .ZN(n3510) );
  TPOAI21D2BWP12T U1315 ( .A1(n4200), .A2(n4707), .B(n3969), .ZN(n3758) );
  OR2D2BWP12T U1316 ( .A1(n1512), .A2(n4625), .Z(n1346) );
  INVD2BWP12T U1317 ( .I(n1512), .ZN(n1513) );
  XNR2D2BWP12T U1318 ( .A1(b[22]), .A2(n2742), .ZN(n2321) );
  TPNR2D2BWP12T U1319 ( .A1(n1073), .A2(n1072), .ZN(n1069) );
  INVD2BWP12T U1320 ( .I(n1050), .ZN(n717) );
  ND2XD8BWP12T U1321 ( .A1(n1307), .A2(n533), .ZN(n2263) );
  CKND0BWP12T U1322 ( .I(n1097), .ZN(n1068) );
  XNR2D2BWP12T U1323 ( .A1(n2619), .A2(n2688), .ZN(n2552) );
  XNR2XD2BWP12T U1324 ( .A1(n2619), .A2(n2679), .ZN(n2090) );
  XNR2XD8BWP12T U1325 ( .A1(n2619), .A2(n2746), .ZN(n1239) );
  XNR2XD4BWP12T U1326 ( .A1(n2096), .A2(n2679), .ZN(n654) );
  TPND2D2BWP12T U1327 ( .A1(n2085), .A2(n2084), .ZN(n1991) );
  INVD1BWP12T U1328 ( .I(n2085), .ZN(n1990) );
  XNR2D2BWP12T U1329 ( .A1(n2072), .A2(n4699), .ZN(n2097) );
  XNR2D2BWP12T U1330 ( .A1(n2072), .A2(n653), .ZN(n747) );
  XOR2XD2BWP12T U1331 ( .A1(n2072), .A2(n431), .Z(n484) );
  XOR3XD4BWP12T U1332 ( .A1(n2188), .A2(n2187), .A3(n2186), .Z(n2208) );
  TPOAI22D1BWP12T U1333 ( .A1(n1348), .A2(n2263), .B1(n1518), .B2(n2265), .ZN(
        n1460) );
  XNR2XD4BWP12T U1334 ( .A1(n4686), .A2(n866), .ZN(n568) );
  DCCKBD4BWP12T U1335 ( .I(n1932), .Z(n1709) );
  DCCKND4BWP12T U1336 ( .I(n1932), .ZN(n4686) );
  DCCKND4BWP12T U1337 ( .I(a[11]), .ZN(n866) );
  TPOAI22D1BWP12T U1338 ( .A1(n423), .A2(n2648), .B1(n430), .B2(n2647), .ZN(
        n445) );
  IOA21D1BWP12T U1339 ( .A1(n1876), .A2(n1875), .B(n1996), .ZN(n1878) );
  TPND2D2BWP12T U1340 ( .A1(n601), .A2(n600), .ZN(n1687) );
  OR2D4BWP12T U1341 ( .A1(n601), .A2(n600), .Z(n1688) );
  XNR2XD2BWP12T U1342 ( .A1(n4754), .A2(n2679), .ZN(n1557) );
  XOR3XD4BWP12T U1343 ( .A1(n2213), .A2(n2212), .A3(n2211), .Z(n2361) );
  RCOAI21D1BWP12T U1344 ( .A1(n2176), .A2(n2175), .B(n2174), .ZN(n2213) );
  TPOAI22D1BWP12T U1345 ( .A1(n1109), .A2(n4257), .B1(n1048), .B2(n2646), .ZN(
        n1084) );
  OAI21D1BWP12T U1346 ( .A1(n2150), .A2(n2151), .B(n2149), .ZN(n2101) );
  TPND2D2BWP12T U1347 ( .A1(n2151), .A2(n2150), .ZN(n2100) );
  BUFFD8BWP12T U1348 ( .I(b[15]), .Z(n2551) );
  XNR2D2BWP12T U1349 ( .A1(n2098), .A2(n2688), .ZN(n2168) );
  INVD2BWP12T U1350 ( .I(n2214), .ZN(n2176) );
  ND2D3BWP12T U1351 ( .A1(n3085), .A2(n4146), .ZN(n2437) );
  XNR2XD4BWP12T U1352 ( .A1(n4628), .A2(n288), .ZN(n554) );
  INVD12BWP12T U1353 ( .I(n853), .ZN(n4628) );
  BUFFXD16BWP12T U1354 ( .I(n1421), .Z(n2691) );
  INR2D2BWP12T U1355 ( .A1(n953), .B1(n5082), .ZN(n4561) );
  INVD8BWP12T U1356 ( .I(n4738), .ZN(n992) );
  TPAOI31D1BWP12T U1357 ( .A1(n1720), .A2(n4573), .A3(n1719), .B(n5100), .ZN(
        n4878) );
  ND2XD4BWP12T U1358 ( .A1(n4283), .A2(n5085), .ZN(n1855) );
  XNR2XD2BWP12T U1359 ( .A1(b[10]), .A2(n4924), .ZN(n1934) );
  DCCKND4BWP12T U1360 ( .I(b[10]), .ZN(n506) );
  TPND2D2BWP12T U1361 ( .A1(n4009), .A2(n4005), .ZN(n1024) );
  CKND0BWP12T U1362 ( .I(n3097), .ZN(n2916) );
  AOI22D1BWP12T U1363 ( .A1(n3107), .A2(n3098), .B1(n3097), .B2(n3096), .ZN(
        n3102) );
  TPNR2D2BWP12T U1364 ( .A1(n1491), .A2(n1490), .ZN(n3020) );
  BUFFXD12BWP12T U1365 ( .I(n3107), .Z(n3941) );
  NR2D4BWP12T U1366 ( .A1(n3436), .A2(n3005), .ZN(n3107) );
  CKND2D2BWP12T U1367 ( .A1(n618), .A2(n349), .ZN(n621) );
  TPND2D3BWP12T U1368 ( .A1(n4083), .A2(n4082), .ZN(result[14]) );
  XOR2XD2BWP12T U1369 ( .A1(n3171), .A2(n3170), .Z(n4278) );
  ND2D4BWP12T U1370 ( .A1(n1855), .A2(n1854), .ZN(result[18]) );
  TPOAI21D1BWP12T U1371 ( .A1(n975), .A2(n4227), .B(n4108), .ZN(n1786) );
  TPOAI22D4BWP12T U1372 ( .A1(n1109), .A2(n2646), .B1(n1187), .B2(n4257), .ZN(
        n1170) );
  TPAOI21D1BWP12T U1373 ( .A1(n3866), .A2(n318), .B(n3864), .ZN(n3871) );
  BUFFXD0BWP12T U1374 ( .I(n4924), .Z(n3771) );
  BUFFD8BWP12T U1375 ( .I(a[11]), .Z(n5014) );
  INVD3BWP12T U1376 ( .I(n4699), .ZN(n2169) );
  BUFFXD0BWP12T U1377 ( .I(n4699), .Z(n2792) );
  BUFFXD0BWP12T U1378 ( .I(n4699), .Z(n2818) );
  BUFFD6BWP12T U1379 ( .I(a[2]), .Z(n4912) );
  INVD2BWP12T U1380 ( .I(n4912), .ZN(n373) );
  INVD6BWP12T U1381 ( .I(n4627), .ZN(n2746) );
  INVD1BWP12T U1382 ( .I(n848), .ZN(n3455) );
  INVD4BWP12T U1383 ( .I(a[15]), .ZN(n1058) );
  BUFFXD0BWP12T U1384 ( .I(n5014), .Z(n4449) );
  BUFFXD0BWP12T U1385 ( .I(n4699), .Z(n3847) );
  OA21D2BWP12T U1386 ( .A1(n2743), .A2(n570), .B(n538), .Z(n349) );
  INVD6BWP12T U1387 ( .I(n1058), .ZN(n2666) );
  INVD3BWP12T U1388 ( .I(n3523), .ZN(n4906) );
  BUFFD2BWP12T U1389 ( .I(n480), .Z(n3523) );
  INVD1BWP12T U1390 ( .I(n5063), .ZN(n5099) );
  INVD1BWP12T U1391 ( .I(n4103), .ZN(n4489) );
  NR2D1BWP12T U1392 ( .A1(n833), .A2(n911), .ZN(n4103) );
  OA211D1BWP12T U1393 ( .A1(n4954), .A2(n942), .B(n941), .C(n940), .Z(n350) );
  INVD1BWP12T U1394 ( .I(n4954), .ZN(n5093) );
  ND2D1BWP12T U1395 ( .A1(n909), .A2(n933), .ZN(n4954) );
  AN2D1BWP12T U1396 ( .A1(n4743), .A2(n1785), .Z(n1770) );
  ND2D1BWP12T U1397 ( .A1(n904), .A2(n765), .ZN(n4260) );
  INVD1BWP12T U1398 ( .I(n5094), .ZN(n5040) );
  INR2D1BWP12T U1399 ( .A1(n933), .B1(n860), .ZN(n5094) );
  ND2D1BWP12T U1400 ( .A1(n4765), .A2(n3523), .ZN(n351) );
  AN2D1BWP12T U1401 ( .A1(n2495), .A2(n2494), .Z(n352) );
  INVD2BWP12T U1402 ( .I(n4260), .ZN(n5085) );
  INVD1BWP12T U1403 ( .I(n2792), .ZN(n4649) );
  INVD1BWP12T U1404 ( .I(n848), .ZN(n4624) );
  AN2D1BWP12T U1405 ( .A1(n3926), .A2(n3925), .Z(n353) );
  OR2D2BWP12T U1406 ( .A1(n2263), .A2(n866), .Z(n355) );
  AN2D1BWP12T U1407 ( .A1(n2170), .A2(n5014), .Z(n356) );
  CKBD1BWP12T U1408 ( .I(n4914), .Z(n3053) );
  INVD1BWP12T U1409 ( .I(n4914), .ZN(n4625) );
  INVD1BWP12T U1410 ( .I(n4910), .ZN(n5079) );
  INVD1BWP12T U1411 ( .I(n2666), .ZN(n710) );
  CKBD1BWP12T U1412 ( .I(n861), .Z(n4653) );
  OR2XD1BWP12T U1413 ( .A1(n3604), .A2(n3292), .Z(n357) );
  CKBD1BWP12T U1414 ( .I(n289), .Z(n4125) );
  INVD1BWP12T U1415 ( .I(n2450), .ZN(n2429) );
  ND2D1BWP12T U1416 ( .A1(n300), .A2(n3548), .ZN(n358) );
  ND2D1BWP12T U1417 ( .A1(n616), .A2(n615), .ZN(n359) );
  TPOAI22D1BWP12T U1418 ( .A1(n1443), .A2(n2747), .B1(n1349), .B2(n2748), .ZN(
        n1458) );
  TPOAI22D2BWP12T U1419 ( .A1(n569), .A2(n2747), .B1(n535), .B2(n2748), .ZN(
        n541) );
  INVD6BWP12T U1420 ( .I(a[5]), .ZN(n4627) );
  XNR2D1BWP12T U1421 ( .A1(n4316), .A2(n2746), .ZN(n362) );
  BUFFD6BWP12T U1422 ( .I(a[4]), .Z(n4921) );
  AN2XD2BWP12T U1423 ( .A1(n4627), .A2(n4921), .Z(n361) );
  INVD3BWP12T U1424 ( .I(a[3]), .ZN(n871) );
  INVD8BWP12T U1425 ( .I(n871), .ZN(n4913) );
  INVD12BWP12T U1426 ( .I(n4913), .ZN(n374) );
  TPOAI21D8BWP12T U1427 ( .A1(n361), .A2(n374), .B(n360), .ZN(n2748) );
  INVD6BWP12T U1428 ( .I(n605), .ZN(n4738) );
  XNR2D1BWP12T U1429 ( .A1(n4738), .A2(n2746), .ZN(n395) );
  INVD18BWP12T U1430 ( .I(n374), .ZN(n2742) );
  XNR2XD8BWP12T U1431 ( .A1(n2742), .A2(n4921), .ZN(n2747) );
  OAI22D1BWP12T U1432 ( .A1(n362), .A2(n2748), .B1(n395), .B2(n2747), .ZN(n402) );
  BUFFXD4BWP12T U1433 ( .I(b[0]), .Z(n1512) );
  IND2D1BWP12T U1434 ( .A1(n1512), .B1(n2746), .ZN(n363) );
  OAI22D1BWP12T U1435 ( .A1(n363), .A2(n2747), .B1(n2748), .B2(n4627), .ZN(
        n401) );
  BUFFXD12BWP12T U1436 ( .I(b[2]), .Z(n2072) );
  XNR2D1BWP12T U1437 ( .A1(n2742), .A2(n2072), .ZN(n367) );
  INVD3BWP12T U1438 ( .I(n4913), .ZN(n4626) );
  TPND2D1BWP12T U1439 ( .A1(a[1]), .A2(n4626), .ZN(n372) );
  INVD1P75BWP12T U1440 ( .I(n4626), .ZN(n365) );
  TPNR2D3BWP12T U1441 ( .A1(a[1]), .A2(n4912), .ZN(n364) );
  TPND2D2BWP12T U1442 ( .A1(n365), .A2(n364), .ZN(n371) );
  OA21D2BWP12T U1443 ( .A1(n373), .A2(n372), .B(n371), .Z(n536) );
  XNR2D1BWP12T U1444 ( .A1(n2742), .A2(b[3]), .ZN(n398) );
  XNR2D2BWP12T U1445 ( .A1(n4912), .A2(a[1]), .ZN(n471) );
  OAI22D1BWP12T U1446 ( .A1(n367), .A2(n536), .B1(n398), .B2(n2743), .ZN(n397)
         );
  INVD4BWP12T U1447 ( .I(a[1]), .ZN(n4644) );
  INVD9BWP12T U1448 ( .I(n4644), .ZN(n2593) );
  XNR2XD0BWP12T U1449 ( .A1(n2071), .A2(n2593), .ZN(n369) );
  INVD1P75BWP12T U1450 ( .I(a[0]), .ZN(n366) );
  ND2D3BWP12T U1451 ( .A1(a[1]), .A2(n366), .ZN(n607) );
  BUFFXD8BWP12T U1452 ( .I(n607), .Z(n2646) );
  BUFFXD3BWP12T U1453 ( .I(a[1]), .Z(n4214) );
  XNR2D1BWP12T U1454 ( .A1(n4214), .A2(n4628), .ZN(n399) );
  INVD12BWP12T U1455 ( .I(n4910), .ZN(n4257) );
  TPOAI22D1BWP12T U1456 ( .A1(n369), .A2(n2646), .B1(n399), .B2(n4257), .ZN(
        n396) );
  INVD12BWP12T U1457 ( .I(n605), .ZN(n1932) );
  XNR2D1BWP12T U1458 ( .A1(n1932), .A2(n2742), .ZN(n377) );
  OAI22D1BWP12T U1459 ( .A1(n367), .A2(n2743), .B1(n377), .B2(n536), .ZN(n387)
         );
  INR2D1BWP12T U1460 ( .A1(n4316), .B1(n2747), .ZN(n386) );
  BUFFXD12BWP12T U1461 ( .I(b[3]), .Z(n2555) );
  CKND1BWP12T U1462 ( .I(n4644), .ZN(n368) );
  XNR2D1BWP12T U1463 ( .A1(n2555), .A2(n368), .ZN(n376) );
  OAI22D1BWP12T U1464 ( .A1(n376), .A2(n2646), .B1(n369), .B2(n4257), .ZN(n385) );
  IND2XD2BWP12T U1465 ( .A1(n393), .B1(n370), .ZN(n3341) );
  IND2D1BWP12T U1466 ( .A1(n1512), .B1(n2742), .ZN(n375) );
  OA21XD4BWP12T U1467 ( .A1(n373), .A2(n372), .B(n371), .Z(n2744) );
  OAI22D1BWP12T U1468 ( .A1(n375), .A2(n2743), .B1(n2744), .B2(n374), .ZN(n389) );
  BUFFXD8BWP12T U1469 ( .I(n2072), .Z(n3748) );
  XNR2D1BWP12T U1470 ( .A1(n3748), .A2(n2593), .ZN(n378) );
  TPOAI22D1BWP12T U1471 ( .A1(n376), .A2(n4257), .B1(n378), .B2(n2646), .ZN(
        n388) );
  TPNR2D2BWP12T U1472 ( .A1(n383), .A2(n382), .ZN(n4095) );
  XNR2D1BWP12T U1473 ( .A1(n2593), .A2(n4738), .ZN(n379) );
  OAI22D1BWP12T U1474 ( .A1(n378), .A2(n4257), .B1(n379), .B2(n2646), .ZN(n381) );
  INVD1BWP12T U1475 ( .I(n4316), .ZN(n4225) );
  NR2D1BWP12T U1476 ( .A1(n4225), .A2(n2743), .ZN(n380) );
  TPOAI22D1BWP12T U1477 ( .A1(n2646), .A2(n1512), .B1(n379), .B2(n4257), .ZN(
        n4238) );
  ND2D1BWP12T U1478 ( .A1(n4238), .A2(n4237), .ZN(n4239) );
  ND2D1BWP12T U1479 ( .A1(n381), .A2(n380), .ZN(n997) );
  TPOAI21D1BWP12T U1480 ( .A1(n996), .A2(n4239), .B(n997), .ZN(n4098) );
  CKND2D2BWP12T U1481 ( .A1(n383), .A2(n382), .ZN(n4096) );
  FA1D2BWP12T U1482 ( .A(n387), .B(n386), .CI(n385), .CO(n392), .S(n391) );
  HA1D2BWP12T U1483 ( .A(n389), .B(n388), .CO(n390), .S(n383) );
  NR2XD2BWP12T U1484 ( .A1(n391), .A2(n390), .ZN(n1753) );
  CKND2D2BWP12T U1485 ( .A1(n391), .A2(n390), .ZN(n1754) );
  TPOAI21D2BWP12T U1486 ( .A1(n1755), .A2(n1753), .B(n1754), .ZN(n3342) );
  INVD1P75BWP12T U1487 ( .I(n3340), .ZN(n394) );
  TPAOI21D2BWP12T U1488 ( .A1(n3341), .A2(n3342), .B(n394), .ZN(n3663) );
  XNR2D1BWP12T U1489 ( .A1(n3748), .A2(n2746), .ZN(n437) );
  OAI22D1BWP12T U1490 ( .A1(n437), .A2(n2747), .B1(n395), .B2(n2748), .ZN(n457) );
  HA1D2BWP12T U1491 ( .A(n397), .B(n396), .CO(n458), .S(n400) );
  BUFFD6BWP12T U1492 ( .I(a[6]), .Z(n4931) );
  XNR2XD8BWP12T U1493 ( .A1(n4627), .A2(n4931), .ZN(n411) );
  TPOAI22D2BWP12T U1494 ( .A1(n435), .A2(n2743), .B1(n2744), .B2(n398), .ZN(
        n438) );
  OAI22D1BWP12T U1495 ( .A1(n399), .A2(n607), .B1(n417), .B2(n4257), .ZN(n439)
         );
  XOR3D2BWP12T U1496 ( .A1(n440), .A2(n438), .A3(n439), .Z(n456) );
  CKND3BWP12T U1497 ( .I(n406), .ZN(n404) );
  FA1D2BWP12T U1498 ( .A(n402), .B(n401), .CI(n400), .CO(n405), .S(n393) );
  INVD1BWP12T U1499 ( .I(n405), .ZN(n403) );
  TPND2D2BWP12T U1500 ( .A1(n404), .A2(n403), .ZN(n3662) );
  CKND2BWP12T U1501 ( .I(n3662), .ZN(n407) );
  ND2D1BWP12T U1502 ( .A1(n406), .A2(n405), .ZN(n3661) );
  TPOAI21D2BWP12T U1503 ( .A1(n3663), .A2(n407), .B(n3661), .ZN(n3249) );
  XNR2XD4BWP12T U1504 ( .A1(a[7]), .A2(a[8]), .ZN(n467) );
  BUFFXD6BWP12T U1505 ( .I(n467), .Z(n2704) );
  INR2D2BWP12T U1506 ( .A1(n4316), .B1(n2704), .ZN(n491) );
  INVD1BWP12T U1507 ( .I(n471), .ZN(n1114) );
  INR2D2BWP12T U1508 ( .A1(n1114), .B1(n470), .ZN(n409) );
  XNR2D1BWP12T U1509 ( .A1(n4628), .A2(n2742), .ZN(n434) );
  TPNR2D2BWP12T U1510 ( .A1(n434), .A2(n536), .ZN(n408) );
  TPNR2D2BWP12T U1511 ( .A1(n409), .A2(n408), .ZN(n486) );
  XNR2D1BWP12T U1512 ( .A1(n2746), .A2(n2071), .ZN(n482) );
  XNR2XD4BWP12T U1513 ( .A1(n2746), .A2(n2555), .ZN(n436) );
  XNR3XD4BWP12T U1514 ( .A1(n485), .A2(n486), .A3(n487), .ZN(n495) );
  IND2D1BWP12T U1515 ( .A1(n1512), .B1(n288), .ZN(n415) );
  INVD3BWP12T U1516 ( .I(n4931), .ZN(n410) );
  XOR2XD4BWP12T U1517 ( .A1(n410), .A2(n414), .Z(n413) );
  BUFFXD1BWP12T U1518 ( .I(n414), .Z(n431) );
  INVD1P25BWP12T U1519 ( .I(n447), .ZN(n422) );
  DCCKND4BWP12T U1520 ( .I(b[7]), .ZN(n416) );
  XNR2D2BWP12T U1521 ( .A1(n2593), .A2(n2094), .ZN(n429) );
  CKND3BWP12T U1522 ( .I(n429), .ZN(n421) );
  CKND2BWP12T U1523 ( .I(n417), .ZN(n419) );
  CKND1BWP12T U1524 ( .I(n607), .ZN(n418) );
  RCAOI22D2BWP12T U1525 ( .A1(n421), .A2(n420), .B1(n419), .B2(n418), .ZN(n446) );
  XNR2D1BWP12T U1526 ( .A1(n4316), .A2(n288), .ZN(n423) );
  BUFFXD16BWP12T U1527 ( .I(n1442), .Z(n2648) );
  XNR2D1BWP12T U1528 ( .A1(n1709), .A2(n288), .ZN(n430) );
  CKND2D2BWP12T U1529 ( .A1(n425), .A2(n447), .ZN(n426) );
  CKND2D2BWP12T U1530 ( .A1(n427), .A2(n426), .ZN(n497) );
  INVD9BWP12T U1531 ( .I(n428), .ZN(n2167) );
  NR2D2BWP12T U1532 ( .A1(n2648), .A2(n430), .ZN(n433) );
  NR2D1BWP12T U1533 ( .A1(n2647), .A2(n484), .ZN(n432) );
  TPNR2D2BWP12T U1534 ( .A1(n433), .A2(n432), .ZN(n475) );
  OAI22D1BWP12T U1535 ( .A1(n435), .A2(n2744), .B1(n434), .B2(n2743), .ZN(n444) );
  AN2XD2BWP12T U1536 ( .A1(n444), .A2(n443), .Z(n473) );
  XNR3XD4BWP12T U1537 ( .A1(n476), .A2(n475), .A3(n473), .ZN(n493) );
  XNR3XD4BWP12T U1538 ( .A1(n495), .A2(n497), .A3(n493), .ZN(n464) );
  OAI21D1BWP12T U1539 ( .A1(n440), .A2(n439), .B(n438), .ZN(n442) );
  CKND2D1BWP12T U1540 ( .A1(n440), .A2(n439), .ZN(n441) );
  XNR2D2BWP12T U1541 ( .A1(n444), .A2(n443), .ZN(n452) );
  INVD1BWP12T U1542 ( .I(n452), .ZN(n450) );
  INVD1BWP12T U1543 ( .I(n453), .ZN(n448) );
  XNR3XD4BWP12T U1544 ( .A1(n447), .A2(n446), .A3(n445), .ZN(n451) );
  IOA21D2BWP12T U1545 ( .A1(n448), .A2(n452), .B(n451), .ZN(n449) );
  IOA21D2BWP12T U1546 ( .A1(n453), .A2(n450), .B(n449), .ZN(n463) );
  TPNR2D3BWP12T U1547 ( .A1(n464), .A2(n463), .ZN(n3378) );
  XNR3XD4BWP12T U1548 ( .A1(n453), .A2(n452), .A3(n451), .ZN(n462) );
  CKND1BWP12T U1549 ( .I(n457), .ZN(n454) );
  ND2D1BWP12T U1550 ( .A1(n458), .A2(n457), .ZN(n459) );
  NR2D2BWP12T U1551 ( .A1(n462), .A2(n461), .ZN(n3376) );
  TPNR2D1BWP12T U1552 ( .A1(n3378), .A2(n3376), .ZN(n466) );
  TPND2D2BWP12T U1553 ( .A1(n462), .A2(n461), .ZN(n3375) );
  TPOAI21D1BWP12T U1554 ( .A1(n3378), .A2(n3375), .B(n3379), .ZN(n465) );
  TPAOI21D2BWP12T U1555 ( .A1(n3249), .A2(n466), .B(n465), .ZN(n3496) );
  INVD4BWP12T U1556 ( .I(a[9]), .ZN(n480) );
  IND2D1BWP12T U1557 ( .A1(n1512), .B1(n4906), .ZN(n469) );
  BUFFD6BWP12T U1558 ( .I(n467), .Z(n2319) );
  XNR2XD2BWP12T U1559 ( .A1(n480), .A2(a[8]), .ZN(n468) );
  ND2XD8BWP12T U1560 ( .A1(n468), .A2(n467), .ZN(n2702) );
  TPOAI22D2BWP12T U1561 ( .A1(n469), .A2(n2319), .B1(n3523), .B2(n2702), .ZN(
        n520) );
  XNR2XD2BWP12T U1562 ( .A1(n2094), .A2(n2742), .ZN(n505) );
  OAI22D2BWP12T U1563 ( .A1(n505), .A2(n471), .B1(n536), .B2(n470), .ZN(n519)
         );
  XNR2D1BWP12T U1564 ( .A1(n2098), .A2(n2593), .ZN(n507) );
  OAI22D1BWP12T U1565 ( .A1(n472), .A2(n2646), .B1(n507), .B2(n4257), .ZN(n518) );
  INVD1BWP12T U1566 ( .I(n476), .ZN(n474) );
  IOA21D1BWP12T U1567 ( .A1(n475), .A2(n474), .B(n473), .ZN(n479) );
  INVD1BWP12T U1568 ( .I(n475), .ZN(n477) );
  ND2D1BWP12T U1569 ( .A1(n477), .A2(n476), .ZN(n478) );
  CKAN2D2BWP12T U1570 ( .A1(n479), .A2(n478), .Z(n524) );
  INVD12BWP12T U1571 ( .I(n480), .ZN(n2701) );
  OAI22D1BWP12T U1572 ( .A1(n481), .A2(n2702), .B1(n504), .B2(n2319), .ZN(n509) );
  INVD1BWP12T U1573 ( .I(n509), .ZN(n492) );
  XNR2D1BWP12T U1574 ( .A1(n4628), .A2(n2746), .ZN(n516) );
  TPOAI22D1BWP12T U1575 ( .A1(n482), .A2(n2748), .B1(n516), .B2(n2747), .ZN(
        n515) );
  XNR2XD1BWP12T U1576 ( .A1(n2555), .A2(n288), .ZN(n517) );
  TPOAI22D2BWP12T U1577 ( .A1(n517), .A2(n2647), .B1(n484), .B2(n483), .ZN(
        n514) );
  ND2D1BWP12T U1578 ( .A1(n486), .A2(n485), .ZN(n488) );
  ND2D1BWP12T U1579 ( .A1(n487), .A2(n488), .ZN(n489) );
  IOA21D2BWP12T U1580 ( .A1(n491), .A2(n490), .B(n489), .ZN(n508) );
  XOR3XD4BWP12T U1581 ( .A1(n492), .A2(n508), .A3(n510), .Z(n526) );
  XNR3XD4BWP12T U1582 ( .A1(n522), .A2(n524), .A3(n526), .ZN(n502) );
  INVD1BWP12T U1583 ( .I(n497), .ZN(n494) );
  IOA21D1BWP12T U1584 ( .A1(n495), .A2(n494), .B(n493), .ZN(n499) );
  INVD1BWP12T U1585 ( .I(n495), .ZN(n496) );
  ND2D1BWP12T U1586 ( .A1(n497), .A2(n496), .ZN(n498) );
  TPND2D2BWP12T U1587 ( .A1(n502), .A2(n501), .ZN(n500) );
  INVD3BWP12T U1588 ( .I(n500), .ZN(n3493) );
  TPNR2D2BWP12T U1589 ( .A1(n502), .A2(n501), .ZN(n3495) );
  INVD1P75BWP12T U1590 ( .I(n3495), .ZN(n503) );
  TPOAI21D2BWP12T U1591 ( .A1(n3496), .A2(n3493), .B(n503), .ZN(n3267) );
  OAI22D1BWP12T U1592 ( .A1(n537), .A2(n2743), .B1(n2744), .B2(n505), .ZN(n549) );
  INVD8BWP12T U1593 ( .I(n506), .ZN(n4754) );
  OAI22D1BWP12T U1594 ( .A1(n561), .A2(n4257), .B1(n507), .B2(n2646), .ZN(n547) );
  XOR3XD4BWP12T U1595 ( .A1(n548), .A2(n549), .A3(n547), .Z(n592) );
  INVD1P75BWP12T U1596 ( .I(n508), .ZN(n513) );
  NR2D2BWP12T U1597 ( .A1(n510), .A2(n509), .ZN(n512) );
  ND2D1BWP12T U1598 ( .A1(n510), .A2(n509), .ZN(n511) );
  OAI21D2BWP12T U1599 ( .A1(n513), .A2(n512), .B(n511), .ZN(n593) );
  HA1D2BWP12T U1600 ( .A(n515), .B(n514), .CO(n577), .S(n510) );
  BUFFD6BWP12T U1601 ( .I(a[10]), .Z(n4904) );
  XNR2XD8BWP12T U1602 ( .A1(n2701), .A2(n4904), .ZN(n1307) );
  INVD6BWP12T U1603 ( .I(n610), .ZN(n2739) );
  NR2XD2BWP12T U1604 ( .A1(n2739), .A2(n4225), .ZN(n543) );
  XNR2XD2BWP12T U1605 ( .A1(n2172), .A2(n2746), .ZN(n535) );
  TPOAI22D2BWP12T U1606 ( .A1(n516), .A2(n2748), .B1(n535), .B2(n2747), .ZN(
        n544) );
  XNR2XD2BWP12T U1607 ( .A1(n2071), .A2(n288), .ZN(n532) );
  TPOAI22D2BWP12T U1608 ( .A1(n517), .A2(n2648), .B1(n532), .B2(n2647), .ZN(
        n542) );
  XOR3XD4BWP12T U1609 ( .A1(n543), .A2(n544), .A3(n542), .Z(n576) );
  XOR3D2BWP12T U1610 ( .A1(n577), .A2(n576), .A3(n578), .Z(n589) );
  XOR3D2BWP12T U1611 ( .A1(n592), .A2(n593), .A3(n589), .Z(n530) );
  INVD2BWP12T U1612 ( .I(n530), .ZN(n528) );
  INVD1BWP12T U1613 ( .I(n524), .ZN(n521) );
  NR2D1BWP12T U1614 ( .A1(n522), .A2(n521), .ZN(n525) );
  INVD1BWP12T U1615 ( .I(n522), .ZN(n523) );
  OAI22D1BWP12T U1616 ( .A1(n526), .A2(n525), .B1(n524), .B2(n523), .ZN(n529)
         );
  INVD1BWP12T U1617 ( .I(n529), .ZN(n527) );
  TPND2D2BWP12T U1618 ( .A1(n528), .A2(n527), .ZN(n3266) );
  TPND2D3BWP12T U1619 ( .A1(n530), .A2(n529), .ZN(n3265) );
  INVD2P3BWP12T U1620 ( .I(n3265), .ZN(n1684) );
  TPAOI21D1BWP12T U1621 ( .A1(n3267), .A2(n3266), .B(n1684), .ZN(n1023) );
  BUFFD8BWP12T U1622 ( .I(b[11]), .Z(n2575) );
  XNR2XD4BWP12T U1623 ( .A1(n2575), .A2(n2593), .ZN(n560) );
  OAI22D2BWP12T U1624 ( .A1(n560), .A2(n607), .B1(n608), .B2(n4257), .ZN(n622)
         );
  XNR2XD0BWP12T U1625 ( .A1(b[3]), .A2(n2701), .ZN(n558) );
  TPOAI22D1BWP12T U1626 ( .A1(n532), .A2(n1442), .B1(n554), .B2(n2647), .ZN(
        n563) );
  DCCKND4BWP12T U1627 ( .I(n1512), .ZN(n2170) );
  XNR2XD4BWP12T U1628 ( .A1(n866), .A2(n4904), .ZN(n533) );
  XNR2XD2BWP12T U1629 ( .A1(n2094), .A2(n2746), .ZN(n569) );
  TPNR2D1BWP12T U1630 ( .A1(n540), .A2(n541), .ZN(n619) );
  OR2D4BWP12T U1631 ( .A1(n537), .A2(n536), .Z(n538) );
  OAI21D1BWP12T U1632 ( .A1(n619), .A2(n349), .B(n618), .ZN(n539) );
  XNR3XD4BWP12T U1633 ( .A1(n541), .A2(n540), .A3(n349), .ZN(n573) );
  OAI21D1BWP12T U1634 ( .A1(n543), .A2(n544), .B(n542), .ZN(n546) );
  ND2D1BWP12T U1635 ( .A1(n544), .A2(n543), .ZN(n545) );
  CKND2D2BWP12T U1636 ( .A1(n546), .A2(n545), .ZN(n575) );
  OAI21D1BWP12T U1637 ( .A1(n549), .A2(n548), .B(n547), .ZN(n551) );
  TPOAI21D1BWP12T U1638 ( .A1(n573), .A2(n575), .B(n574), .ZN(n553) );
  TPND2D1BWP12T U1639 ( .A1(n573), .A2(n575), .ZN(n552) );
  INR2D4BWP12T U1640 ( .A1(a[12]), .B1(n866), .ZN(n603) );
  TPNR2D3BWP12T U1641 ( .A1(a[12]), .A2(a[11]), .ZN(n604) );
  OR2D8BWP12T U1642 ( .A1(n603), .A2(n604), .Z(n2682) );
  INR2D1BWP12T U1643 ( .A1(n4316), .B1(n2682), .ZN(n665) );
  OR2D2BWP12T U1644 ( .A1(n629), .A2(n2647), .Z(n557) );
  ND2D2BWP12T U1645 ( .A1(n631), .A2(n555), .ZN(n556) );
  TPND2D2BWP12T U1646 ( .A1(n557), .A2(n556), .ZN(n666) );
  XNR2XD4BWP12T U1647 ( .A1(n2071), .A2(n2701), .ZN(n609) );
  XNR3XD4BWP12T U1648 ( .A1(n665), .A2(n666), .A3(n559), .ZN(n677) );
  XNR2D1BWP12T U1649 ( .A1(n4316), .A2(n5014), .ZN(n562) );
  TPOAI22D2BWP12T U1650 ( .A1(n562), .A2(n2263), .B1(n568), .B2(n296), .ZN(
        n582) );
  HA1D2BWP12T U1651 ( .A(n563), .B(n564), .CO(n623), .S(n581) );
  NR2XD2BWP12T U1652 ( .A1(n582), .A2(n583), .ZN(n565) );
  INVD1P75BWP12T U1653 ( .I(n565), .ZN(n566) );
  ND2D2BWP12T U1654 ( .A1(n581), .A2(n566), .ZN(n567) );
  IOA21D2BWP12T U1655 ( .A1(n583), .A2(n582), .B(n567), .ZN(n678) );
  XNR2D2BWP12T U1656 ( .A1(n2072), .A2(n5014), .ZN(n611) );
  OA22D4BWP12T U1657 ( .A1(n569), .A2(n2748), .B1(n637), .B2(n2747), .Z(n614)
         );
  XNR2D1BWP12T U1658 ( .A1(n4754), .A2(n2742), .ZN(n669) );
  OAI22D1BWP12T U1659 ( .A1(n570), .A2(n2744), .B1(n669), .B2(n2743), .ZN(n612) );
  INVD1BWP12T U1660 ( .I(n612), .ZN(n571) );
  XNR3XD4BWP12T U1661 ( .A1(n616), .A2(n614), .A3(n571), .ZN(n680) );
  INVD3BWP12T U1662 ( .I(n680), .ZN(n572) );
  XOR3XD4BWP12T U1663 ( .A1(n677), .A2(n678), .A3(n572), .Z(n689) );
  XOR3XD4BWP12T U1664 ( .A1(n690), .A2(n691), .A3(n689), .Z(n601) );
  XNR3XD4BWP12T U1665 ( .A1(n575), .A2(n574), .A3(n573), .ZN(n586) );
  RCOAI21D2BWP12T U1666 ( .A1(n578), .A2(n577), .B(n576), .ZN(n580) );
  ND2D3BWP12T U1667 ( .A1(n578), .A2(n577), .ZN(n579) );
  TPND2D2BWP12T U1668 ( .A1(n580), .A2(n579), .ZN(n587) );
  XOR3D2BWP12T U1669 ( .A1(n583), .A2(n582), .A3(n581), .Z(n588) );
  XNR3XD4BWP12T U1670 ( .A1(n588), .A2(n587), .A3(n586), .ZN(n599) );
  INVD2BWP12T U1671 ( .I(n599), .ZN(n597) );
  INVD1BWP12T U1672 ( .I(n592), .ZN(n591) );
  INVD1BWP12T U1673 ( .I(n593), .ZN(n590) );
  ND2D1BWP12T U1674 ( .A1(n593), .A2(n592), .ZN(n594) );
  INVD1BWP12T U1675 ( .I(n598), .ZN(n596) );
  TPND2D2BWP12T U1676 ( .A1(n597), .A2(n596), .ZN(n4271) );
  TPND2D2BWP12T U1677 ( .A1(n1688), .A2(n4271), .ZN(n1022) );
  INVD1P75BWP12T U1678 ( .I(n1687), .ZN(n602) );
  TPAOI21D2BWP12T U1679 ( .A1(n1688), .A2(n4272), .B(n602), .ZN(n1021) );
  TPOAI21D1BWP12T U1680 ( .A1(n4270), .A2(n1022), .B(n1021), .ZN(n3171) );
  INVD6BWP12T U1681 ( .I(a[13]), .ZN(n861) );
  INVD15BWP12T U1682 ( .I(n4926), .ZN(n1164) );
  INVD9BWP12T U1683 ( .I(n1164), .ZN(n2679) );
  XNR2D1BWP12T U1684 ( .A1(n4316), .A2(n2679), .ZN(n606) );
  INVD2BWP12T U1685 ( .I(n605), .ZN(n2096) );
  BUFFXD8BWP12T U1686 ( .I(b[13]), .Z(n4753) );
  XNR2XD4BWP12T U1687 ( .A1(n4753), .A2(n2593), .ZN(n657) );
  XNR2XD4BWP12T U1688 ( .A1(n4628), .A2(n2701), .ZN(n642) );
  INVD2BWP12T U1689 ( .I(n610), .ZN(n2265) );
  XOR3XD4BWP12T U1690 ( .A1(n648), .A2(n649), .A3(n646), .Z(n682) );
  IND2XD1BWP12T U1691 ( .A1(n616), .B1(n614), .ZN(n613) );
  TPND2D2BWP12T U1692 ( .A1(n613), .A2(n612), .ZN(n617) );
  ND2D4BWP12T U1693 ( .A1(n617), .A2(n359), .ZN(n684) );
  INVD1P75BWP12T U1694 ( .I(n619), .ZN(n620) );
  ND2D2BWP12T U1695 ( .A1(n621), .A2(n620), .ZN(n626) );
  TPNR2D2BWP12T U1696 ( .A1(n623), .A2(n622), .ZN(n625) );
  TPND2D1BWP12T U1697 ( .A1(n623), .A2(n622), .ZN(n624) );
  RCOAI21D2BWP12T U1698 ( .A1(n626), .A2(n625), .B(n624), .ZN(n685) );
  TPND2D2BWP12T U1699 ( .A1(n628), .A2(n627), .ZN(n756) );
  INVD1BWP12T U1700 ( .I(n629), .ZN(n630) );
  CKND2D2BWP12T U1701 ( .A1(n631), .A2(n630), .ZN(n632) );
  TPND2D2BWP12T U1702 ( .A1(n633), .A2(n632), .ZN(n662) );
  INVD2P3BWP12T U1703 ( .I(n2682), .ZN(n635) );
  TPNR2D2BWP12T U1704 ( .A1(n1512), .A2(n653), .ZN(n634) );
  CKND2D2BWP12T U1705 ( .A1(n635), .A2(n634), .ZN(n636) );
  TPOAI21D2BWP12T U1706 ( .A1(n2680), .A2(n653), .B(n636), .ZN(n660) );
  NR2D1BWP12T U1707 ( .A1(n662), .A2(n660), .ZN(n641) );
  XNR2D1BWP12T U1708 ( .A1(n2098), .A2(n2746), .ZN(n656) );
  NR2D1BWP12T U1709 ( .A1(n656), .A2(n2747), .ZN(n639) );
  NR2D1BWP12T U1710 ( .A1(n637), .A2(n2748), .ZN(n638) );
  TPND2D1BWP12T U1711 ( .A1(n662), .A2(n660), .ZN(n640) );
  TPOAI21D2BWP12T U1712 ( .A1(n641), .A2(n661), .B(n640), .ZN(n751) );
  INVD1BWP12T U1713 ( .I(n4316), .ZN(n971) );
  XNR2XD4BWP12T U1714 ( .A1(n4926), .A2(a[14]), .ZN(n2669) );
  TPNR2D1BWP12T U1715 ( .A1(n971), .A2(n2669), .ZN(n738) );
  XNR2XD4BWP12T U1716 ( .A1(n341), .A2(n2701), .ZN(n713) );
  XNR2XD2BWP12T U1717 ( .A1(n2071), .A2(n5014), .ZN(n743) );
  XOR3D2BWP12T U1718 ( .A1(n738), .A2(n737), .A3(n736), .Z(n750) );
  INVD1BWP12T U1719 ( .I(n648), .ZN(n644) );
  CKND2D2BWP12T U1720 ( .A1(n647), .A2(n646), .ZN(n651) );
  ND2XD1BWP12T U1721 ( .A1(n649), .A2(n648), .ZN(n650) );
  TPND2D2BWP12T U1722 ( .A1(n651), .A2(n650), .ZN(n749) );
  XOR3XD4BWP12T U1723 ( .A1(n751), .A2(n750), .A3(n749), .Z(n757) );
  XNR2XD4BWP12T U1724 ( .A1(n2167), .A2(n288), .ZN(n716) );
  TPOAI22D2BWP12T U1725 ( .A1(n652), .A2(n1442), .B1(n716), .B2(n2647), .ZN(
        n705) );
  INVD1P75BWP12T U1726 ( .I(n747), .ZN(n655) );
  TPOAI22D2BWP12T U1727 ( .A1(n655), .A2(n2682), .B1(n654), .B2(n2680), .ZN(
        n704) );
  XNR2XD2BWP12T U1728 ( .A1(n4754), .A2(n2746), .ZN(n732) );
  TPOAI22D1BWP12T U1729 ( .A1(n656), .A2(n2748), .B1(n732), .B2(n2747), .ZN(
        n702) );
  XOR3D2BWP12T U1730 ( .A1(n705), .A2(n704), .A3(n702), .Z(n728) );
  XNR2XD8BWP12T U1731 ( .A1(n2619), .A2(n2593), .ZN(n742) );
  TPOAI22D4BWP12T U1732 ( .A1(n657), .A2(n2646), .B1(n742), .B2(n4257), .ZN(
        n719) );
  XNR2D1BWP12T U1733 ( .A1(n2575), .A2(n2742), .ZN(n670) );
  XNR2XD4BWP12T U1734 ( .A1(n2623), .A2(n2742), .ZN(n733) );
  HA1D2BWP12T U1735 ( .A(n659), .B(n658), .CO(n718), .S(n646) );
  XOR3D2BWP12T U1736 ( .A1(n719), .A2(n720), .A3(n718), .Z(n729) );
  INVD1P75BWP12T U1737 ( .I(n660), .ZN(n663) );
  XNR3XD4BWP12T U1738 ( .A1(n663), .A2(n662), .A3(n661), .ZN(n674) );
  OAI21D1BWP12T U1739 ( .A1(n665), .A2(n666), .B(n664), .ZN(n668) );
  TPND2D1BWP12T U1740 ( .A1(n666), .A2(n665), .ZN(n667) );
  TPND2D2BWP12T U1741 ( .A1(n668), .A2(n667), .ZN(n675) );
  OAI22D1BWP12T U1742 ( .A1(n670), .A2(n2743), .B1(n669), .B2(n2744), .ZN(n676) );
  TPNR2D1BWP12T U1743 ( .A1(n675), .A2(n676), .ZN(n673) );
  INVD1BWP12T U1744 ( .I(n676), .ZN(n672) );
  INVD2BWP12T U1745 ( .I(n675), .ZN(n671) );
  XOR3XD4BWP12T U1746 ( .A1(n728), .A2(n729), .A3(n726), .Z(n755) );
  XNR3XD4BWP12T U1747 ( .A1(n756), .A2(n757), .A3(n755), .ZN(n701) );
  NR2D1BWP12T U1748 ( .A1(n678), .A2(n677), .ZN(n681) );
  ND2D1BWP12T U1749 ( .A1(n678), .A2(n677), .ZN(n679) );
  TPOAI21D2BWP12T U1750 ( .A1(n681), .A2(n680), .B(n679), .ZN(n695) );
  INR2D4BWP12T U1751 ( .A1(n696), .B1(n695), .ZN(n687) );
  XOR3XD4BWP12T U1752 ( .A1(n684), .A2(n685), .A3(n683), .Z(n694) );
  IND2D2BWP12T U1753 ( .A1(n696), .B1(n695), .ZN(n686) );
  TPOAI21D2BWP12T U1754 ( .A1(n687), .A2(n694), .B(n686), .ZN(n699) );
  ND2XD4BWP12T U1755 ( .A1(n701), .A2(n688), .ZN(n4009) );
  OAI21D1BWP12T U1756 ( .A1(n690), .A2(n691), .B(n689), .ZN(n693) );
  ND2D1BWP12T U1757 ( .A1(n691), .A2(n690), .ZN(n692) );
  AN2XD2BWP12T U1758 ( .A1(n693), .A2(n692), .Z(n697) );
  XNR3XD4BWP12T U1759 ( .A1(n696), .A2(n695), .A3(n694), .ZN(n698) );
  ND2D3BWP12T U1760 ( .A1(n697), .A2(n698), .ZN(n4005) );
  NR2XD2BWP12T U1761 ( .A1(n698), .A2(n697), .ZN(n3169) );
  TPNR2D3BWP12T U1762 ( .A1(n701), .A2(n700), .ZN(n4011) );
  RCAOI21D4BWP12T U1763 ( .A1(n3169), .A2(n4009), .B(n4011), .ZN(n1027) );
  OAI21D1BWP12T U1764 ( .A1(n704), .A2(n705), .B(n702), .ZN(n703) );
  IOA21D2BWP12T U1765 ( .A1(n705), .A2(n704), .B(n703), .ZN(n1072) );
  TPND2D2BWP12T U1766 ( .A1(n706), .A2(n2170), .ZN(n711) );
  TPAOI21D1BWP12T U1767 ( .A1(n1058), .A2(a[14]), .B(n1164), .ZN(n709) );
  INVD4BWP12T U1768 ( .I(n707), .ZN(n708) );
  OR2D8BWP12T U1769 ( .A1(n709), .A2(n708), .Z(n2667) );
  DCCKND4BWP12T U1770 ( .I(n2704), .ZN(n712) );
  INR2D4BWP12T U1771 ( .A1(n712), .B1(n329), .ZN(n715) );
  TPNR2D3BWP12T U1772 ( .A1(n713), .A2(n2702), .ZN(n714) );
  XOR3XD4BWP12T U1773 ( .A1(n1054), .A2(n1052), .A3(n717), .Z(n1073) );
  INVD1BWP12T U1774 ( .I(n718), .ZN(n722) );
  ND2D1BWP12T U1775 ( .A1(n720), .A2(n719), .ZN(n721) );
  INVD1BWP12T U1776 ( .I(n729), .ZN(n725) );
  INVD1BWP12T U1777 ( .I(n728), .ZN(n724) );
  CKND2D2BWP12T U1778 ( .A1(n727), .A2(n726), .ZN(n731) );
  ND2D1BWP12T U1779 ( .A1(n729), .A2(n728), .ZN(n730) );
  TPND2D2BWP12T U1780 ( .A1(n731), .A2(n730), .ZN(n1140) );
  XNR2XD4BWP12T U1781 ( .A1(n2575), .A2(n2746), .ZN(n1064) );
  TPOAI22D2BWP12T U1782 ( .A1(n733), .A2(n2744), .B1(n1067), .B2(n2743), .ZN(
        n1042) );
  INVD1BWP12T U1783 ( .I(n738), .ZN(n734) );
  IND2XD2BWP12T U1784 ( .A1(n737), .B1(n734), .ZN(n735) );
  TPND2D1BWP12T U1785 ( .A1(n738), .A2(n737), .ZN(n739) );
  TPND2D2BWP12T U1786 ( .A1(n740), .A2(n739), .ZN(n1040) );
  XNR2D1BWP12T U1787 ( .A1(n4316), .A2(n2666), .ZN(n741) );
  XNR2D1BWP12T U1788 ( .A1(n2551), .A2(n2593), .ZN(n1048) );
  NR2D2BWP12T U1789 ( .A1(n2263), .A2(n743), .ZN(n745) );
  XNR2D1BWP12T U1790 ( .A1(n4628), .A2(n5014), .ZN(n1061) );
  TPNR2D2BWP12T U1791 ( .A1(n1061), .A2(n2739), .ZN(n744) );
  NR2D2BWP12T U1792 ( .A1(n745), .A2(n744), .ZN(n1066) );
  XOR2XD2BWP12T U1793 ( .A1(b[3]), .A2(n1164), .Z(n1060) );
  TPNR2D2BWP12T U1794 ( .A1(n1060), .A2(n2682), .ZN(n746) );
  TPAOI21D2BWP12T U1795 ( .A1(n748), .A2(n747), .B(n746), .ZN(n1065) );
  XNR2XD4BWP12T U1796 ( .A1(n1066), .A2(n1065), .ZN(n1039) );
  XNR3XD4BWP12T U1797 ( .A1(n1035), .A2(n1036), .A3(n1039), .ZN(n1125) );
  TPNR2D1BWP12T U1798 ( .A1(n751), .A2(n750), .ZN(n754) );
  INVD1BWP12T U1799 ( .I(n749), .ZN(n753) );
  TPOAI21D2BWP12T U1800 ( .A1(n754), .A2(n753), .B(n752), .ZN(n1122) );
  XNR3XD4BWP12T U1801 ( .A1(n1124), .A2(n1125), .A3(n1122), .ZN(n1144) );
  XNR3XD4BWP12T U1802 ( .A1(n1139), .A2(n1140), .A3(n1144), .ZN(n761) );
  OAI21D1BWP12T U1803 ( .A1(n757), .A2(n756), .B(n755), .ZN(n759) );
  ND2D1BWP12T U1804 ( .A1(n757), .A2(n756), .ZN(n758) );
  NR2XD2BWP12T U1805 ( .A1(n761), .A2(n760), .ZN(n1026) );
  INVD1BWP12T U1806 ( .I(n1026), .ZN(n762) );
  CKND2D2BWP12T U1807 ( .A1(n761), .A2(n760), .ZN(n1025) );
  ND2D1BWP12T U1808 ( .A1(n762), .A2(n1025), .ZN(n763) );
  ND2XD3BWP12T U1809 ( .A1(n4282), .A2(n5085), .ZN(n943) );
  INR2D1BWP12T U1810 ( .A1(op[1]), .B1(op[0]), .ZN(n909) );
  BUFFD6BWP12T U1811 ( .I(b[2]), .Z(n4742) );
  INVD4BWP12T U1812 ( .I(b[3]), .ZN(n4685) );
  INVD8BWP12T U1813 ( .I(n4685), .ZN(n4743) );
  CKBD1BWP12T U1814 ( .I(n4913), .Z(n817) );
  INR2D1BWP12T U1815 ( .A1(n4109), .B1(n1770), .ZN(n767) );
  INVD1BWP12T U1816 ( .I(n2096), .ZN(n983) );
  TPNR2D1BWP12T U1817 ( .A1(n983), .A2(n4911), .ZN(n4226) );
  CKND2D1BWP12T U1818 ( .A1(n4910), .A2(c_in), .ZN(n4951) );
  ND2D1BWP12T U1819 ( .A1(n983), .A2(n4911), .ZN(n4227) );
  OAI21D1BWP12T U1820 ( .A1(n4226), .A2(n4951), .B(n4227), .ZN(n4110) );
  INVD1P25BWP12T U1821 ( .I(n4742), .ZN(n4848) );
  ND2D1BWP12T U1822 ( .A1(n4848), .A2(n4912), .ZN(n4108) );
  ND2D1BWP12T U1823 ( .A1(n4685), .A2(n817), .ZN(n4112) );
  OAI21D1BWP12T U1824 ( .A1(n1770), .A2(n4108), .B(n4112), .ZN(n766) );
  INVD1BWP12T U1825 ( .I(b[4]), .ZN(n768) );
  BUFFD12BWP12T U1826 ( .I(n768), .Z(n4707) );
  NR2D1BWP12T U1827 ( .A1(n4707), .A2(n4921), .ZN(n3357) );
  BUFFD2BWP12T U1828 ( .I(n4628), .Z(n4741) );
  INVD1BWP12T U1829 ( .I(n4741), .ZN(n4684) );
  NR2D1BWP12T U1830 ( .A1(n4684), .A2(n2746), .ZN(n3346) );
  NR2D1BWP12T U1831 ( .A1(n3357), .A2(n3346), .ZN(n3651) );
  CKBD1BWP12T U1832 ( .I(n2094), .Z(n3234) );
  INVD1BWP12T U1833 ( .I(n3234), .ZN(n769) );
  TPNR2D1BWP12T U1834 ( .A1(n769), .A2(n288), .ZN(n3412) );
  INVD2BWP12T U1835 ( .I(n4748), .ZN(n4706) );
  NR2D1BWP12T U1836 ( .A1(n4706), .A2(n4931), .ZN(n3602) );
  TPNR2D1BWP12T U1837 ( .A1(n3412), .A2(n3602), .ZN(n771) );
  CKND2D1BWP12T U1838 ( .A1(n4707), .A2(n4921), .ZN(n3360) );
  CKND2D1BWP12T U1839 ( .A1(n4684), .A2(n2746), .ZN(n3599) );
  OAI21D1BWP12T U1840 ( .A1(n3360), .A2(n3346), .B(n3599), .ZN(n3650) );
  ND2D1BWP12T U1841 ( .A1(n4706), .A2(n4931), .ZN(n3603) );
  ND2D1BWP12T U1842 ( .A1(n769), .A2(n288), .ZN(n3411) );
  OAI21D1BWP12T U1843 ( .A1(n3412), .A2(n3603), .B(n3411), .ZN(n770) );
  AOI21D1BWP12T U1844 ( .A1(n3650), .A2(n771), .B(n770), .ZN(n772) );
  OAI21D1BWP12T U1845 ( .A1(n3358), .A2(n773), .B(n772), .ZN(n776) );
  CKBD1BWP12T U1846 ( .I(n5075), .Z(n4486) );
  NR2D1BWP12T U1847 ( .A1(n773), .A2(n4486), .ZN(n774) );
  NR2D1BWP12T U1848 ( .A1(n4910), .A2(c_in), .ZN(n4224) );
  NR2D1BWP12T U1849 ( .A1(n4226), .A2(n4224), .ZN(n1769) );
  ND2D1BWP12T U1850 ( .A1(n1769), .A2(n4109), .ZN(n4111) );
  NR2D1BWP12T U1851 ( .A1(n4111), .A2(n1770), .ZN(n3649) );
  AN2D1BWP12T U1852 ( .A1(n774), .A2(n3649), .Z(n775) );
  INVD2BWP12T U1853 ( .I(n1614), .ZN(n4971) );
  BUFFD3BWP12T U1854 ( .I(n2167), .Z(n4749) );
  CKBD1BWP12T U1855 ( .I(a[8]), .Z(n4905) );
  NR2D1BWP12T U1856 ( .A1(n4705), .A2(n4905), .ZN(n796) );
  INVD1BWP12T U1857 ( .I(n796), .ZN(n3528) );
  ND2D1BWP12T U1858 ( .A1(n3528), .A2(n351), .ZN(n4965) );
  CKBD1BWP12T U1859 ( .I(n4754), .Z(n3296) );
  INVD1BWP12T U1860 ( .I(n3296), .ZN(n4676) );
  TPNR2D1BWP12T U1861 ( .A1(n4676), .A2(n4904), .ZN(n4967) );
  INVD1BWP12T U1862 ( .I(n4967), .ZN(n3271) );
  CKBD1BWP12T U1863 ( .I(n2575), .Z(n5015) );
  INVD1BWP12T U1864 ( .I(n5014), .ZN(n777) );
  ND2D1BWP12T U1865 ( .A1(n5015), .A2(n777), .ZN(n4973) );
  ND2D1BWP12T U1866 ( .A1(n3271), .A2(n4973), .ZN(n782) );
  NR2D1BWP12T U1867 ( .A1(n4965), .A2(n782), .ZN(n1703) );
  INVD1BWP12T U1868 ( .I(n1703), .ZN(n4014) );
  INVD1BWP12T U1869 ( .I(n2623), .ZN(n4674) );
  CKBD1BWP12T U1870 ( .I(a[12]), .Z(n4925) );
  NR2D1BWP12T U1871 ( .A1(n4674), .A2(n4925), .ZN(n3173) );
  INVD1BWP12T U1872 ( .I(n3173), .ZN(n1697) );
  CKBD1BWP12T U1873 ( .I(n4926), .Z(n783) );
  ND2D1BWP12T U1874 ( .A1(n1697), .A2(n3176), .ZN(n4016) );
  CKND0BWP12T U1875 ( .I(n4016), .ZN(n778) );
  CKBD1BWP12T U1876 ( .I(n2619), .Z(n4752) );
  CKBD1BWP12T U1877 ( .I(a[14]), .Z(n4932) );
  CKND2D1BWP12T U1878 ( .A1(n778), .A2(n4021), .ZN(n786) );
  NR2D1BWP12T U1879 ( .A1(n4014), .A2(n786), .ZN(n788) );
  CKND2D1BWP12T U1880 ( .A1(n4705), .A2(n4905), .ZN(n3383) );
  INVD1BWP12T U1881 ( .I(n3383), .ZN(n3527) );
  INVD1BWP12T U1882 ( .I(n4765), .ZN(n4704) );
  ND2D1BWP12T U1883 ( .A1(n4704), .A2(n4906), .ZN(n3529) );
  INVD1BWP12T U1884 ( .I(n3529), .ZN(n3270) );
  AOI21D1BWP12T U1885 ( .A1(n351), .A2(n3527), .B(n3270), .ZN(n4968) );
  ND2D1BWP12T U1886 ( .A1(n4676), .A2(n4904), .ZN(n4966) );
  INVD0BWP12T U1887 ( .I(n4966), .ZN(n780) );
  CKND0BWP12T U1888 ( .I(n2575), .ZN(n4675) );
  ND2D1BWP12T U1889 ( .A1(n4675), .A2(n4449), .ZN(n4972) );
  INVD1BWP12T U1890 ( .I(n4972), .ZN(n779) );
  AOI21D1BWP12T U1891 ( .A1(n4973), .A2(n780), .B(n779), .ZN(n781) );
  OAI21D1BWP12T U1892 ( .A1(n4968), .A2(n782), .B(n781), .ZN(n1702) );
  INVD1BWP12T U1893 ( .I(n1702), .ZN(n4017) );
  CKND2D1BWP12T U1894 ( .A1(n4674), .A2(n4925), .ZN(n3172) );
  ND2D1BWP12T U1895 ( .A1(n4673), .A2(n783), .ZN(n4071) );
  CKND0BWP12T U1896 ( .I(n4015), .ZN(n784) );
  CKND2D1BWP12T U1897 ( .A1(n803), .A2(n4932), .ZN(n4020) );
  INVD1BWP12T U1898 ( .I(n4020), .ZN(n1606) );
  TPAOI21D0BWP12T U1899 ( .A1(n784), .A2(n4021), .B(n1606), .ZN(n785) );
  OAI21D1BWP12T U1900 ( .A1(n4017), .A2(n786), .B(n785), .ZN(n787) );
  AOI21D1BWP12T U1901 ( .A1(n4971), .A2(n788), .B(n787), .ZN(n789) );
  CKBD1BWP12T U1902 ( .I(n2551), .Z(n4759) );
  ND2D1BWP12T U1903 ( .A1(n4687), .A2(n2666), .ZN(n1588) );
  CKND2D1BWP12T U1904 ( .A1(n1607), .A2(n1588), .ZN(n812) );
  XOR2XD1BWP12T U1905 ( .A1(n789), .A2(n812), .Z(n4949) );
  INVD1BWP12T U1906 ( .I(n4949), .ZN(n942) );
  INVD0BWP12T U1907 ( .I(op[0]), .ZN(n790) );
  IND2XD1BWP12T U1908 ( .A1(op[2]), .B1(op[1]), .ZN(n833) );
  INVD4BWP12T U1909 ( .I(n4318), .ZN(n5090) );
  INVD1BWP12T U1910 ( .I(n4244), .ZN(n1787) );
  NR2D1BWP12T U1911 ( .A1(n796), .A2(n3412), .ZN(n798) );
  NR2D1BWP12T U1912 ( .A1(n3602), .A2(n3346), .ZN(n3409) );
  ND2D1BWP12T U1913 ( .A1(n798), .A2(n3409), .ZN(n800) );
  CKBD1BWP12T U1914 ( .I(n4913), .Z(n4560) );
  ND2D1BWP12T U1915 ( .A1(n4743), .A2(n1785), .ZN(n4134) );
  INVD15BWP12T U1916 ( .I(n4707), .ZN(n4843) );
  ND2D1BWP12T U1917 ( .A1(n4843), .A2(n1765), .ZN(n1784) );
  INVD1BWP12T U1918 ( .I(n4742), .ZN(n3051) );
  TPNR2D1BWP12T U1919 ( .A1(n975), .A2(n4226), .ZN(n4131) );
  CKND2D1BWP12T U1920 ( .A1(n1784), .A2(n4131), .ZN(n791) );
  OR2D2BWP12T U1921 ( .A1(n1770), .A2(n791), .Z(n3345) );
  NR2D1BWP12T U1922 ( .A1(n800), .A2(n3345), .ZN(n802) );
  NR2D0BWP12T U1923 ( .A1(n4743), .A2(n1785), .ZN(n792) );
  CKND2D1BWP12T U1924 ( .A1(n792), .A2(n1784), .ZN(n793) );
  ND2D1BWP12T U1925 ( .A1(n793), .A2(n3360), .ZN(n795) );
  AN3XD1BWP12T U1926 ( .A1(n1786), .A2(n4134), .A3(n1784), .Z(n794) );
  NR2D2BWP12T U1927 ( .A1(n795), .A2(n794), .ZN(n3344) );
  OAI21D1BWP12T U1928 ( .A1(n3602), .A2(n3599), .B(n3603), .ZN(n3410) );
  OAI21D1BWP12T U1929 ( .A1(n796), .A2(n3411), .B(n3383), .ZN(n797) );
  AOI21D1BWP12T U1930 ( .A1(n798), .A2(n3410), .B(n797), .ZN(n799) );
  OAI21D1BWP12T U1931 ( .A1(n800), .A2(n3344), .B(n799), .ZN(n801) );
  INVD1P75BWP12T U1932 ( .I(n1596), .ZN(n4333) );
  NR2D1BWP12T U1933 ( .A1(n4704), .A2(n4906), .ZN(n3269) );
  NR2D1BWP12T U1934 ( .A1(n4967), .A2(n3269), .ZN(n4332) );
  NR2D1BWP12T U1935 ( .A1(n4675), .A2(n4449), .ZN(n4334) );
  NR2D1BWP12T U1936 ( .A1(n4334), .A2(n3173), .ZN(n806) );
  ND2D1BWP12T U1937 ( .A1(n4332), .A2(n806), .ZN(n4070) );
  CKBD1BWP12T U1938 ( .I(n4926), .Z(n804) );
  NR2D1BWP12T U1939 ( .A1(n4673), .A2(n804), .ZN(n4072) );
  NR2D1BWP12T U1940 ( .A1(n807), .A2(n4072), .ZN(n1587) );
  INVD1BWP12T U1941 ( .I(n1587), .ZN(n809) );
  TPNR2D0BWP12T U1942 ( .A1(n4070), .A2(n809), .ZN(n811) );
  OAI21D1BWP12T U1943 ( .A1(n4967), .A2(n3529), .B(n4966), .ZN(n4331) );
  OAI21D1BWP12T U1944 ( .A1(n3173), .A2(n4972), .B(n3172), .ZN(n805) );
  TPAOI21D1BWP12T U1945 ( .A1(n806), .A2(n4331), .B(n805), .ZN(n4073) );
  OAI21D1BWP12T U1946 ( .A1(n807), .A2(n4071), .B(n4020), .ZN(n1589) );
  INVD1BWP12T U1947 ( .I(n1589), .ZN(n808) );
  TPOAI21D0BWP12T U1948 ( .A1(n4073), .A2(n809), .B(n808), .ZN(n810) );
  AOI21D1BWP12T U1949 ( .A1(n4333), .A2(n811), .B(n810), .ZN(n813) );
  XOR2XD1BWP12T U1950 ( .A1(n813), .A2(n812), .Z(n4342) );
  TPNR2D2BWP12T U1951 ( .A1(n4742), .A2(n4912), .ZN(n4114) );
  NR2D1BWP12T U1952 ( .A1(n1709), .A2(n4214), .ZN(n961) );
  CKND1BWP12T U1953 ( .I(n961), .ZN(n4230) );
  IND2XD1BWP12T U1954 ( .A1(n4114), .B1(n4230), .ZN(n816) );
  CKND2D1BWP12T U1955 ( .A1(n4486), .A2(n4910), .ZN(n4487) );
  INVD1BWP12T U1956 ( .I(n992), .ZN(n4645) );
  ND2D1BWP12T U1957 ( .A1(n4645), .A2(n4214), .ZN(n4229) );
  INVD1BWP12T U1958 ( .I(n4229), .ZN(n814) );
  INVD1BWP12T U1959 ( .I(n4114), .ZN(n887) );
  ND2D1BWP12T U1960 ( .A1(n4742), .A2(n4912), .ZN(n963) );
  INVD1BWP12T U1961 ( .I(n963), .ZN(n4116) );
  AOI21D1BWP12T U1962 ( .A1(n814), .A2(n887), .B(n4116), .ZN(n815) );
  OAI21D1BWP12T U1963 ( .A1(n816), .A2(n4487), .B(n815), .ZN(n1774) );
  NR2D4BWP12T U1964 ( .A1(n4743), .A2(n817), .ZN(n1775) );
  INVD1BWP12T U1965 ( .I(n1775), .ZN(n4101) );
  ND2D1BWP12T U1966 ( .A1(n4101), .A2(n3352), .ZN(n3626) );
  OR2D2BWP12T U1967 ( .A1(n4748), .A2(n4931), .Z(n3633) );
  OR2XD1BWP12T U1968 ( .A1(n4741), .A2(n2746), .Z(n3366) );
  ND2D1BWP12T U1969 ( .A1(n3633), .A2(n3366), .ZN(n820) );
  NR2D1BWP12T U1970 ( .A1(n3626), .A2(n820), .ZN(n822) );
  INVD0BWP12T U1971 ( .I(n4100), .ZN(n818) );
  CKND2D1BWP12T U1972 ( .A1(n4843), .A2(n4921), .ZN(n1776) );
  INVD1BWP12T U1973 ( .I(n1776), .ZN(n3351) );
  AOI21D1BWP12T U1974 ( .A1(n3352), .A2(n818), .B(n3351), .ZN(n3629) );
  CKND2D1BWP12T U1975 ( .A1(n4741), .A2(n2746), .ZN(n3627) );
  ND2D1BWP12T U1976 ( .A1(n4748), .A2(n4931), .ZN(n3632) );
  OAI21D1BWP12T U1977 ( .A1(n3629), .A2(n820), .B(n819), .ZN(n821) );
  NR2D1BWP12T U1978 ( .A1(n3296), .A2(n4904), .ZN(n4380) );
  NR2D1BWP12T U1979 ( .A1(n4765), .A2(n4906), .ZN(n3283) );
  NR2D1BWP12T U1980 ( .A1(n4380), .A2(n3283), .ZN(n824) );
  NR2D1BWP12T U1981 ( .A1(n3234), .A2(n288), .ZN(n3214) );
  NR2D1BWP12T U1982 ( .A1(n891), .A2(n3214), .ZN(n3533) );
  ND2D1BWP12T U1983 ( .A1(n824), .A2(n3533), .ZN(n826) );
  ND2D1BWP12T U1984 ( .A1(n3234), .A2(n288), .ZN(n3402) );
  ND2D1BWP12T U1985 ( .A1(n4749), .A2(n4905), .ZN(n3398) );
  OAI21D1BWP12T U1986 ( .A1(n891), .A2(n3402), .B(n3398), .ZN(n3532) );
  ND2D1BWP12T U1987 ( .A1(n4765), .A2(n4906), .ZN(n3535) );
  ND2D1BWP12T U1988 ( .A1(n3296), .A2(n4904), .ZN(n4379) );
  OAI21D1BWP12T U1989 ( .A1(n4380), .A2(n3535), .B(n4379), .ZN(n823) );
  AOI21D1BWP12T U1990 ( .A1(n824), .A2(n3532), .B(n823), .ZN(n825) );
  NR2D1BWP12T U1991 ( .A1(n5015), .A2(n5014), .ZN(n1691) );
  NR2D0BWP12T U1992 ( .A1(n2623), .A2(n4925), .ZN(n3208) );
  NR2D1BWP12T U1993 ( .A1(n1691), .A2(n3208), .ZN(n4023) );
  NR2D1BWP12T U1994 ( .A1(n4752), .A2(n4932), .ZN(n828) );
  CKBD1BWP12T U1995 ( .I(n4926), .Z(n827) );
  ND2D1BWP12T U1996 ( .A1(n4023), .A2(n830), .ZN(n1802) );
  CKND2D1BWP12T U1997 ( .A1(n5015), .A2(n5014), .ZN(n4491) );
  INVD1BWP12T U1998 ( .I(n4674), .ZN(n4760) );
  OAI21D1BWP12T U1999 ( .A1(n3208), .A2(n4491), .B(n3207), .ZN(n4026) );
  CKBD1BWP12T U2000 ( .I(n4926), .Z(n892) );
  ND2XD0BWP12T U2001 ( .A1(n4753), .A2(n892), .ZN(n3200) );
  ND2D1BWP12T U2002 ( .A1(n4752), .A2(n4932), .ZN(n4029) );
  OAI21D1BWP12T U2003 ( .A1(n828), .A2(n3200), .B(n4029), .ZN(n829) );
  AOI21D1BWP12T U2004 ( .A1(n830), .A2(n4026), .B(n829), .ZN(n1803) );
  OAI21D1BWP12T U2005 ( .A1(n4493), .A2(n1802), .B(n1803), .ZN(n832) );
  NR2D1BWP12T U2006 ( .A1(n4759), .A2(n2666), .ZN(n1641) );
  INVD1BWP12T U2007 ( .I(n1641), .ZN(n4183) );
  CKND2D1BWP12T U2008 ( .A1(n4759), .A2(n2666), .ZN(n1642) );
  CKND2D1BWP12T U2009 ( .A1(n4183), .A2(n1642), .ZN(n831) );
  AOI22D1BWP12T U2010 ( .A1(n5090), .A2(n4342), .B1(n4508), .B2(n4103), .ZN(
        n941) );
  NR2D3BWP12T U2011 ( .A1(n992), .A2(n5075), .ZN(n3217) );
  INVD8BWP12T U2012 ( .I(a[17]), .ZN(n1810) );
  CKBD1BWP12T U2013 ( .I(a[16]), .Z(n4927) );
  OAI22D1BWP12T U2014 ( .A1(n3321), .A2(n1810), .B1(n275), .B2(n4638), .ZN(
        n837) );
  IND2XD8BWP12T U2015 ( .A1(n5075), .B1(n4686), .ZN(n3323) );
  INVD4BWP12T U2016 ( .I(n5075), .ZN(n835) );
  NR2D4BWP12T U2017 ( .A1(n835), .A2(n992), .ZN(n3220) );
  INVD3BWP12T U2018 ( .I(n3220), .ZN(n3322) );
  BUFFD6BWP12T U2019 ( .I(a[18]), .Z(n4923) );
  INVD1BWP12T U2020 ( .I(n4923), .ZN(n4637) );
  OAI22D0BWP12T U2021 ( .A1(n3323), .A2(n4930), .B1(n3322), .B2(n4637), .ZN(
        n836) );
  NR2D1BWP12T U2022 ( .A1(n837), .A2(n836), .ZN(n4522) );
  NR2D4BWP12T U2023 ( .A1(n5075), .A2(n4738), .ZN(n3219) );
  DCCKND4BWP12T U2024 ( .I(a[19]), .ZN(n1652) );
  INVD4BWP12T U2025 ( .I(a[21]), .ZN(n838) );
  INVD12BWP12T U2026 ( .I(n838), .ZN(n4914) );
  BUFFD6BWP12T U2027 ( .I(a[20]), .Z(n5051) );
  ND2D1BWP12T U2028 ( .A1(n3218), .A2(n5051), .ZN(n840) );
  BUFFD6BWP12T U2029 ( .I(a[22]), .Z(n4728) );
  TPND2D0BWP12T U2030 ( .A1(n3220), .A2(n4915), .ZN(n839) );
  OAI211D1BWP12T U2031 ( .A1(n3321), .A2(n4625), .B(n840), .C(n839), .ZN(n841)
         );
  AOI21D1BWP12T U2032 ( .A1(n3219), .A2(n3771), .B(n841), .ZN(n4517) );
  MUX2D1BWP12T U2033 ( .I0(n4522), .I1(n4517), .S(n4742), .Z(n3223) );
  INVD4BWP12T U2034 ( .I(a[29]), .ZN(n982) );
  BUFFD6BWP12T U2035 ( .I(a[28]), .Z(n4908) );
  INVD1BWP12T U2036 ( .I(n4908), .ZN(n4665) );
  OAI22D1BWP12T U2037 ( .A1(n3321), .A2(n4664), .B1(n275), .B2(n4665), .ZN(
        n843) );
  BUFFXD3BWP12T U2038 ( .I(a[27]), .Z(n3040) );
  INVD1BWP12T U2039 ( .I(n3040), .ZN(n4667) );
  BUFFD6BWP12T U2040 ( .I(a[30]), .Z(n4933) );
  OAI22D1BWP12T U2041 ( .A1(n3323), .A2(n4667), .B1(n3322), .B2(n4636), .ZN(
        n842) );
  NR2D1BWP12T U2042 ( .A1(n843), .A2(n842), .ZN(n3767) );
  INVD1P75BWP12T U2043 ( .I(n3219), .ZN(n3318) );
  DCCKND4BWP12T U2044 ( .I(a[23]), .ZN(n2981) );
  INVD9BWP12T U2045 ( .I(n2981), .ZN(n4916) );
  CKND3BWP12T U2046 ( .I(n4916), .ZN(n4465) );
  BUFFD6BWP12T U2047 ( .I(a[24]), .Z(n4907) );
  INVD1BWP12T U2048 ( .I(n4907), .ZN(n4650) );
  INVD3BWP12T U2049 ( .I(a[25]), .ZN(n3850) );
  OAI22D1BWP12T U2050 ( .A1(n275), .A2(n4650), .B1(n3321), .B2(n3850), .ZN(
        n846) );
  BUFFD6BWP12T U2051 ( .I(a[26]), .Z(n4922) );
  INVD1BWP12T U2052 ( .I(n4922), .ZN(n4666) );
  INVD0BWP12T U2053 ( .I(n4666), .ZN(n844) );
  INR2D1BWP12T U2054 ( .A1(n844), .B1(n3322), .ZN(n845) );
  NR2D1BWP12T U2055 ( .A1(n846), .A2(n845), .ZN(n847) );
  OA21D1BWP12T U2056 ( .A1(n3318), .A2(n4465), .B(n847), .Z(n4518) );
  IND2D1BWP12T U2057 ( .A1(n4843), .B1(n4743), .ZN(n3968) );
  OAI22D1BWP12T U2058 ( .A1(n3223), .A2(n4611), .B1(n3224), .B2(n3968), .ZN(
        n4528) );
  INVD1BWP12T U2059 ( .I(n4528), .ZN(n849) );
  INR2D8BWP12T U2060 ( .A1(n4848), .B1(n3323), .ZN(n4200) );
  INVD3BWP12T U2061 ( .I(n4200), .ZN(n1673) );
  BUFFD2BWP12T U2062 ( .I(a[31]), .Z(n848) );
  NR3XD0BWP12T U2063 ( .A1(n1673), .A2(n4743), .A3(n4624), .ZN(n4534) );
  CKND2D1BWP12T U2064 ( .A1(n4534), .A2(n4843), .ZN(n4530) );
  ND2D1BWP12T U2065 ( .A1(n849), .A2(n4530), .ZN(n877) );
  BUFFXD4BWP12T U2066 ( .I(b[24]), .Z(n4740) );
  NR2D1BWP12T U2067 ( .A1(n2578), .A2(n4740), .ZN(n921) );
  NR4D0BWP12T U2068 ( .A1(n2575), .A2(n4754), .A3(n2098), .A4(n2167), .ZN(n922) );
  BUFFXD8BWP12T U2069 ( .I(b[21]), .Z(n4726) );
  NR2D1BWP12T U2070 ( .A1(n4726), .A2(n2243), .ZN(n925) );
  BUFFD6BWP12T U2071 ( .I(b[30]), .Z(n4727) );
  NR2D1BWP12T U2072 ( .A1(n4751), .A2(n4727), .ZN(n923) );
  NR4D0BWP12T U2073 ( .A1(n4753), .A2(n2619), .A3(n2623), .A4(n2094), .ZN(n920) );
  ND2D1BWP12T U2074 ( .A1(n923), .A2(n920), .ZN(n850) );
  TPNR2D2BWP12T U2075 ( .A1(n851), .A2(n850), .ZN(n859) );
  BUFFD6BWP12T U2076 ( .I(b[19]), .Z(n4764) );
  BUFFD6BWP12T U2077 ( .I(b[18]), .Z(n2226) );
  NR2D1BWP12T U2078 ( .A1(n336), .A2(n2226), .ZN(n926) );
  NR2D1BWP12T U2079 ( .A1(n280), .A2(n4761), .ZN(n924) );
  BUFFXD4BWP12T U2080 ( .I(b[23]), .Z(n2591) );
  CKND2D0BWP12T U2081 ( .A1(n317), .A2(n347), .ZN(n854) );
  ND3D1BWP12T U2082 ( .A1(n926), .A2(n924), .A3(n919), .ZN(n857) );
  BUFFXD4BWP12T U2083 ( .I(b[29]), .Z(n4730) );
  BUFFD6BWP12T U2084 ( .I(b[28]), .Z(n4733) );
  TPNR2D2BWP12T U2085 ( .A1(n857), .A2(n927), .ZN(n858) );
  CKND2D8BWP12T U2086 ( .A1(n859), .A2(n858), .ZN(n4891) );
  INVD8BWP12T U2087 ( .I(n4891), .ZN(n4573) );
  ND2D1BWP12T U2088 ( .A1(op[0]), .A2(op[1]), .ZN(n860) );
  ND2D1BWP12T U2089 ( .A1(n4573), .A2(n4209), .ZN(n4068) );
  ND2D1BWP12T U2090 ( .A1(n4068), .A2(n5040), .ZN(n5026) );
  XNR2XD8BWP12T U2091 ( .A1(n1673), .A2(n4743), .ZN(n4032) );
  ND2XD4BWP12T U2092 ( .A1(n4032), .A2(n3758), .ZN(n3818) );
  MUX2XD0BWP12T U2093 ( .I0(n4653), .I1(n4652), .S(n5075), .Z(n3120) );
  INVD1BWP12T U2094 ( .I(n3120), .ZN(n3104) );
  INVD1P75BWP12T U2095 ( .I(n3322), .ZN(n862) );
  INR2D4BWP12T U2096 ( .A1(n3318), .B1(n862), .ZN(n3005) );
  ND2D2BWP12T U2097 ( .A1(n3323), .A2(n4742), .ZN(n2887) );
  INVD1BWP12T U2098 ( .I(n2887), .ZN(n863) );
  CKND2D2BWP12T U2099 ( .A1(n3322), .A2(n2887), .ZN(n864) );
  TPNR2D3BWP12T U2100 ( .A1(n864), .A2(n3219), .ZN(n3940) );
  INVD2P3BWP12T U2101 ( .I(n4905), .ZN(n4655) );
  MUX2D1BWP12T U2102 ( .I0(n3523), .I1(n4655), .S(n5075), .Z(n3098) );
  INVD1BWP12T U2103 ( .I(n3098), .ZN(n3112) );
  AOI22D1BWP12T U2104 ( .A1(n3104), .A2(n3939), .B1(n3940), .B2(n3112), .ZN(
        n870) );
  INVD1P75BWP12T U2105 ( .I(n4200), .ZN(n865) );
  ND2D2BWP12T U2106 ( .A1(n865), .A2(n2887), .ZN(n867) );
  TPNR2D3BWP12T U2107 ( .A1(n867), .A2(n3005), .ZN(n3937) );
  MUX2XD0BWP12T U2108 ( .I0(n777), .I1(n4654), .S(n5075), .Z(n3121) );
  INVD1BWP12T U2109 ( .I(n3121), .ZN(n3105) );
  TPND2D0BWP12T U2110 ( .A1(n3937), .A2(n3105), .ZN(n869) );
  INVD2BWP12T U2111 ( .I(n867), .ZN(n3436) );
  MUX2D1BWP12T U2112 ( .I0(n2666), .I1(n4932), .S(n5075), .Z(n3103) );
  CKND2D1BWP12T U2113 ( .A1(n3941), .A2(n3103), .ZN(n868) );
  ND3D1BWP12T U2114 ( .A1(n870), .A2(n869), .A3(n868), .ZN(n1671) );
  MUX2D1BWP12T U2115 ( .I0(n4679), .I1(n4631), .S(n5075), .Z(n3096) );
  INVD1BWP12T U2116 ( .I(n3096), .ZN(n3113) );
  ND2D1BWP12T U2117 ( .A1(n3941), .A2(n3113), .ZN(n876) );
  MUX2XD0BWP12T U2118 ( .I0(n871), .I1(n373), .S(n5075), .Z(n3099) );
  INVD1BWP12T U2119 ( .I(n3099), .ZN(n3115) );
  IND2D1BWP12T U2120 ( .A1(n5075), .B1(n901), .ZN(n872) );
  ND2D1BWP12T U2121 ( .A1(n5075), .A2(n5079), .ZN(n5084) );
  ND2D1BWP12T U2122 ( .A1(n872), .A2(n5084), .ZN(n3061) );
  MUX2D1BWP12T U2123 ( .I0(n4627), .I1(n1765), .S(n5075), .Z(n3100) );
  TPNR2D2BWP12T U2124 ( .A1(n4032), .A2(n4045), .ZN(n4799) );
  AOI22D1BWP12T U2125 ( .A1(n4801), .A2(n1671), .B1(n4779), .B2(n4799), .ZN(
        n4835) );
  MAOI22D1BWP12T U2126 ( .A1(n877), .A2(n5026), .B1(n4835), .B2(n5040), .ZN(
        n939) );
  TPNR2D0BWP12T U2127 ( .A1(n4114), .A2(n1775), .ZN(n880) );
  CKND2D1BWP12T U2128 ( .A1(n4910), .A2(c_in), .ZN(n4394) );
  BUFFD1BWP12T U2129 ( .I(a[1]), .Z(n878) );
  CKND2D2BWP12T U2130 ( .A1(n4645), .A2(n878), .ZN(n4221) );
  OAI21D1BWP12T U2131 ( .A1(n1775), .A2(n963), .B(n4100), .ZN(n879) );
  AOI21D1BWP12T U2132 ( .A1(n880), .A2(n4115), .B(n879), .ZN(n1766) );
  NR2D1BWP12T U2133 ( .A1(n4741), .A2(n2746), .ZN(n3628) );
  TPNR2D1BWP12T U2134 ( .A1(n3214), .A2(n3231), .ZN(n881) );
  ND2D1BWP12T U2135 ( .A1(n3620), .A2(n881), .ZN(n886) );
  NR2D1BWP12T U2136 ( .A1(n1766), .A2(n886), .ZN(n885) );
  OAI21D1BWP12T U2137 ( .A1(n1776), .A2(n3628), .B(n3627), .ZN(n3619) );
  CKND2D1BWP12T U2138 ( .A1(n3619), .A2(n881), .ZN(n883) );
  OA21D1BWP12T U2139 ( .A1(n3214), .A2(n3632), .B(n3402), .Z(n882) );
  CKND2D1BWP12T U2140 ( .A1(n883), .A2(n882), .ZN(n884) );
  TPNR2D1BWP12T U2141 ( .A1(n885), .A2(n884), .ZN(n890) );
  INR2D1BWP12T U2142 ( .A1(n5075), .B1(n886), .ZN(n888) );
  INVD1BWP12T U2143 ( .I(n962), .ZN(n4113) );
  INR3D2BWP12T U2144 ( .A1(n887), .B1(n4113), .B2(n1775), .ZN(n3618) );
  ND2D1BWP12T U2145 ( .A1(n888), .A2(n3618), .ZN(n889) );
  CKND2D2BWP12T U2146 ( .A1(n890), .A2(n889), .ZN(n4384) );
  INVD1BWP12T U2147 ( .I(n891), .ZN(n3515) );
  INVD1BWP12T U2148 ( .I(n3283), .ZN(n3536) );
  ND2D1BWP12T U2149 ( .A1(n3515), .A2(n3536), .ZN(n4378) );
  INVD1BWP12T U2150 ( .I(n4380), .ZN(n3273) );
  INVD1BWP12T U2151 ( .I(n1691), .ZN(n4492) );
  ND2D1BWP12T U2152 ( .A1(n3273), .A2(n4492), .ZN(n895) );
  NR2D1BWP12T U2153 ( .A1(n4378), .A2(n895), .ZN(n3206) );
  CKND0BWP12T U2154 ( .I(n3206), .ZN(n4049) );
  INVD1BWP12T U2155 ( .I(n3208), .ZN(n3205) );
  OR2XD0BWP12T U2156 ( .A1(n4753), .A2(n892), .Z(n4025) );
  ND2D1BWP12T U2157 ( .A1(n3205), .A2(n4025), .ZN(n4051) );
  CKND0BWP12T U2158 ( .I(n4051), .ZN(n893) );
  INVD1BWP12T U2159 ( .I(n3398), .ZN(n3514) );
  INVD1BWP12T U2160 ( .I(n3535), .ZN(n894) );
  AOI21D1BWP12T U2161 ( .A1(n3536), .A2(n3514), .B(n894), .ZN(n4381) );
  INVD1BWP12T U2162 ( .I(n1734), .ZN(n4052) );
  CKND0BWP12T U2163 ( .I(n3207), .ZN(n896) );
  INVD1BWP12T U2164 ( .I(n3200), .ZN(n4024) );
  AOI21D1BWP12T U2165 ( .A1(n4025), .A2(n896), .B(n4024), .ZN(n4050) );
  CKND0BWP12T U2166 ( .I(n4050), .ZN(n897) );
  INVD1BWP12T U2167 ( .I(n4029), .ZN(n1623) );
  INVD1BWP12T U2168 ( .I(n933), .ZN(n899) );
  IND2XD1BWP12T U2169 ( .A1(op[1]), .B1(op[0]), .ZN(n898) );
  TPNR2D2BWP12T U2170 ( .A1(n899), .A2(n898), .ZN(n5088) );
  CKND2D1BWP12T U2171 ( .A1(n4406), .A2(n5088), .ZN(n938) );
  ND2D1BWP12T U2172 ( .A1(n777), .A2(n4654), .ZN(n900) );
  NR2D1BWP12T U2173 ( .A1(n4446), .A2(n900), .ZN(n1721) );
  CKND1BWP12T U2174 ( .I(n1721), .ZN(n4058) );
  CKBD1BWP12T U2175 ( .I(n4926), .Z(n3187) );
  ND2D1BWP12T U2176 ( .A1(n4653), .A2(n4652), .ZN(n4057) );
  INVD1BWP12T U2177 ( .I(n4932), .ZN(n4680) );
  ND2D1BWP12T U2178 ( .A1(n901), .A2(n5079), .ZN(n964) );
  ND2D1BWP12T U2179 ( .A1(n1785), .A2(n373), .ZN(n902) );
  NR2D1BWP12T U2180 ( .A1(n964), .A2(n902), .ZN(n1762) );
  AN2XD1BWP12T U2181 ( .A1(n4679), .A2(n4631), .Z(n903) );
  INVD1BWP12T U2182 ( .I(n3605), .ZN(n3233) );
  AN3XD2BWP12T U2183 ( .A1(n1762), .A2(n903), .A3(n3233), .Z(n4448) );
  NR2D0BWP12T U2184 ( .A1(op[2]), .A2(op[1]), .ZN(n906) );
  ND2D1BWP12T U2185 ( .A1(n904), .A2(n906), .ZN(n4420) );
  INVD4BWP12T U2186 ( .I(n4420), .ZN(n5078) );
  NR2D1BWP12T U2187 ( .A1(op[0]), .A2(op[1]), .ZN(n2870) );
  CKND2D0BWP12T U2188 ( .A1(op[3]), .A2(op[2]), .ZN(n908) );
  INR2D1BWP12T U2189 ( .A1(n2870), .B1(n908), .ZN(n905) );
  CKND0BWP12T U2190 ( .I(op[3]), .ZN(n931) );
  AN3D1BWP12T U2191 ( .A1(n906), .A2(op[0]), .A3(n931), .Z(n4633) );
  NR2D0BWP12T U2192 ( .A1(n2666), .A2(n5083), .ZN(n907) );
  OA21XD0BWP12T U2193 ( .A1(n905), .A2(n907), .B(n4759), .Z(n914) );
  INR2D1BWP12T U2194 ( .A1(n909), .B1(n908), .ZN(n4623) );
  MUX2ND0BWP12T U2195 ( .I0(n5077), .I1(n5076), .S(n4759), .ZN(n910) );
  NR2D0BWP12T U2196 ( .A1(n910), .A2(n905), .ZN(n912) );
  MUX2ND0BWP12T U2197 ( .I0(n912), .I1(n5080), .S(n4930), .ZN(n913) );
  AOI211D1BWP12T U2198 ( .A1(n4439), .A2(n5078), .B(n914), .C(n913), .ZN(n936)
         );
  TPNR2D2BWP12T U2199 ( .A1(n4738), .A2(n4742), .ZN(n3067) );
  INVD4BWP12T U2200 ( .I(n3067), .ZN(n3957) );
  INVD4BWP12T U2201 ( .I(n3957), .ZN(n3125) );
  INVD1BWP12T U2202 ( .I(n3103), .ZN(n3118) );
  AOI22D1BWP12T U2203 ( .A1(n3125), .A2(n3118), .B1(n3120), .B2(n953), .ZN(
        n916) );
  TPND2D1BWP12T U2204 ( .A1(n2096), .A2(n4742), .ZN(n3959) );
  INVD1BWP12T U2205 ( .I(n3959), .ZN(n3122) );
  AOI22D1BWP12T U2206 ( .A1(n3122), .A2(n3098), .B1(n3121), .B2(n3701), .ZN(
        n915) );
  ND2D1BWP12T U2207 ( .A1(n916), .A2(n915), .ZN(n2866) );
  INVD1BWP12T U2208 ( .I(n2866), .ZN(n1655) );
  OAI22D1BWP12T U2209 ( .A1(n3126), .A2(n3959), .B1(n3114), .B2(n3961), .ZN(
        n918) );
  INVD9BWP12T U2210 ( .I(n3701), .ZN(n3963) );
  OAI22D1BWP12T U2211 ( .A1(n3113), .A2(n3957), .B1(n3115), .B2(n3963), .ZN(
        n917) );
  NR2D1BWP12T U2212 ( .A1(n918), .A2(n917), .ZN(n4585) );
  ND4D0BWP12T U2213 ( .A1(n922), .A2(n921), .A3(n920), .A4(n919), .ZN(n929) );
  ND4D1BWP12T U2214 ( .A1(n926), .A2(n925), .A3(n924), .A4(n923), .ZN(n928) );
  NR4D1BWP12T U2215 ( .A1(n929), .A2(n928), .A3(n927), .A4(n4843), .ZN(n930)
         );
  INVD3BWP12T U2216 ( .I(n930), .ZN(n4890) );
  INVD6BWP12T U2217 ( .I(n4890), .ZN(n4605) );
  TPNR2D3BWP12T U2218 ( .A1(n4605), .A2(n4624), .ZN(n3982) );
  TPAOI21D0BWP12T U2219 ( .A1(n4528), .A2(n4573), .B(n3982), .ZN(n4872) );
  ND2D1BWP12T U2220 ( .A1(n933), .A2(n2870), .ZN(n5063) );
  NR2XD0BWP12T U2221 ( .A1(n4872), .A2(n5063), .ZN(n934) );
  INR3XD1BWP12T U2222 ( .A1(n936), .B1(n935), .B2(n934), .ZN(n937) );
  AN3XD2BWP12T U2223 ( .A1(n939), .A2(n938), .A3(n937), .Z(n940) );
  ND2D8BWP12T U2224 ( .A1(n943), .A2(n350), .ZN(result[15]) );
  TPAOI22D0BWP12T U2225 ( .A1(n3218), .A2(n777), .B1(n3217), .B2(n4652), .ZN(
        n945) );
  AOI22D0BWP12T U2226 ( .A1(n3220), .A2(n4653), .B1(n3219), .B2(n4654), .ZN(
        n944) );
  ND2D1BWP12T U2227 ( .A1(n945), .A2(n944), .ZN(n3638) );
  INVD1BWP12T U2228 ( .I(n3638), .ZN(n3274) );
  IND2D2BWP12T U2229 ( .A1(n4742), .B1(n4743), .ZN(n4206) );
  AOI22D0BWP12T U2230 ( .A1(n3218), .A2(n2666), .B1(n3217), .B2(n4927), .ZN(
        n947) );
  AOI22D1BWP12T U2231 ( .A1(n3220), .A2(n2688), .B1(n3219), .B2(n4932), .ZN(
        n946) );
  ND2D3BWP12T U2232 ( .A1(n4743), .A2(n4742), .ZN(n4554) );
  NR3XD0BWP12T U2233 ( .A1(n949), .A2(n948), .A3(n4843), .ZN(n958) );
  OAI21D1BWP12T U2234 ( .A1(n3462), .A2(n289), .B(n3902), .ZN(n950) );
  TPAOI21D0BWP12T U2235 ( .A1(n4200), .A2(n373), .B(n950), .ZN(n956) );
  OAI22D1BWP12T U2236 ( .A1(n3321), .A2(n4655), .B1(n275), .B2(n4679), .ZN(
        n952) );
  OAI22D1BWP12T U2237 ( .A1(n3318), .A2(n4631), .B1(n3322), .B2(n3523), .ZN(
        n951) );
  NR2D1BWP12T U2238 ( .A1(n952), .A2(n951), .ZN(n3636) );
  CKND2D1BWP12T U2239 ( .A1(n3636), .A2(n3748), .ZN(n955) );
  CKND6BWP12T U2240 ( .I(n5075), .ZN(n5082) );
  AOI22D1BWP12T U2241 ( .A1(n4561), .A2(n4627), .B1(n4562), .B2(n1765), .ZN(
        n954) );
  ND3D1BWP12T U2242 ( .A1(n956), .A2(n955), .A3(n954), .ZN(n957) );
  ND2D1BWP12T U2243 ( .A1(n958), .A2(n957), .ZN(n4886) );
  AN3XD1BWP12T U2244 ( .A1(n4886), .A2(n4605), .A3(n4209), .Z(n979) );
  INR2D1BWP12T U2245 ( .A1(n4707), .B1(n5042), .ZN(n3295) );
  CKAN2D1BWP12T U2246 ( .A1(n4685), .A2(n3295), .Z(n959) );
  INR2D2BWP12T U2247 ( .A1(n959), .B1(n4891), .ZN(n4249) );
  INR2D1BWP12T U2248 ( .A1(n4910), .B1(n3321), .ZN(n3469) );
  INVD1BWP12T U2249 ( .I(n3469), .ZN(n1004) );
  ND2D1BWP12T U2250 ( .A1(n2972), .A2(n1004), .ZN(n3468) );
  TPOAI21D0BWP12T U2251 ( .A1(n1004), .A2(n4742), .B(n3957), .ZN(n960) );
  ND2D1BWP12T U2252 ( .A1(n3468), .A2(n960), .ZN(n3292) );
  CKND1BWP12T U2253 ( .I(n964), .ZN(n4124) );
  XNR2D1BWP12T U2254 ( .A1(n4124), .A2(n4912), .ZN(n4418) );
  CKND2D0BWP12T U2255 ( .A1(n4418), .A2(n5078), .ZN(n968) );
  INVD4BWP12T U2256 ( .I(n905), .ZN(n5081) );
  OAI21D1BWP12T U2257 ( .A1(n4912), .A2(n5083), .B(n5081), .ZN(n965) );
  CKND2D0BWP12T U2258 ( .A1(n4742), .A2(n965), .ZN(n966) );
  ND3D1BWP12T U2259 ( .A1(n968), .A2(n967), .A3(n966), .ZN(n969) );
  TPAOI21D0BWP12T U2260 ( .A1(n4395), .A2(n5088), .B(n969), .ZN(n970) );
  IOA21D0BWP12T U2261 ( .A1(n4488), .A2(n4103), .B(n970), .ZN(n974) );
  INVD1BWP12T U2262 ( .I(n4953), .ZN(n972) );
  INR2D1BWP12T U2263 ( .A1(n5093), .B1(n972), .ZN(n973) );
  CKND2D0BWP12T U2264 ( .A1(n4317), .A2(n5090), .ZN(n976) );
  ND3D1BWP12T U2265 ( .A1(n357), .A2(n977), .A3(n976), .ZN(n978) );
  NR2D1BWP12T U2266 ( .A1(n3318), .A2(n4636), .ZN(n981) );
  NR2D1BWP12T U2267 ( .A1(n275), .A2(n4624), .ZN(n980) );
  INVD9BWP12T U2268 ( .I(n982), .ZN(n4909) );
  OAI22D1BWP12T U2269 ( .A1(n3321), .A2(n4908), .B1(n3322), .B2(n4909), .ZN(
        n986) );
  MUX2D1BWP12T U2270 ( .I0(n4922), .I1(a[27]), .S(n5075), .Z(n1710) );
  INVD1BWP12T U2271 ( .I(n1710), .ZN(n984) );
  AN2XD1BWP12T U2272 ( .A1(n984), .A2(n983), .Z(n985) );
  TPNR2D2BWP12T U2273 ( .A1(n986), .A2(n985), .ZN(n4036) );
  CKND0BWP12T U2274 ( .I(n3969), .ZN(n2984) );
  ND2D1BWP12T U2275 ( .A1(n3694), .A2(n2984), .ZN(n4830) );
  ND2D1BWP12T U2276 ( .A1(n5075), .A2(n4924), .ZN(n988) );
  CKND2D0BWP12T U2277 ( .A1(n992), .A2(n4923), .ZN(n987) );
  OA22D1BWP12T U2278 ( .A1(n988), .A2(n4645), .B1(n987), .B2(n5075), .Z(n991)
         );
  CKND2D1BWP12T U2279 ( .A1(n3220), .A2(n4914), .ZN(n990) );
  ND2D1BWP12T U2280 ( .A1(n3217), .A2(n5051), .ZN(n989) );
  ND3D1BWP12T U2281 ( .A1(n991), .A2(n990), .A3(n989), .ZN(n4041) );
  INVD1BWP12T U2282 ( .I(n4041), .ZN(n3639) );
  ND3D1BWP12T U2283 ( .A1(n5082), .A2(n992), .A3(n4728), .ZN(n995) );
  INVD8BWP12T U2284 ( .I(n3850), .ZN(n4699) );
  AOI22D1BWP12T U2285 ( .A1(n3217), .A2(n4907), .B1(n3220), .B2(n4699), .ZN(
        n994) );
  CKND2D1BWP12T U2286 ( .A1(n3218), .A2(n4916), .ZN(n993) );
  ND3D1BWP12T U2287 ( .A1(n995), .A2(n994), .A3(n993), .ZN(n4037) );
  INVD1BWP12T U2288 ( .I(n4037), .ZN(n1009) );
  AOI22D1BWP12T U2289 ( .A1(n3639), .A2(n3051), .B1(n1009), .B2(n4742), .ZN(
        n3277) );
  INR2D1BWP12T U2290 ( .A1(n4843), .B1(n4743), .ZN(n3972) );
  INVD1BWP12T U2291 ( .I(n996), .ZN(n998) );
  CKND2D1BWP12T U2292 ( .A1(n998), .A2(n997), .ZN(n1000) );
  INVD1BWP12T U2293 ( .I(n4239), .ZN(n999) );
  XNR2D1BWP12T U2294 ( .A1(n1000), .A2(n999), .ZN(n4262) );
  INVD1BWP12T U2295 ( .I(n4262), .ZN(n1001) );
  OR2D2BWP12T U2296 ( .A1(n1001), .A2(n4260), .Z(n1003) );
  INR2D8BWP12T U2297 ( .A1(n848), .B1(n4573), .ZN(n5100) );
  ND2D1BWP12T U2298 ( .A1(n5100), .A2(n5099), .ZN(n1002) );
  ND2D1BWP12T U2299 ( .A1(n1003), .A2(n1002), .ZN(n1007) );
  TPNR2D0BWP12T U2300 ( .A1(n3436), .A2(n1004), .ZN(n1005) );
  OAI21D1BWP12T U2301 ( .A1(n3107), .A2(n1005), .B(n3468), .ZN(n1816) );
  INVD1BWP12T U2302 ( .I(n4886), .ZN(n4832) );
  NR2D1BWP12T U2303 ( .A1(n3639), .A2(n4742), .ZN(n1011) );
  NR2D1BWP12T U2304 ( .A1(n1009), .A2(n3051), .ZN(n1010) );
  NR3D1BWP12T U2305 ( .A1(n1011), .A2(n4743), .A3(n1010), .ZN(n1818) );
  NR2D1BWP12T U2306 ( .A1(n4036), .A2(n4206), .ZN(n1012) );
  NR2D1BWP12T U2307 ( .A1(n1818), .A2(n1012), .ZN(n1015) );
  INVD1BWP12T U2308 ( .I(n3456), .ZN(n1013) );
  INVD1BWP12T U2309 ( .I(n4554), .ZN(n3766) );
  CKND2D1BWP12T U2310 ( .A1(n1013), .A2(n3766), .ZN(n1014) );
  ND2D1BWP12T U2311 ( .A1(n1015), .A2(n1014), .ZN(n1846) );
  OAI21D1BWP12T U2312 ( .A1(n1846), .A2(n4891), .B(n4890), .ZN(n4885) );
  IND3D1BWP12T U2313 ( .A1(n4832), .B1(n5099), .B2(n4885), .ZN(n1018) );
  CKND2D1BWP12T U2314 ( .A1(n4886), .A2(n4209), .ZN(n1016) );
  INR2D1BWP12T U2315 ( .A1(n4573), .B1(n4544), .ZN(n4549) );
  IND2XD1BWP12T U2316 ( .A1(n1016), .B1(n4549), .ZN(n1017) );
  TPOAI21D1BWP12T U2317 ( .A1(n1023), .A2(n1022), .B(n1021), .ZN(n1030) );
  TPAOI21D2BWP12T U2318 ( .A1(n1030), .A2(n1029), .B(n1028), .ZN(n3084) );
  TPOAI22D2BWP12T U2319 ( .A1(n1031), .A2(n2667), .B1(n1119), .B2(n2669), .ZN(
        n1102) );
  TPOAI22D2BWP12T U2320 ( .A1(n1108), .A2(n2647), .B1(n2648), .B2(n1032), .ZN(
        n1103) );
  XNR2XD2BWP12T U2321 ( .A1(n2167), .A2(n2701), .ZN(n1094) );
  OAI22D1BWP12T U2322 ( .A1(n1094), .A2(n2319), .B1(n1033), .B2(n2702), .ZN(
        n1104) );
  INVD1BWP12T U2323 ( .I(n1104), .ZN(n1034) );
  XOR3XD4BWP12T U2324 ( .A1(n1102), .A2(n1103), .A3(n1034), .Z(n1130) );
  INVD1BWP12T U2325 ( .I(n1130), .ZN(n1047) );
  NR2D1BWP12T U2326 ( .A1(n1036), .A2(n1035), .ZN(n1038) );
  ND2D1BWP12T U2327 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  TPOAI21D2BWP12T U2328 ( .A1(n1039), .A2(n1038), .B(n1037), .ZN(n1129) );
  OR2XD1BWP12T U2329 ( .A1(n1043), .A2(n1042), .Z(n1041) );
  ND2D1BWP12T U2330 ( .A1(n1041), .A2(n1040), .ZN(n1045) );
  ND2D1BWP12T U2331 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  OAI21D1BWP12T U2332 ( .A1(n1129), .A2(n1047), .B(n1128), .ZN(n1046) );
  TPND2D2BWP12T U2333 ( .A1(n1051), .A2(n1050), .ZN(n1056) );
  ND2D3BWP12T U2334 ( .A1(n1056), .A2(n1055), .ZN(n1083) );
  CKND3BWP12T U2335 ( .I(a[16]), .ZN(n1057) );
  XNR2XD8BWP12T U2336 ( .A1(n1058), .A2(n1057), .ZN(n1421) );
  INVD1BWP12T U2337 ( .I(n1421), .ZN(n1059) );
  INVD1BWP12T U2338 ( .I(n1086), .ZN(n1063) );
  TPOAI22D2BWP12T U2339 ( .A1(n2263), .A2(n1061), .B1(n2739), .B2(n1093), .ZN(
        n1087) );
  INVD1BWP12T U2340 ( .I(n1087), .ZN(n1062) );
  XOR3D2BWP12T U2341 ( .A1(n1063), .A2(n1085), .A3(n1062), .Z(n1079) );
  XNR2XD4BWP12T U2342 ( .A1(n2623), .A2(n2746), .ZN(n1107) );
  OAI22D1BWP12T U2343 ( .A1(n1107), .A2(n2747), .B1(n1064), .B2(n2748), .ZN(
        n1098) );
  TPNR2D1BWP12T U2344 ( .A1(n1066), .A2(n1065), .ZN(n1096) );
  OAI22D1BWP12T U2345 ( .A1(n1067), .A2(n2744), .B1(n1113), .B2(n2743), .ZN(
        n1097) );
  XOR3D2BWP12T U2346 ( .A1(n1098), .A2(n1096), .A3(n1068), .Z(n1133) );
  ND2D3BWP12T U2347 ( .A1(n1131), .A2(n1076), .ZN(n1078) );
  INVD2BWP12T U2348 ( .I(n1069), .ZN(n1071) );
  TPND2D3BWP12T U2349 ( .A1(n1071), .A2(n1070), .ZN(n1075) );
  ND2D3BWP12T U2350 ( .A1(n1073), .A2(n1072), .ZN(n1074) );
  TPOAI21D2BWP12T U2351 ( .A1(n1131), .A2(n1076), .B(n1132), .ZN(n1077) );
  ND2D3BWP12T U2352 ( .A1(n1078), .A2(n1077), .ZN(n1274) );
  IOA21D2BWP12T U2353 ( .A1(n1081), .A2(n1080), .B(n1079), .ZN(n1082) );
  IOA21D2BWP12T U2354 ( .A1(n1084), .A2(n1083), .B(n1082), .ZN(n1255) );
  ND2D1BWP12T U2355 ( .A1(n1087), .A2(n1086), .ZN(n1089) );
  TPND2D2BWP12T U2356 ( .A1(n1089), .A2(n1088), .ZN(n1201) );
  INVD1BWP12T U2357 ( .I(a[16]), .ZN(n1090) );
  XNR2XD4BWP12T U2358 ( .A1(n1090), .A2(a[17]), .ZN(n1091) );
  ND2D8BWP12T U2359 ( .A1(n1421), .A2(n1091), .ZN(n2689) );
  TPOAI22D2BWP12T U2360 ( .A1(n1092), .A2(n2691), .B1(n2689), .B2(n1810), .ZN(
        n1191) );
  XNR2XD4BWP12T U2361 ( .A1(n2098), .A2(n2701), .ZN(n1176) );
  TPOAI22D2BWP12T U2362 ( .A1(n1176), .A2(n2319), .B1(n1094), .B2(n2702), .ZN(
        n1189) );
  INVD2BWP12T U2363 ( .I(n1189), .ZN(n1095) );
  XOR3XD4BWP12T U2364 ( .A1(n1191), .A2(n1190), .A3(n1095), .Z(n1202) );
  INVD1BWP12T U2365 ( .I(n1096), .ZN(n1100) );
  ND2D1BWP12T U2366 ( .A1(n1098), .A2(n1097), .ZN(n1099) );
  TPOAI21D2BWP12T U2367 ( .A1(n1101), .A2(n1100), .B(n1099), .ZN(n1204) );
  XNR3XD4BWP12T U2368 ( .A1(n1201), .A2(n1202), .A3(n1204), .ZN(n1256) );
  OAI21D1BWP12T U2369 ( .A1(n1104), .A2(n1103), .B(n1102), .ZN(n1106) );
  ND2D1BWP12T U2370 ( .A1(n1104), .A2(n1103), .ZN(n1105) );
  XNR2XD4BWP12T U2371 ( .A1(n4753), .A2(n2746), .ZN(n1150) );
  TPOAI22D4BWP12T U2372 ( .A1(n1107), .A2(n2748), .B1(n1150), .B2(n2747), .ZN(
        n1171) );
  XNR2XD4BWP12T U2373 ( .A1(n2575), .A2(n288), .ZN(n1151) );
  XNR2XD4BWP12T U2374 ( .A1(n279), .A2(n2593), .ZN(n1187) );
  INVD1P75BWP12T U2375 ( .I(n1170), .ZN(n1110) );
  XNR3XD4BWP12T U2376 ( .A1(n1171), .A2(n1172), .A3(n1110), .ZN(n1196) );
  XNR2XD4BWP12T U2377 ( .A1(n1932), .A2(n2688), .ZN(n1175) );
  IND2D2BWP12T U2378 ( .A1(n1175), .B1(n1059), .ZN(n1111) );
  OAI21D1BWP12T U2379 ( .A1(n2689), .A2(n1112), .B(n1111), .ZN(n1219) );
  OR2XD4BWP12T U2380 ( .A1(n2744), .A2(n1113), .Z(n1117) );
  XNR2D1BWP12T U2381 ( .A1(n2551), .A2(n2742), .ZN(n1185) );
  INR2D1BWP12T U2382 ( .A1(n1114), .B1(n1185), .ZN(n1115) );
  INVD1BWP12T U2383 ( .I(n1115), .ZN(n1116) );
  TPND2D3BWP12T U2384 ( .A1(n1117), .A2(n1116), .ZN(n1220) );
  XNR2D1BWP12T U2385 ( .A1(n4628), .A2(n2679), .ZN(n1160) );
  OAI22D2BWP12T U2386 ( .A1(n1118), .A2(n2680), .B1(n2682), .B2(n1160), .ZN(
        n1155) );
  XNR2XD2BWP12T U2387 ( .A1(n2555), .A2(n2666), .ZN(n1161) );
  TPOAI22D2BWP12T U2388 ( .A1(n1119), .A2(n2667), .B1(n1161), .B2(n2669), .ZN(
        n1154) );
  XOR3D2BWP12T U2389 ( .A1(n1219), .A2(n1220), .A3(n1218), .Z(n1194) );
  XOR3XD4BWP12T U2390 ( .A1(n1195), .A2(n1196), .A3(n1194), .Z(n1253) );
  XOR3XD4BWP12T U2391 ( .A1(n1255), .A2(n1256), .A3(n1253), .Z(n1270) );
  CKND2D2BWP12T U2392 ( .A1(n1121), .A2(n1120), .ZN(n1123) );
  ND2D3BWP12T U2393 ( .A1(n1123), .A2(n1122), .ZN(n1127) );
  ND2D1BWP12T U2394 ( .A1(n1125), .A2(n1124), .ZN(n1126) );
  TPND2D2BWP12T U2395 ( .A1(n1127), .A2(n1126), .ZN(n1137) );
  XNR3XD4BWP12T U2396 ( .A1(n1130), .A2(n1129), .A3(n1128), .ZN(n1138) );
  NR2D1BWP12T U2397 ( .A1(n1137), .A2(n1138), .ZN(n1135) );
  XOR3XD4BWP12T U2398 ( .A1(n1133), .A2(n1132), .A3(n1131), .Z(n1136) );
  ND2D1BWP12T U2399 ( .A1(n1137), .A2(n1138), .ZN(n1134) );
  OA21XD2BWP12T U2400 ( .A1(n1135), .A2(n1136), .B(n1134), .Z(n1148) );
  TPND2D3BWP12T U2401 ( .A1(n1149), .A2(n1148), .ZN(n3085) );
  XNR3XD4BWP12T U2402 ( .A1(n1138), .A2(n1137), .A3(n1136), .ZN(n1147) );
  NR2D1BWP12T U2403 ( .A1(n1140), .A2(n1139), .ZN(n1143) );
  INVD1BWP12T U2404 ( .I(n1139), .ZN(n1142) );
  CKND0BWP12T U2405 ( .I(n1140), .ZN(n1141) );
  OAI22D1BWP12T U2406 ( .A1(n1144), .A2(n1143), .B1(n1142), .B2(n1141), .ZN(
        n1145) );
  INR2D4BWP12T U2407 ( .A1(n1147), .B1(n1146), .ZN(n4144) );
  NR2D2BWP12T U2408 ( .A1(n1149), .A2(n1148), .ZN(n3086) );
  TPAOI21D2BWP12T U2409 ( .A1(n3085), .A2(n4144), .B(n3086), .ZN(n2436) );
  TPOAI21D1BWP12T U2410 ( .A1(n3084), .A2(n2437), .B(n2436), .ZN(n1795) );
  INVD1BWP12T U2411 ( .I(n1229), .ZN(n1156) );
  HA1D2BWP12T U2412 ( .A(n1155), .B(n1154), .CO(n1227), .S(n1218) );
  IND2XD1BWP12T U2413 ( .A1(n1228), .B1(n1229), .ZN(n1157) );
  DCCKBD4BWP12T U2414 ( .I(n2701), .Z(n1347) );
  XNR2XD4BWP12T U2415 ( .A1(n2575), .A2(n1347), .ZN(n1351) );
  XNR2D1BWP12T U2416 ( .A1(n280), .A2(n2742), .ZN(n1282) );
  OAI22D2BWP12T U2417 ( .A1(n2648), .A2(n1159), .B1(n1352), .B2(n2647), .ZN(
        n1296) );
  XOR3D2BWP12T U2418 ( .A1(n1295), .A2(n1293), .A3(n1296), .Z(n1325) );
  XNR2D2BWP12T U2419 ( .A1(n2226), .A2(n2593), .ZN(n1188) );
  XNR2D2BWP12T U2420 ( .A1(n2172), .A2(n4926), .ZN(n1166) );
  TPOAI22D2BWP12T U2421 ( .A1(n1160), .A2(n2680), .B1(n1166), .B2(n2682), .ZN(
        n1225) );
  XOR2XD8BWP12T U2422 ( .A1(n1810), .A2(n4923), .Z(n2220) );
  BUFFXD12BWP12T U2423 ( .I(n2220), .Z(n2620) );
  NR2XD2BWP12T U2424 ( .A1(n2620), .A2(n5082), .ZN(n1226) );
  ND2D1BWP12T U2425 ( .A1(n1225), .A2(n1226), .ZN(n1163) );
  XNR2XD4BWP12T U2426 ( .A1(n2071), .A2(n2666), .ZN(n1241) );
  TPOAI22D2BWP12T U2427 ( .A1(n1161), .A2(n2667), .B1(n1241), .B2(n2669), .ZN(
        n1224) );
  INVD1BWP12T U2428 ( .I(n1164), .ZN(n1165) );
  XNR2XD4BWP12T U2429 ( .A1(n2094), .A2(n1165), .ZN(n1304) );
  TPOAI22D2BWP12T U2430 ( .A1(n1304), .A2(n2682), .B1(n1166), .B2(n2680), .ZN(
        n1290) );
  IND2XD1BWP12T U2431 ( .A1(n1512), .B1(n4924), .ZN(n1169) );
  INVD2BWP12T U2432 ( .I(n4923), .ZN(n1167) );
  XNR2XD4BWP12T U2433 ( .A1(n1167), .A2(n4924), .ZN(n1168) );
  ND2XD16BWP12T U2434 ( .A1(n1168), .A2(n2220), .ZN(n2218) );
  TPOAI22D2BWP12T U2435 ( .A1(n1169), .A2(n2220), .B1(n2218), .B2(n1342), .ZN(
        n1289) );
  XNR2D1BWP12T U2436 ( .A1(n2098), .A2(n5014), .ZN(n1306) );
  TPOAI22D2BWP12T U2437 ( .A1(n1306), .A2(n2739), .B1(n2263), .B2(n1180), .ZN(
        n1287) );
  XOR3XD4BWP12T U2438 ( .A1(n1290), .A2(n1289), .A3(n1287), .Z(n1380) );
  XOR3D2BWP12T U2439 ( .A1(n1378), .A2(n1379), .A3(n1380), .Z(n1323) );
  XOR3D2BWP12T U2440 ( .A1(n1324), .A2(n1325), .A3(n1323), .Z(n1412) );
  OAI21D1BWP12T U2441 ( .A1(n1172), .A2(n1171), .B(n1170), .ZN(n1174) );
  TPOAI22D1BWP12T U2442 ( .A1(n1242), .A2(n2691), .B1(n1175), .B2(n2689), .ZN(
        n1235) );
  TPNR2D2BWP12T U2443 ( .A1(n1177), .A2(n2319), .ZN(n1178) );
  TPNR2D2BWP12T U2444 ( .A1(n1179), .A2(n1178), .ZN(n1232) );
  NR2D3BWP12T U2445 ( .A1(n1180), .A2(n2739), .ZN(n1183) );
  NR2D1BWP12T U2446 ( .A1(n1181), .A2(n2263), .ZN(n1182) );
  NR2D2BWP12T U2447 ( .A1(n1183), .A2(n1182), .ZN(n1236) );
  INVD1BWP12T U2448 ( .I(n1236), .ZN(n1184) );
  XOR3XD4BWP12T U2449 ( .A1(n1235), .A2(n1232), .A3(n1184), .Z(n1213) );
  TPOAI22D1BWP12T U2450 ( .A1(n1186), .A2(n2743), .B1(n2744), .B2(n1185), .ZN(
        n1248) );
  OAI21D0BWP12T U2451 ( .A1(n1191), .A2(n1190), .B(n1189), .ZN(n1193) );
  CKND2D0BWP12T U2452 ( .A1(n1191), .A2(n1190), .ZN(n1192) );
  ND2D1BWP12T U2453 ( .A1(n1196), .A2(n1195), .ZN(n1197) );
  TPOAI21D2BWP12T U2454 ( .A1(n1199), .A2(n1198), .B(n1197), .ZN(n1261) );
  INVD1BWP12T U2455 ( .I(n1202), .ZN(n1200) );
  ND2D1BWP12T U2456 ( .A1(n1200), .A2(n1201), .ZN(n1207) );
  INVD1BWP12T U2457 ( .I(n1201), .ZN(n1203) );
  ND2D1BWP12T U2458 ( .A1(n1203), .A2(n1202), .ZN(n1205) );
  ND2D1BWP12T U2459 ( .A1(n1205), .A2(n1204), .ZN(n1206) );
  TPNR2D1BWP12T U2460 ( .A1(n1261), .A2(n1262), .ZN(n1210) );
  INVD1BWP12T U2461 ( .I(n1261), .ZN(n1209) );
  INVD1BWP12T U2462 ( .I(n1262), .ZN(n1208) );
  TPOAI22D2BWP12T U2463 ( .A1(n1260), .A2(n1210), .B1(n1209), .B2(n1208), .ZN(
        n1413) );
  INVD1BWP12T U2464 ( .I(n1214), .ZN(n1212) );
  IOA21D2BWP12T U2465 ( .A1(n1212), .A2(n1213), .B(n1211), .ZN(n1217) );
  ND2D1BWP12T U2466 ( .A1(n1215), .A2(n1214), .ZN(n1216) );
  TPND2D2BWP12T U2467 ( .A1(n1217), .A2(n1216), .ZN(n1396) );
  INVD1BWP12T U2468 ( .I(n1218), .ZN(n1223) );
  TPNR2D1BWP12T U2469 ( .A1(n1220), .A2(n1219), .ZN(n1222) );
  ND2D1BWP12T U2470 ( .A1(n1220), .A2(n1219), .ZN(n1221) );
  TPOAI21D2BWP12T U2471 ( .A1(n1223), .A2(n1222), .B(n1221), .ZN(n1249) );
  XOR3XD4BWP12T U2472 ( .A1(n1226), .A2(n1225), .A3(n1224), .Z(n1252) );
  ND2D1BWP12T U2473 ( .A1(n1249), .A2(n1252), .ZN(n1231) );
  XNR3XD4BWP12T U2474 ( .A1(n1229), .A2(n1228), .A3(n1227), .ZN(n1251) );
  OAI21D2BWP12T U2475 ( .A1(n1249), .A2(n1252), .B(n1251), .ZN(n1230) );
  ND2D2BWP12T U2476 ( .A1(n1231), .A2(n1230), .ZN(n1397) );
  INVD1BWP12T U2477 ( .I(n1235), .ZN(n1234) );
  XNR2D1BWP12T U2478 ( .A1(n2551), .A2(n2746), .ZN(n1281) );
  TPOAI22D2BWP12T U2479 ( .A1(n1239), .A2(n2748), .B1(n1281), .B2(n2747), .ZN(
        n1303) );
  XNR2XD2BWP12T U2480 ( .A1(n1932), .A2(n4924), .ZN(n1305) );
  TPOAI22D1BWP12T U2481 ( .A1(n1240), .A2(n2218), .B1(n1305), .B2(n2220), .ZN(
        n1302) );
  XNR2XD4BWP12T U2482 ( .A1(n4628), .A2(n2666), .ZN(n1284) );
  TPOAI22D2BWP12T U2483 ( .A1(n1241), .A2(n2667), .B1(n1284), .B2(n2669), .ZN(
        n1356) );
  XNR2XD4BWP12T U2484 ( .A1(n2555), .A2(n2688), .ZN(n1285) );
  TPOAI22D2BWP12T U2485 ( .A1(n1285), .A2(n2691), .B1(n1242), .B2(n2689), .ZN(
        n1355) );
  INVD1BWP12T U2486 ( .I(n1247), .ZN(n1245) );
  INVD1BWP12T U2487 ( .I(n1248), .ZN(n1244) );
  IOA21D1BWP12T U2488 ( .A1(n1245), .A2(n1244), .B(n1243), .ZN(n1246) );
  IOA21D1BWP12T U2489 ( .A1(n1248), .A2(n1247), .B(n1246), .ZN(n1319) );
  XOR3XD4BWP12T U2490 ( .A1(n1322), .A2(n1321), .A3(n1319), .Z(n1398) );
  XOR3XD4BWP12T U2491 ( .A1(n1396), .A2(n1397), .A3(n1398), .Z(n1410) );
  XOR3XD4BWP12T U2492 ( .A1(n1412), .A2(n1413), .A3(n1410), .Z(n1279) );
  XNR3XD4BWP12T U2493 ( .A1(n1252), .A2(n1251), .A3(n1250), .ZN(n1264) );
  TPND2D2BWP12T U2494 ( .A1(n1254), .A2(n1253), .ZN(n1258) );
  ND2D1BWP12T U2495 ( .A1(n1256), .A2(n1255), .ZN(n1257) );
  TPND2D2BWP12T U2496 ( .A1(n1258), .A2(n1257), .ZN(n1268) );
  INR2D2BWP12T U2497 ( .A1(n1269), .B1(n1268), .ZN(n1259) );
  INVD1BWP12T U2498 ( .I(n1259), .ZN(n1263) );
  XNR3XD4BWP12T U2499 ( .A1(n1262), .A2(n1261), .A3(n1260), .ZN(n1267) );
  ND2D1BWP12T U2500 ( .A1(n1263), .A2(n1267), .ZN(n1266) );
  ND2D1BWP12T U2501 ( .A1(n1268), .A2(n1264), .ZN(n1265) );
  TPND2D1BWP12T U2502 ( .A1(n1266), .A2(n1265), .ZN(n1278) );
  XNR3XD4BWP12T U2503 ( .A1(n1269), .A2(n1268), .A3(n1267), .ZN(n1277) );
  INVD1BWP12T U2504 ( .I(n1274), .ZN(n1272) );
  IOA21D1BWP12T U2505 ( .A1(n1272), .A2(n1271), .B(n1270), .ZN(n1273) );
  ND2D2BWP12T U2506 ( .A1(n1277), .A2(n1276), .ZN(n3730) );
  AO21D1BWP12T U2507 ( .A1(n1795), .A2(n2439), .B(n2438), .Z(n3866) );
  XNR2XD8BWP12T U2508 ( .A1(n4761), .A2(n2746), .ZN(n1349) );
  TPOAI22D1BWP12T U2509 ( .A1(n1349), .A2(n2747), .B1(n1281), .B2(n2748), .ZN(
        n1309) );
  XNR2D1BWP12T U2510 ( .A1(n2226), .A2(n2742), .ZN(n1368) );
  OAI22D1BWP12T U2511 ( .A1(n1282), .A2(n2744), .B1(n1368), .B2(n2743), .ZN(
        n1308) );
  CKND3BWP12T U2512 ( .I(n1478), .ZN(n1474) );
  XNR2XD4BWP12T U2513 ( .A1(n4924), .A2(n5051), .ZN(n2624) );
  XNR2XD4BWP12T U2514 ( .A1(n341), .A2(n2666), .ZN(n1339) );
  TPOAI22D4BWP12T U2515 ( .A1(n1284), .A2(n2667), .B1(n1339), .B2(n2669), .ZN(
        n1371) );
  XNR2XD8BWP12T U2516 ( .A1(n2071), .A2(n2688), .ZN(n1365) );
  TPOAI22D2BWP12T U2517 ( .A1(n1285), .A2(n2689), .B1(n1365), .B2(n2691), .ZN(
        n1370) );
  XOR3XD4BWP12T U2518 ( .A1(n1373), .A2(n1371), .A3(n1370), .Z(n1388) );
  TPNR2D1BWP12T U2519 ( .A1(n1290), .A2(n1289), .ZN(n1286) );
  INVD1BWP12T U2520 ( .I(n1286), .ZN(n1288) );
  TPND2D2BWP12T U2521 ( .A1(n1288), .A2(n1287), .ZN(n1292) );
  ND2D1BWP12T U2522 ( .A1(n1290), .A2(n1289), .ZN(n1291) );
  TPND2D2BWP12T U2523 ( .A1(n1292), .A2(n1291), .ZN(n1387) );
  INVD1BWP12T U2524 ( .I(n1293), .ZN(n1385) );
  TPNR2D1BWP12T U2525 ( .A1(n1385), .A2(n1384), .ZN(n1294) );
  TPOAI21D1BWP12T U2526 ( .A1(n1388), .A2(n1387), .B(n1294), .ZN(n1300) );
  TPND2D1BWP12T U2527 ( .A1(n1296), .A2(n1295), .ZN(n1383) );
  INVD1BWP12T U2528 ( .I(n1383), .ZN(n1297) );
  TPOAI21D1BWP12T U2529 ( .A1(n1297), .A2(n1388), .B(n1387), .ZN(n1299) );
  ND2D1BWP12T U2530 ( .A1(n1388), .A2(n1297), .ZN(n1298) );
  ND3XD3BWP12T U2531 ( .A1(n1300), .A2(n1299), .A3(n1298), .ZN(n1479) );
  FA1D2BWP12T U2532 ( .A(n1303), .B(n1302), .CI(n1301), .CO(n1315), .S(n1321)
         );
  XNR2D2BWP12T U2533 ( .A1(n2072), .A2(n4924), .ZN(n1366) );
  TPOAI22D2BWP12T U2534 ( .A1(n1305), .A2(n2218), .B1(n1366), .B2(n2620), .ZN(
        n1335) );
  TPOAI22D1BWP12T U2535 ( .A1(n1348), .A2(n296), .B1(n1306), .B2(n2263), .ZN(
        n1333) );
  XOR3XD4BWP12T U2536 ( .A1(n1334), .A2(n1335), .A3(n1333), .Z(n1316) );
  FA1D2BWP12T U2537 ( .A(n1309), .B(n1310), .CI(n1308), .CO(n1478), .S(n1314)
         );
  TPOAI21D1BWP12T U2538 ( .A1(n1315), .A2(n1311), .B(n1314), .ZN(n1313) );
  TPND2D1BWP12T U2539 ( .A1(n1311), .A2(n1315), .ZN(n1312) );
  TPND2D2BWP12T U2540 ( .A1(n1313), .A2(n1312), .ZN(n1477) );
  XOR3XD4BWP12T U2541 ( .A1(n1474), .A2(n1479), .A3(n1477), .Z(n1484) );
  XOR3D2BWP12T U2542 ( .A1(n1316), .A2(n1315), .A3(n1314), .Z(n1394) );
  INVD1BWP12T U2543 ( .I(n1322), .ZN(n1317) );
  TPND2D1BWP12T U2544 ( .A1(n1318), .A2(n1317), .ZN(n1320) );
  TPND2D2BWP12T U2545 ( .A1(n1320), .A2(n1319), .ZN(n1330) );
  ND2D1BWP12T U2546 ( .A1(n1322), .A2(n1321), .ZN(n1329) );
  INVD1BWP12T U2547 ( .I(n1323), .ZN(n1328) );
  NR2D2BWP12T U2548 ( .A1(n1325), .A2(n1324), .ZN(n1327) );
  ND2D1BWP12T U2549 ( .A1(n1325), .A2(n1324), .ZN(n1326) );
  TPOAI21D1BWP12T U2550 ( .A1(n1328), .A2(n1327), .B(n1326), .ZN(n1392) );
  TPOAI21D1BWP12T U2551 ( .A1(n1394), .A2(n1395), .B(n1392), .ZN(n1332) );
  TPND2D2BWP12T U2552 ( .A1(n1332), .A2(n1331), .ZN(n1485) );
  INVD1BWP12T U2553 ( .I(n1333), .ZN(n1338) );
  NR2D1BWP12T U2554 ( .A1(n1335), .A2(n312), .ZN(n1337) );
  ND2XD0BWP12T U2555 ( .A1(n1335), .A2(n312), .ZN(n1336) );
  XNR2XD4BWP12T U2556 ( .A1(n2094), .A2(n2666), .ZN(n1438) );
  TPOAI22D2BWP12T U2557 ( .A1(n1438), .A2(n2669), .B1(n1339), .B2(n2667), .ZN(
        n1416) );
  XNR2XD4BWP12T U2558 ( .A1(n2098), .A2(n2679), .ZN(n1439) );
  CKND4BWP12T U2559 ( .I(n5051), .ZN(n1341) );
  CKND2D2BWP12T U2560 ( .A1(n4914), .A2(n1341), .ZN(n1343) );
  INVD1P75BWP12T U2561 ( .I(n5051), .ZN(n1658) );
  TPOAI21D2BWP12T U2562 ( .A1(n4914), .A2(n1658), .B(n4924), .ZN(n1344) );
  TPOAI22D2BWP12T U2563 ( .A1(n1346), .A2(n2624), .B1(n2625), .B2(n4625), .ZN(
        n1417) );
  XOR3XD4BWP12T U2564 ( .A1(n1416), .A2(n1415), .A3(n1417), .Z(n1426) );
  XNR2XD4BWP12T U2565 ( .A1(n4753), .A2(n2701), .ZN(n1464) );
  XNR2XD8BWP12T U2566 ( .A1(n2623), .A2(n1347), .ZN(n1350) );
  XNR2D1BWP12T U2567 ( .A1(n279), .A2(n2746), .ZN(n1443) );
  XOR3XD4BWP12T U2568 ( .A1(n1459), .A2(n1460), .A3(n1458), .Z(n1427) );
  XOR3XD4BWP12T U2569 ( .A1(n1425), .A2(n1426), .A3(n1427), .Z(n1449) );
  TPOAI22D2BWP12T U2570 ( .A1(n2702), .A2(n1351), .B1(n1350), .B2(n2319), .ZN(
        n1376) );
  ND2D1BWP12T U2571 ( .A1(n1357), .A2(n1375), .ZN(n1359) );
  ND2D1BWP12T U2572 ( .A1(n1376), .A2(n1377), .ZN(n1358) );
  TPND2D2BWP12T U2573 ( .A1(n1359), .A2(n1358), .ZN(n1454) );
  XNR2D2BWP12T U2574 ( .A1(n2551), .A2(n288), .ZN(n1441) );
  TPOAI22D4BWP12T U2575 ( .A1(n1360), .A2(n2648), .B1(n1441), .B2(n2647), .ZN(
        n1433) );
  XNR2XD4BWP12T U2576 ( .A1(n1932), .A2(n4914), .ZN(n1437) );
  OR2D2BWP12T U2577 ( .A1(n1437), .A2(n2624), .Z(n1364) );
  XNR2XD4BWP12T U2578 ( .A1(n4316), .A2(n4914), .ZN(n1361) );
  INVD1P75BWP12T U2579 ( .I(n1362), .ZN(n1363) );
  TPND2D3BWP12T U2580 ( .A1(n1364), .A2(n1363), .ZN(n1434) );
  XNR2XD4BWP12T U2581 ( .A1(n4628), .A2(n2688), .ZN(n1420) );
  TPOAI22D2BWP12T U2582 ( .A1(n1365), .A2(n2689), .B1(n1420), .B2(n2691), .ZN(
        n1466) );
  XNR2XD4BWP12T U2583 ( .A1(b[3]), .A2(n4924), .ZN(n1422) );
  TPOAI22D2BWP12T U2584 ( .A1(n1366), .A2(n2218), .B1(n2620), .B2(n1422), .ZN(
        n1465) );
  XOR3XD4BWP12T U2585 ( .A1(n1433), .A2(n1434), .A3(n1432), .Z(n1455) );
  TPOAI22D1BWP12T U2586 ( .A1(n1367), .A2(n2646), .B1(n1440), .B2(n4257), .ZN(
        n1470) );
  XNR2XD8BWP12T U2587 ( .A1(n4764), .A2(n2742), .ZN(n1414) );
  INVD1BWP12T U2588 ( .I(n1371), .ZN(n1369) );
  INVD1BWP12T U2589 ( .I(n1369), .ZN(n1374) );
  OAI21D0BWP12T U2590 ( .A1(n1373), .A2(n1371), .B(n1370), .ZN(n1372) );
  XOR3XD4BWP12T U2591 ( .A1(n1470), .A2(n1471), .A3(n1469), .Z(n1453) );
  XNR3XD4BWP12T U2592 ( .A1(n1454), .A2(n1455), .A3(n1453), .ZN(n1448) );
  XOR3D2BWP12T U2593 ( .A1(n1377), .A2(n1376), .A3(n1375), .Z(n1403) );
  OAI21D1BWP12T U2594 ( .A1(n1385), .A2(n1384), .B(n1383), .ZN(n1386) );
  XOR3XD4BWP12T U2595 ( .A1(n1388), .A2(n1387), .A3(n1386), .Z(n1401) );
  ND2D1BWP12T U2596 ( .A1(n1402), .A2(n1403), .ZN(n1389) );
  CKND3BWP12T U2597 ( .I(n1446), .ZN(n1391) );
  XOR3XD4BWP12T U2598 ( .A1(n1449), .A2(n1448), .A3(n1391), .Z(n1483) );
  XNR3XD4BWP12T U2599 ( .A1(n1484), .A2(n1485), .A3(n1483), .ZN(n1493) );
  XNR3XD4BWP12T U2600 ( .A1(n1395), .A2(n1394), .A3(n1393), .ZN(n1407) );
  INVD2BWP12T U2601 ( .I(n1407), .ZN(n1406) );
  ND2D1BWP12T U2602 ( .A1(n1398), .A2(n1397), .ZN(n1400) );
  TPOAI21D1BWP12T U2603 ( .A1(n1398), .A2(n1397), .B(n1396), .ZN(n1399) );
  TPND2D2BWP12T U2604 ( .A1(n1399), .A2(n1400), .ZN(n1408) );
  XOR3D2BWP12T U2605 ( .A1(n1403), .A2(n1402), .A3(n1401), .Z(n1409) );
  NR2D2BWP12T U2606 ( .A1(n1408), .A2(n1409), .ZN(n1405) );
  ND2D1BWP12T U2607 ( .A1(n1408), .A2(n1409), .ZN(n1404) );
  TPNR2D3BWP12T U2608 ( .A1(n1493), .A2(n1492), .ZN(n3022) );
  XOR3XD4BWP12T U2609 ( .A1(n1409), .A2(n1408), .A3(n1407), .Z(n1491) );
  OAI21D1BWP12T U2610 ( .A1(n1413), .A2(n1412), .B(n1410), .ZN(n1411) );
  INVD1BWP12T U2611 ( .I(n3865), .ZN(n1489) );
  TPOAI22D2BWP12T U2612 ( .A1(n1414), .A2(n2744), .B1(n1550), .B2(n2743), .ZN(
        n1563) );
  INVD1P75BWP12T U2613 ( .I(n1563), .ZN(n1423) );
  OAI21D1BWP12T U2614 ( .A1(n1416), .A2(n1417), .B(n1415), .ZN(n1419) );
  ND2D1BWP12T U2615 ( .A1(n1417), .A2(n1416), .ZN(n1418) );
  CKND4BWP12T U2616 ( .I(n4316), .ZN(n1868) );
  TPNR2D1BWP12T U2617 ( .A1(n1868), .A2(n2643), .ZN(n1508) );
  XNR2XD4BWP12T U2618 ( .A1(n2172), .A2(n2688), .ZN(n1516) );
  TPOAI22D2BWP12T U2619 ( .A1(n1516), .A2(n1421), .B1(n1420), .B2(n2689), .ZN(
        n1509) );
  BUFFXD8BWP12T U2620 ( .I(n2218), .Z(n2621) );
  TPOAI22D2BWP12T U2621 ( .A1(n2621), .A2(n1422), .B1(n1548), .B2(n2620), .ZN(
        n1506) );
  XOR3XD4BWP12T U2622 ( .A1(n1508), .A2(n1509), .A3(n1506), .Z(n1562) );
  XOR3XD4BWP12T U2623 ( .A1(n1423), .A2(n1564), .A3(n1562), .Z(n1571) );
  TPNR2D2BWP12T U2624 ( .A1(n1426), .A2(n337), .ZN(n1424) );
  CKND3BWP12T U2625 ( .I(n1424), .ZN(n1428) );
  RCAOI21D4BWP12T U2626 ( .A1(n1428), .A2(n1427), .B(n354), .ZN(n1570) );
  INVD2BWP12T U2627 ( .I(n1433), .ZN(n1429) );
  TPND2D2BWP12T U2628 ( .A1(n1430), .A2(n1429), .ZN(n1431) );
  TPND2D2BWP12T U2629 ( .A1(n1432), .A2(n1431), .ZN(n1436) );
  ND2D1BWP12T U2630 ( .A1(n1434), .A2(n1433), .ZN(n1435) );
  XNR2D2BWP12T U2631 ( .A1(n2072), .A2(n4914), .ZN(n1549) );
  TPOAI22D2BWP12T U2632 ( .A1(n1549), .A2(n2624), .B1(n1437), .B2(n2625), .ZN(
        n1542) );
  TPOAI22D2BWP12T U2633 ( .A1(n1517), .A2(n2669), .B1(n1438), .B2(n2667), .ZN(
        n1543) );
  XOR3XD4BWP12T U2634 ( .A1(n1542), .A2(n1543), .A3(n1540), .Z(n1501) );
  TPOAI22D4BWP12T U2635 ( .A1(n1551), .A2(n4257), .B1(n1440), .B2(n2646), .ZN(
        n1554) );
  XNR2XD4BWP12T U2636 ( .A1(n4761), .A2(n288), .ZN(n1561) );
  TPOAI22D1BWP12T U2637 ( .A1(n1443), .A2(n2748), .B1(n1552), .B2(n2747), .ZN(
        n1556) );
  XOR3XD4BWP12T U2638 ( .A1(n1554), .A2(n1553), .A3(n1556), .Z(n1499) );
  CKND3BWP12T U2639 ( .I(n1499), .ZN(n1444) );
  XNR3XD4BWP12T U2640 ( .A1(n1500), .A2(n1501), .A3(n1444), .ZN(n1569) );
  XOR3XD4BWP12T U2641 ( .A1(n1571), .A2(n1570), .A3(n1569), .Z(n1576) );
  CKND3BWP12T U2642 ( .I(n1449), .ZN(n1445) );
  TPND2D2BWP12T U2643 ( .A1(n1448), .A2(n1445), .ZN(n1447) );
  CKND2D2BWP12T U2644 ( .A1(n1450), .A2(n1449), .ZN(n1451) );
  OAI21D1BWP12T U2645 ( .A1(n1455), .A2(n1454), .B(n1453), .ZN(n1457) );
  ND2D1BWP12T U2646 ( .A1(n1455), .A2(n1454), .ZN(n1456) );
  NR2D1BWP12T U2647 ( .A1(n1460), .A2(n1459), .ZN(n1463) );
  INVD1P75BWP12T U2648 ( .I(n1458), .ZN(n1462) );
  ND2XD1BWP12T U2649 ( .A1(n1460), .A2(n1459), .ZN(n1461) );
  TPOAI21D1BWP12T U2650 ( .A1(n1463), .A2(n1462), .B(n1461), .ZN(n1530) );
  XNR2XD4BWP12T U2651 ( .A1(n2619), .A2(n2701), .ZN(n1547) );
  XNR2XD4BWP12T U2652 ( .A1(n2623), .A2(n5014), .ZN(n1558) );
  TPOAI22D1BWP12T U2653 ( .A1(n1558), .A2(n2265), .B1(n1518), .B2(n2263), .ZN(
        n1525) );
  HA1D2BWP12T U2654 ( .A(n1466), .B(n1465), .CO(n1523), .S(n1432) );
  XOR3D2BWP12T U2655 ( .A1(n1524), .A2(n1525), .A3(n1523), .Z(n1529) );
  CKND2BWP12T U2656 ( .I(n1470), .ZN(n1467) );
  IND2D2BWP12T U2657 ( .A1(n1471), .B1(n1467), .ZN(n1468) );
  TPND2D2BWP12T U2658 ( .A1(n1473), .A2(n1472), .ZN(n1528) );
  XOR3XD4BWP12T U2659 ( .A1(n1530), .A2(n1529), .A3(n1528), .Z(n1536) );
  INVD2P3BWP12T U2660 ( .I(n1479), .ZN(n1475) );
  TPND2D2BWP12T U2661 ( .A1(n1475), .A2(n1474), .ZN(n1476) );
  ND2D1BWP12T U2662 ( .A1(n1479), .A2(n1478), .ZN(n1480) );
  TPND2D3BWP12T U2663 ( .A1(n1481), .A2(n1480), .ZN(n1534) );
  XOR3XD4BWP12T U2664 ( .A1(n1535), .A2(n1536), .A3(n1534), .Z(n1577) );
  XOR3XD4BWP12T U2665 ( .A1(n1576), .A2(n1579), .A3(n1577), .Z(n1495) );
  IND2D2BWP12T U2666 ( .A1(n1485), .B1(n1484), .ZN(n1482) );
  ND2D3BWP12T U2667 ( .A1(n1483), .A2(n1482), .ZN(n1488) );
  ND2D1BWP12T U2668 ( .A1(n1486), .A2(n1485), .ZN(n1487) );
  TPND2D2BWP12T U2669 ( .A1(n1488), .A2(n1487), .ZN(n1494) );
  TPNR2D3BWP12T U2670 ( .A1(n1495), .A2(n1494), .ZN(n3867) );
  TPND2D2BWP12T U2671 ( .A1(n1491), .A2(n1490), .ZN(n4291) );
  TPOAI21D4BWP12T U2672 ( .A1(n3022), .A2(n4291), .B(n3023), .ZN(n3864) );
  TPAOI21D1BWP12T U2673 ( .A1(n3866), .A2(n1498), .B(n1497), .ZN(n1586) );
  CKND2D2BWP12T U2674 ( .A1(n1501), .A2(n332), .ZN(n1502) );
  ND2XD3BWP12T U2675 ( .A1(n1503), .A2(n1502), .ZN(n2459) );
  CKND3BWP12T U2676 ( .I(n1509), .ZN(n1505) );
  INVD1BWP12T U2677 ( .I(n1508), .ZN(n1504) );
  TPND2D2BWP12T U2678 ( .A1(n1505), .A2(n1504), .ZN(n1507) );
  ND2D1BWP12T U2679 ( .A1(n1509), .A2(n1508), .ZN(n1510) );
  ND2D3BWP12T U2680 ( .A1(n1511), .A2(n1510), .ZN(n2329) );
  ND2D3BWP12T U2681 ( .A1(n1513), .A2(n4916), .ZN(n1515) );
  XOR2XD4BWP12T U2682 ( .A1(n4916), .A2(n4728), .Z(n1514) );
  ND2XD16BWP12T U2683 ( .A1(n2643), .A2(n1514), .ZN(n1894) );
  TPOAI22D4BWP12T U2684 ( .A1(n2233), .A2(n2691), .B1(n1516), .B2(n2689), .ZN(
        n2257) );
  XNR2XD4BWP12T U2685 ( .A1(n2098), .A2(n2666), .ZN(n2237) );
  XOR3XD4BWP12T U2686 ( .A1(n2261), .A2(n2257), .A3(n2258), .Z(n2328) );
  TPNR2D1BWP12T U2687 ( .A1(n1520), .A2(n1519), .ZN(n1521) );
  TPND2D1BWP12T U2688 ( .A1(n340), .A2(n1521), .ZN(n1522) );
  ND2D1BWP12T U2689 ( .A1(n1523), .A2(n1522), .ZN(n1527) );
  ND2D1BWP12T U2690 ( .A1(n1525), .A2(n1524), .ZN(n1526) );
  AN2D4BWP12T U2691 ( .A1(n1527), .A2(n1526), .Z(n2331) );
  XOR3XD4BWP12T U2692 ( .A1(n2329), .A2(n2328), .A3(n2331), .Z(n2458) );
  OAI21D1BWP12T U2693 ( .A1(n1529), .A2(n1530), .B(n1528), .ZN(n1532) );
  ND2D1BWP12T U2694 ( .A1(n1530), .A2(n1529), .ZN(n1531) );
  TPND2D2BWP12T U2695 ( .A1(n1532), .A2(n1531), .ZN(n2456) );
  INVD1P75BWP12T U2696 ( .I(n2456), .ZN(n1533) );
  XOR3XD4BWP12T U2697 ( .A1(n2459), .A2(n2458), .A3(n1533), .Z(n2499) );
  DCCKND4BWP12T U2698 ( .I(n1534), .ZN(n1538) );
  TPOAI21D2BWP12T U2699 ( .A1(n1539), .A2(n1538), .B(n1537), .ZN(n2498) );
  IND2XD1BWP12T U2700 ( .A1(n1541), .B1(n1540), .ZN(n1545) );
  ND2D1BWP12T U2701 ( .A1(n1543), .A2(n1542), .ZN(n1544) );
  CKND2D2BWP12T U2702 ( .A1(n1545), .A2(n1544), .ZN(n2410) );
  XNR2D1BWP12T U2703 ( .A1(n4316), .A2(n4916), .ZN(n1546) );
  XNR2D1BWP12T U2704 ( .A1(n1932), .A2(n4916), .ZN(n2236) );
  XNR2D1BWP12T U2705 ( .A1(n2551), .A2(n2701), .ZN(n2318) );
  TPOAI22D2BWP12T U2706 ( .A1(n1547), .A2(n2702), .B1(n2318), .B2(n2319), .ZN(
        n2377) );
  XNR2XD4BWP12T U2707 ( .A1(n4628), .A2(n4924), .ZN(n2219) );
  TPOAI22D4BWP12T U2708 ( .A1(n1548), .A2(n2218), .B1(n2220), .B2(n2219), .ZN(
        n2270) );
  TPOAI22D2BWP12T U2709 ( .A1(n1549), .A2(n306), .B1(n2624), .B2(n2222), .ZN(
        n2269) );
  XOR3XD4BWP12T U2710 ( .A1(n2378), .A2(n2377), .A3(n2373), .Z(n2411) );
  XNR2XD4BWP12T U2711 ( .A1(n4726), .A2(n2742), .ZN(n2322) );
  XNR2XD2BWP12T U2712 ( .A1(n2591), .A2(n2593), .ZN(n2323) );
  XNR2D1BWP12T U2713 ( .A1(n4764), .A2(n2746), .ZN(n2255) );
  OAI22D1BWP12T U2714 ( .A1(n1552), .A2(n2748), .B1(n2255), .B2(n2747), .ZN(
        n2325) );
  XOR3XD4BWP12T U2715 ( .A1(n2410), .A2(n2411), .A3(n2409), .Z(n2483) );
  ND2D1BWP12T U2716 ( .A1(n1554), .A2(n335), .ZN(n1555) );
  IOA21D2BWP12T U2717 ( .A1(n1556), .A2(n316), .B(n1555), .ZN(n2416) );
  TPOAI22D1BWP12T U2718 ( .A1(n1557), .A2(n2680), .B1(n2267), .B2(n2682), .ZN(
        n2338) );
  NR2D2BWP12T U2719 ( .A1(n2263), .A2(n1558), .ZN(n1560) );
  TPNR2D1BWP12T U2720 ( .A1(n2264), .A2(n2739), .ZN(n1559) );
  TPNR2D2BWP12T U2721 ( .A1(n1560), .A2(n1559), .ZN(n2340) );
  XNR2D1BWP12T U2722 ( .A1(n280), .A2(n288), .ZN(n2254) );
  OAI22D1BWP12T U2723 ( .A1(n2648), .A2(n1561), .B1(n2254), .B2(n2647), .ZN(
        n2343) );
  XOR3D2BWP12T U2724 ( .A1(n2338), .A2(n2340), .A3(n2343), .Z(n2418) );
  NR2D1BWP12T U2725 ( .A1(n1564), .A2(n1563), .ZN(n1566) );
  ND2D1BWP12T U2726 ( .A1(n1564), .A2(n1563), .ZN(n1565) );
  OAI21D2BWP12T U2727 ( .A1(n1567), .A2(n1566), .B(n1565), .ZN(n2414) );
  XNR3XD4BWP12T U2728 ( .A1(n2416), .A2(n2418), .A3(n2414), .ZN(n2484) );
  INVD1BWP12T U2729 ( .I(n1570), .ZN(n1573) );
  INVD1BWP12T U2730 ( .I(n1571), .ZN(n1572) );
  ND2D1BWP12T U2731 ( .A1(n1573), .A2(n1572), .ZN(n1574) );
  TPND2D2BWP12T U2732 ( .A1(n1575), .A2(n1574), .ZN(n2480) );
  XOR3XD4BWP12T U2733 ( .A1(n2483), .A2(n2484), .A3(n2480), .Z(n2497) );
  XOR3XD4BWP12T U2734 ( .A1(n2499), .A2(n2498), .A3(n2497), .Z(n1583) );
  BUFFXD3BWP12T U2735 ( .I(n1576), .Z(n1578) );
  TPOAI21D2BWP12T U2736 ( .A1(n1579), .A2(n1578), .B(n1577), .ZN(n1581) );
  TPND2D2BWP12T U2737 ( .A1(n1581), .A2(n1580), .ZN(n1582) );
  ND2D3BWP12T U2738 ( .A1(n1583), .A2(n1582), .ZN(n2441) );
  INVD1BWP12T U2739 ( .I(n304), .ZN(n1584) );
  AN2XD2BWP12T U2740 ( .A1(n2441), .A2(n1584), .Z(n1585) );
  XNR2XD4BWP12T U2741 ( .A1(n1586), .A2(n1585), .ZN(n4294) );
  ND2XD8BWP12T U2742 ( .A1(n4294), .A2(n5085), .ZN(n1683) );
  NR2D1BWP12T U2743 ( .A1(n4716), .A2(n4927), .ZN(n4189) );
  NR2D1BWP12T U2744 ( .A1(n4717), .A2(n2688), .ZN(n3089) );
  NR2D1BWP12T U2745 ( .A1(n4189), .A2(n3089), .ZN(n1593) );
  ND2D1BWP12T U2746 ( .A1(n1587), .A2(n1607), .ZN(n1591) );
  NR2D1BWP12T U2747 ( .A1(n4070), .A2(n1591), .ZN(n4192) );
  CKND2D1BWP12T U2748 ( .A1(n1593), .A2(n4192), .ZN(n1595) );
  INVD1BWP12T U2749 ( .I(n1588), .ZN(n1605) );
  AOI21D1BWP12T U2750 ( .A1(n1589), .A2(n1607), .B(n1605), .ZN(n1590) );
  OAI21D1BWP12T U2751 ( .A1(n4073), .A2(n1591), .B(n1590), .ZN(n4191) );
  ND2D1BWP12T U2752 ( .A1(n4716), .A2(n4927), .ZN(n4190) );
  ND2D1BWP12T U2753 ( .A1(n4717), .A2(n2688), .ZN(n3090) );
  OAI21D1BWP12T U2754 ( .A1(n3089), .A2(n4190), .B(n3090), .ZN(n1592) );
  AOI21D1BWP12T U2755 ( .A1(n1593), .A2(n4191), .B(n1592), .ZN(n1594) );
  INVD3BWP12T U2756 ( .I(n3788), .ZN(n4353) );
  BUFFD3BWP12T U2757 ( .I(n2226), .Z(n4762) );
  NR2D1BWP12T U2758 ( .A1(n4714), .A2(n4923), .ZN(n1800) );
  CKBD1BWP12T U2759 ( .I(n4924), .Z(n1597) );
  NR2D1BWP12T U2760 ( .A1(n4715), .A2(n1597), .ZN(n3743) );
  NR2D1BWP12T U2761 ( .A1(n1800), .A2(n3743), .ZN(n4349) );
  BUFFXD8BWP12T U2762 ( .I(n2243), .Z(n5053) );
  NR2D1BWP12T U2763 ( .A1(n4713), .A2(n5051), .ZN(n3026) );
  NR2D1BWP12T U2764 ( .A1(n4712), .A2(n4914), .ZN(n3029) );
  NR2D1BWP12T U2765 ( .A1(n3026), .A2(n3029), .ZN(n1599) );
  ND2D1BWP12T U2766 ( .A1(n4349), .A2(n1599), .ZN(n3873) );
  CKBD1BWP12T U2767 ( .I(b[22]), .Z(n4729) );
  NR2D1BWP12T U2768 ( .A1(n4683), .A2(n4728), .ZN(n2941) );
  INVD1BWP12T U2769 ( .I(n2941), .ZN(n3875) );
  ND2XD0BWP12T U2770 ( .A1(n3930), .A2(n3875), .ZN(n1601) );
  ND2D1BWP12T U2771 ( .A1(n4714), .A2(n4923), .ZN(n3739) );
  ND2D1BWP12T U2772 ( .A1(n4715), .A2(n1597), .ZN(n3744) );
  OAI21D1BWP12T U2773 ( .A1(n3743), .A2(n3739), .B(n3744), .ZN(n4350) );
  ND2D1BWP12T U2774 ( .A1(n4713), .A2(n5051), .ZN(n4354) );
  ND2D1BWP12T U2775 ( .A1(n4712), .A2(n1598), .ZN(n3030) );
  ND2D1BWP12T U2776 ( .A1(n4683), .A2(n4728), .ZN(n3874) );
  CKND0BWP12T U2777 ( .I(n3874), .ZN(n2954) );
  AOI21D1BWP12T U2778 ( .A1(n3933), .A2(n3875), .B(n2954), .ZN(n1600) );
  OAI21D1BWP12T U2779 ( .A1(n4353), .A2(n1601), .B(n1600), .ZN(n1604) );
  BUFFXD4BWP12T U2780 ( .I(n2591), .Z(n4732) );
  CKND0BWP12T U2781 ( .I(n4732), .ZN(n4688) );
  CKBD1BWP12T U2782 ( .I(n4916), .Z(n1663) );
  NR2D1BWP12T U2783 ( .A1(n4688), .A2(n1663), .ZN(n2943) );
  INVD1BWP12T U2784 ( .I(n2943), .ZN(n2953) );
  CKBD1BWP12T U2785 ( .I(n4916), .Z(n1602) );
  ND2D1BWP12T U2786 ( .A1(n4688), .A2(n1602), .ZN(n2942) );
  CKND2D1BWP12T U2787 ( .A1(n2953), .A2(n2942), .ZN(n1603) );
  ND2D1BWP12T U2788 ( .A1(n4021), .A2(n1607), .ZN(n1609) );
  NR2D1BWP12T U2789 ( .A1(n4016), .A2(n1609), .ZN(n1611) );
  ND2D1BWP12T U2790 ( .A1(n1703), .A2(n1611), .ZN(n1613) );
  AOI21D1BWP12T U2791 ( .A1(n1607), .A2(n1606), .B(n1605), .ZN(n1608) );
  OAI21D1BWP12T U2792 ( .A1(n4015), .A2(n1609), .B(n1608), .ZN(n1610) );
  AOI21D1BWP12T U2793 ( .A1(n1702), .A2(n1611), .B(n1610), .ZN(n1612) );
  NR2D1BWP12T U2794 ( .A1(n4189), .A2(n3089), .ZN(n3738) );
  NR2D1BWP12T U2795 ( .A1(n1800), .A2(n3743), .ZN(n1616) );
  ND2D1BWP12T U2796 ( .A1(n3738), .A2(n1616), .ZN(n4984) );
  INVD1BWP12T U2797 ( .I(n4984), .ZN(n3876) );
  NR2D1BWP12T U2798 ( .A1(n3026), .A2(n3029), .ZN(n3878) );
  INVD1BWP12T U2799 ( .I(n3878), .ZN(n2951) );
  NR2XD0BWP12T U2800 ( .A1(n2951), .A2(n2941), .ZN(n1618) );
  TPND2D0BWP12T U2801 ( .A1(n3876), .A2(n1618), .ZN(n1620) );
  OAI21D1BWP12T U2802 ( .A1(n3089), .A2(n4190), .B(n3090), .ZN(n3740) );
  OAI21D1BWP12T U2803 ( .A1(n3743), .A2(n3739), .B(n3744), .ZN(n1615) );
  AOI21D1BWP12T U2804 ( .A1(n1616), .A2(n3740), .B(n1615), .ZN(n4983) );
  INVD1BWP12T U2805 ( .I(n4983), .ZN(n3879) );
  OAI21D1BWP12T U2806 ( .A1(n3029), .A2(n4354), .B(n3030), .ZN(n3877) );
  CKND0BWP12T U2807 ( .I(n3877), .ZN(n2957) );
  OAI21D0BWP12T U2808 ( .A1(n2957), .A2(n2941), .B(n3874), .ZN(n1617) );
  AOI21D1BWP12T U2809 ( .A1(n3879), .A2(n1618), .B(n1617), .ZN(n1619) );
  OAI21D1BWP12T U2810 ( .A1(n4985), .A2(n1620), .B(n1619), .ZN(n1622) );
  ND2D1BWP12T U2811 ( .A1(n2953), .A2(n2942), .ZN(n1621) );
  XNR2XD1BWP12T U2812 ( .A1(n1622), .A2(n1621), .ZN(n4988) );
  INVD1BWP12T U2813 ( .I(n4384), .ZN(n1630) );
  ND2D1BWP12T U2814 ( .A1(n4030), .A2(n4183), .ZN(n1625) );
  NR2D1BWP12T U2815 ( .A1(n4051), .A2(n1625), .ZN(n1627) );
  ND2D1BWP12T U2816 ( .A1(n3206), .A2(n1627), .ZN(n1629) );
  INVD1BWP12T U2817 ( .I(n1642), .ZN(n4182) );
  AOI21D1BWP12T U2818 ( .A1(n4183), .A2(n1623), .B(n4182), .ZN(n1624) );
  OAI21D1BWP12T U2819 ( .A1(n4050), .A2(n1625), .B(n1624), .ZN(n1626) );
  AOI21D1BWP12T U2820 ( .A1(n1734), .A2(n1627), .B(n1626), .ZN(n1628) );
  TPOAI21D1BWP12T U2821 ( .A1(n1630), .A2(n1629), .B(n1628), .ZN(n2791) );
  INVD2BWP12T U2822 ( .I(n2791), .ZN(n4367) );
  NR2D1BWP12T U2823 ( .A1(n4761), .A2(n4927), .ZN(n4149) );
  NR2D1BWP12T U2824 ( .A1(n279), .A2(n2688), .ZN(n1808) );
  NR2D1BWP12T U2825 ( .A1(n4149), .A2(n1808), .ZN(n3781) );
  NR2D1BWP12T U2826 ( .A1(n4762), .A2(n4923), .ZN(n1809) );
  NR2D1BWP12T U2827 ( .A1(n3771), .A2(n4764), .ZN(n4475) );
  NR2D1BWP12T U2828 ( .A1(n1809), .A2(n4475), .ZN(n1633) );
  ND2D1BWP12T U2829 ( .A1(n3781), .A2(n1633), .ZN(n4366) );
  INVD1BWP12T U2830 ( .I(n4366), .ZN(n3907) );
  NR2D1BWP12T U2831 ( .A1(n5053), .A2(n5051), .ZN(n3072) );
  NR2D1BWP12T U2832 ( .A1(n4726), .A2(n1631), .ZN(n3039) );
  NR2D1BWP12T U2833 ( .A1(n3072), .A2(n3039), .ZN(n3909) );
  INVD0BWP12T U2834 ( .I(n3909), .ZN(n2965) );
  NR2D1BWP12T U2835 ( .A1(n4729), .A2(n4728), .ZN(n2964) );
  NR2XD0BWP12T U2836 ( .A1(n2965), .A2(n2964), .ZN(n1636) );
  TPND2D0BWP12T U2837 ( .A1(n3907), .A2(n1636), .ZN(n1638) );
  ND2D1BWP12T U2838 ( .A1(n4761), .A2(n4927), .ZN(n4150) );
  ND2D1BWP12T U2839 ( .A1(n279), .A2(n2688), .ZN(n3093) );
  OAI21D1BWP12T U2840 ( .A1(n1808), .A2(n4150), .B(n3093), .ZN(n3784) );
  ND2D1BWP12T U2841 ( .A1(n4762), .A2(n4923), .ZN(n3782) );
  ND2D1BWP12T U2842 ( .A1(n336), .A2(n3771), .ZN(n4474) );
  TPOAI21D0BWP12T U2843 ( .A1(n4475), .A2(n3782), .B(n4474), .ZN(n1632) );
  AOI21D1BWP12T U2844 ( .A1(n1633), .A2(n3784), .B(n1632), .ZN(n4365) );
  INVD1BWP12T U2845 ( .I(n4365), .ZN(n3910) );
  ND2D1BWP12T U2846 ( .A1(n5053), .A2(n5051), .ZN(n4368) );
  ND2D1BWP12T U2847 ( .A1(n4726), .A2(n1634), .ZN(n3884) );
  OAI21D1BWP12T U2848 ( .A1(n3039), .A2(n4368), .B(n3884), .ZN(n3908) );
  CKND0BWP12T U2849 ( .I(n3908), .ZN(n2966) );
  ND2D1BWP12T U2850 ( .A1(n4729), .A2(n4728), .ZN(n3888) );
  OAI21D0BWP12T U2851 ( .A1(n2966), .A2(n2964), .B(n3888), .ZN(n1635) );
  TPAOI21D0BWP12T U2852 ( .A1(n3910), .A2(n1636), .B(n1635), .ZN(n1637) );
  OAI21D1BWP12T U2853 ( .A1(n4367), .A2(n1638), .B(n1637), .ZN(n1640) );
  NR2D1BWP12T U2854 ( .A1(n4732), .A2(n1639), .ZN(n2795) );
  INVD1BWP12T U2855 ( .I(n2795), .ZN(n2970) );
  CKBD1BWP12T U2856 ( .I(n4916), .Z(n4648) );
  ND2D1BWP12T U2857 ( .A1(n4732), .A2(n4648), .ZN(n2798) );
  CKND2D0BWP12T U2858 ( .A1(n2970), .A2(n2798), .ZN(n1651) );
  XNR2D1BWP12T U2859 ( .A1(n1640), .A2(n1651), .ZN(n4371) );
  NR2D1BWP12T U2860 ( .A1(n1808), .A2(n1809), .ZN(n1644) );
  NR2D1BWP12T U2861 ( .A1(n4149), .A2(n1641), .ZN(n1805) );
  CKND2D1BWP12T U2862 ( .A1(n1644), .A2(n1805), .ZN(n1646) );
  NR2D1BWP12T U2863 ( .A1(n1646), .A2(n1802), .ZN(n1648) );
  OAI21D1BWP12T U2864 ( .A1(n4149), .A2(n1642), .B(n4150), .ZN(n1804) );
  OAI21D0BWP12T U2865 ( .A1(n1809), .A2(n3093), .B(n3782), .ZN(n1643) );
  AOI21D1BWP12T U2866 ( .A1(n1644), .A2(n1804), .B(n1643), .ZN(n1645) );
  OAI21D1BWP12T U2867 ( .A1(n1646), .A2(n1803), .B(n1645), .ZN(n1647) );
  TPAOI21D2BWP12T U2868 ( .A1(n3199), .A2(n1648), .B(n1647), .ZN(n4476) );
  TPNR2D0BWP12T U2869 ( .A1(n3072), .A2(n4475), .ZN(n3037) );
  NR2D1BWP12T U2870 ( .A1(n3039), .A2(n2964), .ZN(n1650) );
  ND2D1BWP12T U2871 ( .A1(n3037), .A2(n1650), .ZN(n2796) );
  OAI21D1BWP12T U2872 ( .A1(n3072), .A2(n4474), .B(n4368), .ZN(n3038) );
  TPOAI21D0BWP12T U2873 ( .A1(n2964), .A2(n3884), .B(n3888), .ZN(n1649) );
  AOI21D1BWP12T U2874 ( .A1(n1650), .A2(n3038), .B(n1649), .ZN(n2801) );
  XNR2XD1BWP12T U2875 ( .A1(n3830), .A2(n1651), .ZN(n4511) );
  NR2D1BWP12T U2876 ( .A1(n3224), .A2(n4743), .ZN(n1674) );
  TPAOI21D0BWP12T U2877 ( .A1(n4889), .A2(n1674), .B(n3843), .ZN(n4851) );
  INVD3BWP12T U2878 ( .I(n4611), .ZN(n4158) );
  MUX2D1BWP12T U2879 ( .I0(n4465), .I1(n4651), .S(n5075), .Z(n2918) );
  INVD1BWP12T U2880 ( .I(n5051), .ZN(n5047) );
  MUX2D1BWP12T U2881 ( .I0(n4625), .I1(n5047), .S(n5075), .Z(n3810) );
  AOI22D1BWP12T U2882 ( .A1(n3125), .A2(n2918), .B1(n3810), .B2(n953), .ZN(
        n1654) );
  MUX2XD0BWP12T U2883 ( .I0(n1810), .I1(n4638), .S(n5075), .Z(n3119) );
  MUX2XD0BWP12T U2884 ( .I0(n1342), .I1(n4637), .S(n5075), .Z(n3811) );
  AOI22D1BWP12T U2885 ( .A1(n3122), .A2(n3119), .B1(n3811), .B2(n3701), .ZN(
        n1653) );
  ND2D1BWP12T U2886 ( .A1(n1654), .A2(n1653), .ZN(n2867) );
  OAI22D1BWP12T U2887 ( .A1(n1655), .A2(n4685), .B1(n4585), .B2(n4707), .ZN(
        n1656) );
  CKND2D2BWP12T U2888 ( .A1(n4573), .A2(n3969), .ZN(n4156) );
  AOI211D1BWP12T U2889 ( .A1(n4158), .A2(n2867), .B(n1656), .C(n4156), .ZN(
        n4603) );
  AN2XD2BWP12T U2890 ( .A1(n4448), .A2(n3142), .Z(n4426) );
  ND2D1BWP12T U2891 ( .A1(n1810), .A2(n4638), .ZN(n3770) );
  CKND0BWP12T U2892 ( .I(n4923), .ZN(n1833) );
  CKND2D1BWP12T U2893 ( .A1(n1342), .A2(n1833), .ZN(n1657) );
  NR2D1BWP12T U2894 ( .A1(n3770), .A2(n1657), .ZN(n4425) );
  CKND1BWP12T U2895 ( .I(n4425), .ZN(n3892) );
  ND2D1BWP12T U2896 ( .A1(n4625), .A2(n1658), .ZN(n3891) );
  CKND0BWP12T U2897 ( .I(n3891), .ZN(n1659) );
  CKND2D0BWP12T U2898 ( .A1(n1659), .A2(n4651), .ZN(n1660) );
  NR2D1BWP12T U2899 ( .A1(n3892), .A2(n1660), .ZN(n1661) );
  CKND2D1BWP12T U2900 ( .A1(n4426), .A2(n1661), .ZN(n1662) );
  CKBD1BWP12T U2901 ( .I(n4916), .Z(n2781) );
  XOR2D1BWP12T U2902 ( .A1(n1662), .A2(n2781), .Z(n4442) );
  OAI21D0BWP12T U2903 ( .A1(n1663), .A2(n5083), .B(n5081), .ZN(n1667) );
  MUX2ND0BWP12T U2904 ( .I0(n5077), .I1(n5076), .S(n4732), .ZN(n1664) );
  NR2D0BWP12T U2905 ( .A1(n1664), .A2(n905), .ZN(n1665) );
  MUX2ND0BWP12T U2906 ( .I0(n1665), .I1(n5080), .S(n1856), .ZN(n1666) );
  RCAOI21D0BWP12T U2907 ( .A1(n4732), .A2(n1667), .B(n1666), .ZN(n1668) );
  IOA21D1BWP12T U2908 ( .A1(n4442), .A2(n5078), .B(n1668), .ZN(n1669) );
  TPAOI21D0BWP12T U2909 ( .A1(n4167), .A2(n4603), .B(n1669), .ZN(n1670) );
  OAI21D0BWP12T U2910 ( .A1(n4851), .A2(n5063), .B(n1670), .ZN(n1677) );
  INVD1BWP12T U2911 ( .I(n1671), .ZN(n2858) );
  AOI22D1BWP12T U2912 ( .A1(n4801), .A2(n2859), .B1(n2858), .B2(n3754), .ZN(
        n1672) );
  NR2D1BWP12T U2913 ( .A1(n4032), .A2(n3758), .ZN(n3947) );
  ND2D1BWP12T U2914 ( .A1(n4200), .A2(n4158), .ZN(n3817) );
  INVD1BWP12T U2915 ( .I(n3817), .ZN(n3690) );
  NR2D1BWP12T U2916 ( .A1(n3947), .A2(n3690), .ZN(n3756) );
  OAI211D1BWP12T U2917 ( .A1(n3758), .A2(n4779), .B(n1672), .C(n3756), .ZN(
        n4807) );
  NR2D1BWP12T U2918 ( .A1(n4807), .A2(n5040), .ZN(n1676) );
  TPNR2D0BWP12T U2919 ( .A1(n3899), .A2(n4540), .ZN(n1675) );
  NR3XD0BWP12T U2920 ( .A1(n1677), .A2(n1676), .A3(n1675), .ZN(n1678) );
  IOA21D1BWP12T U2921 ( .A1(n4511), .A2(n4103), .B(n1678), .ZN(n1679) );
  AOI21D1BWP12T U2922 ( .A1(n5088), .A2(n4371), .B(n1679), .ZN(n1680) );
  TPAOI21D4BWP12T U2923 ( .A1(n5090), .A2(n4357), .B(n1681), .ZN(n1682) );
  TPND2D8BWP12T U2924 ( .A1(n1683), .A2(n1682), .ZN(result[23]) );
  TPAOI21D1BWP12T U2925 ( .A1(n3267), .A2(n3266), .B(n1684), .ZN(n4270) );
  INVD1BWP12T U2926 ( .I(n4271), .ZN(n1686) );
  ND2D1BWP12T U2927 ( .A1(n1688), .A2(n1687), .ZN(n1689) );
  XNR2XD4BWP12T U2928 ( .A1(n1690), .A2(n1689), .ZN(n4275) );
  ND2D4BWP12T U2929 ( .A1(n4275), .A2(n5085), .ZN(n1743) );
  OAI21D1BWP12T U2930 ( .A1(n4493), .A2(n1691), .B(n4491), .ZN(n1692) );
  CKND2D1BWP12T U2931 ( .A1(n3205), .A2(n3207), .ZN(n1735) );
  XNR2D1BWP12T U2932 ( .A1(n1692), .A2(n1735), .ZN(n4481) );
  CKND0BWP12T U2933 ( .I(n4332), .ZN(n1693) );
  NR2D0BWP12T U2934 ( .A1(n1693), .A2(n4334), .ZN(n1696) );
  CKND0BWP12T U2935 ( .I(n4331), .ZN(n1694) );
  OAI21D0BWP12T U2936 ( .A1(n1694), .A2(n4334), .B(n4972), .ZN(n1695) );
  AOI21D1BWP12T U2937 ( .A1(n4333), .A2(n1696), .B(n1695), .ZN(n1698) );
  CKND2D0BWP12T U2938 ( .A1(n1697), .A2(n3172), .ZN(n1704) );
  XOR2XD1BWP12T U2939 ( .A1(n1698), .A2(n1704), .Z(n4339) );
  MUX2XD0BWP12T U2940 ( .I0(n4631), .I1(n4627), .S(n5075), .Z(n1822) );
  MUX2XD0BWP12T U2941 ( .I0(n4652), .I1(n777), .S(n5075), .Z(n2999) );
  AOI22D1BWP12T U2942 ( .A1(n3122), .A2(n1822), .B1(n2999), .B2(n3125), .ZN(
        n1700) );
  MUX2XD0BWP12T U2943 ( .I0(n4654), .I1(n3523), .S(n5075), .Z(n3447) );
  MUX2D1BWP12T U2944 ( .I0(n4655), .I1(n4679), .S(n5075), .Z(n1821) );
  AOI22D1BWP12T U2945 ( .A1(n953), .A2(n3447), .B1(n1821), .B2(n3701), .ZN(
        n1699) );
  ND2D1BWP12T U2946 ( .A1(n1700), .A2(n1699), .ZN(n4608) );
  ND2D1BWP12T U2947 ( .A1(n3219), .A2(n4910), .ZN(n4567) );
  MUX2D1BWP12T U2948 ( .I0(n4921), .I1(n289), .S(n5075), .Z(n3471) );
  INVD1BWP12T U2949 ( .I(n3471), .ZN(n3004) );
  MUX2ND0BWP12T U2950 ( .I0(n4608), .I1(n4607), .S(n4743), .ZN(n1701) );
  CKND2D1BWP12T U2951 ( .A1(n1701), .A2(n4605), .ZN(n4593) );
  AOI21D1BWP12T U2952 ( .A1(n4971), .A2(n1703), .B(n1702), .ZN(n1705) );
  XOR2XD1BWP12T U2953 ( .A1(n1705), .A2(n1704), .Z(n4976) );
  MOAI22D1BWP12T U2954 ( .A1(n5042), .A2(n4593), .B1(n4976), .B2(n5093), .ZN(
        n1732) );
  CKND0BWP12T U2955 ( .I(n4173), .ZN(n4535) );
  OR2XD4BWP12T U2956 ( .A1(n4743), .A2(n4742), .Z(n4566) );
  ND2XD0BWP12T U2957 ( .A1(n4535), .A2(n4039), .ZN(n1717) );
  OAI22D1BWP12T U2958 ( .A1(n3323), .A2(n5047), .B1(n3321), .B2(n4651), .ZN(
        n1707) );
  OAI22D1BWP12T U2959 ( .A1(n3322), .A2(n4465), .B1(n275), .B2(n4625), .ZN(
        n1706) );
  NR2D1BWP12T U2960 ( .A1(n1707), .A2(n1706), .ZN(n4170) );
  INR2D1BWP12T U2961 ( .A1(n3051), .B1(n4170), .ZN(n1708) );
  INVD1BWP12T U2962 ( .I(n4171), .ZN(n1711) );
  OAI22D1BWP12T U2963 ( .A1(n3321), .A2(n4680), .B1(n275), .B2(n4653), .ZN(
        n1713) );
  OAI22D1BWP12T U2964 ( .A1(n3323), .A2(n4652), .B1(n3322), .B2(n4930), .ZN(
        n1712) );
  NR2D1BWP12T U2965 ( .A1(n1713), .A2(n1712), .ZN(n4555) );
  OAI22D1BWP12T U2966 ( .A1(n3323), .A2(n4638), .B1(n275), .B2(n1810), .ZN(
        n1715) );
  OAI22D1BWP12T U2967 ( .A1(n3321), .A2(n4637), .B1(n3322), .B2(n1342), .ZN(
        n1714) );
  NR2D1BWP12T U2968 ( .A1(n1715), .A2(n1714), .ZN(n4172) );
  INVD1BWP12T U2969 ( .I(n1720), .ZN(n1716) );
  AOI21D1BWP12T U2970 ( .A1(n4843), .A2(n1717), .B(n1716), .ZN(n4552) );
  INVD1BWP12T U2971 ( .I(n4068), .ZN(n3186) );
  CKND2D1BWP12T U2972 ( .A1(n4552), .A2(n3186), .ZN(n1730) );
  MUX2NXD0BWP12T U2973 ( .I0(n4173), .I1(n4624), .S(n4566), .ZN(n3983) );
  CKND0BWP12T U2974 ( .I(n3983), .ZN(n1718) );
  CKND2D0BWP12T U2975 ( .A1(n1718), .A2(n4843), .ZN(n1719) );
  CKND2D0BWP12T U2976 ( .A1(n4448), .A2(n1721), .ZN(n1722) );
  XOR2XD1BWP12T U2977 ( .A1(n1722), .A2(n4925), .Z(n4451) );
  MUX2ND0BWP12T U2978 ( .I0(n5077), .I1(n5076), .S(n4760), .ZN(n1723) );
  NR2D0BWP12T U2979 ( .A1(n1723), .A2(n905), .ZN(n1724) );
  MUX2ND0BWP12T U2980 ( .I0(n1724), .I1(n5080), .S(n4652), .ZN(n1727) );
  NR2D0BWP12T U2981 ( .A1(n4925), .A2(n5083), .ZN(n1725) );
  OA21XD0BWP12T U2982 ( .A1(n905), .A2(n1725), .B(n4760), .Z(n1726) );
  AOI211D1BWP12T U2983 ( .A1(n4451), .A2(n5078), .B(n1727), .C(n1726), .ZN(
        n1728) );
  OA21D1BWP12T U2984 ( .A1(n4878), .A2(n5063), .B(n1728), .Z(n1729) );
  CKND2D1BWP12T U2985 ( .A1(n1730), .A2(n1729), .ZN(n1731) );
  TPNR2D1BWP12T U2986 ( .A1(n1732), .A2(n1731), .ZN(n1733) );
  IOA21D1BWP12T U2987 ( .A1(n4339), .A2(n5090), .B(n1733), .ZN(n1739) );
  INVD1BWP12T U2988 ( .I(n4392), .ZN(n1737) );
  INVD3BWP12T U2989 ( .I(n3937), .ZN(n3945) );
  INVD1BWP12T U2990 ( .I(n2999), .ZN(n3458) );
  MUX2NXD0BWP12T U2991 ( .I0(n3946), .I1(n3938), .S(n4032), .ZN(n1736) );
  AOI21D1BWP12T U2992 ( .A1(n3758), .A2(n1736), .B(n4552), .ZN(n4828) );
  TPOAI22D1BWP12T U2993 ( .A1(n1737), .A2(n4396), .B1(n4828), .B2(n5040), .ZN(
        n1738) );
  TPNR2D1BWP12T U2994 ( .A1(n1739), .A2(n1738), .ZN(n1740) );
  IOA21D2BWP12T U2995 ( .A1(n4481), .A2(n4103), .B(n1740), .ZN(n1741) );
  INVD3BWP12T U2996 ( .I(n1741), .ZN(n1742) );
  ND2D8BWP12T U2997 ( .A1(n1743), .A2(n1742), .ZN(result[12]) );
  OAI22D0BWP12T U2998 ( .A1(n3321), .A2(n4631), .B1(n275), .B2(n4627), .ZN(
        n1745) );
  OAI22D1BWP12T U2999 ( .A1(n3318), .A2(n1765), .B1(n3322), .B2(n4679), .ZN(
        n1744) );
  NR2D1BWP12T U3000 ( .A1(n1745), .A2(n1744), .ZN(n4553) );
  OAI22D1BWP12T U3001 ( .A1(n4555), .A2(n4206), .B1(n4553), .B2(n4566), .ZN(
        n1750) );
  AOI22D0BWP12T U3002 ( .A1(n3218), .A2(n3523), .B1(n3217), .B2(n4654), .ZN(
        n1747) );
  AOI22D0BWP12T U3003 ( .A1(n3220), .A2(n777), .B1(n3219), .B2(n4655), .ZN(
        n1746) );
  ND2D1BWP12T U3004 ( .A1(n1747), .A2(n1746), .ZN(n4558) );
  INVD3BWP12T U3005 ( .I(n4556), .ZN(n4521) );
  OAI21D1BWP12T U3006 ( .A1(n4558), .A2(n4521), .B(n4707), .ZN(n1749) );
  NR2D1BWP12T U3007 ( .A1(n4172), .A2(n4554), .ZN(n1748) );
  TPNR3D2BWP12T U3008 ( .A1(n1750), .A2(n1749), .A3(n1748), .ZN(n4819) );
  NR2D1BWP12T U3009 ( .A1(n4173), .A2(n4206), .ZN(n1751) );
  AOI21D1BWP12T U3010 ( .A1(n1752), .A2(n4685), .B(n1751), .ZN(n4541) );
  OAI22D1BWP12T U3011 ( .A1(n4819), .A2(n4541), .B1(n3946), .B2(n3818), .ZN(
        n4837) );
  XNR2D1BWP12T U3012 ( .A1(n1756), .A2(n1755), .ZN(n4264) );
  CKND2D1BWP12T U3013 ( .A1(n4264), .A2(n5085), .ZN(n1757) );
  IOA21D1BWP12T U3014 ( .A1(n5094), .A2(n4837), .B(n1757), .ZN(n1761) );
  INVD1BWP12T U3015 ( .I(n3509), .ZN(n3408) );
  AOI21D0BWP12T U3016 ( .A1(n4742), .A2(n3408), .B(n4707), .ZN(n1758) );
  AOI211D1BWP12T U3017 ( .A1(n4541), .A2(n1758), .B(n4819), .C(n4891), .ZN(
        n1759) );
  INR2D1BWP12T U3018 ( .A1(n4046), .B1(n1759), .ZN(n4867) );
  INR2D1BWP12T U3019 ( .A1(n5099), .B1(n4867), .ZN(n1760) );
  INVD1BWP12T U3020 ( .I(n1762), .ZN(n3606) );
  XOR2XD1BWP12T U3021 ( .A1(n3606), .A2(n4921), .Z(n4422) );
  INVD1BWP12T U3022 ( .I(n5076), .ZN(n5044) );
  MUX2ND0BWP12T U3023 ( .I0(n5045), .I1(n5044), .S(n4843), .ZN(n1763) );
  CKND2D1BWP12T U3024 ( .A1(n1763), .A2(n5081), .ZN(n1764) );
  CKND1BWP12T U3025 ( .I(n1766), .ZN(n3621) );
  CKND2D1BWP12T U3026 ( .A1(n3352), .A2(n1776), .ZN(n1767) );
  XOR2XD1BWP12T U3027 ( .A1(n1768), .A2(n1767), .Z(n4401) );
  CKND1BWP12T U3028 ( .I(n3357), .ZN(n3359) );
  CKND2D1BWP12T U3029 ( .A1(n3359), .A2(n3360), .ZN(n1772) );
  XOR2XD1BWP12T U3030 ( .A1(n1773), .A2(n1772), .Z(n4958) );
  AOI22D1BWP12T U3031 ( .A1(n5088), .A2(n4401), .B1(n4958), .B2(n5093), .ZN(
        n1781) );
  OAI21D1BWP12T U3032 ( .A1(n4102), .A2(n1775), .B(n4100), .ZN(n1778) );
  CKND2D1BWP12T U3033 ( .A1(n3352), .A2(n1776), .ZN(n1777) );
  XNR2XD1BWP12T U3034 ( .A1(n1778), .A2(n1777), .ZN(n4496) );
  ND2XD0BWP12T U3035 ( .A1(n4496), .A2(n4103), .ZN(n1780) );
  OR2XD1BWP12T U3036 ( .A1(n3604), .A2(n4607), .Z(n1779) );
  ND3D1BWP12T U3037 ( .A1(n1781), .A2(n1780), .A3(n1779), .ZN(n1791) );
  OAI21D1BWP12T U3038 ( .A1(n4541), .A2(n4891), .B(n4890), .ZN(n1783) );
  INVD1BWP12T U3039 ( .I(n4819), .ZN(n1782) );
  ND2D1BWP12T U3040 ( .A1(n1783), .A2(n1782), .ZN(n4576) );
  INR2D1BWP12T U3041 ( .A1(n4209), .B1(n4576), .ZN(n1790) );
  OR2XD1BWP12T U3042 ( .A1(n4743), .A2(n1785), .Z(n4133) );
  INVD1BWP12T U3043 ( .I(n1786), .ZN(n4132) );
  CKND2D0BWP12T U3044 ( .A1(n4131), .A2(n1787), .ZN(n1788) );
  INVD1BWP12T U3045 ( .I(n1795), .ZN(n3732) );
  INVD1BWP12T U3046 ( .I(n3731), .ZN(n1796) );
  TPND2D1BWP12T U3047 ( .A1(n1796), .A2(n3730), .ZN(n1797) );
  XOR2XD4BWP12T U3048 ( .A1(n3732), .A2(n1797), .Z(n4283) );
  CKND0BWP12T U3049 ( .I(n3738), .ZN(n1799) );
  INVD1BWP12T U3050 ( .I(n3740), .ZN(n1798) );
  OAI21D1BWP12T U3051 ( .A1(n4985), .A2(n1799), .B(n1798), .ZN(n1801) );
  INVD1BWP12T U3052 ( .I(n1800), .ZN(n3787) );
  CKND2D0BWP12T U3053 ( .A1(n3787), .A2(n3739), .ZN(n1845) );
  INVD1BWP12T U3054 ( .I(n1802), .ZN(n4181) );
  CKND2D1BWP12T U3055 ( .A1(n4181), .A2(n1805), .ZN(n1807) );
  INVD1BWP12T U3056 ( .I(n1803), .ZN(n4184) );
  AOI21D1BWP12T U3057 ( .A1(n4184), .A2(n1805), .B(n1804), .ZN(n1806) );
  INVD0BWP12T U3058 ( .I(n1808), .ZN(n3094) );
  INVD1BWP12T U3059 ( .I(n1809), .ZN(n3783) );
  CKND2D1BWP12T U3060 ( .A1(n3783), .A2(n3782), .ZN(n1844) );
  ND2D1BWP12T U3061 ( .A1(n4502), .A2(n4103), .ZN(n1852) );
  MUX2XD0BWP12T U3062 ( .I0(n4637), .I1(n1810), .S(n5075), .Z(n3444) );
  MUX2XD0BWP12T U3063 ( .I0(n4932), .I1(n4926), .S(n5075), .Z(n3954) );
  NR2D0BWP12T U3064 ( .A1(n3945), .A2(n3954), .ZN(n1812) );
  MUX2XD0BWP12T U3065 ( .I0(n4927), .I1(n2666), .S(n5075), .Z(n3953) );
  OAI22D1BWP12T U3066 ( .A1(n3813), .A2(n3458), .B1(n3812), .B2(n3953), .ZN(
        n1811) );
  AOI211D1BWP12T U3067 ( .A1(n3941), .A2(n3444), .B(n1812), .C(n1811), .ZN(
        n3687) );
  INVD1BWP12T U3068 ( .I(n1821), .ZN(n3459) );
  TPND2D0BWP12T U3069 ( .A1(n3107), .A2(n3447), .ZN(n1813) );
  TPOAI21D0BWP12T U3070 ( .A1(n2916), .A2(n3459), .B(n1813), .ZN(n1815) );
  INVD1BWP12T U3071 ( .I(n1822), .ZN(n3470) );
  OAI22D1BWP12T U3072 ( .A1(n3945), .A2(n3470), .B1(n3471), .B2(n3813), .ZN(
        n1814) );
  NR2D1BWP12T U3073 ( .A1(n1815), .A2(n1814), .ZN(n3289) );
  OAI22D0BWP12T U3074 ( .A1(n3687), .A2(n3818), .B1(n3289), .B2(n4032), .ZN(
        n1820) );
  INVD1BWP12T U3075 ( .I(n1816), .ZN(n3290) );
  OAI21D0BWP12T U3076 ( .A1(n3290), .A2(n3758), .B(n3756), .ZN(n1819) );
  INVD1BWP12T U3077 ( .I(n3694), .ZN(n4789) );
  AOI21D0BWP12T U3078 ( .A1(n4707), .A2(n4789), .B(n4158), .ZN(n1817) );
  OAI22D1BWP12T U3079 ( .A1(n1820), .A2(n1819), .B1(n1818), .B2(n1817), .ZN(
        n4841) );
  INVD0BWP12T U3080 ( .I(n3849), .ZN(n3716) );
  INVD1BWP12T U3081 ( .I(n3968), .ZN(n3761) );
  NR2XD0BWP12T U3082 ( .A1(n3292), .A2(n4743), .ZN(n4606) );
  AOI21D0BWP12T U3083 ( .A1(n4573), .A2(n4606), .B(n4605), .ZN(n1826) );
  INVD1BWP12T U3084 ( .I(n3444), .ZN(n3952) );
  AOI22D1BWP12T U3085 ( .A1(n3125), .A2(n3952), .B1(n3953), .B2(n953), .ZN(
        n3703) );
  INVD1BWP12T U3086 ( .I(n3703), .ZN(n1824) );
  AOI22D1BWP12T U3087 ( .A1(n3122), .A2(n3458), .B1(n3954), .B2(n3701), .ZN(
        n3702) );
  INVD1BWP12T U3088 ( .I(n3702), .ZN(n1823) );
  NR3XD0BWP12T U3089 ( .A1(n1824), .A2(n1823), .A3(n4611), .ZN(n1825) );
  AOI211D1BWP12T U3090 ( .A1(n3761), .A2(n3291), .B(n1826), .C(n1825), .ZN(
        n4597) );
  MUX2ND0BWP12T U3091 ( .I0(n5045), .I1(n5044), .S(n4762), .ZN(n1827) );
  TPND2D0BWP12T U3092 ( .A1(n1827), .A2(n5081), .ZN(n1828) );
  MUX2NXD0BWP12T U3093 ( .I0(n1828), .I1(n5048), .S(n4637), .ZN(n1840) );
  ND2XD0BWP12T U3094 ( .A1(n1829), .A2(n1833), .ZN(n1832) );
  INVD1BWP12T U3095 ( .I(n4448), .ZN(n1834) );
  INR2D1BWP12T U3096 ( .A1(n1830), .B1(n1834), .ZN(n1831) );
  INR2D1BWP12T U3097 ( .A1(n1832), .B1(n1831), .ZN(n1836) );
  CKND2D1BWP12T U3098 ( .A1(n1834), .A2(n1833), .ZN(n1835) );
  ND2D1BWP12T U3099 ( .A1(n1836), .A2(n1835), .ZN(n4428) );
  CKND2D1BWP12T U3100 ( .A1(n4428), .A2(n5078), .ZN(n1839) );
  OAI21D1BWP12T U3101 ( .A1(n4923), .A2(n5083), .B(n5081), .ZN(n1837) );
  ND2D1BWP12T U3102 ( .A1(n4762), .A2(n1837), .ZN(n1838) );
  ND3D1BWP12T U3103 ( .A1(n1840), .A2(n1839), .A3(n1838), .ZN(n1841) );
  AOI21D1BWP12T U3104 ( .A1(n4597), .A2(n4167), .B(n1841), .ZN(n1842) );
  OAI21D1BWP12T U3105 ( .A1(n4544), .A2(n3716), .B(n1842), .ZN(n1843) );
  AO21D1BWP12T U3106 ( .A1(n5094), .A2(n4841), .B(n1843), .Z(n1850) );
  ND2XD0BWP12T U3107 ( .A1(n4411), .A2(n5088), .ZN(n1848) );
  XOR2XD1BWP12T U3108 ( .A1(n4353), .A2(n1845), .Z(n4327) );
  INVD1BWP12T U3109 ( .I(n3982), .ZN(n4847) );
  OAI21D1BWP12T U3110 ( .A1(n1846), .A2(n3566), .B(n4847), .ZN(n4899) );
  AOI22D1BWP12T U3111 ( .A1(n4327), .A2(n5090), .B1(n4899), .B2(n5099), .ZN(
        n1847) );
  CKND2D1BWP12T U3112 ( .A1(n1848), .A2(n1847), .ZN(n1849) );
  NR2D1BWP12T U3113 ( .A1(n1850), .A2(n1849), .ZN(n1851) );
  ND2D1BWP12T U3114 ( .A1(n1852), .A2(n1851), .ZN(n1853) );
  TPAOI21D2BWP12T U3115 ( .A1(n5093), .A2(n4980), .B(n1853), .ZN(n1854) );
  XNR2XD4BWP12T U3116 ( .A1(n4628), .A2(n4916), .ZN(n1895) );
  BUFFXD8BWP12T U3117 ( .I(n1894), .Z(n1982) );
  XNR2XD4BWP12T U3118 ( .A1(n341), .A2(n1856), .ZN(n1871) );
  TPND2D3BWP12T U3119 ( .A1(n1871), .A2(n1870), .ZN(n1857) );
  TPOAI21D4BWP12T U3120 ( .A1(n1895), .A2(n1982), .B(n1857), .ZN(n1880) );
  INVD4BWP12T U3121 ( .I(a[27]), .ZN(n2631) );
  INVD8BWP12T U3122 ( .I(n4908), .ZN(n1858) );
  XNR2XD8BWP12T U3123 ( .A1(n2631), .A2(n1858), .ZN(n2686) );
  INR2D8BWP12T U3124 ( .A1(n4316), .B1(n2686), .ZN(n1863) );
  CKND2D2BWP12T U3125 ( .A1(n1859), .A2(n1881), .ZN(n1862) );
  INVD1BWP12T U3126 ( .I(n4907), .ZN(n1860) );
  XOR2D2BWP12T U3127 ( .A1(n2169), .A2(n1860), .Z(n1861) );
  XNR2XD4BWP12T U3128 ( .A1(n4916), .A2(n4907), .ZN(n2678) );
  ND2XD8BWP12T U3129 ( .A1(n1861), .A2(n2678), .ZN(n2676) );
  TPOAI22D2BWP12T U3130 ( .A1(n1896), .A2(n2676), .B1(n1929), .B2(n2678), .ZN(
        n1879) );
  ND2D1BWP12T U3131 ( .A1(n1863), .A2(n1880), .ZN(n1864) );
  TPND2D2BWP12T U3132 ( .A1(n1865), .A2(n1864), .ZN(n1917) );
  INVD8BWP12T U3133 ( .I(n4909), .ZN(n2017) );
  XNR2D2BWP12T U3134 ( .A1(n2017), .A2(n4908), .ZN(n1866) );
  CKND2D4BWP12T U3135 ( .A1(n1866), .A2(n2686), .ZN(n2685) );
  CKND3BWP12T U3136 ( .I(n2017), .ZN(n1867) );
  TPND2D2BWP12T U3137 ( .A1(n1868), .A2(n1867), .ZN(n1869) );
  TPOAI22D4BWP12T U3138 ( .A1(n2685), .A2(n2017), .B1(n1869), .B2(n2686), .ZN(
        n2044) );
  ND2D4BWP12T U3139 ( .A1(n2035), .A2(n1870), .ZN(n1874) );
  INVD1BWP12T U3140 ( .I(n1894), .ZN(n1872) );
  CKND2D2BWP12T U3141 ( .A1(n1872), .A2(n1871), .ZN(n1873) );
  XNR2D1BWP12T U3142 ( .A1(n2098), .A2(n4914), .ZN(n2037) );
  XNR3XD4BWP12T U3143 ( .A1(n2044), .A2(n2043), .A3(n2041), .ZN(n1918) );
  XNR2XD8BWP12T U3144 ( .A1(n2623), .A2(n2688), .ZN(n1909) );
  XNR2XD8BWP12T U3145 ( .A1(n2575), .A2(n2688), .ZN(n2000) );
  TPOAI22D2BWP12T U3146 ( .A1(n1909), .A2(n2691), .B1(n2000), .B2(n2689), .ZN(
        n1997) );
  CKND3BWP12T U3147 ( .I(n1997), .ZN(n1876) );
  XNR2XD4BWP12T U3148 ( .A1(n2619), .A2(n2666), .ZN(n1925) );
  XNR2XD4BWP12T U3149 ( .A1(n4753), .A2(n2666), .ZN(n1999) );
  TPOAI22D4BWP12T U3150 ( .A1(n1925), .A2(n2669), .B1(n1999), .B2(n2667), .ZN(
        n1998) );
  XNR2D1BWP12T U3151 ( .A1(b[26]), .A2(n2742), .ZN(n1905) );
  OAI22D1BWP12T U3152 ( .A1(n2001), .A2(n2744), .B1(n1905), .B2(n2743), .ZN(
        n1996) );
  ND2D3BWP12T U3153 ( .A1(n1998), .A2(n1997), .ZN(n1877) );
  ND2D3BWP12T U3154 ( .A1(n1878), .A2(n1877), .ZN(n1916) );
  XOR3XD4BWP12T U3155 ( .A1(n1917), .A2(n1918), .A3(n1916), .Z(n1974) );
  XNR3XD4BWP12T U3156 ( .A1(n1881), .A2(n1880), .A3(n1879), .ZN(n1977) );
  INVD1P75BWP12T U3157 ( .I(n1977), .ZN(n1891) );
  XNR2D1BWP12T U3158 ( .A1(b[24]), .A2(n2746), .ZN(n1910) );
  OAI22D1BWP12T U3159 ( .A1(n1910), .A2(n2747), .B1(n1994), .B2(n2748), .ZN(
        n1979) );
  XNR2XD4BWP12T U3160 ( .A1(n2094), .A2(n4914), .ZN(n1931) );
  XNR2XD4BWP12T U3161 ( .A1(n341), .A2(n4914), .ZN(n2177) );
  TPOAI22D2BWP12T U3162 ( .A1(n1931), .A2(n2624), .B1(n306), .B2(n2177), .ZN(
        n2105) );
  OR2D2BWP12T U3163 ( .A1(n4316), .A2(n2631), .Z(n1886) );
  CKND3BWP12T U3164 ( .I(n4922), .ZN(n1882) );
  NR2XD2BWP12T U3165 ( .A1(n1883), .A2(n1882), .ZN(n1927) );
  TPNR2D2BWP12T U3166 ( .A1(n4699), .A2(n4922), .ZN(n1926) );
  OR2XD4BWP12T U3167 ( .A1(n1927), .A2(n1926), .Z(n2634) );
  CKND0BWP12T U3168 ( .I(n4922), .ZN(n1884) );
  TPOAI21D1BWP12T U3169 ( .A1(n1886), .A2(n2634), .B(n1885), .ZN(n2104) );
  XNR2XD4BWP12T U3170 ( .A1(n2098), .A2(n4924), .ZN(n1935) );
  TPOAI21D1BWP12T U3171 ( .A1(n2105), .A2(n2104), .B(n2102), .ZN(n1888) );
  TPND2D1BWP12T U3172 ( .A1(n2104), .A2(n2105), .ZN(n1887) );
  NR2D1BWP12T U3173 ( .A1(n1979), .A2(n330), .ZN(n1890) );
  ND2D1BWP12T U3174 ( .A1(n1979), .A2(n330), .ZN(n1889) );
  TPOAI21D1BWP12T U3175 ( .A1(n1891), .A2(n1890), .B(n1889), .ZN(n1975) );
  XNR2XD4BWP12T U3176 ( .A1(n4764), .A2(n4906), .ZN(n1980) );
  XNR2XD2BWP12T U3177 ( .A1(n279), .A2(n5014), .ZN(n1981) );
  TPNR2D1BWP12T U3178 ( .A1(n1981), .A2(n2740), .ZN(n1893) );
  XNR2XD2BWP12T U3179 ( .A1(n2226), .A2(n5014), .ZN(n1936) );
  TPNR2D2BWP12T U3180 ( .A1(n1936), .A2(n2739), .ZN(n1892) );
  TPNR2D2BWP12T U3181 ( .A1(n1893), .A2(n1892), .ZN(n1966) );
  IND2XD2BWP12T U3182 ( .A1(n293), .B1(n1966), .ZN(n1897) );
  XNR2XD2BWP12T U3183 ( .A1(n2071), .A2(n4916), .ZN(n1983) );
  BUFFXD6BWP12T U3184 ( .I(n1894), .Z(n2641) );
  TPND2D1BWP12T U3185 ( .A1(n1897), .A2(n1964), .ZN(n1900) );
  INVD1BWP12T U3186 ( .I(n1966), .ZN(n1898) );
  CKND2D2BWP12T U3187 ( .A1(n1898), .A2(n293), .ZN(n1899) );
  TPND2D2BWP12T U3188 ( .A1(n1900), .A2(n1899), .ZN(n1976) );
  NR2D1BWP12T U3189 ( .A1(n1975), .A2(n1976), .ZN(n1903) );
  INVD1BWP12T U3190 ( .I(n1976), .ZN(n1902) );
  INVD1BWP12T U3191 ( .I(n1975), .ZN(n1901) );
  TPOAI22D1BWP12T U3192 ( .A1(n1904), .A2(n2702), .B1(n1921), .B2(n2319), .ZN(
        n2052) );
  XNR2D1BWP12T U3193 ( .A1(n2591), .A2(n288), .ZN(n2039) );
  OAI22D1BWP12T U3194 ( .A1(n1906), .A2(n2648), .B1(n2647), .B2(n2039), .ZN(
        n2053) );
  XNR2D1BWP12T U3195 ( .A1(n4731), .A2(n2742), .ZN(n1922) );
  OAI22D1BWP12T U3196 ( .A1(n1922), .A2(n2743), .B1(n2744), .B2(n1905), .ZN(
        n2051) );
  XOR3XD4BWP12T U3197 ( .A1(n2052), .A2(n2053), .A3(n2051), .Z(n1945) );
  INVD1BWP12T U3198 ( .I(n1945), .ZN(n1914) );
  XNR2XD4BWP12T U3199 ( .A1(n2551), .A2(n2679), .ZN(n1953) );
  TPOAI22D2BWP12T U3200 ( .A1(n1937), .A2(n2682), .B1(n2680), .B2(n1953), .ZN(
        n2006) );
  XNR2XD4BWP12T U3201 ( .A1(n4726), .A2(n288), .ZN(n1993) );
  ND2D1BWP12T U3202 ( .A1(n2006), .A2(n2007), .ZN(n1908) );
  XNR2XD4BWP12T U3203 ( .A1(n4731), .A2(n2593), .ZN(n1995) );
  XNR2XD4BWP12T U3204 ( .A1(n4214), .A2(n4733), .ZN(n1940) );
  TPOAI22D2BWP12T U3205 ( .A1(n2646), .A2(n1995), .B1(n1940), .B2(n4257), .ZN(
        n2005) );
  XNR2XD4BWP12T U3206 ( .A1(n2575), .A2(n4924), .ZN(n2026) );
  TPOAI22D2BWP12T U3207 ( .A1(n2026), .A2(n2620), .B1(n1934), .B2(n2218), .ZN(
        n2033) );
  XNR2XD4BWP12T U3208 ( .A1(n4753), .A2(n2688), .ZN(n2027) );
  XNR2XD4BWP12T U3209 ( .A1(n2578), .A2(n2746), .ZN(n2028) );
  XOR3D2BWP12T U3210 ( .A1(n2033), .A2(n2034), .A3(n2029), .Z(n1947) );
  NR2D0BWP12T U3211 ( .A1(n1946), .A2(n1947), .ZN(n1913) );
  INVD1BWP12T U3212 ( .I(n1946), .ZN(n1912) );
  INVD1BWP12T U3213 ( .I(n1947), .ZN(n1911) );
  ND2D1BWP12T U3214 ( .A1(n1916), .A2(n1915), .ZN(n1920) );
  OAI22D1BWP12T U3215 ( .A1(n1921), .A2(n2702), .B1(n2592), .B2(n2704), .ZN(
        n2597) );
  XNR2D1BWP12T U3216 ( .A1(n2666), .A2(n4761), .ZN(n2546) );
  XNR2D1BWP12T U3217 ( .A1(n4733), .A2(n2742), .ZN(n2564) );
  OAI22D1BWP12T U3218 ( .A1(n1922), .A2(n2744), .B1(n2564), .B2(n2743), .ZN(
        n2596) );
  XNR2XD8BWP12T U3219 ( .A1(n4316), .A2(n4909), .ZN(n1923) );
  XNR2XD4BWP12T U3220 ( .A1(n1932), .A2(n4909), .ZN(n2038) );
  TPOAI22D2BWP12T U3221 ( .A1(n1923), .A2(n2685), .B1(n2686), .B2(n2038), .ZN(
        n2022) );
  TPOAI22D2BWP12T U3222 ( .A1(n1927), .A2(a[27]), .B1(n1926), .B2(n2631), .ZN(
        n2632) );
  CKND3BWP12T U3223 ( .I(n2631), .ZN(n1928) );
  XNR2XD4BWP12T U3224 ( .A1(b[3]), .A2(n1928), .ZN(n2018) );
  XNR2XD2BWP12T U3225 ( .A1(n4628), .A2(n4699), .ZN(n2019) );
  TPOAI22D2BWP12T U3226 ( .A1(n1929), .A2(n2676), .B1(n2019), .B2(n2678), .ZN(
        n2059) );
  XOR3XD4BWP12T U3227 ( .A1(n2022), .A2(n2023), .A3(n2021), .Z(n1949) );
  XNR2XD4BWP12T U3228 ( .A1(n1932), .A2(n3040), .ZN(n1951) );
  OAI22D1BWP12T U3229 ( .A1(n1935), .A2(n2621), .B1(n1934), .B2(n2620), .ZN(
        n1959) );
  INVD1BWP12T U3230 ( .I(n1950), .ZN(n1941) );
  XNR2XD4BWP12T U3231 ( .A1(n4764), .A2(n5014), .ZN(n2058) );
  NR2D2BWP12T U3232 ( .A1(n1937), .A2(n2680), .ZN(n1939) );
  XNR2D1BWP12T U3233 ( .A1(n4763), .A2(n2679), .ZN(n2057) );
  NR2D2BWP12T U3234 ( .A1(n2057), .A2(n2682), .ZN(n1938) );
  XOR3XD4BWP12T U3235 ( .A1(n2047), .A2(n2045), .A3(n2050), .Z(n1948) );
  IOA21D1BWP12T U3236 ( .A1(n1949), .A2(n1950), .B(n1943), .ZN(n2531) );
  XOR3XD4BWP12T U3237 ( .A1(n1947), .A2(n1946), .A3(n1945), .Z(n2061) );
  INVD1P75BWP12T U3238 ( .I(n2061), .ZN(n1973) );
  XNR2D1BWP12T U3239 ( .A1(n4316), .A2(n3040), .ZN(n1952) );
  OAI22D1BWP12T U3240 ( .A1(n1952), .A2(n2632), .B1(n1951), .B2(n2634), .ZN(
        n2087) );
  INVD1BWP12T U3241 ( .I(n2087), .ZN(n1957) );
  INVD2BWP12T U3242 ( .I(n2088), .ZN(n1956) );
  HA1D2BWP12T U3243 ( .A(n1955), .B(n1954), .CO(n1964), .S(n2086) );
  INVD2BWP12T U3244 ( .I(n2127), .ZN(n1963) );
  CKND2BWP12T U3245 ( .I(n2126), .ZN(n1962) );
  TPND2D2BWP12T U3246 ( .A1(n1963), .A2(n1962), .ZN(n1968) );
  INVD1P75BWP12T U3247 ( .I(n1964), .ZN(n1965) );
  XOR3XD4BWP12T U3248 ( .A1(n1967), .A2(n1966), .A3(n1965), .Z(n2125) );
  ND2D1BWP12T U3249 ( .A1(n2126), .A2(n2127), .ZN(n1969) );
  TPOAI21D1BWP12T U3250 ( .A1(n1973), .A2(n1972), .B(n1971), .ZN(n2526) );
  XNR3XD4BWP12T U3251 ( .A1(n1976), .A2(n1975), .A3(n1974), .ZN(n2121) );
  XOR3XD4BWP12T U3252 ( .A1(n1979), .A2(n1978), .A3(n1977), .Z(n2132) );
  XNR2XD4BWP12T U3253 ( .A1(n2226), .A2(n4906), .ZN(n2063) );
  TPOAI22D2BWP12T U3254 ( .A1(n1980), .A2(n2704), .B1(n2063), .B2(n2702), .ZN(
        n2085) );
  XNR2D2BWP12T U3255 ( .A1(n5014), .A2(n4761), .ZN(n2069) );
  CKND3BWP12T U3256 ( .I(n2084), .ZN(n1989) );
  ND2D1BWP12T U3257 ( .A1(n1985), .A2(n1984), .ZN(n1988) );
  XNR2D2BWP12T U3258 ( .A1(n2555), .A2(n4916), .ZN(n2073) );
  INVD2BWP12T U3259 ( .I(n1984), .ZN(n2181) );
  IND2D2BWP12T U3260 ( .A1(n1985), .B1(n2181), .ZN(n1986) );
  ND2D2BWP12T U3261 ( .A1(n2179), .A2(n1986), .ZN(n1987) );
  ND2D2BWP12T U3262 ( .A1(n1988), .A2(n1987), .ZN(n2083) );
  IOA21D2BWP12T U3263 ( .A1(n1990), .A2(n1989), .B(n2083), .ZN(n1992) );
  ND2D3BWP12T U3264 ( .A1(n1992), .A2(n1991), .ZN(n2133) );
  XNR2XD2BWP12T U3265 ( .A1(b[20]), .A2(n288), .ZN(n2064) );
  TPOAI22D2BWP12T U3266 ( .A1(n1993), .A2(n2647), .B1(n2648), .B2(n2064), .ZN(
        n2079) );
  XNR2XD1BWP12T U3267 ( .A1(b[26]), .A2(n2593), .ZN(n2091) );
  OAI22D1BWP12T U3268 ( .A1(n2091), .A2(n2646), .B1(n1995), .B2(n4257), .ZN(
        n2077) );
  RCOAI21D2BWP12T U3269 ( .A1(n2132), .A2(n2133), .B(n2134), .ZN(n2120) );
  TPND2D3BWP12T U3270 ( .A1(n2133), .A2(n2132), .ZN(n2119) );
  TPND2D2BWP12T U3271 ( .A1(n2120), .A2(n2119), .ZN(n2013) );
  INVD2BWP12T U3272 ( .I(n2013), .ZN(n2011) );
  XNR2XD2BWP12T U3273 ( .A1(n2623), .A2(n2666), .ZN(n2089) );
  TPOAI22D1BWP12T U3274 ( .A1(n2089), .A2(n2667), .B1(n1999), .B2(n2669), .ZN(
        n2108) );
  INVD1P25BWP12T U3275 ( .I(n2108), .ZN(n2003) );
  XNR2D1BWP12T U3276 ( .A1(n4740), .A2(n2742), .ZN(n2066) );
  OAI22D1BWP12T U3277 ( .A1(n2066), .A2(n2744), .B1(n2001), .B2(n2743), .ZN(
        n2106) );
  IOA21D2BWP12T U3278 ( .A1(n2003), .A2(n2002), .B(n2106), .ZN(n2004) );
  IOA21D2BWP12T U3279 ( .A1(n2108), .A2(n2107), .B(n2004), .ZN(n2131) );
  ND2D1BWP12T U3280 ( .A1(n2131), .A2(n2130), .ZN(n2008) );
  TPND2D2BWP12T U3281 ( .A1(n2011), .A2(n2010), .ZN(n2012) );
  ND2D1BWP12T U3282 ( .A1(n2122), .A2(n2013), .ZN(n2014) );
  TPND2D2BWP12T U3283 ( .A1(n2015), .A2(n2014), .ZN(n2527) );
  CKND1BWP12T U3284 ( .I(n4933), .ZN(n2016) );
  XNR2D2BWP12T U3285 ( .A1(n2017), .A2(n2016), .ZN(n2629) );
  TPNR2D3BWP12T U3286 ( .A1(n2629), .A2(n5082), .ZN(n2545) );
  XNR2XD2BWP12T U3287 ( .A1(n2071), .A2(n3040), .ZN(n2554) );
  TPOAI22D1BWP12T U3288 ( .A1(n2554), .A2(n2634), .B1(n2018), .B2(n2632), .ZN(
        n2542) );
  OAI22D1BWP12T U3289 ( .A1(n2019), .A2(n2676), .B1(n2678), .B2(n2550), .ZN(
        n2544) );
  XOR3XD4BWP12T U3290 ( .A1(n2545), .A2(n2542), .A3(n2544), .Z(n2538) );
  OR2D2BWP12T U3291 ( .A1(n2023), .A2(n2022), .Z(n2020) );
  CKND2D2BWP12T U3292 ( .A1(n2023), .A2(n284), .ZN(n2024) );
  CKND2D2BWP12T U3293 ( .A1(n2025), .A2(n2024), .ZN(n2539) );
  RCOAI22D1BWP12T U3294 ( .A1(n2552), .A2(n2691), .B1(n2689), .B2(n2027), .ZN(
        n2581) );
  XNR2D1BWP12T U3295 ( .A1(b[26]), .A2(n2746), .ZN(n2595) );
  XOR3XD4BWP12T U3296 ( .A1(n2538), .A2(n2539), .A3(n2537), .Z(n2569) );
  CKND0BWP12T U3297 ( .I(n2033), .ZN(n2031) );
  IOA21D1BWP12T U3298 ( .A1(n2034), .A2(n2033), .B(n2032), .ZN(n2588) );
  CKND3BWP12T U3299 ( .I(n2035), .ZN(n2036) );
  TPOAI22D2BWP12T U3300 ( .A1(n2036), .A2(n2641), .B1(n2643), .B2(n2549), .ZN(
        n2558) );
  TPOAI22D1BWP12T U3301 ( .A1(n2037), .A2(n305), .B1(n2576), .B2(n2624), .ZN(
        n2557) );
  XNR2D1BWP12T U3302 ( .A1(n3748), .A2(n4909), .ZN(n2556) );
  XOR3XD4BWP12T U3303 ( .A1(n2558), .A2(n2557), .A3(n2559), .Z(n2587) );
  XNR2D1BWP12T U3304 ( .A1(b[24]), .A2(n288), .ZN(n2579) );
  TPOAI22D1BWP12T U3305 ( .A1(n2579), .A2(n2647), .B1(n2039), .B2(n2648), .ZN(
        n2585) );
  XNR2D1BWP12T U3306 ( .A1(n4727), .A2(n2593), .ZN(n2594) );
  TPOAI22D1BWP12T U3307 ( .A1(n2040), .A2(n2646), .B1(n2594), .B2(n4257), .ZN(
        n2584) );
  OAI21D1BWP12T U3308 ( .A1(n281), .A2(n2044), .B(n290), .ZN(n2042) );
  IOA21D1BWP12T U3309 ( .A1(n2044), .A2(n281), .B(n2042), .ZN(n2583) );
  XOR3XD4BWP12T U3310 ( .A1(n2588), .A2(n2587), .A3(n2586), .Z(n2568) );
  INVD2P3BWP12T U3311 ( .I(n2045), .ZN(n2046) );
  TPOAI21D1BWP12T U3312 ( .A1(n2050), .A2(n2049), .B(n2048), .ZN(n2536) );
  CKND2D1BWP12T U3313 ( .A1(n2053), .A2(n2052), .ZN(n2054) );
  TPOAI21D1BWP12T U3314 ( .A1(n2056), .A2(n2055), .B(n2054), .ZN(n2535) );
  XNR2D1BWP12T U3315 ( .A1(n2226), .A2(n2679), .ZN(n2562) );
  OAI22D1BWP12T U3316 ( .A1(n2562), .A2(n2682), .B1(n2680), .B2(n2057), .ZN(
        n2604) );
  TPOAI22D2BWP12T U3317 ( .A1(n2563), .A2(n2739), .B1(n2740), .B2(n2058), .ZN(
        n2603) );
  HA1D2BWP12T U3318 ( .A(n2060), .B(n2059), .CO(n2602), .S(n2021) );
  XOR3XD4BWP12T U3319 ( .A1(n2569), .A2(n2568), .A3(n2567), .Z(n2528) );
  XNR3XD4BWP12T U3320 ( .A1(n2526), .A2(n2527), .A3(n2528), .ZN(n2605) );
  XOR3XD4BWP12T U3321 ( .A1(n2062), .A2(n326), .A3(n2061), .Z(n2197) );
  TPOAI22D1BWP12T U3322 ( .A1(n2242), .A2(n2702), .B1(n2063), .B2(n2319), .ZN(
        n2148) );
  XNR2XD4BWP12T U3323 ( .A1(n4764), .A2(n288), .ZN(n2227) );
  XNR2D1BWP12T U3324 ( .A1(n2591), .A2(n2742), .ZN(n2241) );
  OR2XD1BWP12T U3325 ( .A1(n2241), .A2(n2744), .Z(n2065) );
  OAI21D1BWP12T U3326 ( .A1(n2066), .A2(n2743), .B(n2065), .ZN(n2145) );
  OAI21D1BWP12T U3327 ( .A1(n2148), .A2(n2147), .B(n2145), .ZN(n2068) );
  XNR2D1BWP12T U3328 ( .A1(n2551), .A2(n5014), .ZN(n2152) );
  OAI22D1BWP12T U3329 ( .A1(n2740), .A2(n2152), .B1(n2069), .B2(n2739), .ZN(
        n2290) );
  XNR2XD2BWP12T U3330 ( .A1(n4726), .A2(n2746), .ZN(n2244) );
  OAI22D1BWP12T U3331 ( .A1(n2223), .A2(n306), .B1(n2178), .B2(n2624), .ZN(
        n2156) );
  TPOAI22D1BWP12T U3332 ( .A1(n2235), .A2(n2641), .B1(n2073), .B2(n2643), .ZN(
        n2155) );
  TPOAI21D1BWP12T U3333 ( .A1(n2290), .A2(n2074), .B(n2289), .ZN(n2076) );
  CKND2D2BWP12T U3334 ( .A1(n2290), .A2(n2074), .ZN(n2075) );
  TPND2D1BWP12T U3335 ( .A1(n2076), .A2(n2075), .ZN(n2304) );
  FA1D1BWP12T U3336 ( .A(n2079), .B(n2078), .CI(n2077), .CO(n2134), .S(n2302)
         );
  OAI21D1BWP12T U3337 ( .A1(n2303), .A2(n2304), .B(n2302), .ZN(n2082) );
  INVD1BWP12T U3338 ( .I(n2303), .ZN(n2080) );
  XOR3XD4BWP12T U3339 ( .A1(n2085), .A2(n2084), .A3(n2083), .Z(n2186) );
  XOR3XD4BWP12T U3340 ( .A1(n2088), .A2(n2087), .A3(n2086), .Z(n2187) );
  XNR2XD4BWP12T U3341 ( .A1(n2575), .A2(n2666), .ZN(n2165) );
  TPOAI22D1BWP12T U3342 ( .A1(n2165), .A2(n2667), .B1(n2089), .B2(n2669), .ZN(
        n2287) );
  TPOAI22D1BWP12T U3343 ( .A1(n2090), .A2(n2682), .B1(n2164), .B2(n2680), .ZN(
        n2288) );
  OAI22D1BWP12T U3344 ( .A1(n2166), .A2(n2646), .B1(n2091), .B2(n4257), .ZN(
        n2286) );
  OAI21D1BWP12T U3345 ( .A1(n2287), .A2(n2288), .B(n2286), .ZN(n2093) );
  ND2D1BWP12T U3346 ( .A1(n2287), .A2(n2288), .ZN(n2092) );
  CKND2D2BWP12T U3347 ( .A1(n2093), .A2(n2092), .ZN(n2188) );
  TPNR2D2BWP12T U3348 ( .A1(n2187), .A2(n2188), .ZN(n2113) );
  TPND2D2BWP12T U3349 ( .A1(n2187), .A2(n2188), .ZN(n2112) );
  TPOAI21D2BWP12T U3350 ( .A1(n2114), .A2(n2113), .B(n2112), .ZN(n2143) );
  XNR2XD4BWP12T U3351 ( .A1(n2094), .A2(n4924), .ZN(n2173) );
  TPOAI22D2BWP12T U3352 ( .A1(n2095), .A2(n2620), .B1(n2173), .B2(n2218), .ZN(
        n2150) );
  TPOAI22D2BWP12T U3353 ( .A1(n2153), .A2(n2676), .B1(n2097), .B2(n2678), .ZN(
        n2151) );
  OAI22D1BWP12T U3354 ( .A1(n2168), .A2(n2689), .B1(n2099), .B2(n2691), .ZN(
        n2149) );
  TPND2D2BWP12T U3355 ( .A1(n2101), .A2(n2100), .ZN(n2295) );
  INVD1BWP12T U3356 ( .I(n2102), .ZN(n2103) );
  XOR3D2BWP12T U3357 ( .A1(n2105), .A2(n2104), .A3(n2103), .Z(n2298) );
  IND2D2BWP12T U3358 ( .A1(n2295), .B1(n2298), .ZN(n2110) );
  XOR3D2BWP12T U3359 ( .A1(n2108), .A2(n2107), .A3(n2106), .Z(n2296) );
  CKND3BWP12T U3360 ( .I(n2298), .ZN(n2109) );
  CKND3BWP12T U3361 ( .I(n2144), .ZN(n2111) );
  OA21D1BWP12T U3362 ( .A1(n2114), .A2(n2113), .B(n2112), .Z(n2115) );
  INVD1BWP12T U3363 ( .I(n2197), .ZN(n2118) );
  INVD1BWP12T U3364 ( .I(n2198), .ZN(n2117) );
  TPND2D1BWP12T U3365 ( .A1(n2118), .A2(n2117), .ZN(n2123) );
  ND2D1BWP12T U3366 ( .A1(n2123), .A2(n2196), .ZN(n2124) );
  XOR3D2BWP12T U3367 ( .A1(n2127), .A2(n2126), .A3(n2125), .Z(n2140) );
  INVD1P75BWP12T U3368 ( .I(n2128), .ZN(n2129) );
  XNR3XD4BWP12T U3369 ( .A1(n2131), .A2(n2130), .A3(n2129), .ZN(n2141) );
  XNR3D2BWP12T U3370 ( .A1(n2134), .A2(n2133), .A3(n2132), .ZN(n2139) );
  OAI21D1BWP12T U3371 ( .A1(n2138), .A2(n2139), .B(n2137), .ZN(n2201) );
  XNR3XD4BWP12T U3372 ( .A1(n2141), .A2(n2140), .A3(n2139), .ZN(n2205) );
  XOR3XD4BWP12T U3373 ( .A1(n2144), .A2(n2143), .A3(n2142), .Z(n2206) );
  DCCKND4BWP12T U3374 ( .I(n2206), .ZN(n2193) );
  XNR3XD4BWP12T U3375 ( .A1(n2148), .A2(n2147), .A3(n2146), .ZN(n2277) );
  CKND3BWP12T U3376 ( .I(n2277), .ZN(n2163) );
  XOR3XD4BWP12T U3377 ( .A1(n2151), .A2(n2150), .A3(n2149), .Z(n2279) );
  TPOAI22D2BWP12T U3378 ( .A1(n2266), .A2(n2263), .B1(n2739), .B2(n2152), .ZN(
        n2231) );
  INVD1BWP12T U3379 ( .I(n2231), .ZN(n2158) );
  XNR2D1BWP12T U3380 ( .A1(n4316), .A2(n4699), .ZN(n2154) );
  TPOAI22D1BWP12T U3381 ( .A1(n2676), .A2(n2154), .B1(n2153), .B2(n2678), .ZN(
        n2232) );
  CKND3BWP12T U3382 ( .I(n2232), .ZN(n2157) );
  IOA21D2BWP12T U3383 ( .A1(n2158), .A2(n2157), .B(n2230), .ZN(n2160) );
  ND2XD1BWP12T U3384 ( .A1(n2232), .A2(n2231), .ZN(n2159) );
  TPND2D2BWP12T U3385 ( .A1(n2160), .A2(n2159), .ZN(n2278) );
  NR2D1BWP12T U3386 ( .A1(n2279), .A2(n2278), .ZN(n2162) );
  ND2D1BWP12T U3387 ( .A1(n2279), .A2(n2278), .ZN(n2161) );
  TPOAI21D2BWP12T U3388 ( .A1(n2163), .A2(n2162), .B(n2161), .ZN(n2209) );
  XNR2XD4BWP12T U3389 ( .A1(n2623), .A2(n2679), .ZN(n2268) );
  TPOAI22D2BWP12T U3390 ( .A1(n2268), .A2(n2680), .B1(n2164), .B2(n2682), .ZN(
        n2273) );
  TPOAI22D2BWP12T U3391 ( .A1(n2238), .A2(n2667), .B1(n2165), .B2(n2669), .ZN(
        n2272) );
  TPOAI22D2BWP12T U3392 ( .A1(n2234), .A2(n2689), .B1(n2168), .B2(n2691), .ZN(
        n2214) );
  CKND2D2BWP12T U3393 ( .A1(n2170), .A2(n4699), .ZN(n2171) );
  TPOAI22D2BWP12T U3394 ( .A1(n2676), .A2(n4649), .B1(n2171), .B2(n2678), .ZN(
        n2216) );
  XNR2D2BWP12T U3395 ( .A1(n341), .A2(n4924), .ZN(n2221) );
  TPNR2D1BWP12T U3396 ( .A1(n2216), .A2(n2215), .ZN(n2175) );
  ND2D1BWP12T U3397 ( .A1(n2215), .A2(n2216), .ZN(n2174) );
  XOR3XD4BWP12T U3398 ( .A1(n2181), .A2(n2180), .A3(n2179), .Z(n2212) );
  IND2D1BWP12T U3399 ( .A1(n2213), .B1(n2212), .ZN(n2182) );
  ND2D1BWP12T U3400 ( .A1(n2182), .A2(n2211), .ZN(n2184) );
  IND2D1BWP12T U3401 ( .A1(n2212), .B1(n2213), .ZN(n2183) );
  CKND2D2BWP12T U3402 ( .A1(n2184), .A2(n2183), .ZN(n2210) );
  INVD1BWP12T U3403 ( .I(n2210), .ZN(n2185) );
  IND2D2BWP12T U3404 ( .A1(n2209), .B1(n2185), .ZN(n2189) );
  CKND2D2BWP12T U3405 ( .A1(n2189), .A2(n2208), .ZN(n2191) );
  ND2D1BWP12T U3406 ( .A1(n2209), .A2(n2210), .ZN(n2190) );
  TPND2D2BWP12T U3407 ( .A1(n2191), .A2(n2190), .ZN(n2207) );
  INVD1P75BWP12T U3408 ( .I(n2207), .ZN(n2192) );
  TPND2D2BWP12T U3409 ( .A1(n2193), .A2(n2192), .ZN(n2195) );
  TPNR2D3BWP12T U3410 ( .A1(n2193), .A2(n2192), .ZN(n2194) );
  CKND1BWP12T U3411 ( .I(n2203), .ZN(n2200) );
  XOR3XD4BWP12T U3412 ( .A1(n2198), .A2(n2197), .A3(n2196), .Z(n2202) );
  IOA21D2BWP12T U3413 ( .A1(n2201), .A2(n2200), .B(n2199), .ZN(n2520) );
  NR2XD2BWP12T U3414 ( .A1(n2521), .A2(n2520), .ZN(n3424) );
  XOR3XD4BWP12T U3415 ( .A1(n2204), .A2(n2203), .A3(n2202), .Z(n2519) );
  XOR3XD4BWP12T U3416 ( .A1(n2207), .A2(n2206), .A3(n2205), .Z(n2309) );
  XOR3XD4BWP12T U3417 ( .A1(n2210), .A2(n2209), .A3(n2208), .Z(n2313) );
  XNR3XD4BWP12T U3418 ( .A1(n2216), .A2(n2215), .A3(n2214), .ZN(n2364) );
  INVD1BWP12T U3419 ( .I(n4316), .ZN(n2217) );
  TPNR2D1BWP12T U3420 ( .A1(n2678), .A2(n2217), .ZN(n2381) );
  TPOAI22D2BWP12T U3421 ( .A1(n2221), .A2(n2220), .B1(n2219), .B2(n2218), .ZN(
        n2379) );
  TPOAI22D2BWP12T U3422 ( .A1(n2223), .A2(n2624), .B1(n2222), .B2(n305), .ZN(
        n2382) );
  TPOAI21D1BWP12T U3423 ( .A1(n2381), .A2(n2379), .B(n2382), .ZN(n2225) );
  TPND2D2BWP12T U3424 ( .A1(n2225), .A2(n2224), .ZN(n2366) );
  XNR2D1BWP12T U3425 ( .A1(n2226), .A2(n288), .ZN(n2253) );
  TPOAI22D1BWP12T U3426 ( .A1(n2253), .A2(n2648), .B1(n2227), .B2(n2647), .ZN(
        n2363) );
  NR2D1BWP12T U3427 ( .A1(n2366), .A2(n2363), .ZN(n2229) );
  ND2D1BWP12T U3428 ( .A1(n2366), .A2(n2363), .ZN(n2228) );
  TPOAI22D1BWP12T U3429 ( .A1(n2234), .A2(n2691), .B1(n2233), .B2(n2689), .ZN(
        n2346) );
  OAI22D1BWP12T U3430 ( .A1(n2641), .A2(n2236), .B1(n2643), .B2(n2235), .ZN(
        n2344) );
  ND2D1BWP12T U3431 ( .A1(n2346), .A2(n2344), .ZN(n2240) );
  OAI22D1BWP12T U3432 ( .A1(n2238), .A2(n2669), .B1(n2237), .B2(n2667), .ZN(
        n2345) );
  ND2D3BWP12T U3433 ( .A1(n2240), .A2(n2239), .ZN(n2353) );
  ND2D1BWP12T U3434 ( .A1(n2354), .A2(n2353), .ZN(n2248) );
  TPOAI22D2BWP12T U3435 ( .A1(n2241), .A2(n2743), .B1(n2744), .B2(n2321), .ZN(
        n2284) );
  XNR2XD4BWP12T U3436 ( .A1(n4761), .A2(n2701), .ZN(n2320) );
  TPOAI22D2BWP12T U3437 ( .A1(n2320), .A2(n2702), .B1(n2242), .B2(n2704), .ZN(
        n2280) );
  XNR2XD2BWP12T U3438 ( .A1(n2243), .A2(n2746), .ZN(n2256) );
  OAI22D2BWP12T U3439 ( .A1(n2256), .A2(n2748), .B1(n2244), .B2(n2747), .ZN(
        n2245) );
  CKND3BWP12T U3440 ( .I(n2245), .ZN(n2281) );
  XOR3XD4BWP12T U3441 ( .A1(n2284), .A2(n2280), .A3(n2281), .Z(n2355) );
  ND2D1BWP12T U3442 ( .A1(n2248), .A2(n2247), .ZN(n2360) );
  ND2D1BWP12T U3443 ( .A1(n2249), .A2(n2360), .ZN(n2252) );
  INR2D1BWP12T U3444 ( .A1(n2362), .B1(n2361), .ZN(n2250) );
  INVD0BWP12T U3445 ( .I(n2250), .ZN(n2251) );
  TPND2D2BWP12T U3446 ( .A1(n2252), .A2(n2251), .ZN(n2314) );
  TPOAI22D1BWP12T U3447 ( .A1(n2254), .A2(n2648), .B1(n2647), .B2(n2253), .ZN(
        n2349) );
  TPOAI22D1BWP12T U3448 ( .A1(n2256), .A2(n2747), .B1(n2255), .B2(n2748), .ZN(
        n2348) );
  INVD1BWP12T U3449 ( .I(n2257), .ZN(n2259) );
  CKND0BWP12T U3450 ( .I(n2259), .ZN(n2262) );
  TPOAI22D2BWP12T U3451 ( .A1(n2268), .A2(n2682), .B1(n2267), .B2(n2680), .ZN(
        n2371) );
  HA1D2BWP12T U3452 ( .A(n2270), .B(n2269), .CO(n2370), .S(n2373) );
  FA1D2BWP12T U3453 ( .A(n2273), .B(n2272), .CI(n2271), .CO(n2211), .S(n2405)
         );
  TPOAI21D2BWP12T U3454 ( .A1(n2276), .A2(n2275), .B(n2274), .ZN(n2426) );
  XOR3D2BWP12T U3455 ( .A1(n2279), .A2(n2278), .A3(n2277), .Z(n2427) );
  CKND0BWP12T U3456 ( .I(n2281), .ZN(n2285) );
  CKND0BWP12T U3457 ( .I(n2284), .ZN(n2282) );
  IOA21D1BWP12T U3458 ( .A1(n2282), .A2(n2281), .B(n2280), .ZN(n2283) );
  XOR3D2BWP12T U3459 ( .A1(n2288), .A2(n2287), .A3(n2286), .Z(n2300) );
  XNR3XD4BWP12T U3460 ( .A1(n2291), .A2(n2290), .A3(n2289), .ZN(n2299) );
  OAI21D1BWP12T U3461 ( .A1(n2426), .A2(n2427), .B(n2424), .ZN(n2292) );
  IOA21D2BWP12T U3462 ( .A1(n2426), .A2(n2427), .B(n2292), .ZN(n2312) );
  ND2D3BWP12T U3463 ( .A1(n2313), .A2(n2314), .ZN(n2293) );
  TPND2D2BWP12T U3464 ( .A1(n2294), .A2(n2293), .ZN(n2310) );
  INVD1BWP12T U3465 ( .I(n2295), .ZN(n2297) );
  XOR3D2BWP12T U3466 ( .A1(n2298), .A2(n2297), .A3(n2296), .Z(n2317) );
  FA1D2BWP12T U3467 ( .A(n2301), .B(n2300), .CI(n2299), .CO(n2316), .S(n2424)
         );
  IND2D2BWP12T U3468 ( .A1(n2310), .B1(n2305), .ZN(n2306) );
  ND2D3BWP12T U3469 ( .A1(n2309), .A2(n2306), .ZN(n2308) );
  ND2XD4BWP12T U3470 ( .A1(n2308), .A2(n2307), .ZN(n2518) );
  XOR3XD4BWP12T U3471 ( .A1(n2311), .A2(n2310), .A3(n2309), .Z(n2517) );
  XOR3XD4BWP12T U3472 ( .A1(n2314), .A2(n2313), .A3(n2312), .Z(n2432) );
  TPOAI22D2BWP12T U3473 ( .A1(n2322), .A2(n2744), .B1(n2743), .B2(n2321), .ZN(
        n2368) );
  OAI22D1BWP12T U3474 ( .A1(n2324), .A2(n4257), .B1(n2323), .B2(n2646), .ZN(
        n2367) );
  NR2XD2BWP12T U3475 ( .A1(n2464), .A2(n2465), .ZN(n2337) );
  INVD3BWP12T U3476 ( .I(n2328), .ZN(n2332) );
  RCOAI21D2BWP12T U3477 ( .A1(n2331), .A2(n2332), .B(n2330), .ZN(n2334) );
  ND2D3BWP12T U3478 ( .A1(n2332), .A2(n2331), .ZN(n2333) );
  TPND2D3BWP12T U3479 ( .A1(n2334), .A2(n2333), .ZN(n2463) );
  CKND3BWP12T U3480 ( .I(n2465), .ZN(n2335) );
  TPOAI22D4BWP12T U3481 ( .A1(n2337), .A2(n2463), .B1(n2336), .B2(n2335), .ZN(
        n2454) );
  INVD1P75BWP12T U3482 ( .I(n2454), .ZN(n2359) );
  INVD1BWP12T U3483 ( .I(n2338), .ZN(n2339) );
  CKND2D1BWP12T U3484 ( .A1(n2340), .A2(n2339), .ZN(n2342) );
  NR2D1BWP12T U3485 ( .A1(n2339), .A2(n2340), .ZN(n2341) );
  XNR3XD4BWP12T U3486 ( .A1(n2346), .A2(n2345), .A3(n2344), .ZN(n2467) );
  FA1D2BWP12T U3487 ( .A(n2349), .B(n2348), .CI(n2347), .CO(n2403), .S(n2466)
         );
  IOA21D2BWP12T U3488 ( .A1(n2468), .A2(n2467), .B(n2466), .ZN(n2352) );
  INVD1BWP12T U3489 ( .I(n2467), .ZN(n2350) );
  IND2XD1BWP12T U3490 ( .A1(n2468), .B1(n2350), .ZN(n2351) );
  CKND2D2BWP12T U3491 ( .A1(n2352), .A2(n2351), .ZN(n2453) );
  INVD1P75BWP12T U3492 ( .I(n2353), .ZN(n2356) );
  XOR3XD4BWP12T U3493 ( .A1(n2356), .A2(n2355), .A3(n2354), .Z(n2451) );
  TPNR2D1BWP12T U3494 ( .A1(n2453), .A2(n2451), .ZN(n2358) );
  ND2D1BWP12T U3495 ( .A1(n2451), .A2(n2453), .ZN(n2357) );
  OAI21D2BWP12T U3496 ( .A1(n2359), .A2(n2358), .B(n2357), .ZN(n2397) );
  INVD1BWP12T U3497 ( .I(n2397), .ZN(n2392) );
  XNR3XD4BWP12T U3498 ( .A1(n2362), .A2(n2361), .A3(n2360), .ZN(n2398) );
  INVD1P75BWP12T U3499 ( .I(n2363), .ZN(n2365) );
  XOR3XD4BWP12T U3500 ( .A1(n2366), .A2(n2365), .A3(n2364), .Z(n2401) );
  FA1D2BWP12T U3501 ( .A(n2369), .B(n2368), .CI(n2367), .CO(n2387), .S(n2464)
         );
  INVD1P75BWP12T U3502 ( .I(n2387), .ZN(n2402) );
  FA1D2BWP12T U3503 ( .A(n2372), .B(n2371), .CI(n2370), .CO(n2404), .S(n2406)
         );
  INVD1BWP12T U3504 ( .I(n2406), .ZN(n2385) );
  INVD1BWP12T U3505 ( .I(n2377), .ZN(n2375) );
  INVD1BWP12T U3506 ( .I(n2378), .ZN(n2374) );
  IOA21D1BWP12T U3507 ( .A1(n2375), .A2(n2374), .B(n2373), .ZN(n2376) );
  IOA21D2BWP12T U3508 ( .A1(n2378), .A2(n2377), .B(n2376), .ZN(n2407) );
  INVD1BWP12T U3509 ( .I(n2379), .ZN(n2380) );
  XNR3XD4BWP12T U3510 ( .A1(n2382), .A2(n2381), .A3(n2380), .ZN(n2408) );
  TPNR2D1BWP12T U3511 ( .A1(n2407), .A2(n2408), .ZN(n2384) );
  ND2D1BWP12T U3512 ( .A1(n2407), .A2(n2408), .ZN(n2383) );
  TPOAI21D1BWP12T U3513 ( .A1(n2385), .A2(n2384), .B(n2383), .ZN(n2400) );
  IOA21D1BWP12T U3514 ( .A1(n2386), .A2(n2402), .B(n2400), .ZN(n2389) );
  ND2D1BWP12T U3515 ( .A1(n2401), .A2(n2387), .ZN(n2388) );
  CKND2D2BWP12T U3516 ( .A1(n2389), .A2(n2388), .ZN(n2399) );
  TPNR2D1BWP12T U3517 ( .A1(n2398), .A2(n2399), .ZN(n2391) );
  ND2D1BWP12T U3518 ( .A1(n2398), .A2(n2399), .ZN(n2390) );
  TPOAI21D2BWP12T U3519 ( .A1(n2392), .A2(n2391), .B(n2390), .ZN(n2433) );
  TPNR2D1BWP12T U3520 ( .A1(n2434), .A2(n2433), .ZN(n2393) );
  INVD1P75BWP12T U3521 ( .I(n2393), .ZN(n2394) );
  ND2D3BWP12T U3522 ( .A1(n2432), .A2(n2394), .ZN(n2396) );
  ND2D1BWP12T U3523 ( .A1(n2433), .A2(n2434), .ZN(n2395) );
  TPND2D2BWP12T U3524 ( .A1(n2396), .A2(n2395), .ZN(n2516) );
  TPNR2D3BWP12T U3525 ( .A1(n2517), .A2(n2516), .ZN(n3924) );
  XOR3XD4BWP12T U3526 ( .A1(n2399), .A2(n2398), .A3(n2397), .Z(n2448) );
  XNR3XD4BWP12T U3527 ( .A1(n2402), .A2(n2401), .A3(n2400), .ZN(n2472) );
  XOR3XD4BWP12T U3528 ( .A1(n2405), .A2(n2404), .A3(n2403), .Z(n2473) );
  OAI21D1BWP12T U3529 ( .A1(n2410), .A2(n338), .B(n2409), .ZN(n2413) );
  ND2D1BWP12T U3530 ( .A1(n338), .A2(n2410), .ZN(n2412) );
  TPNR2D1BWP12T U3531 ( .A1(n2489), .A2(n2490), .ZN(n2422) );
  INVD1BWP12T U3532 ( .I(n2414), .ZN(n2420) );
  INVD1BWP12T U3533 ( .I(n2418), .ZN(n2415) );
  NR2D1BWP12T U3534 ( .A1(n2415), .A2(n2416), .ZN(n2419) );
  CKND0BWP12T U3535 ( .I(n2416), .ZN(n2417) );
  OA22D2BWP12T U3536 ( .A1(n2420), .A2(n2419), .B1(n2418), .B2(n2417), .Z(
        n2487) );
  TPND2D1BWP12T U3537 ( .A1(n2489), .A2(n2490), .ZN(n2421) );
  TPOAI21D1BWP12T U3538 ( .A1(n2422), .A2(n2487), .B(n2421), .ZN(n2471) );
  OAI21D1BWP12T U3539 ( .A1(n2473), .A2(n2472), .B(n2471), .ZN(n2423) );
  IOA21D2BWP12T U3540 ( .A1(n2472), .A2(n2473), .B(n2423), .ZN(n2449) );
  CKND3BWP12T U3541 ( .I(n2424), .ZN(n2425) );
  XNR3XD4BWP12T U3542 ( .A1(n2426), .A2(n2427), .A3(n2425), .ZN(n2450) );
  IND2D2BWP12T U3543 ( .A1(n2449), .B1(n2429), .ZN(n2428) );
  ND2D2BWP12T U3544 ( .A1(n2448), .A2(n2428), .ZN(n2431) );
  ND2D1BWP12T U3545 ( .A1(n2449), .A2(n2450), .ZN(n2430) );
  TPND2D2BWP12T U3546 ( .A1(n2431), .A2(n2430), .ZN(n2514) );
  INVD1P75BWP12T U3547 ( .I(n2514), .ZN(n2435) );
  XOR3XD4BWP12T U3548 ( .A1(n2434), .A2(n2433), .A3(n2432), .Z(n2515) );
  INR2D4BWP12T U3549 ( .A1(n2435), .B1(n327), .ZN(n3922) );
  TPNR2D1BWP12T U3550 ( .A1(n3924), .A2(n3922), .ZN(n3419) );
  CKND2D1BWP12T U3551 ( .A1(n2523), .A2(n3419), .ZN(n2525) );
  TPOAI21D1BWP12T U3552 ( .A1(n3084), .A2(n2437), .B(n2436), .ZN(n2440) );
  TPAOI21D2BWP12T U3553 ( .A1(n2440), .A2(n2439), .B(n2438), .ZN(n4293) );
  TPNR2D2BWP12T U3554 ( .A1(n304), .A2(n3867), .ZN(n2445) );
  TPND2D1BWP12T U3555 ( .A1(n2445), .A2(n3865), .ZN(n2447) );
  TPOAI21D1BWP12T U3556 ( .A1(n2443), .A2(n2442), .B(n2441), .ZN(n2444) );
  TPAOI21D2BWP12T U3557 ( .A1(n3864), .A2(n2445), .B(n2444), .ZN(n2446) );
  XOR3XD4BWP12T U3558 ( .A1(n2450), .A2(n2449), .A3(n2448), .Z(n2511) );
  CKND3BWP12T U3559 ( .I(n2451), .ZN(n2452) );
  XNR3XD4BWP12T U3560 ( .A1(n2454), .A2(n2453), .A3(n2452), .ZN(n2507) );
  INVD1BWP12T U3561 ( .I(n2459), .ZN(n2455) );
  ND2D1BWP12T U3562 ( .A1(n2455), .A2(n2458), .ZN(n2457) );
  ND2D1BWP12T U3563 ( .A1(n2457), .A2(n2456), .ZN(n2462) );
  ND2D1BWP12T U3564 ( .A1(n2460), .A2(n2459), .ZN(n2461) );
  AN2XD2BWP12T U3565 ( .A1(n2462), .A2(n2461), .Z(n2477) );
  XNR3XD4BWP12T U3566 ( .A1(n2465), .A2(n2464), .A3(n2463), .ZN(n2478) );
  XOR3D2BWP12T U3567 ( .A1(n2468), .A2(n2467), .A3(n2466), .Z(n2479) );
  NR2D2BWP12T U3568 ( .A1(n2478), .A2(n2479), .ZN(n2470) );
  CKND2D2BWP12T U3569 ( .A1(n2478), .A2(n2479), .ZN(n2469) );
  INVD1BWP12T U3570 ( .I(n2506), .ZN(n2475) );
  XOR3XD4BWP12T U3571 ( .A1(n2473), .A2(n2472), .A3(n2471), .Z(n2505) );
  IOA21D0BWP12T U3572 ( .A1(n2475), .A2(n2474), .B(n2505), .ZN(n2476) );
  IOA21D2BWP12T U3573 ( .A1(n2507), .A2(n282), .B(n2476), .ZN(n2510) );
  XNR3XD4BWP12T U3574 ( .A1(n2507), .A2(n282), .A3(n2505), .ZN(n2492) );
  XNR3XD4BWP12T U3575 ( .A1(n2479), .A2(n2478), .A3(n2477), .ZN(n2493) );
  CKND2BWP12T U3576 ( .I(n2484), .ZN(n2481) );
  ND2D1BWP12T U3577 ( .A1(n315), .A2(n343), .ZN(n2485) );
  INVD1P75BWP12T U3578 ( .I(n2487), .ZN(n2488) );
  XOR3XD4BWP12T U3579 ( .A1(n2490), .A2(n2489), .A3(n2488), .Z(n2494) );
  OR2D2BWP12T U3580 ( .A1(n2495), .A2(n2494), .Z(n2491) );
  RCAOI21D4BWP12T U3581 ( .A1(n2493), .A2(n2491), .B(n352), .ZN(n2508) );
  ND2XD4BWP12T U3582 ( .A1(n2492), .A2(n2508), .ZN(n3797) );
  XNR3XD4BWP12T U3583 ( .A1(n2495), .A2(n2494), .A3(n2493), .ZN(n2503) );
  OR2XD1BWP12T U3584 ( .A1(n2499), .A2(n333), .Z(n2496) );
  ND2D1BWP12T U3585 ( .A1(n2496), .A2(n2497), .ZN(n2501) );
  CKND2D0BWP12T U3586 ( .A1(n2499), .A2(n334), .ZN(n2500) );
  TPND2D2BWP12T U3587 ( .A1(n2501), .A2(n2500), .ZN(n2504) );
  INVD1P75BWP12T U3588 ( .I(n2504), .ZN(n2502) );
  ND2D3BWP12T U3589 ( .A1(n2503), .A2(n2502), .ZN(n3795) );
  TPNR2D2BWP12T U3590 ( .A1(n273), .A2(n3667), .ZN(n2513) );
  XNR3XD4BWP12T U3591 ( .A1(n2507), .A2(n2506), .A3(n2505), .ZN(n2509) );
  RCAOI21D2BWP12T U3592 ( .A1(n3794), .A2(n3797), .B(n3798), .ZN(n3669) );
  TPAOI21D2BWP12T U3593 ( .A1(n3796), .A2(n2513), .B(n2512), .ZN(n3923) );
  TPOAI21D2BWP12T U3594 ( .A1(n3924), .A2(n3921), .B(n3925), .ZN(n3420) );
  TPOAI21D2BWP12T U3595 ( .A1(n3424), .A2(n3549), .B(n3425), .ZN(n2522) );
  TPAOI21D2BWP12T U3596 ( .A1(n3420), .A2(n2523), .B(n2522), .ZN(n2524) );
  TPOAI21D1BWP12T U3597 ( .A1(n2525), .A2(n3923), .B(n2524), .ZN(n2847) );
  ND2D1BWP12T U3598 ( .A1(n331), .A2(n301), .ZN(n2530) );
  OAI21D1BWP12T U3599 ( .A1(n301), .A2(n331), .B(n2526), .ZN(n2529) );
  FA1D2BWP12T U3600 ( .A(n2533), .B(n2532), .CI(n2531), .CO(n2763), .S(n2572)
         );
  FA1D2BWP12T U3601 ( .A(n2536), .B(n2535), .CI(n2534), .CO(n2762), .S(n2567)
         );
  ND2D1BWP12T U3602 ( .A1(n2539), .A2(n2538), .ZN(n2541) );
  OAI21D1BWP12T U3603 ( .A1(n2539), .A2(n2538), .B(n2537), .ZN(n2540) );
  ND2D1BWP12T U3604 ( .A1(n2541), .A2(n2540), .ZN(n2618) );
  IOA21D1BWP12T U3605 ( .A1(n2545), .A2(n2544), .B(n2543), .ZN(n2655) );
  XNR2D1BWP12T U3606 ( .A1(n279), .A2(n2666), .ZN(n2668) );
  OAI22D1BWP12T U3607 ( .A1(n2546), .A2(n2667), .B1(n2668), .B2(n2669), .ZN(
        n2654) );
  IND2D1BWP12T U3608 ( .A1(n4258), .B1(n848), .ZN(n2548) );
  XOR2XD1BWP12T U3609 ( .A1(n4933), .A2(n848), .Z(n2547) );
  XNR2D1BWP12T U3610 ( .A1(n4765), .A2(n4916), .ZN(n2642) );
  OAI22D1BWP12T U3611 ( .A1(n2642), .A2(n2643), .B1(n2549), .B2(n2641), .ZN(
        n2706) );
  OAI22D1BWP12T U3612 ( .A1(n2677), .A2(n2678), .B1(n2550), .B2(n2676), .ZN(
        n2709) );
  XOR3D2BWP12T U3613 ( .A1(n2708), .A2(n2706), .A3(n2709), .Z(n2653) );
  OAI22D1BWP12T U3614 ( .A1(n2552), .A2(n2689), .B1(n2690), .B2(n2691), .ZN(
        n2712) );
  XNR2D1BWP12T U3615 ( .A1(n4258), .A2(n848), .ZN(n2553) );
  XNR2D1BWP12T U3616 ( .A1(n848), .A2(n4738), .ZN(n2628) );
  OAI22D1BWP12T U3617 ( .A1(n2553), .A2(n2627), .B1(n2628), .B2(n2629), .ZN(
        n2711) );
  TPOAI22D1BWP12T U3618 ( .A1(n2554), .A2(n2632), .B1(n2633), .B2(n2634), .ZN(
        n2665) );
  XNR2D1BWP12T U3619 ( .A1(n2555), .A2(n4909), .ZN(n2684) );
  OAI22D1BWP12T U3620 ( .A1(n2684), .A2(n2686), .B1(n2556), .B2(n2685), .ZN(
        n2664) );
  OAI21D1BWP12T U3621 ( .A1(n2559), .A2(n2558), .B(n2557), .ZN(n2561) );
  ND2D1BWP12T U3622 ( .A1(n2559), .A2(n2558), .ZN(n2560) );
  ND2D1BWP12T U3623 ( .A1(n2561), .A2(n2560), .ZN(n2731) );
  XNR2D1BWP12T U3624 ( .A1(n2679), .A2(n4764), .ZN(n2681) );
  OAI22D1BWP12T U3625 ( .A1(n2562), .A2(n2680), .B1(n2682), .B2(n2681), .ZN(
        n2738) );
  OAI22D1BWP12T U3626 ( .A1(n2740), .A2(n2563), .B1(n2741), .B2(n2739), .ZN(
        n2737) );
  XNR2D1BWP12T U3627 ( .A1(n4730), .A2(n2742), .ZN(n2745) );
  OAI22D1BWP12T U3628 ( .A1(n2564), .A2(n2744), .B1(n2745), .B2(n2743), .ZN(
        n2736) );
  INVD1BWP12T U3629 ( .I(n2568), .ZN(n2565) );
  IND2XD1BWP12T U3630 ( .A1(n2569), .B1(n2565), .ZN(n2566) );
  ND2D1BWP12T U3631 ( .A1(n2567), .A2(n2566), .ZN(n2571) );
  ND2D1BWP12T U3632 ( .A1(n2569), .A2(n2568), .ZN(n2570) );
  ND2D1BWP12T U3633 ( .A1(n2571), .A2(n2570), .ZN(n2726) );
  FA1D2BWP12T U3634 ( .A(n2574), .B(n2573), .CI(n2572), .CO(n2725), .S(n1944)
         );
  XNR2D1BWP12T U3635 ( .A1(n2575), .A2(n4914), .ZN(n2626) );
  OAI22D1BWP12T U3636 ( .A1(n2576), .A2(n306), .B1(n2626), .B2(n2624), .ZN(
        n2675) );
  XNR2XD0BWP12T U3637 ( .A1(n4753), .A2(n4924), .ZN(n2622) );
  TPOAI22D1BWP12T U3638 ( .A1(n2577), .A2(n2621), .B1(n2622), .B2(n2620), .ZN(
        n2674) );
  XNR2D1BWP12T U3639 ( .A1(n4739), .A2(n288), .ZN(n2649) );
  FA1D2BWP12T U3640 ( .A(n2582), .B(n2581), .CI(n2580), .CO(n2660), .S(n2537)
         );
  FA1D2BWP12T U3641 ( .A(n2585), .B(n2584), .CI(n2583), .CO(n2659), .S(n2586)
         );
  ND2D1BWP12T U3642 ( .A1(n2588), .A2(n2587), .ZN(n2589) );
  ND2D1BWP12T U3643 ( .A1(n2590), .A2(n2589), .ZN(n2759) );
  OAI22D1BWP12T U3644 ( .A1(n2592), .A2(n2702), .B1(n2703), .B2(n2704), .ZN(
        n2735) );
  OAI22D1BWP12T U3645 ( .A1(n2594), .A2(n2646), .B1(n2645), .B2(n4257), .ZN(
        n2734) );
  XNR2D1BWP12T U3646 ( .A1(n4731), .A2(n2746), .ZN(n2749) );
  OAI22D1BWP12T U3647 ( .A1(n2595), .A2(n2748), .B1(n2749), .B2(n2747), .ZN(
        n2733) );
  CKND1BWP12T U3648 ( .I(n2596), .ZN(n2601) );
  NR2D1BWP12T U3649 ( .A1(n2598), .A2(n2597), .ZN(n2600) );
  CKND2D1BWP12T U3650 ( .A1(n2598), .A2(n2597), .ZN(n2599) );
  OAI21D1BWP12T U3651 ( .A1(n2601), .A2(n2600), .B(n2599), .ZN(n2717) );
  FA1D2BWP12T U3652 ( .A(n2604), .B(n2603), .CI(n2602), .CO(n2716), .S(n2534)
         );
  XNR3XD4BWP12T U3653 ( .A1(n2726), .A2(n2725), .A3(n2727), .ZN(n2774) );
  XNR3XD4BWP12T U3654 ( .A1(n2770), .A2(n2771), .A3(n2774), .ZN(n2614) );
  CKBD1BWP12T U3655 ( .I(n2605), .Z(n2608) );
  INVD1BWP12T U3656 ( .I(n2606), .ZN(n2610) );
  OR2D2BWP12T U3657 ( .A1(n2608), .A2(n2607), .Z(n2609) );
  TPOAI21D2BWP12T U3658 ( .A1(n2611), .A2(n2610), .B(n2609), .ZN(n2613) );
  TPNR2D3BWP12T U3659 ( .A1(n2614), .A2(n2613), .ZN(n2612) );
  INVD2BWP12T U3660 ( .I(n2612), .ZN(n2845) );
  INVD1BWP12T U3661 ( .I(n2844), .ZN(n2615) );
  TPAOI21D1BWP12T U3662 ( .A1(n2847), .A2(n2845), .B(n2615), .ZN(n2780) );
  FA1D2BWP12T U3663 ( .A(n2618), .B(n2617), .CI(n2616), .CO(n2724), .S(n2761)
         );
  OAI22D1BWP12T U3664 ( .A1(n2630), .A2(n2629), .B1(n2628), .B2(n2627), .ZN(
        n2637) );
  CKXOR2D0BWP12T U3665 ( .A1(n4748), .A2(n2631), .Z(n2635) );
  OAI22D1BWP12T U3666 ( .A1(n2635), .A2(n2634), .B1(n2633), .B2(n2632), .ZN(
        n2636) );
  XNR2XD1BWP12T U3667 ( .A1(n2637), .A2(n2636), .ZN(n2638) );
  XOR3D1BWP12T U3668 ( .A1(n2640), .A2(n2639), .A3(n2638), .Z(n2658) );
  XNR2D1BWP12T U3669 ( .A1(n3296), .A2(n4916), .ZN(n2644) );
  OAI22D1BWP12T U3670 ( .A1(n2644), .A2(n2643), .B1(n2642), .B2(n2641), .ZN(
        n2652) );
  AO21D1BWP12T U3671 ( .A1(n2646), .A2(n4257), .B(n2645), .Z(n2651) );
  XOR3D1BWP12T U3672 ( .A1(n2652), .A2(n2651), .A3(n2650), .Z(n2657) );
  FA1D2BWP12T U3673 ( .A(n2655), .B(n2654), .CI(n2653), .CO(n2656), .S(n2617)
         );
  XOR3D2BWP12T U3674 ( .A1(n2658), .A2(n2657), .A3(n2656), .Z(n2663) );
  FA1D2BWP12T U3675 ( .A(n2661), .B(n2660), .CI(n2659), .CO(n2662), .S(n2760)
         );
  XOR2D2BWP12T U3676 ( .A1(n2663), .A2(n2662), .Z(n2723) );
  HA1D1BWP12T U3677 ( .A(n2665), .B(n2664), .CO(n2672), .S(n2710) );
  FA1D2BWP12T U3678 ( .A(n2674), .B(n2675), .CI(n2673), .CO(n2699), .S(n2661)
         );
  XNR2D1BWP12T U3679 ( .A1(n5053), .A2(n2679), .ZN(n2683) );
  OAI22D1BWP12T U3680 ( .A1(n2683), .A2(n2682), .B1(n2681), .B2(n2680), .ZN(
        n2696) );
  OAI22D1BWP12T U3681 ( .A1(n2692), .A2(n2691), .B1(n2690), .B2(n2689), .ZN(
        n2693) );
  OAI22D1BWP12T U3682 ( .A1(n2705), .A2(n2704), .B1(n2703), .B2(n2702), .ZN(
        n2715) );
  IOA21D1BWP12T U3683 ( .A1(n2709), .A2(n2708), .B(n2707), .ZN(n2714) );
  FA1D1BWP12T U3684 ( .A(n2712), .B(n2711), .CI(n2710), .CO(n2713), .S(n2732)
         );
  XOR3D1BWP12T U3685 ( .A1(n2715), .A2(n2714), .A3(n2713), .Z(n2720) );
  XOR3XD4BWP12T U3686 ( .A1(n2721), .A2(n2720), .A3(n2719), .Z(n2722) );
  XOR3XD4BWP12T U3687 ( .A1(n2724), .A2(n2723), .A3(n2722), .Z(n2769) );
  FA1D2BWP12T U3688 ( .A(n2732), .B(n2731), .CI(n2730), .CO(n2757), .S(n2616)
         );
  FA1D0BWP12T U3689 ( .A(n2735), .B(n2734), .CI(n2733), .CO(n2755), .S(n2718)
         );
  FA1D1BWP12T U3690 ( .A(n2738), .B(n2737), .CI(n2736), .CO(n2754), .S(n2730)
         );
  XOR3D1BWP12T U3691 ( .A1(n2752), .A2(n2751), .A3(n2750), .Z(n2753) );
  XOR3D1BWP12T U3692 ( .A1(n2755), .A2(n2754), .A3(n2753), .Z(n2756) );
  XNR2D1BWP12T U3693 ( .A1(n2757), .A2(n2756), .ZN(n2766) );
  FA1D2BWP12T U3694 ( .A(n2760), .B(n2759), .CI(n2758), .CO(n2765), .S(n2727)
         );
  FA1D2BWP12T U3695 ( .A(n2763), .B(n2762), .CI(n2761), .CO(n2764), .S(n2771)
         );
  XOR3D2BWP12T U3696 ( .A1(n2766), .A2(n2765), .A3(n2764), .Z(n2767) );
  XNR3XD4BWP12T U3697 ( .A1(n2769), .A2(n2768), .A3(n2767), .ZN(n2776) );
  CKND2D1BWP12T U3698 ( .A1(n321), .A2(n2770), .ZN(n2772) );
  OR2XD4BWP12T U3699 ( .A1(n2776), .A2(n2775), .Z(n2778) );
  ND2D1BWP12T U3700 ( .A1(n2776), .A2(n2775), .ZN(n2777) );
  AN2D4BWP12T U3701 ( .A1(n2778), .A2(n2777), .Z(n2779) );
  XNR2XD4BWP12T U3702 ( .A1(n2780), .A2(n2779), .ZN(n3486) );
  INVD1BWP12T U3703 ( .I(n3486), .ZN(n2843) );
  ND2D1BWP12T U3704 ( .A1(n4649), .A2(n4650), .ZN(n3707) );
  NR2D1BWP12T U3705 ( .A1(n3707), .A2(n4922), .ZN(n2901) );
  CKND2D1BWP12T U3706 ( .A1(n2901), .A2(n4667), .ZN(n2782) );
  NR2D1BWP12T U3707 ( .A1(n3708), .A2(n2782), .ZN(n2783) );
  ND2D1BWP12T U3708 ( .A1(n2783), .A2(n4426), .ZN(n3973) );
  NR2D1BWP12T U3709 ( .A1(n2851), .A2(n848), .ZN(n3488) );
  OR2XD1BWP12T U3710 ( .A1(n4740), .A2(n4907), .Z(n2968) );
  ND2D1BWP12T U3711 ( .A1(n2968), .A2(n2970), .ZN(n2784) );
  NR2D1BWP12T U3712 ( .A1(n2964), .A2(n2784), .ZN(n2786) );
  CKND2D1BWP12T U3713 ( .A1(n3909), .A2(n2786), .ZN(n2788) );
  NR2D1BWP12T U3714 ( .A1(n4366), .A2(n2788), .ZN(n2790) );
  INVD1BWP12T U3715 ( .I(n2798), .ZN(n2969) );
  ND2D1BWP12T U3716 ( .A1(n4740), .A2(n4907), .ZN(n2967) );
  TPAOI21D0BWP12T U3717 ( .A1(n2786), .A2(n3908), .B(n2785), .ZN(n2787) );
  OAI21D1BWP12T U3718 ( .A1(n4365), .A2(n2788), .B(n2787), .ZN(n2789) );
  TPAOI21D1BWP12T U3719 ( .A1(n2791), .A2(n2790), .B(n2789), .ZN(n3997) );
  NR2D1BWP12T U3720 ( .A1(n4739), .A2(n2792), .ZN(n3683) );
  NR2D1BWP12T U3721 ( .A1(b[26]), .A2(n4922), .ZN(n2797) );
  NR2D1BWP12T U3722 ( .A1(n3683), .A2(n2797), .ZN(n3993) );
  ND2D1BWP12T U3723 ( .A1(n4739), .A2(n2792), .ZN(n3831) );
  ND2D1BWP12T U3724 ( .A1(b[26]), .A2(n4922), .ZN(n3684) );
  OAI21D1BWP12T U3725 ( .A1(n2797), .A2(n3831), .B(n3684), .ZN(n3996) );
  OR2XD1BWP12T U3726 ( .A1(n4731), .A2(a[27]), .Z(n3995) );
  NR2D1BWP12T U3727 ( .A1(n4733), .A2(n4908), .ZN(n2805) );
  INVD0BWP12T U3728 ( .I(n2805), .ZN(n3999) );
  CKND2D0BWP12T U3729 ( .A1(n4731), .A2(a[27]), .ZN(n2930) );
  INVD1BWP12T U3730 ( .I(n2930), .ZN(n3994) );
  CKBD1BWP12T U3731 ( .I(n4909), .Z(n2793) );
  NR2D1BWP12T U3732 ( .A1(n4730), .A2(n2793), .ZN(n2806) );
  ND2D1BWP12T U3733 ( .A1(n4730), .A2(n2793), .ZN(n3589) );
  TPOAI21D1BWP12T U3734 ( .A1(n3555), .A2(n2806), .B(n3589), .ZN(n3480) );
  INVD1BWP12T U3735 ( .I(n4751), .ZN(n2853) );
  NR2D1BWP12T U3736 ( .A1(n4740), .A2(n4907), .ZN(n2799) );
  NR2D1BWP12T U3737 ( .A1(n2799), .A2(n2795), .ZN(n3829) );
  ND2D1BWP12T U3738 ( .A1(n3829), .A2(n3832), .ZN(n2800) );
  NR2D1BWP12T U3739 ( .A1(n2800), .A2(n2796), .ZN(n3696) );
  INVD0BWP12T U3740 ( .I(n2797), .ZN(n3685) );
  TPND2D0BWP12T U3741 ( .A1(n3696), .A2(n3685), .ZN(n2804) );
  TPOAI21D0BWP12T U3742 ( .A1(n2799), .A2(n2798), .B(n2967), .ZN(n3828) );
  CKND0BWP12T U3743 ( .I(n3684), .ZN(n2802) );
  TPAOI21D0BWP12T U3744 ( .A1(n3695), .A2(n3685), .B(n2802), .ZN(n2803) );
  CKND0BWP12T U3745 ( .I(n2806), .ZN(n3590) );
  INVD1BWP12T U3746 ( .I(n3589), .ZN(n2807) );
  AOI21D1BWP12T U3747 ( .A1(n3591), .A2(n3590), .B(n2807), .ZN(n3434) );
  NR2D1BWP12T U3748 ( .A1(n4727), .A2(n4933), .ZN(n3432) );
  ND2D1BWP12T U3749 ( .A1(n4727), .A2(n4933), .ZN(n3433) );
  OAI21D1BWP12T U3750 ( .A1(n3434), .A2(n3432), .B(n3433), .ZN(n2852) );
  OR2XD1BWP12T U3751 ( .A1(n4697), .A2(n4907), .Z(n2949) );
  ND2D1BWP12T U3752 ( .A1(n2949), .A2(n2953), .ZN(n2810) );
  NR2D1BWP12T U3753 ( .A1(n2941), .A2(n2810), .ZN(n2812) );
  ND2D1BWP12T U3754 ( .A1(n3878), .A2(n2812), .ZN(n2814) );
  NR2D1BWP12T U3755 ( .A1(n4984), .A2(n2814), .ZN(n2816) );
  INVD1BWP12T U3756 ( .I(n2942), .ZN(n2952) );
  ND2D1BWP12T U3757 ( .A1(n4697), .A2(n4907), .ZN(n2948) );
  INVD1BWP12T U3758 ( .I(n2948), .ZN(n2826) );
  AOI21D1BWP12T U3759 ( .A1(n2949), .A2(n2952), .B(n2826), .ZN(n2809) );
  TPOAI21D0BWP12T U3760 ( .A1(n3874), .A2(n2810), .B(n2809), .ZN(n2811) );
  AOI21D1BWP12T U3761 ( .A1(n2812), .A2(n3877), .B(n2811), .ZN(n2813) );
  OAI21D1BWP12T U3762 ( .A1(n4983), .A2(n2814), .B(n2813), .ZN(n2815) );
  NR2D1BWP12T U3763 ( .A1(n4695), .A2(n4922), .ZN(n2819) );
  NR2D1BWP12T U3764 ( .A1(n3723), .A2(n2819), .ZN(n3987) );
  INVD1BWP12T U3765 ( .I(n3987), .ZN(n2821) );
  ND2D1BWP12T U3766 ( .A1(n4698), .A2(n2818), .ZN(n3805) );
  ND2D1BWP12T U3767 ( .A1(n4695), .A2(n4922), .ZN(n3680) );
  OAI21D1BWP12T U3768 ( .A1(n2819), .A2(n3805), .B(n3680), .ZN(n3990) );
  INVD1BWP12T U3769 ( .I(n3990), .ZN(n2820) );
  CKBD1BWP12T U3770 ( .I(a[27]), .Z(n2885) );
  OR2XD0BWP12T U3771 ( .A1(n4696), .A2(n2885), .Z(n3989) );
  CKBD1BWP12T U3772 ( .I(a[27]), .Z(n2822) );
  ND2D1BWP12T U3773 ( .A1(n4696), .A2(n2822), .ZN(n2928) );
  INVD1BWP12T U3774 ( .I(n2928), .ZN(n3988) );
  ND2D1BWP12T U3775 ( .A1(n4694), .A2(n4908), .ZN(n3934) );
  INVD1BWP12T U3776 ( .I(n3934), .ZN(n2829) );
  CKBD1BWP12T U3777 ( .I(n4909), .Z(n2823) );
  NR2D1BWP12T U3778 ( .A1(n4693), .A2(n2823), .ZN(n3551) );
  ND2D1BWP12T U3779 ( .A1(n4693), .A2(n2823), .ZN(n3552) );
  OR2D1BWP12T U3780 ( .A1(n4711), .A2(n4933), .Z(n3429) );
  ND2D1BWP12T U3781 ( .A1(n4711), .A2(n4933), .ZN(n3428) );
  INVD1BWP12T U3782 ( .I(n3428), .ZN(n2824) );
  TPAOI21D0BWP12T U3783 ( .A1(n3430), .A2(n3429), .B(n2824), .ZN(n2850) );
  INVD1BWP12T U3784 ( .I(n2825), .ZN(n2840) );
  ND2D1BWP12T U3785 ( .A1(n2949), .A2(n2953), .ZN(n2828) );
  INVD1BWP12T U3786 ( .I(n3723), .ZN(n3806) );
  ND2D1BWP12T U3787 ( .A1(n3806), .A2(n3681), .ZN(n3928) );
  ND2D1BWP12T U3788 ( .A1(n3989), .A2(n3935), .ZN(n2831) );
  NR2D1BWP12T U3789 ( .A1(n3928), .A2(n2831), .ZN(n2833) );
  CKND2D1BWP12T U3790 ( .A1(n3802), .A2(n2833), .ZN(n2835) );
  OR2XD1BWP12T U3791 ( .A1(n3873), .A2(n2835), .Z(n2837) );
  AOI21D1BWP12T U3792 ( .A1(n2949), .A2(n2952), .B(n2826), .ZN(n2827) );
  OAI21D1BWP12T U3793 ( .A1(n3874), .A2(n2828), .B(n2827), .ZN(n3801) );
  AOI21D1BWP12T U3794 ( .A1(n3935), .A2(n3988), .B(n2829), .ZN(n2830) );
  OAI21D1BWP12T U3795 ( .A1(n3931), .A2(n2831), .B(n2830), .ZN(n2832) );
  TPAOI21D0BWP12T U3796 ( .A1(n3801), .A2(n2833), .B(n2832), .ZN(n2834) );
  OA21D1BWP12T U3797 ( .A1(n3872), .A2(n2835), .B(n2834), .Z(n2836) );
  INVD1BWP12T U3798 ( .I(n2838), .ZN(n2839) );
  AOI22D1BWP12T U3799 ( .A1(n2840), .A2(n5093), .B1(n5090), .B2(n2839), .ZN(
        n3487) );
  AN2XD2BWP12T U3800 ( .A1(n2841), .A2(n3487), .Z(n2842) );
  TPOAI21D1BWP12T U3801 ( .A1(n2843), .A2(n4260), .B(n2842), .ZN(c_out) );
  TPND2D3BWP12T U3802 ( .A1(n2845), .A2(n2844), .ZN(n2846) );
  XNR2XD4BWP12T U3803 ( .A1(n2847), .A2(n2846), .ZN(n4300) );
  ND2D4BWP12T U3804 ( .A1(n4300), .A2(n5085), .ZN(n2883) );
  FA1D0BWP12T U3805 ( .A(n4751), .B(n848), .CI(n2848), .CO(n2794), .S(n4472)
         );
  INVD1BWP12T U3806 ( .I(n4472), .ZN(n2849) );
  OR2XD1BWP12T U3807 ( .A1(n2849), .A2(n4396), .Z(n2881) );
  FICIND1BWP12T U3808 ( .CIN(n2850), .B(n3455), .A(n4751), .CO(n2825), .S(
        n4998) );
  ND2D1BWP12T U3809 ( .A1(n4998), .A2(n5093), .ZN(n2879) );
  XNR2D1BWP12T U3810 ( .A1(n2851), .A2(n848), .ZN(n4458) );
  INVD1BWP12T U3811 ( .I(n4458), .ZN(n2875) );
  INVD1BWP12T U3812 ( .I(n4799), .ZN(n3558) );
  CKND2D1BWP12T U3813 ( .A1(n3817), .A2(n4045), .ZN(n2854) );
  INVD1BWP12T U3814 ( .I(n4797), .ZN(n3108) );
  MUX2D1BWP12T U3815 ( .I0(n4667), .I1(n4666), .S(n5075), .Z(n2919) );
  TPNR2D0BWP12T U3816 ( .A1(n3945), .A2(n2919), .ZN(n2856) );
  MUX2D1BWP12T U3817 ( .I0(n3850), .I1(n4650), .S(n5075), .Z(n3816) );
  MUX2D1BWP12T U3818 ( .I0(n4664), .I1(n4665), .S(n5075), .Z(n2861) );
  OAI22D0BWP12T U3819 ( .A1(n3813), .A2(n3816), .B1(n3812), .B2(n2861), .ZN(
        n2855) );
  AOI211D0BWP12T U3820 ( .A1(n3941), .A2(n4933), .B(n2856), .C(n2855), .ZN(
        n2857) );
  OAI222D1BWP12T U3821 ( .A1(n3558), .A2(n2859), .B1(n3108), .B2(n2858), .C1(
        n3818), .C2(n2857), .ZN(n4840) );
  RCAOI21D0BWP12T U3822 ( .A1(n3947), .A2(n4779), .B(n4840), .ZN(n2860) );
  NR2XD0BWP12T U3823 ( .A1(n2860), .A2(n5040), .ZN(n2872) );
  INVD1BWP12T U3824 ( .I(n2861), .ZN(n3569) );
  INVD1BWP12T U3825 ( .I(n3816), .ZN(n3834) );
  OAI22D1BWP12T U3826 ( .A1(n3569), .A2(n3961), .B1(n3834), .B2(n3959), .ZN(
        n2863) );
  INVD1BWP12T U3827 ( .I(n2919), .ZN(n3570) );
  OAI22D1BWP12T U3828 ( .A1(n3570), .A2(n3963), .B1(n4933), .B2(n3462), .ZN(
        n2862) );
  NR2D1BWP12T U3829 ( .A1(n2863), .A2(n2862), .ZN(n2864) );
  OAI22D0BWP12T U3830 ( .A1(n2864), .A2(n4611), .B1(n848), .B2(n3817), .ZN(
        n2865) );
  AOI211D1BWP12T U3831 ( .A1(n3972), .A2(n2866), .B(n4891), .C(n2865), .ZN(
        n2869) );
  CKND2D0BWP12T U3832 ( .A1(n2867), .A2(n3761), .ZN(n2868) );
  OAI211D1BWP12T U3833 ( .A1(n4585), .A2(n3969), .B(n2869), .C(n2868), .ZN(
        n4616) );
  XNR2D1BWP12T U3834 ( .A1(n4751), .A2(n4624), .ZN(n4668) );
  RCAOI211D0BWP12T U3835 ( .A1(n4534), .A2(n5038), .B(n2872), .C(n2871), .ZN(
        n2873) );
  OAI211D1BWP12T U3836 ( .A1(n2875), .A2(n4420), .B(n2874), .C(n2873), .ZN(
        n2878) );
  FA1D0BWP12T U3837 ( .A(n4751), .B(n3455), .CI(n2876), .CO(n2838), .S(n4364)
         );
  INR3XD1BWP12T U3838 ( .A1(n2879), .B1(n2878), .B2(n2877), .ZN(n2880) );
  TPND2D2BWP12T U3839 ( .A1(n2881), .A2(n2880), .ZN(n4084) );
  INVD3BWP12T U3840 ( .I(n4084), .ZN(n2882) );
  ND2D4BWP12T U3841 ( .A1(n2883), .A2(n2882), .ZN(result[31]) );
  INR2D2BWP12T U3842 ( .A1(n3921), .B1(n3922), .ZN(n2884) );
  XNR2XD4BWP12T U3843 ( .A1(n3923), .A2(n2884), .ZN(n4301) );
  ND2XD8BWP12T U3844 ( .A1(n4301), .A2(n5085), .ZN(n2937) );
  INVD1BWP12T U3845 ( .I(n3802), .ZN(n3929) );
  INVD1BWP12T U3846 ( .I(n3801), .ZN(n3932) );
  ND2D1BWP12T U3847 ( .A1(n4315), .A2(n5090), .ZN(n2935) );
  IOA21D0BWP12T U3848 ( .A1(n4624), .A2(n3748), .B(n2887), .ZN(n2888) );
  AOI21D1BWP12T U3849 ( .A1(n3767), .A2(n3051), .B(n2888), .ZN(n3752) );
  TPND2D0BWP12T U3850 ( .A1(n3752), .A2(n4685), .ZN(n4821) );
  CKND0BWP12T U3851 ( .I(n3767), .ZN(n2890) );
  OAI21D0BWP12T U3852 ( .A1(n4521), .A2(n4624), .B(n3509), .ZN(n2889) );
  AOI21D0BWP12T U3853 ( .A1(n2890), .A2(n4039), .B(n2889), .ZN(n4892) );
  TPNR2D0BWP12T U3854 ( .A1(n3566), .A2(n4892), .ZN(n4887) );
  AOI22D1BWP12T U3855 ( .A1(n3125), .A2(n3121), .B1(n3098), .B2(n953), .ZN(
        n2892) );
  TPND2D0BWP12T U3856 ( .A1(n3096), .A2(n3701), .ZN(n2891) );
  OAI211D1BWP12T U3857 ( .A1(n3114), .A2(n3959), .B(n2892), .C(n2891), .ZN(
        n3762) );
  OAI22D1BWP12T U3858 ( .A1(n3099), .A2(n3957), .B1(n3061), .B2(n3961), .ZN(
        n4583) );
  AOI22D1BWP12T U3859 ( .A1(n3125), .A2(n3811), .B1(n3119), .B2(n953), .ZN(
        n2894) );
  TPND2D0BWP12T U3860 ( .A1(n3118), .A2(n3701), .ZN(n2893) );
  OAI211D1BWP12T U3861 ( .A1(n3104), .A2(n3959), .B(n2894), .C(n2893), .ZN(
        n3760) );
  AOI22D0BWP12T U3862 ( .A1(n3125), .A2(n2919), .B1(n3816), .B2(n953), .ZN(
        n2896) );
  AOI22D0BWP12T U3863 ( .A1(n3122), .A2(n3810), .B1(n2918), .B2(n3701), .ZN(
        n2895) );
  AOI21D0BWP12T U3864 ( .A1(n2896), .A2(n2895), .B(n4611), .ZN(n2897) );
  AOI211D1BWP12T U3865 ( .A1(n3760), .A2(n3761), .B(n2897), .C(n4891), .ZN(
        n2898) );
  TPOAI21D0BWP12T U3866 ( .A1(n5020), .A2(n4707), .B(n2898), .ZN(n4617) );
  NR2XD0BWP12T U3867 ( .A1(n4617), .A2(n5042), .ZN(n2899) );
  ND2D2BWP12T U3868 ( .A1(n3982), .A2(n5099), .ZN(n4165) );
  AOI211XD0BWP12T U3869 ( .A1(n5099), .A2(n4887), .B(n2899), .C(n3763), .ZN(
        n2908) );
  INVD1BWP12T U3870 ( .I(n3708), .ZN(n2900) );
  ND2D1BWP12T U3871 ( .A1(n4426), .A2(n2900), .ZN(n3846) );
  MUX2ND0BWP12T U3872 ( .I0(n5077), .I1(n5076), .S(n4731), .ZN(n2902) );
  NR2D0BWP12T U3873 ( .A1(n2902), .A2(n905), .ZN(n2903) );
  MUX2NXD0BWP12T U3874 ( .I0(n2903), .I1(n5080), .S(n4667), .ZN(n2906) );
  NR2D1BWP12T U3875 ( .A1(a[27]), .A2(n5083), .ZN(n2904) );
  OA21XD0BWP12T U3876 ( .A1(n905), .A2(n2904), .B(n4731), .Z(n2905) );
  AOI211D1BWP12T U3877 ( .A1(n4438), .A2(n5078), .B(n2906), .C(n2905), .ZN(
        n2907) );
  OAI211D1BWP12T U3878 ( .A1(n3899), .A2(n4821), .B(n2908), .C(n2907), .ZN(
        n2927) );
  AOI22D1BWP12T U3879 ( .A1(n3939), .A2(n3119), .B1(n3940), .B2(n3120), .ZN(
        n2911) );
  TPND2D0BWP12T U3880 ( .A1(n3937), .A2(n3118), .ZN(n2910) );
  TPND2D0BWP12T U3881 ( .A1(n3941), .A2(n3811), .ZN(n2909) );
  ND3D1BWP12T U3882 ( .A1(n2911), .A2(n2910), .A3(n2909), .ZN(n3753) );
  INVD1BWP12T U3883 ( .I(n3753), .ZN(n2925) );
  AOI22D1BWP12T U3884 ( .A1(n3941), .A2(n3121), .B1(n3940), .B2(n3100), .ZN(
        n2915) );
  ND2XD0BWP12T U3885 ( .A1(n3097), .A2(n3098), .ZN(n2913) );
  INR2XD0BWP12T U3886 ( .A1(n3096), .B1(n3945), .ZN(n2912) );
  INR2D1BWP12T U3887 ( .A1(n2913), .B1(n2912), .ZN(n2914) );
  ND2D1BWP12T U3888 ( .A1(n2915), .A2(n2914), .ZN(n3755) );
  AO21D1BWP12T U3889 ( .A1(n3755), .A2(n4032), .B(n2917), .Z(n5023) );
  CKND2D1BWP12T U3890 ( .A1(n5023), .A2(n4045), .ZN(n2924) );
  INVD1BWP12T U3891 ( .I(n2918), .ZN(n3835) );
  TPND2D0BWP12T U3892 ( .A1(n3941), .A2(n2919), .ZN(n2921) );
  AOI22D0BWP12T U3893 ( .A1(n3940), .A2(n3810), .B1(n3939), .B2(n3816), .ZN(
        n2920) );
  OAI211D1BWP12T U3894 ( .A1(n3835), .A2(n3945), .B(n2921), .C(n2920), .ZN(
        n2922) );
  AOI21D1BWP12T U3895 ( .A1(n2922), .A2(n4801), .B(n3690), .ZN(n2923) );
  OAI211D1BWP12T U3896 ( .A1(n2925), .A2(n3558), .B(n2924), .C(n2923), .ZN(
        n4813) );
  NR2D1BWP12T U3897 ( .A1(n4813), .A2(n5040), .ZN(n2926) );
  AOI211D1BWP12T U3898 ( .A1(n4503), .A2(n4103), .B(n2927), .C(n2926), .ZN(
        n2934) );
  ND2D1BWP12T U3899 ( .A1(n4945), .A2(n5093), .ZN(n2933) );
  ND2D1BWP12T U3900 ( .A1(n4413), .A2(n5088), .ZN(n2932) );
  AN4D4BWP12T U3901 ( .A1(n2935), .A2(n2934), .A3(n2933), .A4(n2932), .Z(n2936) );
  TPND2D8BWP12T U3902 ( .A1(n2937), .A2(n2936), .ZN(result[27]) );
  INVD1BWP12T U3903 ( .I(n291), .ZN(n2940) );
  INVD0BWP12T U3904 ( .I(n302), .ZN(n2938) );
  AN2XD2BWP12T U3905 ( .A1(n3795), .A2(n2938), .Z(n2939) );
  XNR2XD4BWP12T U3906 ( .A1(n2940), .A2(n2939), .ZN(n4289) );
  TPNR2D0BWP12T U3907 ( .A1(n2941), .A2(n2943), .ZN(n2945) );
  CKND2D1BWP12T U3908 ( .A1(n3930), .A2(n2945), .ZN(n2947) );
  TPOAI21D0BWP12T U3909 ( .A1(n3874), .A2(n2943), .B(n2942), .ZN(n2944) );
  AOI21D1BWP12T U3910 ( .A1(n3933), .A2(n2945), .B(n2944), .ZN(n2946) );
  OAI21D1BWP12T U3911 ( .A1(n4353), .A2(n2947), .B(n2946), .ZN(n2950) );
  ND2D1BWP12T U3912 ( .A1(n2949), .A2(n2948), .ZN(n2962) );
  CKND2D1BWP12T U3913 ( .A1(n3875), .A2(n2953), .ZN(n2956) );
  NR2D1BWP12T U3914 ( .A1(n2951), .A2(n2956), .ZN(n2959) );
  CKND2D1BWP12T U3915 ( .A1(n3876), .A2(n2959), .ZN(n2961) );
  TPAOI21D0BWP12T U3916 ( .A1(n2954), .A2(n2953), .B(n2952), .ZN(n2955) );
  OAI21D1BWP12T U3917 ( .A1(n2957), .A2(n2956), .B(n2955), .ZN(n2958) );
  TPAOI21D0BWP12T U3918 ( .A1(n3879), .A2(n2959), .B(n2958), .ZN(n2960) );
  OAI21D1BWP12T U3919 ( .A1(n4985), .A2(n2961), .B(n2960), .ZN(n2963) );
  INVD1BWP12T U3920 ( .I(n2964), .ZN(n3889) );
  CKND2D1BWP12T U3921 ( .A1(n2968), .A2(n2967), .ZN(n2971) );
  INVD1BWP12T U3922 ( .I(n4412), .ZN(n3016) );
  ND2D1BWP12T U3923 ( .A1(n4510), .A2(n4103), .ZN(n3015) );
  INVD1BWP12T U3924 ( .I(n2972), .ZN(n3435) );
  OAI22D1BWP12T U3925 ( .A1(n3435), .A2(n3959), .B1(n3471), .B2(n3963), .ZN(
        n2974) );
  INVD0BWP12T U3926 ( .I(n4154), .ZN(n2990) );
  INVD0BWP12T U3927 ( .I(n3953), .ZN(n2976) );
  INVD0BWP12T U3928 ( .I(n3954), .ZN(n2975) );
  AOI22D1BWP12T U3929 ( .A1(n3125), .A2(n2976), .B1(n2975), .B2(n953), .ZN(
        n2980) );
  CKND2D0BWP12T U3930 ( .A1(n2999), .A2(n3701), .ZN(n2978) );
  INVD1BWP12T U3931 ( .I(n3447), .ZN(n3457) );
  NR2D1BWP12T U3932 ( .A1(n3457), .A2(n3959), .ZN(n2977) );
  INR2XD0BWP12T U3933 ( .A1(n2978), .B1(n2977), .ZN(n2979) );
  ND2D1BWP12T U3934 ( .A1(n2980), .A2(n2979), .ZN(n4157) );
  CKND1BWP12T U3935 ( .I(n4157), .ZN(n2988) );
  MUX2XD0BWP12T U3936 ( .I0(n5051), .I1(n4924), .S(n5075), .Z(n3951) );
  OAI22D1BWP12T U3937 ( .A1(n3952), .A2(n3959), .B1(n3951), .B2(n3963), .ZN(
        n2983) );
  MUX2XD0BWP12T U3938 ( .I0(n4650), .I1(n2981), .S(n5075), .Z(n3944) );
  INVD1BWP12T U3939 ( .I(n3944), .ZN(n3964) );
  MUX2XD0BWP12T U3940 ( .I0(n4728), .I1(n4914), .S(n5075), .Z(n3960) );
  OAI22D1BWP12T U3941 ( .A1(n3964), .A2(n3957), .B1(n3960), .B2(n3961), .ZN(
        n2982) );
  TPOAI21D0BWP12T U3942 ( .A1(n2983), .A2(n2982), .B(n4158), .ZN(n2986) );
  NR2D1BWP12T U3943 ( .A1(n4567), .A2(n4742), .ZN(n4153) );
  IND2D0BWP12T U3944 ( .A1(n4153), .B1(n2984), .ZN(n2985) );
  AN2XD1BWP12T U3945 ( .A1(n2986), .A2(n2985), .Z(n2987) );
  OAI21D1BWP12T U3946 ( .A1(n2988), .A2(n3968), .B(n2987), .ZN(n2989) );
  AOI211D1BWP12T U3947 ( .A1(n3972), .A2(n2990), .B(n2989), .C(n4891), .ZN(
        n4591) );
  INVD1BWP12T U3948 ( .I(n4591), .ZN(n2996) );
  XOR2XD1BWP12T U3949 ( .A1(n3846), .A2(n4907), .Z(n4424) );
  OAI21D1BWP12T U3950 ( .A1(n4907), .A2(n5083), .B(n5081), .ZN(n2991) );
  AOI22D1BWP12T U3951 ( .A1(n4424), .A2(n5078), .B1(n4740), .B2(n2991), .ZN(
        n2995) );
  MUX2ND0BWP12T U3952 ( .I0(n5045), .I1(n5044), .S(n4740), .ZN(n2992) );
  TPND2D0BWP12T U3953 ( .A1(n2992), .A2(n5081), .ZN(n2993) );
  MUX2NXD0BWP12T U3954 ( .I0(n2993), .I1(n5048), .S(n4650), .ZN(n2994) );
  OAI211D1BWP12T U3955 ( .A1(n5042), .A2(n2996), .B(n2995), .C(n2994), .ZN(
        n3013) );
  NR2D1BWP12T U3956 ( .A1(n5038), .A2(n3903), .ZN(n4176) );
  OAI22D1BWP12T U3957 ( .A1(n4171), .A2(n4566), .B1(n4173), .B2(n4521), .ZN(
        n4888) );
  INVD1BWP12T U3958 ( .I(n4888), .ZN(n4539) );
  AOI22D0BWP12T U3959 ( .A1(n3954), .A2(n3939), .B1(n3940), .B2(n3457), .ZN(
        n2998) );
  CKND2D1BWP12T U3960 ( .A1(n3941), .A2(n3953), .ZN(n2997) );
  OAI211D1BWP12T U3961 ( .A1(n3945), .A2(n2999), .B(n2998), .C(n2997), .ZN(
        n4152) );
  CKND1BWP12T U3962 ( .I(n3960), .ZN(n3700) );
  AOI22D0BWP12T U3963 ( .A1(n3939), .A2(n3700), .B1(n3940), .B2(n3444), .ZN(
        n3001) );
  CKND2D0BWP12T U3964 ( .A1(n3941), .A2(n3944), .ZN(n3000) );
  OAI211D0BWP12T U3965 ( .A1(n3951), .A2(n3945), .B(n3001), .C(n3000), .ZN(
        n3003) );
  INVD1BWP12T U3966 ( .I(n3947), .ZN(n3556) );
  NR2XD0BWP12T U3967 ( .A1(n3556), .A2(n4153), .ZN(n3002) );
  AOI211D1BWP12T U3968 ( .A1(n3003), .A2(n4801), .B(n3690), .C(n3002), .ZN(
        n3011) );
  MAOI22D1BWP12T U3969 ( .A1(n3097), .A2(n3470), .B1(n3945), .B2(n3004), .ZN(
        n3008) );
  ND2D1BWP12T U3970 ( .A1(n3941), .A2(n3459), .ZN(n3007) );
  ND3D1BWP12T U3971 ( .A1(n3436), .A2(n3435), .A3(n3005), .ZN(n3006) );
  ND3D2BWP12T U3972 ( .A1(n3008), .A2(n3007), .A3(n3006), .ZN(n4151) );
  INVD1BWP12T U3973 ( .I(n4151), .ZN(n3009) );
  TPND3D0BWP12T U3974 ( .A1(n3009), .A2(n4045), .A3(n4032), .ZN(n3010) );
  OAI211D1BWP12T U3975 ( .A1(n3558), .A2(n4152), .B(n3011), .C(n3010), .ZN(
        n4795) );
  OAI22D1BWP12T U3976 ( .A1(n4176), .A2(n4539), .B1(n4795), .B2(n5040), .ZN(
        n3012) );
  OAI211D1BWP12T U3977 ( .A1(n3016), .A2(n4396), .B(n3015), .C(n3014), .ZN(
        n3017) );
  AOI21D1BWP12T U3978 ( .A1(n5093), .A2(n4978), .B(n3017), .ZN(n3018) );
  INVD1BWP12T U3979 ( .I(n3020), .ZN(n4290) );
  INVD1BWP12T U3980 ( .I(n311), .ZN(n3021) );
  TPAOI21D1BWP12T U3981 ( .A1(n3866), .A2(n4290), .B(n3021), .ZN(n3025) );
  AN2XD2BWP12T U3982 ( .A1(n3023), .A2(n277), .Z(n3024) );
  XNR2XD4BWP12T U3983 ( .A1(n3025), .A2(n3024), .ZN(n4296) );
  ND2D3BWP12T U3984 ( .A1(n4296), .A2(n5085), .ZN(n3083) );
  INVD1BWP12T U3985 ( .I(n3026), .ZN(n4355) );
  CKND2D0BWP12T U3986 ( .A1(n4349), .A2(n4355), .ZN(n3028) );
  INVD1BWP12T U3987 ( .I(n4354), .ZN(n3032) );
  TPAOI21D0BWP12T U3988 ( .A1(n4350), .A2(n4355), .B(n3032), .ZN(n3027) );
  OAI21D1BWP12T U3989 ( .A1(n4353), .A2(n3028), .B(n3027), .ZN(n3031) );
  XNR2XD1BWP12T U3990 ( .A1(n3031), .A2(n3035), .ZN(n4359) );
  CKND2D1BWP12T U3991 ( .A1(n4359), .A2(n5090), .ZN(n3081) );
  TPND2D0BWP12T U3992 ( .A1(n3876), .A2(n4355), .ZN(n3034) );
  AOI21D1BWP12T U3993 ( .A1(n3879), .A2(n4355), .B(n3032), .ZN(n3033) );
  OAI21D1BWP12T U3994 ( .A1(n4985), .A2(n3034), .B(n3033), .ZN(n3036) );
  XNR2XD1BWP12T U3995 ( .A1(n3036), .A2(n3035), .ZN(n4990) );
  CKND2D1BWP12T U3996 ( .A1(n4990), .A2(n5093), .ZN(n3080) );
  INVD0BWP12T U3997 ( .I(n3039), .ZN(n3886) );
  CKND2D1BWP12T U3998 ( .A1(n3886), .A2(n3884), .ZN(n3076) );
  XNR2XD1BWP12T U3999 ( .A1(n3887), .A2(n3076), .ZN(n4504) );
  INVD1BWP12T U4000 ( .I(n4665), .ZN(n4459) );
  CKND2D1BWP12T U4001 ( .A1(n3220), .A2(n4459), .ZN(n3042) );
  CKND2D1BWP12T U4002 ( .A1(n3217), .A2(n3040), .ZN(n3041) );
  ND2D1BWP12T U4003 ( .A1(n3042), .A2(n3041), .ZN(n3044) );
  AN2D1BWP12T U4004 ( .A1(n3219), .A2(n3847), .Z(n3043) );
  NR2D1BWP12T U4005 ( .A1(n275), .A2(n4666), .ZN(n3045) );
  INR2D2BWP12T U4006 ( .A1(n3046), .B1(n3045), .ZN(n3824) );
  TPOAI22D1BWP12T U4007 ( .A1(n3321), .A2(n4465), .B1(n275), .B2(n4651), .ZN(
        n3048) );
  OAI22D1BWP12T U4008 ( .A1(n3323), .A2(n4625), .B1(n3322), .B2(n4650), .ZN(
        n3047) );
  NR2D2BWP12T U4009 ( .A1(n3048), .A2(n3047), .ZN(n3502) );
  OAI22D1BWP12T U4010 ( .A1(n3824), .A2(n4521), .B1(n3502), .B2(n4566), .ZN(
        n3052) );
  CKND2D1BWP12T U4011 ( .A1(n3218), .A2(n4933), .ZN(n3050) );
  CKND2D1BWP12T U4012 ( .A1(n3219), .A2(n4909), .ZN(n3049) );
  ND2D1BWP12T U4013 ( .A1(n3050), .A2(n3049), .ZN(n3128) );
  INVD1BWP12T U4014 ( .I(n3823), .ZN(n4536) );
  TPND2D0BWP12T U4015 ( .A1(n5038), .A2(n4542), .ZN(n3060) );
  MUX2ND0BWP12T U4016 ( .I0(n5077), .I1(n5076), .S(n4726), .ZN(n3054) );
  NR2D0BWP12T U4017 ( .A1(n3054), .A2(n905), .ZN(n3055) );
  MUX2NXD0BWP12T U4018 ( .I0(n3055), .I1(n5080), .S(n4625), .ZN(n3058) );
  NR2D0BWP12T U4019 ( .A1(n4914), .A2(n5083), .ZN(n3056) );
  AOI211D1BWP12T U4020 ( .A1(n4430), .A2(n5078), .B(n3058), .C(n3057), .ZN(
        n3059) );
  OAI211D1BWP12T U4021 ( .A1(n4859), .A2(n3777), .B(n3060), .C(n3059), .ZN(
        n3071) );
  INVD1BWP12T U4022 ( .I(n3203), .ZN(n3565) );
  AOI22D1BWP12T U4023 ( .A1(n4801), .A2(n3559), .B1(n3557), .B2(n4045), .ZN(
        n3062) );
  OAI211D1BWP12T U4024 ( .A1(n4032), .A2(n3565), .B(n3062), .C(n3756), .ZN(
        n4794) );
  AOI22D1BWP12T U4025 ( .A1(n3125), .A2(n3810), .B1(n3811), .B2(n953), .ZN(
        n3064) );
  AOI22D1BWP12T U4026 ( .A1(n3122), .A2(n3118), .B1(n3119), .B2(n3701), .ZN(
        n3063) );
  ND2D1BWP12T U4027 ( .A1(n3064), .A2(n3063), .ZN(n3568) );
  OAI22D1BWP12T U4028 ( .A1(n3105), .A2(n3961), .B1(n3104), .B2(n3957), .ZN(
        n3066) );
  OAI22D1BWP12T U4029 ( .A1(n3113), .A2(n3959), .B1(n3112), .B2(n3963), .ZN(
        n3065) );
  NR2D1BWP12T U4030 ( .A1(n3066), .A2(n3065), .ZN(n3178) );
  OAI22D1BWP12T U4031 ( .A1(n3178), .A2(n4685), .B1(n3575), .B2(n4707), .ZN(
        n3068) );
  AOI211D1BWP12T U4032 ( .A1(n4158), .A2(n3568), .B(n4156), .C(n3068), .ZN(
        n4602) );
  CKND2D1BWP12T U4033 ( .A1(n4602), .A2(n4167), .ZN(n3069) );
  OAI211D1BWP12T U4034 ( .A1(n5040), .A2(n4794), .B(n4165), .C(n3069), .ZN(
        n3070) );
  AOI211D1BWP12T U4035 ( .A1(n4504), .A2(n4103), .B(n3071), .C(n3070), .ZN(
        n3079) );
  INVD1BWP12T U4036 ( .I(n3072), .ZN(n4369) );
  ND2XD0BWP12T U4037 ( .A1(n3907), .A2(n4369), .ZN(n3075) );
  INVD0BWP12T U4038 ( .I(n4368), .ZN(n3073) );
  AOI21D1BWP12T U4039 ( .A1(n3910), .A2(n4369), .B(n3073), .ZN(n3074) );
  OAI21D1BWP12T U4040 ( .A1(n4367), .A2(n3075), .B(n3074), .ZN(n3077) );
  XNR2D1BWP12T U4041 ( .A1(n3077), .A2(n3076), .ZN(n4373) );
  CKND2D1BWP12T U4042 ( .A1(n4373), .A2(n5088), .ZN(n3078) );
  AN4D2BWP12T U4043 ( .A1(n3081), .A2(n3080), .A3(n3079), .A4(n3078), .Z(n3082) );
  TPND2D3BWP12T U4044 ( .A1(n3083), .A2(n3082), .ZN(result[21]) );
  INVD1BWP12T U4045 ( .I(n3084), .ZN(n4148) );
  TPAOI21D1BWP12T U4046 ( .A1(n4148), .A2(n4146), .B(n4144), .ZN(n3088) );
  IND2D1BWP12T U4047 ( .A1(n3086), .B1(n3085), .ZN(n3087) );
  OAI21D1BWP12T U4048 ( .A1(n4985), .A2(n4189), .B(n4190), .ZN(n3092) );
  INVD1BWP12T U4049 ( .I(n3089), .ZN(n3091) );
  ND2D1BWP12T U4050 ( .A1(n3091), .A2(n3090), .ZN(n3158) );
  OAI21D1BWP12T U4051 ( .A1(n4367), .A2(n4149), .B(n4150), .ZN(n3095) );
  CKND2D1BWP12T U4052 ( .A1(n3094), .A2(n3093), .ZN(n3160) );
  INVD1BWP12T U4053 ( .I(n4409), .ZN(n3166) );
  AOI22D0BWP12T U4054 ( .A1(n3937), .A2(n3100), .B1(n3940), .B2(n3099), .ZN(
        n3101) );
  INVD1BWP12T U4055 ( .I(n3499), .ZN(n3111) );
  AOI22D1BWP12T U4056 ( .A1(n3937), .A2(n3104), .B1(n3103), .B2(n3939), .ZN(
        n3821) );
  INVD0BWP12T U4057 ( .I(n3119), .ZN(n3106) );
  AOI22D1BWP12T U4058 ( .A1(n3941), .A2(n3106), .B1(n3105), .B2(n3940), .ZN(
        n3822) );
  TPAOI21D0BWP12T U4059 ( .A1(n3821), .A2(n3822), .B(n3818), .ZN(n3110) );
  ND2D1BWP12T U4060 ( .A1(n3107), .A2(n3126), .ZN(n4251) );
  NR2D1BWP12T U4061 ( .A1(n3108), .A2(n4251), .ZN(n3109) );
  AOI211D1BWP12T U4062 ( .A1(n4799), .A2(n3111), .B(n3110), .C(n3109), .ZN(
        n4793) );
  OAI22D1BWP12T U4063 ( .A1(n3113), .A2(n3961), .B1(n3112), .B2(n3957), .ZN(
        n3117) );
  OAI22D1BWP12T U4064 ( .A1(n3115), .A2(n3959), .B1(n3114), .B2(n3963), .ZN(
        n3116) );
  NR2D1BWP12T U4065 ( .A1(n3117), .A2(n3116), .ZN(n3520) );
  INVD1BWP12T U4066 ( .I(n4156), .ZN(n4610) );
  AOI22D1BWP12T U4067 ( .A1(n3125), .A2(n3119), .B1(n3118), .B2(n953), .ZN(
        n3124) );
  AOI22D1BWP12T U4068 ( .A1(n3122), .A2(n3121), .B1(n3120), .B2(n3701), .ZN(
        n3123) );
  ND2D1BWP12T U4069 ( .A1(n3124), .A2(n3123), .ZN(n3833) );
  ND2D1BWP12T U4070 ( .A1(n3126), .A2(n3125), .ZN(n4248) );
  AOI22D1BWP12T U4071 ( .A1(n3833), .A2(n4158), .B1(n4843), .B2(n4248), .ZN(
        n3127) );
  OAI211D1BWP12T U4072 ( .A1(n3520), .A2(n3968), .B(n4610), .C(n3127), .ZN(
        n4613) );
  NR2D1BWP12T U4073 ( .A1(n3824), .A2(n4742), .ZN(n3132) );
  NR2D1BWP12T U4074 ( .A1(n3959), .A2(n4624), .ZN(n3130) );
  NR2XD0BWP12T U4075 ( .A1(n3130), .A2(n3129), .ZN(n3131) );
  OR2D2BWP12T U4076 ( .A1(n3502), .A2(n4521), .Z(n3141) );
  INVD0BWP12T U4077 ( .I(n4637), .ZN(n3133) );
  CKND2D1BWP12T U4078 ( .A1(n3218), .A2(n3133), .ZN(n3134) );
  OAI21D1BWP12T U4079 ( .A1(n3323), .A2(n1810), .B(n3134), .ZN(n3137) );
  ND2D1BWP12T U4080 ( .A1(n3220), .A2(n5051), .ZN(n3135) );
  OAI21D1BWP12T U4081 ( .A1(n3321), .A2(n1342), .B(n3135), .ZN(n3136) );
  NR2D1BWP12T U4082 ( .A1(n3137), .A2(n3136), .ZN(n3503) );
  NR2D1BWP12T U4083 ( .A1(n3503), .A2(n4566), .ZN(n3140) );
  INVD1BWP12T U4084 ( .I(n3140), .ZN(n3138) );
  ND2D1BWP12T U4085 ( .A1(n3141), .A2(n3138), .ZN(n3139) );
  OA22D1BWP12T U4086 ( .A1(n4613), .A2(n5042), .B1(n4861), .B2(n3777), .Z(
        n3153) );
  INVD1BWP12T U4087 ( .I(n4788), .ZN(n4822) );
  AO21D1BWP12T U4088 ( .A1(n4638), .A2(n3142), .B(n2688), .Z(n3145) );
  ND4D0BWP12T U4089 ( .A1(n4448), .A2(n3142), .A3(n2688), .A4(n4638), .ZN(
        n3144) );
  OR2XD1BWP12T U4090 ( .A1(n4448), .A2(n2688), .Z(n3143) );
  ND3D1BWP12T U4091 ( .A1(n3145), .A2(n3144), .A3(n3143), .ZN(n4429) );
  OAI21D0BWP12T U4092 ( .A1(n2688), .A2(n5083), .B(n5081), .ZN(n3146) );
  AOI22D1BWP12T U4093 ( .A1(n4429), .A2(n5078), .B1(n279), .B2(n3146), .ZN(
        n3150) );
  MUX2ND0BWP12T U4094 ( .I0(n5045), .I1(n5044), .S(n280), .ZN(n3147) );
  TPND2D0BWP12T U4095 ( .A1(n3147), .A2(n5081), .ZN(n3148) );
  MUX2NXD0BWP12T U4096 ( .I0(n3148), .I1(n5048), .S(n1810), .ZN(n3149) );
  CKND2D1BWP12T U4097 ( .A1(n3150), .A2(n3149), .ZN(n3151) );
  AOI211D1BWP12T U4098 ( .A1(n4822), .A2(n5038), .B(n3763), .C(n3151), .ZN(
        n3152) );
  OA211D1BWP12T U4099 ( .A1(n4793), .A2(n5040), .B(n3153), .C(n3152), .Z(n3165) );
  CKND0BWP12T U4100 ( .I(n4192), .ZN(n3154) );
  NR2XD0BWP12T U4101 ( .A1(n3154), .A2(n4189), .ZN(n3157) );
  CKND1BWP12T U4102 ( .I(n4191), .ZN(n3155) );
  TPOAI21D0BWP12T U4103 ( .A1(n3155), .A2(n4189), .B(n4190), .ZN(n3156) );
  AOI21D1BWP12T U4104 ( .A1(n4333), .A2(n3157), .B(n3156), .ZN(n3159) );
  XOR2XD1BWP12T U4105 ( .A1(n3159), .A2(n3158), .Z(n4325) );
  ND2D1BWP12T U4106 ( .A1(n4325), .A2(n5090), .ZN(n3163) );
  XNR2D1BWP12T U4107 ( .A1(n3161), .A2(n3160), .ZN(n4512) );
  AN2XD2BWP12T U4108 ( .A1(n4512), .A2(n4103), .Z(n3162) );
  INR2D2BWP12T U4109 ( .A1(n3163), .B1(n3162), .ZN(n3164) );
  OAI211D1BWP12T U4110 ( .A1(n4396), .A2(n3166), .B(n3165), .C(n3164), .ZN(
        n3167) );
  AOI21D2BWP12T U4111 ( .A1(n5093), .A2(n4947), .B(n3167), .ZN(n3168) );
  INVD1BWP12T U4112 ( .I(n3169), .ZN(n4006) );
  ND2D1BWP12T U4113 ( .A1(n4005), .A2(n4006), .ZN(n3170) );
  NR2D0BWP12T U4114 ( .A1(n4014), .A2(n3173), .ZN(n3175) );
  OAI21D0BWP12T U4115 ( .A1(n4017), .A2(n3173), .B(n3172), .ZN(n3174) );
  TPAOI21D0BWP12T U4116 ( .A1(n4971), .A2(n3175), .B(n3174), .ZN(n3177) );
  CKND2D1BWP12T U4117 ( .A1(n3176), .A2(n4071), .ZN(n3197) );
  XOR2XD1BWP12T U4118 ( .A1(n3177), .A2(n3197), .Z(n4977) );
  INVD1BWP12T U4119 ( .I(n4977), .ZN(n3194) );
  INVD1BWP12T U4120 ( .I(n3178), .ZN(n3578) );
  INVD1BWP12T U4121 ( .I(n3575), .ZN(n4588) );
  MUX2NXD0BWP12T U4122 ( .I0(n3578), .I1(n4588), .S(n4743), .ZN(n3179) );
  CKND2D1BWP12T U4123 ( .A1(n3179), .A2(n4605), .ZN(n4594) );
  CKND2D1BWP12T U4124 ( .A1(n4536), .A2(n4039), .ZN(n3185) );
  OAI22D1BWP12T U4125 ( .A1(n3824), .A2(n4554), .B1(n3503), .B2(n4521), .ZN(
        n3184) );
  OAI21D0BWP12T U4126 ( .A1(n3502), .A2(n4206), .B(n4707), .ZN(n3183) );
  OAI22D1BWP12T U4127 ( .A1(n3321), .A2(n4930), .B1(n275), .B2(n4680), .ZN(
        n3181) );
  OAI22D1BWP12T U4128 ( .A1(n3323), .A2(n4653), .B1(n3322), .B2(n4638), .ZN(
        n3180) );
  NR2D1BWP12T U4129 ( .A1(n3181), .A2(n3180), .ZN(n4208) );
  NR2D1BWP12T U4130 ( .A1(n4208), .A2(n4566), .ZN(n3182) );
  NR3D1BWP12T U4131 ( .A1(n3184), .A2(n3183), .A3(n3182), .ZN(n3191) );
  AOI21D1BWP12T U4132 ( .A1(n4843), .A2(n3185), .B(n3191), .ZN(n4551) );
  CKND2D1BWP12T U4133 ( .A1(n3186), .A2(n4551), .ZN(n3189) );
  OA211D1BWP12T U4134 ( .A1(n5042), .A2(n4594), .B(n3189), .C(n3188), .Z(n3193) );
  NR2D0BWP12T U4135 ( .A1(n3190), .A2(n4743), .ZN(n3567) );
  CKND2D1BWP12T U4136 ( .A1(n4896), .A2(n5099), .ZN(n3192) );
  OAI211D1BWP12T U4137 ( .A1(n4954), .A2(n3194), .B(n3193), .C(n3192), .ZN(
        n3202) );
  CKND0BWP12T U4138 ( .I(n4070), .ZN(n3196) );
  INVD1BWP12T U4139 ( .I(n4073), .ZN(n3195) );
  AOI21D1BWP12T U4140 ( .A1(n4333), .A2(n3196), .B(n3195), .ZN(n3198) );
  XOR2XD1BWP12T U4141 ( .A1(n3198), .A2(n3197), .Z(n4338) );
  AN2XD1BWP12T U4142 ( .A1(n4025), .A2(n3200), .Z(n3209) );
  AOI22D1BWP12T U4143 ( .A1(n5090), .A2(n4338), .B1(n4480), .B2(n4103), .ZN(
        n3201) );
  MUX2ND0BWP12T U4144 ( .I0(n3203), .I1(n3557), .S(n3754), .ZN(n3204) );
  AOI21D1BWP12T U4145 ( .A1(n3204), .A2(n3758), .B(n4551), .ZN(n4826) );
  TPOAI21D2BWP12T U4146 ( .A1(n4278), .A2(n4260), .B(n3212), .ZN(result[13])
         );
  CKND0BWP12T U4147 ( .I(n3214), .ZN(n3404) );
  CKND2D1BWP12T U4148 ( .A1(n3404), .A2(n3402), .ZN(n3232) );
  XNR2D1BWP12T U4149 ( .A1(n3534), .A2(n3232), .ZN(n4498) );
  CKND2D1BWP12T U4150 ( .A1(n4498), .A2(n4103), .ZN(n3247) );
  AOI22D0BWP12T U4151 ( .A1(n3218), .A2(n4925), .B1(n3217), .B2(n4926), .ZN(
        n3216) );
  AOI22D0BWP12T U4152 ( .A1(n3220), .A2(n4932), .B1(n3219), .B2(n5014), .ZN(
        n3215) );
  ND2D1BWP12T U4153 ( .A1(n3216), .A2(n3215), .ZN(n4089) );
  INVD1BWP12T U4154 ( .I(n4089), .ZN(n4520) );
  AOI22D0BWP12T U4155 ( .A1(n3218), .A2(n4905), .B1(n4906), .B2(n3217), .ZN(
        n3222) );
  AOI22D0BWP12T U4156 ( .A1(n3220), .A2(n4904), .B1(n3219), .B2(n288), .ZN(
        n3221) );
  CKND2D1BWP12T U4157 ( .A1(n3222), .A2(n3221), .ZN(n4088) );
  TPOAI21D0BWP12T U4158 ( .A1(n4540), .A2(n5040), .B(n5098), .ZN(n3229) );
  CKND1BWP12T U4159 ( .I(n3224), .ZN(n3225) );
  TPOAI21D0BWP12T U4160 ( .A1(n3225), .A2(n4707), .B(n3969), .ZN(n3226) );
  ND2D0BWP12T U4161 ( .A1(n3226), .A2(n3509), .ZN(n3227) );
  TPAOI31D0BWP12T U4162 ( .A1(n3227), .A2(n4573), .A3(n4823), .B(n5100), .ZN(
        n4879) );
  OR2D0BWP12T U4163 ( .A1(n4879), .A2(n5063), .Z(n3228) );
  IOA21D1BWP12T U4164 ( .A1(n4823), .A2(n3229), .B(n3228), .ZN(n3246) );
  NR2D1BWP12T U4165 ( .A1(n4540), .A2(n4891), .ZN(n3230) );
  OAI21D1BWP12T U4166 ( .A1(n3230), .A2(n4605), .B(n4823), .ZN(n4577) );
  NR2D1BWP12T U4167 ( .A1(n3818), .A2(n5040), .ZN(n4094) );
  AN2XD1BWP12T U4168 ( .A1(n4094), .A2(n4779), .Z(n3243) );
  INVD1BWP12T U4169 ( .I(n4585), .ZN(n3241) );
  MUX2ND0BWP12T U4170 ( .I0(n5077), .I1(n5076), .S(n4750), .ZN(n3235) );
  NR2XD0BWP12T U4171 ( .A1(n3235), .A2(n905), .ZN(n3236) );
  MUX2NXD0BWP12T U4172 ( .I0(n3236), .I1(n5080), .S(n4679), .ZN(n3239) );
  NR2D0BWP12T U4173 ( .A1(n288), .A2(n5083), .ZN(n3237) );
  OA21XD1BWP12T U4174 ( .A1(n905), .A2(n3237), .B(n4750), .Z(n3238) );
  AOI211XD0BWP12T U4175 ( .A1(n4431), .A2(n5078), .B(n3239), .C(n3238), .ZN(
        n3240) );
  TPOAI21D0BWP12T U4176 ( .A1(n3604), .A2(n3241), .B(n3240), .ZN(n3242) );
  AOI211D1BWP12T U4177 ( .A1(n4389), .A2(n5088), .B(n3243), .C(n3242), .ZN(
        n3244) );
  OAI21D1BWP12T U4178 ( .A1(n4577), .A2(n5102), .B(n3244), .ZN(n3245) );
  INVD1BWP12T U4179 ( .I(n3376), .ZN(n3248) );
  ND2D1BWP12T U4180 ( .A1(n3248), .A2(n3375), .ZN(n3250) );
  XOR2XD1BWP12T U4181 ( .A1(n3250), .A2(n3377), .Z(n4269) );
  INVD0BWP12T U4182 ( .I(n3651), .ZN(n3251) );
  NR2XD0BWP12T U4183 ( .A1(n3251), .A2(n3602), .ZN(n3254) );
  ND2XD0BWP12T U4184 ( .A1(n3254), .A2(n3649), .ZN(n3256) );
  CKND0BWP12T U4185 ( .I(n3650), .ZN(n3252) );
  TPOAI21D0BWP12T U4186 ( .A1(n3252), .A2(n3602), .B(n3603), .ZN(n3253) );
  AOI21D1BWP12T U4187 ( .A1(n3652), .A2(n3254), .B(n3253), .ZN(n3255) );
  OAI21D1BWP12T U4188 ( .A1(n4486), .A2(n3256), .B(n3255), .ZN(n3257) );
  XNR2D1BWP12T U4189 ( .A1(n3257), .A2(n3260), .ZN(n4961) );
  INVD1BWP12T U4190 ( .I(n3345), .ZN(n3598) );
  ND2XD0BWP12T U4191 ( .A1(n3598), .A2(n3409), .ZN(n3259) );
  INVD1BWP12T U4192 ( .I(n3344), .ZN(n3601) );
  AOI21D1BWP12T U4193 ( .A1(n3601), .A2(n3409), .B(n3410), .ZN(n3258) );
  OAI21D1BWP12T U4194 ( .A1(n4244), .A2(n3259), .B(n3258), .ZN(n3261) );
  XNR2D1BWP12T U4195 ( .A1(n3261), .A2(n3260), .ZN(n4329) );
  AO22D1BWP12T U4196 ( .A1(n5093), .A2(n4961), .B1(n4329), .B2(n5090), .Z(
        n3262) );
  CKND2D2BWP12T U4197 ( .A1(n4276), .A2(n5085), .ZN(n3317) );
  INVD1BWP12T U4198 ( .I(n3269), .ZN(n3498) );
  AOI21D1BWP12T U4199 ( .A1(n4333), .A2(n3498), .B(n3270), .ZN(n3272) );
  CKND2D1BWP12T U4200 ( .A1(n3271), .A2(n4966), .ZN(n3309) );
  XOR2XD1BWP12T U4201 ( .A1(n3272), .A2(n3309), .Z(n4340) );
  CKND2D0BWP12T U4202 ( .A1(n3273), .A2(n4379), .ZN(n3287) );
  CKND2D1BWP12T U4203 ( .A1(n4789), .A2(n4685), .ZN(n4543) );
  TPAOI21D0BWP12T U4204 ( .A1(n3274), .A2(n4039), .B(n4843), .ZN(n3275) );
  OAI21D1BWP12T U4205 ( .A1(n3637), .A2(n4521), .B(n3275), .ZN(n3276) );
  AOI21D1BWP12T U4206 ( .A1(n4743), .A2(n3277), .B(n3276), .ZN(n4836) );
  INVD1BWP12T U4207 ( .I(n4836), .ZN(n3278) );
  TPOAI21D0BWP12T U4208 ( .A1(n4543), .A2(n4891), .B(n4890), .ZN(n3279) );
  ND2D1BWP12T U4209 ( .A1(n3279), .A2(n3278), .ZN(n4550) );
  NR2D1BWP12T U4210 ( .A1(n4550), .A2(n5102), .ZN(n3280) );
  CKND0BWP12T U4211 ( .I(n3533), .ZN(n3282) );
  NR2D0BWP12T U4212 ( .A1(n3282), .A2(n3283), .ZN(n3286) );
  CKND0BWP12T U4213 ( .I(n3532), .ZN(n3284) );
  OAI21D0BWP12T U4214 ( .A1(n3284), .A2(n3283), .B(n3535), .ZN(n3285) );
  TPAOI21D0BWP12T U4215 ( .A1(n3534), .A2(n3286), .B(n3285), .ZN(n3288) );
  XOR2XD1BWP12T U4216 ( .A1(n3288), .A2(n3287), .Z(n4497) );
  MUX2NXD0BWP12T U4217 ( .I0(n3290), .I1(n3289), .S(n4032), .ZN(n4806) );
  CKND2D1BWP12T U4218 ( .A1(n3758), .A2(n5094), .ZN(n5024) );
  TPND2D0BWP12T U4219 ( .A1(n3292), .A2(n4743), .ZN(n3293) );
  INR2D1BWP12T U4220 ( .A1(n3295), .B1(n4891), .ZN(n5097) );
  INVD1BWP12T U4221 ( .I(n5097), .ZN(n3526) );
  OAI21D1BWP12T U4222 ( .A1(n4904), .A2(n5083), .B(n5081), .ZN(n3300) );
  MUX2ND0BWP12T U4223 ( .I0(n5077), .I1(n5076), .S(n3296), .ZN(n3297) );
  NR2D0BWP12T U4224 ( .A1(n3297), .A2(n905), .ZN(n3298) );
  MUX2NXD0BWP12T U4225 ( .I0(n3298), .I1(n5080), .S(n4654), .ZN(n3299) );
  AOI21D1BWP12T U4226 ( .A1(n342), .A2(n3300), .B(n3299), .ZN(n3302) );
  CKND2D1BWP12T U4227 ( .A1(n4443), .A2(n5078), .ZN(n3301) );
  OAI211D1BWP12T U4228 ( .A1(n4580), .A2(n3526), .B(n3302), .C(n3301), .ZN(
        n3303) );
  CKND0BWP12T U4229 ( .I(n4965), .ZN(n3308) );
  INVD1BWP12T U4230 ( .I(n4968), .ZN(n3307) );
  AOI21D1BWP12T U4231 ( .A1(n4971), .A2(n3308), .B(n3307), .ZN(n3310) );
  XOR2XD1BWP12T U4232 ( .A1(n3310), .A2(n3309), .Z(n4962) );
  MUX2D1BWP12T U4233 ( .I0(n4036), .I1(n3456), .S(n4742), .Z(n3311) );
  TPAOI21D0BWP12T U4234 ( .A1(n3311), .A2(n4685), .B(n3408), .ZN(n4877) );
  CKND0BWP12T U4235 ( .I(n4877), .ZN(n3312) );
  AOI21D0BWP12T U4236 ( .A1(n3312), .A2(n4573), .B(n4605), .ZN(n3313) );
  OAI21D1BWP12T U4237 ( .A1(n3313), .A2(n4836), .B(n4046), .ZN(n4898) );
  AOI211XD1BWP12T U4238 ( .A1(n5090), .A2(n4340), .B(n3315), .C(n3314), .ZN(
        n3316) );
  TPND2D2BWP12T U4239 ( .A1(n3317), .A2(n3316), .ZN(result[10]) );
  TPOAI21D0BWP12T U4240 ( .A1(n4208), .A2(n4206), .B(n4707), .ZN(n3329) );
  TPNR2D0BWP12T U4241 ( .A1(n3503), .A2(n4554), .ZN(n3328) );
  OAI22D1BWP12T U4242 ( .A1(n3321), .A2(n777), .B1(n275), .B2(n4654), .ZN(
        n3320) );
  OAI22D1BWP12T U4243 ( .A1(n3318), .A2(n3523), .B1(n3322), .B2(n4652), .ZN(
        n3319) );
  NR2D1BWP12T U4244 ( .A1(n3320), .A2(n3319), .ZN(n4207) );
  TPNR2D0BWP12T U4245 ( .A1(n4207), .A2(n4521), .ZN(n3327) );
  OAI22D1BWP12T U4246 ( .A1(n3321), .A2(n4679), .B1(n275), .B2(n4631), .ZN(
        n3325) );
  OAI22D0BWP12T U4247 ( .A1(n3323), .A2(n4627), .B1(n3322), .B2(n4655), .ZN(
        n3324) );
  NR2D1BWP12T U4248 ( .A1(n3325), .A2(n3324), .ZN(n4199) );
  TPNR2D0BWP12T U4249 ( .A1(n4199), .A2(n4566), .ZN(n3326) );
  NR4D0BWP12T U4250 ( .A1(n3329), .A2(n3328), .A3(n3327), .A4(n3326), .ZN(
        n3332) );
  INVD1BWP12T U4251 ( .I(n3337), .ZN(n4546) );
  INR2D1BWP12T U4252 ( .A1(n4209), .B1(n4546), .ZN(n3330) );
  ND2D1BWP12T U4253 ( .A1(n4785), .A2(n3330), .ZN(n3335) );
  ND2XD0BWP12T U4254 ( .A1(n4542), .A2(n5094), .ZN(n3331) );
  CKND2D1BWP12T U4255 ( .A1(n3331), .A2(n5098), .ZN(n3333) );
  INVD1BWP12T U4256 ( .I(n3332), .ZN(n4786) );
  ND2D1BWP12T U4257 ( .A1(n3333), .A2(n4786), .ZN(n3334) );
  ND2D1BWP12T U4258 ( .A1(n3335), .A2(n3334), .ZN(n3339) );
  CKND2D1BWP12T U4259 ( .A1(n4859), .A2(n4843), .ZN(n3336) );
  AOI21D1BWP12T U4260 ( .A1(n3337), .A2(n3336), .B(n5100), .ZN(n4852) );
  TPNR2D2BWP12T U4261 ( .A1(n3339), .A2(n3338), .ZN(n3374) );
  ND2D1BWP12T U4262 ( .A1(n3341), .A2(n278), .ZN(n3343) );
  XNR2D1BWP12T U4263 ( .A1(n3343), .A2(n3342), .ZN(n4265) );
  OAI21D1BWP12T U4264 ( .A1(n4244), .A2(n3345), .B(n3344), .ZN(n3348) );
  CKND0BWP12T U4265 ( .I(n3346), .ZN(n3600) );
  CKND2D1BWP12T U4266 ( .A1(n3600), .A2(n3599), .ZN(n3347) );
  XNR2D1BWP12T U4267 ( .A1(n3348), .A2(n3347), .ZN(n4321) );
  INVD1BWP12T U4268 ( .I(n3557), .ZN(n4778) );
  TPND2D0BWP12T U4269 ( .A1(n3618), .A2(n3352), .ZN(n3354) );
  AOI21D1BWP12T U4270 ( .A1(n3621), .A2(n3352), .B(n3351), .ZN(n3353) );
  OAI21D1BWP12T U4271 ( .A1(n5082), .A2(n3354), .B(n3353), .ZN(n3356) );
  CKND2D1BWP12T U4272 ( .A1(n3366), .A2(n3627), .ZN(n3355) );
  XNR2XD1BWP12T U4273 ( .A1(n3356), .A2(n3355), .ZN(n4398) );
  CKND2D1BWP12T U4274 ( .A1(n4398), .A2(n5088), .ZN(n3369) );
  TPNR2D0BWP12T U4275 ( .A1(n3358), .A2(n3357), .ZN(n3363) );
  CKND2D0BWP12T U4276 ( .A1(n3649), .A2(n3359), .ZN(n3361) );
  TPOAI21D0BWP12T U4277 ( .A1(n3361), .A2(n4486), .B(n3360), .ZN(n3362) );
  NR2D1BWP12T U4278 ( .A1(n3363), .A2(n3362), .ZN(n3365) );
  AN2XD1BWP12T U4279 ( .A1(n3600), .A2(n3599), .Z(n3364) );
  XNR2XD1BWP12T U4280 ( .A1(n3365), .A2(n3364), .ZN(n4956) );
  CKND2D1BWP12T U4281 ( .A1(n4956), .A2(n5093), .ZN(n3368) );
  CKND2D1BWP12T U4282 ( .A1(n4485), .A2(n4103), .ZN(n3367) );
  ND3D1BWP12T U4283 ( .A1(n3369), .A2(n3368), .A3(n3367), .ZN(n3370) );
  TPNR2D2BWP12T U4284 ( .A1(n3371), .A2(n3370), .ZN(n3372) );
  ND3D4BWP12T U4285 ( .A1(n3374), .A2(n3373), .A3(n3372), .ZN(result[5]) );
  OAI21D1BWP12T U4286 ( .A1(n3377), .A2(n3376), .B(n3375), .ZN(n3382) );
  INVD1BWP12T U4287 ( .I(n3378), .ZN(n3380) );
  ND2D1BWP12T U4288 ( .A1(n3380), .A2(n3379), .ZN(n3381) );
  TPND2D0BWP12T U4289 ( .A1(n3528), .A2(n3383), .ZN(n3414) );
  XNR2D1BWP12T U4290 ( .A1(n4971), .A2(n3414), .ZN(n4959) );
  CKND2D1BWP12T U4291 ( .A1(n4959), .A2(n5093), .ZN(n3401) );
  MUX2ND0BWP12T U4292 ( .I0(n4154), .I1(n4153), .S(n4743), .ZN(n3384) );
  OR2XD1BWP12T U4293 ( .A1(n3384), .A2(n4890), .Z(n4595) );
  CKND2D1BWP12T U4294 ( .A1(n4573), .A2(n4888), .ZN(n3388) );
  OAI22D1BWP12T U4295 ( .A1(n4558), .A2(n4566), .B1(n4170), .B2(n4554), .ZN(
        n3387) );
  OAI21D1BWP12T U4296 ( .A1(n4555), .A2(n4521), .B(n4707), .ZN(n3386) );
  NR2D1BWP12T U4297 ( .A1(n4172), .A2(n4206), .ZN(n3385) );
  NR3D1BWP12T U4298 ( .A1(n3387), .A2(n3386), .A3(n3385), .ZN(n3396) );
  AOI21D1BWP12T U4299 ( .A1(n4890), .A2(n3388), .B(n3396), .ZN(n4547) );
  CKND2D1BWP12T U4300 ( .A1(n4547), .A2(n4209), .ZN(n3395) );
  XNR2D0BWP12T U4301 ( .A1(n4448), .A2(n4905), .ZN(n4437) );
  MUX2ND0BWP12T U4302 ( .I0(n5077), .I1(n5076), .S(n4749), .ZN(n3389) );
  NR2D0BWP12T U4303 ( .A1(n3389), .A2(n905), .ZN(n3390) );
  MUX2NXD0BWP12T U4304 ( .I0(n3390), .I1(n5080), .S(n4655), .ZN(n3393) );
  NR2D0BWP12T U4305 ( .A1(n4905), .A2(n5083), .ZN(n3391) );
  OA21XD0BWP12T U4306 ( .A1(n905), .A2(n3391), .B(n4749), .Z(n3392) );
  AOI211D1BWP12T U4307 ( .A1(n4437), .A2(n5078), .B(n3393), .C(n3392), .ZN(
        n3394) );
  OAI211D1BWP12T U4308 ( .A1(n5042), .A2(n4595), .B(n3395), .C(n3394), .ZN(
        n3400) );
  CKND2D1BWP12T U4309 ( .A1(n4539), .A2(n4843), .ZN(n3397) );
  INVD1BWP12T U4310 ( .I(n3396), .ZN(n3407) );
  AOI222D2BWP12T U4311 ( .A1(n3397), .A2(n3407), .B1(n4153), .B2(n4799), .C1(
        n4151), .C2(n4801), .ZN(n4796) );
  ND2D0BWP12T U4312 ( .A1(n3515), .A2(n3398), .ZN(n3405) );
  XNR2XD1BWP12T U4313 ( .A1(n4384), .A2(n3405), .ZN(n4403) );
  MOAI22D1BWP12T U4314 ( .A1(n4796), .A2(n5040), .B1(n4403), .B2(n5088), .ZN(
        n3399) );
  INR3XD1BWP12T U4315 ( .A1(n3401), .B1(n3400), .B2(n3399), .ZN(n3417) );
  INVD1BWP12T U4316 ( .I(n3402), .ZN(n3403) );
  AOI21D1BWP12T U4317 ( .A1(n3534), .A2(n3404), .B(n3403), .ZN(n3406) );
  XOR2XD1BWP12T U4318 ( .A1(n3406), .A2(n3405), .Z(n4484) );
  AOI211D1BWP12T U4319 ( .A1(n3408), .A2(n3407), .B(n4547), .C(n5100), .ZN(
        n4873) );
  MAOI22D2BWP12T U4320 ( .A1(n4484), .A2(n4103), .B1(n4873), .B2(n5063), .ZN(
        n3416) );
  CKND0BWP12T U4321 ( .I(n3410), .ZN(n3413) );
  CKND2D1BWP12T U4322 ( .A1(n4328), .A2(n5090), .ZN(n3415) );
  ND3D1BWP12T U4323 ( .A1(n3417), .A2(n3416), .A3(n3415), .ZN(n3418) );
  INVD1BWP12T U4324 ( .I(n3923), .ZN(n3423) );
  INVD1BWP12T U4325 ( .I(n3419), .ZN(n3546) );
  TPNR2D1BWP12T U4326 ( .A1(n3546), .A2(n3547), .ZN(n3422) );
  TPOAI21D1BWP12T U4327 ( .A1(n3545), .A2(n3547), .B(n300), .ZN(n3421) );
  TPAOI21D2BWP12T U4328 ( .A1(n3423), .A2(n3422), .B(n3421), .ZN(n3427) );
  AN2D1BWP12T U4329 ( .A1(n3425), .A2(n274), .Z(n3426) );
  XNR2XD4BWP12T U4330 ( .A1(n3427), .A2(n3426), .ZN(n5009) );
  ND2D1BWP12T U4331 ( .A1(n5038), .A2(n4039), .ZN(n3984) );
  ND2D1BWP12T U4332 ( .A1(n3937), .A2(n3435), .ZN(n3439) );
  AOI22D1BWP12T U4333 ( .A1(n3939), .A2(n3471), .B1(n3436), .B2(n3469), .ZN(
        n3438) );
  ND2D1BWP12T U4334 ( .A1(n3941), .A2(n3470), .ZN(n3437) );
  ND3D1BWP12T U4335 ( .A1(n3439), .A2(n3438), .A3(n3437), .ZN(n4034) );
  CKND1BWP12T U4336 ( .I(n4034), .ZN(n4781) );
  MUX2D1BWP12T U4337 ( .I0(n4922), .I1(n2818), .S(n5075), .Z(n3962) );
  INVD1BWP12T U4338 ( .I(n3962), .ZN(n3688) );
  MUX2D1BWP12T U4339 ( .I0(n4908), .I1(a[27]), .S(n5075), .Z(n3958) );
  RCAOI22D0BWP12T U4340 ( .A1(n3958), .A2(n3939), .B1(n3940), .B2(n3964), .ZN(
        n3441) );
  CKND2D0BWP12T U4341 ( .A1(n3941), .A2(n4909), .ZN(n3440) );
  OAI211D1BWP12T U4342 ( .A1(n3945), .A2(n3688), .B(n3441), .C(n3440), .ZN(
        n3448) );
  AOI22D1BWP12T U4343 ( .A1(n3951), .A2(n3939), .B1(n3940), .B2(n3953), .ZN(
        n3443) );
  CKND2D1BWP12T U4344 ( .A1(n3941), .A2(n3960), .ZN(n3442) );
  OAI211D1BWP12T U4345 ( .A1(n3945), .A2(n3444), .B(n3443), .C(n3442), .ZN(
        n3900) );
  AOI22D1BWP12T U4346 ( .A1(n3458), .A2(n3939), .B1(n3940), .B2(n3459), .ZN(
        n3446) );
  CKND2D1BWP12T U4347 ( .A1(n3941), .A2(n3954), .ZN(n3445) );
  OAI211D1BWP12T U4348 ( .A1(n3945), .A2(n3447), .B(n3446), .C(n3445), .ZN(
        n4033) );
  AOI222D1BWP12T U4349 ( .A1(n3448), .A2(n4801), .B1(n3900), .B2(n4799), .C1(
        n4033), .C2(n4797), .ZN(n4804) );
  OAI21D1BWP12T U4350 ( .A1(n4781), .A2(n3556), .B(n4804), .ZN(n3449) );
  HA1D1BWP12T U4351 ( .A(n4636), .B(n3450), .CO(n2851), .S(n4457) );
  INVD1BWP12T U4352 ( .I(n4457), .ZN(n3477) );
  OAI21D0BWP12T U4353 ( .A1(n4933), .A2(n5083), .B(n5081), .ZN(n3454) );
  MUX2ND0BWP12T U4354 ( .I0(n5077), .I1(n5076), .S(n4727), .ZN(n3451) );
  NR2D0BWP12T U4355 ( .A1(n3451), .A2(n905), .ZN(n3452) );
  MUX2ND0BWP12T U4356 ( .I0(n3452), .I1(n5080), .S(n4636), .ZN(n3453) );
  AOI211XD0BWP12T U4357 ( .A1(n4727), .A2(n3454), .B(n3763), .C(n3453), .ZN(
        n3476) );
  OAI21D1BWP12T U4358 ( .A1(n3643), .A2(n4743), .B(n3509), .ZN(n4864) );
  OAI22D1BWP12T U4359 ( .A1(n3954), .A2(n3957), .B1(n3457), .B2(n3963), .ZN(
        n3461) );
  OAI22D1BWP12T U4360 ( .A1(n3459), .A2(n3959), .B1(n3458), .B2(n3961), .ZN(
        n3460) );
  NR2D1BWP12T U4361 ( .A1(n3461), .A2(n3460), .ZN(n4064) );
  OAI22D1BWP12T U4362 ( .A1(n3964), .A2(n3959), .B1(n3962), .B2(n3963), .ZN(
        n3464) );
  OAI22D0BWP12T U4363 ( .A1(n3958), .A2(n3961), .B1(n4909), .B2(n3462), .ZN(
        n3463) );
  TPNR2D0BWP12T U4364 ( .A1(n3817), .A2(n4933), .ZN(n4470) );
  OAI22D1BWP12T U4365 ( .A1(n3952), .A2(n3963), .B1(n3951), .B2(n3961), .ZN(
        n3466) );
  OAI22D1BWP12T U4366 ( .A1(n3953), .A2(n3959), .B1(n3960), .B2(n3957), .ZN(
        n3465) );
  NR2D1BWP12T U4367 ( .A1(n3466), .A2(n3465), .ZN(n3901) );
  INVD0BWP12T U4368 ( .I(n3901), .ZN(n3467) );
  NR2D1BWP12T U4369 ( .A1(n3468), .A2(n4848), .ZN(n3474) );
  OAI22D1BWP12T U4370 ( .A1(n3470), .A2(n3957), .B1(n3469), .B2(n3959), .ZN(
        n3473) );
  NR2D1BWP12T U4371 ( .A1(n3471), .A2(n3961), .ZN(n3472) );
  TPNR3D2BWP12T U4372 ( .A1(n3474), .A2(n3473), .A3(n3472), .ZN(n4586) );
  AOI22D1BWP12T U4373 ( .A1(n3903), .A2(n4864), .B1(n4600), .B2(n4167), .ZN(
        n3475) );
  OAI211D1BWP12T U4374 ( .A1(n4420), .A2(n3477), .B(n3476), .C(n3475), .ZN(
        n3478) );
  FA1D2BWP12T U4375 ( .A(n4727), .B(n4933), .CI(n3480), .CO(n2848), .S(n4374)
         );
  XNR2D2BWP12T U4376 ( .A1(n3486), .A2(n4300), .ZN(n3492) );
  AOI21D1BWP12T U4377 ( .A1(n4668), .A2(n3490), .B(n3489), .ZN(n3491) );
  RCOAI21D2BWP12T U4378 ( .A1(n3492), .A2(n4260), .B(n3491), .ZN(v) );
  INVD1BWP12T U4379 ( .I(n3493), .ZN(n3494) );
  IND2XD1BWP12T U4380 ( .A1(n3495), .B1(n3494), .ZN(n3497) );
  XOR2D2BWP12T U4381 ( .A1(n3497), .A2(n3496), .Z(n4268) );
  CKND2D1BWP12T U4382 ( .A1(n3499), .A2(n4032), .ZN(n3501) );
  TPND2D0BWP12T U4383 ( .A1(n4251), .A2(n3754), .ZN(n3500) );
  ND2D1BWP12T U4384 ( .A1(n3501), .A2(n3500), .ZN(n3809) );
  OAI22D1BWP12T U4385 ( .A1(n3502), .A2(n4554), .B1(n4208), .B2(n4521), .ZN(
        n3506) );
  OAI21D1BWP12T U4386 ( .A1(n3503), .A2(n4206), .B(n4707), .ZN(n3505) );
  NR2D1BWP12T U4387 ( .A1(n4207), .A2(n4566), .ZN(n3504) );
  OAI22D1BWP12T U4388 ( .A1(n3823), .A2(n4521), .B1(n3824), .B2(n4566), .ZN(
        n4532) );
  NR2D1BWP12T U4389 ( .A1(n4532), .A2(n4707), .ZN(n3507) );
  OR2XD1BWP12T U4390 ( .A1(n3518), .A2(n3507), .Z(n3508) );
  OAI21D1BWP12T U4391 ( .A1(n3809), .A2(n4045), .B(n3508), .ZN(n4842) );
  TPOAI21D1BWP12T U4392 ( .A1(n3510), .A2(n4156), .B(n3509), .ZN(n3512) );
  INVD0BWP12T U4393 ( .I(n3518), .ZN(n3511) );
  AOI21D1BWP12T U4394 ( .A1(n3512), .A2(n3511), .B(n5100), .ZN(n4868) );
  OR2D0BWP12T U4395 ( .A1(n4868), .A2(n5063), .Z(n3513) );
  AOI21D1BWP12T U4396 ( .A1(n4384), .A2(n3515), .B(n3514), .ZN(n3517) );
  CKND2D1BWP12T U4397 ( .A1(n3536), .A2(n3535), .ZN(n3516) );
  XOR2XD1BWP12T U4398 ( .A1(n3517), .A2(n3516), .Z(n4388) );
  CKND2D1BWP12T U4399 ( .A1(n4573), .A2(n4532), .ZN(n3519) );
  AOI21D1BWP12T U4400 ( .A1(n4890), .A2(n3519), .B(n3518), .ZN(n4574) );
  MUX2ND0BWP12T U4401 ( .I0(n5077), .I1(n5076), .S(n4765), .ZN(n3521) );
  NR2D0BWP12T U4402 ( .A1(n3521), .A2(n905), .ZN(n3522) );
  MUX2ND0BWP12T U4403 ( .I0(n3522), .I1(n5080), .S(n3523), .ZN(n3525) );
  AOI21D0BWP12T U4404 ( .A1(n3523), .A2(n4633), .B(n905), .ZN(n3524) );
  AOI21D1BWP12T U4405 ( .A1(n4971), .A2(n3528), .B(n3527), .ZN(n3531) );
  ND2D1BWP12T U4406 ( .A1(n351), .A2(n3529), .ZN(n3530) );
  XOR2XD1BWP12T U4407 ( .A1(n3531), .A2(n3530), .Z(n4963) );
  CKND2D1BWP12T U4408 ( .A1(n4963), .A2(n5093), .ZN(n3540) );
  AOI21D1BWP12T U4409 ( .A1(n3534), .A2(n3533), .B(n3532), .ZN(n3538) );
  ND2D1BWP12T U4410 ( .A1(n3536), .A2(n3535), .ZN(n3537) );
  XOR2XD1BWP12T U4411 ( .A1(n3538), .A2(n3537), .Z(n4483) );
  CKND2D1BWP12T U4412 ( .A1(n4483), .A2(n4103), .ZN(n3539) );
  OAI21D1BWP12T U4413 ( .A1(n3923), .A2(n3546), .B(n3545), .ZN(n3550) );
  INVD1BWP12T U4414 ( .I(n3547), .ZN(n3548) );
  XNR2XD4BWP12T U4415 ( .A1(n3550), .A2(n358), .ZN(n4299) );
  ND2D4BWP12T U4416 ( .A1(n4299), .A2(n5085), .ZN(n3597) );
  ND2D1BWP12T U4417 ( .A1(n4946), .A2(n5093), .ZN(n3595) );
  ND2D1BWP12T U4418 ( .A1(n4362), .A2(n5090), .ZN(n3594) );
  OAI22D1BWP12T U4419 ( .A1(n3559), .A2(n3558), .B1(n3557), .B2(n3556), .ZN(
        n3564) );
  AOI22D0BWP12T U4420 ( .A1(n3570), .A2(n3939), .B1(n3940), .B2(n3835), .ZN(
        n3562) );
  TPND2D0BWP12T U4421 ( .A1(n3937), .A2(n3834), .ZN(n3561) );
  TPND2D0BWP12T U4422 ( .A1(n3941), .A2(n3569), .ZN(n3560) );
  TPAOI31D0BWP12T U4423 ( .A1(n3562), .A2(n3561), .A3(n3560), .B(n3818), .ZN(
        n3563) );
  AOI211D1BWP12T U4424 ( .A1(n4797), .A2(n3565), .B(n3564), .C(n3563), .ZN(
        n4803) );
  OAI22D1BWP12T U4425 ( .A1(n3984), .A2(n3823), .B1(n4803), .B2(n5040), .ZN(
        n3588) );
  TPOAI21D0BWP12T U4426 ( .A1(n3843), .A2(n3567), .B(n4874), .ZN(n4850) );
  CKND1BWP12T U4427 ( .I(n3568), .ZN(n3574) );
  OAI22D0BWP12T U4428 ( .A1(n3570), .A2(n3961), .B1(n3569), .B2(n3957), .ZN(
        n3572) );
  OAI22D1BWP12T U4429 ( .A1(n3835), .A2(n3959), .B1(n3834), .B2(n3963), .ZN(
        n3571) );
  RCOAI21D0BWP12T U4430 ( .A1(n3572), .A2(n3571), .B(n4158), .ZN(n3573) );
  OAI211D1BWP12T U4431 ( .A1(n3574), .A2(n3968), .B(n4573), .C(n3573), .ZN(
        n3577) );
  NR2D0BWP12T U4432 ( .A1(n3575), .A2(n3969), .ZN(n3576) );
  AOI211D1BWP12T U4433 ( .A1(n3972), .A2(n3578), .B(n3577), .C(n3576), .ZN(
        n4589) );
  MUX2ND0BWP12T U4434 ( .I0(n5077), .I1(n5076), .S(n4730), .ZN(n3579) );
  NR2D0BWP12T U4435 ( .A1(n3579), .A2(n905), .ZN(n3580) );
  MUX2NXD0BWP12T U4436 ( .I0(n3580), .I1(n5080), .S(n4664), .ZN(n3583) );
  NR2D1BWP12T U4437 ( .A1(n4909), .A2(n5083), .ZN(n3581) );
  OA21XD0BWP12T U4438 ( .A1(n905), .A2(n3581), .B(n4730), .Z(n3582) );
  AOI211D1BWP12T U4439 ( .A1(n4589), .A2(n4167), .B(n3583), .C(n3582), .ZN(
        n3586) );
  HA1D1BWP12T U4440 ( .A(n4664), .B(n3584), .CO(n3450), .S(n4434) );
  ND2D1BWP12T U4441 ( .A1(n4434), .A2(n5078), .ZN(n3585) );
  OAI211D1BWP12T U4442 ( .A1(n5063), .A2(n4850), .B(n3586), .C(n3585), .ZN(
        n3587) );
  AOI211D1BWP12T U4443 ( .A1(n4416), .A2(n5088), .B(n3588), .C(n3587), .ZN(
        n3593) );
  ND2D1BWP12T U4444 ( .A1(n4514), .A2(n4103), .ZN(n3592) );
  AN4D2BWP12T U4445 ( .A1(n3595), .A2(n3594), .A3(n3593), .A4(n3592), .Z(n3596) );
  ND2D4BWP12T U4446 ( .A1(n3597), .A2(n3596), .ZN(result[29]) );
  CKND2D1BWP12T U4447 ( .A1(n4034), .A2(n4094), .ZN(n3616) );
  OR2D0BWP12T U4448 ( .A1(n4046), .A2(n5063), .Z(n3615) );
  MUX2ND0BWP12T U4449 ( .I0(n5077), .I1(n5076), .S(n4748), .ZN(n3607) );
  NR2D0BWP12T U4450 ( .A1(n3607), .A2(n905), .ZN(n3608) );
  MUX2NXD0BWP12T U4451 ( .I0(n3608), .I1(n5080), .S(n4631), .ZN(n3611) );
  NR2D1BWP12T U4452 ( .A1(n4931), .A2(n5083), .ZN(n3609) );
  OA21XD0BWP12T U4453 ( .A1(n905), .A2(n3609), .B(n4748), .Z(n3610) );
  AO211D1BWP12T U4454 ( .A1(n4432), .A2(n5078), .B(n3611), .C(n3610), .Z(n3612) );
  NR2D1BWP12T U4455 ( .A1(n3613), .A2(n3612), .ZN(n3614) );
  ND3D1BWP12T U4456 ( .A1(n3616), .A2(n3615), .A3(n3614), .ZN(n3617) );
  AOI21D1BWP12T U4457 ( .A1(n5090), .A2(n4324), .B(n3617), .ZN(n3660) );
  CKND2D0BWP12T U4458 ( .A1(n3618), .A2(n3620), .ZN(n3623) );
  TPAOI21D0BWP12T U4459 ( .A1(n3621), .A2(n3620), .B(n3619), .ZN(n3622) );
  OAI21D1BWP12T U4460 ( .A1(n5082), .A2(n3623), .B(n3622), .ZN(n3625) );
  ND2XD0BWP12T U4461 ( .A1(n3633), .A2(n3632), .ZN(n3624) );
  XNR2XD1BWP12T U4462 ( .A1(n3625), .A2(n3624), .ZN(n4390) );
  TPNR3D0BWP12T U4463 ( .A1(n4102), .A2(n3626), .A3(n3628), .ZN(n3631) );
  OAI21D0BWP12T U4464 ( .A1(n3629), .A2(n3628), .B(n3627), .ZN(n3630) );
  NR2D1BWP12T U4465 ( .A1(n3631), .A2(n3630), .ZN(n3635) );
  CKAN2D1BWP12T U4466 ( .A1(n3633), .A2(n3632), .Z(n3634) );
  XNR2XD1BWP12T U4467 ( .A1(n3635), .A2(n3634), .ZN(n4482) );
  AOI22D1BWP12T U4468 ( .A1(n5088), .A2(n4390), .B1(n4482), .B2(n4103), .ZN(
        n3658) );
  OAI22D1BWP12T U4469 ( .A1(n3637), .A2(n4206), .B1(n3636), .B2(n4566), .ZN(
        n3642) );
  OAI21D0BWP12T U4470 ( .A1(n3638), .A2(n4521), .B(n4707), .ZN(n3641) );
  NR2D1BWP12T U4471 ( .A1(n3639), .A2(n4554), .ZN(n3640) );
  NR3D1BWP12T U4472 ( .A1(n3642), .A2(n3641), .A3(n3640), .ZN(n4853) );
  AOI22D1BWP12T U4473 ( .A1(n4039), .A2(n4037), .B1(n4036), .B2(n4556), .ZN(
        n3644) );
  OAI21D1BWP12T U4474 ( .A1(n3643), .A2(n3902), .B(n3644), .ZN(n4863) );
  AOI21D1BWP12T U4475 ( .A1(n4863), .A2(n4573), .B(n4605), .ZN(n4854) );
  INVD0BWP12T U4476 ( .I(n4538), .ZN(n3646) );
  AO21D1BWP12T U4477 ( .A1(n5094), .A2(n3646), .B(n3645), .Z(n3648) );
  INVD1BWP12T U4478 ( .I(n4853), .ZN(n3647) );
  ND2D1BWP12T U4479 ( .A1(n3648), .A2(n3647), .ZN(n3656) );
  AOI211D1BWP12T U4480 ( .A1(n4843), .A2(n4538), .B(n4853), .C(n4891), .ZN(
        n4575) );
  TPAOI21D0BWP12T U4481 ( .A1(n3652), .A2(n3651), .B(n3650), .ZN(n3653) );
  AOI22D1BWP12T U4482 ( .A1(n4575), .A2(n4209), .B1(n4964), .B2(n5093), .ZN(
        n3655) );
  ND4D1BWP12T U4483 ( .A1(n3658), .A2(n3657), .A3(n3656), .A4(n3655), .ZN(
        n3659) );
  ND2D1BWP12T U4484 ( .A1(n3662), .A2(n3661), .ZN(n3664) );
  INVD1BWP12T U4485 ( .I(n3667), .ZN(n3668) );
  TPND2D1BWP12T U4486 ( .A1(n291), .A2(n3668), .ZN(n3670) );
  TPND2D1BWP12T U4487 ( .A1(n3670), .A2(n292), .ZN(n3675) );
  XNR2XD4BWP12T U4488 ( .A1(n3675), .A2(n3674), .ZN(n4305) );
  NR2XD0BWP12T U4489 ( .A1(n3929), .A2(n3723), .ZN(n3677) );
  TPND2D0BWP12T U4490 ( .A1(n3930), .A2(n3677), .ZN(n3679) );
  TPOAI21D0BWP12T U4491 ( .A1(n3932), .A2(n3723), .B(n3805), .ZN(n3676) );
  AOI21D1BWP12T U4492 ( .A1(n3933), .A2(n3677), .B(n3676), .ZN(n3678) );
  OAI21D1BWP12T U4493 ( .A1(n4353), .A2(n3679), .B(n3678), .ZN(n3682) );
  ND2D1BWP12T U4494 ( .A1(n3681), .A2(n3680), .ZN(n3724) );
  XNR2XD1BWP12T U4495 ( .A1(n3682), .A2(n3724), .ZN(n4311) );
  INVD1BWP12T U4496 ( .I(n4311), .ZN(n3728) );
  OAI21D1BWP12T U4497 ( .A1(n3997), .A2(n3683), .B(n3831), .ZN(n3686) );
  CKND2D1BWP12T U4498 ( .A1(n3685), .A2(n3684), .ZN(n3697) );
  CKND0BWP12T U4499 ( .I(n4806), .ZN(n3693) );
  INVD1BWP12T U4500 ( .I(n3687), .ZN(n3691) );
  AOI211D1BWP12T U4501 ( .A1(n3691), .A2(n4799), .B(n3690), .C(n3689), .ZN(
        n3692) );
  OAI21D1BWP12T U4502 ( .A1(n3693), .A2(n3758), .B(n3692), .ZN(n4814) );
  OA21D1BWP12T U4503 ( .A1(n3694), .A2(n4611), .B(n4814), .Z(n3721) );
  INVD1BWP12T U4504 ( .I(n4476), .ZN(n3746) );
  CKND2D1BWP12T U4505 ( .A1(n4505), .A2(n4103), .ZN(n3720) );
  OAI22D0BWP12T U4506 ( .A1(n3964), .A2(n3961), .B1(n3962), .B2(n3957), .ZN(
        n3699) );
  NR2D0BWP12T U4507 ( .A1(n3951), .A2(n3959), .ZN(n3698) );
  RCAOI211D0BWP12T U4508 ( .A1(n3701), .A2(n3700), .B(n3699), .C(n3698), .ZN(
        n3705) );
  TPND3D0BWP12T U4509 ( .A1(n3703), .A2(n3702), .A3(n3761), .ZN(n3704) );
  OAI211D0BWP12T U4510 ( .A1(n3705), .A2(n4611), .B(n4573), .C(n3704), .ZN(
        n3706) );
  AOI21D1BWP12T U4511 ( .A1(n4580), .A2(n4843), .B(n3706), .ZN(n4620) );
  ND2D1BWP12T U4512 ( .A1(n4874), .A2(n5099), .ZN(n3845) );
  AOI21D1BWP12T U4513 ( .A1(n4877), .A2(n4847), .B(n3845), .ZN(n3718) );
  TPNR2D0BWP12T U4514 ( .A1(n3708), .A2(n3707), .ZN(n3709) );
  CKND2D1BWP12T U4515 ( .A1(n3709), .A2(n4426), .ZN(n3710) );
  XOR2XD1BWP12T U4516 ( .A1(n3710), .A2(n4922), .Z(n4435) );
  OAI21D1BWP12T U4517 ( .A1(n4922), .A2(n5083), .B(n5081), .ZN(n3711) );
  AOI22D1BWP12T U4518 ( .A1(n4435), .A2(n5078), .B1(b[26]), .B2(n3711), .ZN(
        n3715) );
  MUX2ND0BWP12T U4519 ( .I0(n5045), .I1(n5044), .S(b[26]), .ZN(n3712) );
  TPND2D0BWP12T U4520 ( .A1(n3712), .A2(n5081), .ZN(n3713) );
  MUX2NXD0BWP12T U4521 ( .I0(n3713), .I1(n5048), .S(n4666), .ZN(n3714) );
  OAI211D1BWP12T U4522 ( .A1(n4543), .A2(n3716), .B(n3715), .C(n3714), .ZN(
        n3717) );
  AOI211D1BWP12T U4523 ( .A1(n4620), .A2(n4167), .B(n3718), .C(n3717), .ZN(
        n3719) );
  OAI211D1BWP12T U4524 ( .A1(n3721), .A2(n5040), .B(n3720), .C(n3719), .ZN(
        n3722) );
  AOI21D1BWP12T U4525 ( .A1(n5088), .A2(n4377), .B(n3722), .ZN(n3727) );
  TPND2D1BWP12T U4526 ( .A1(n4993), .A2(n5093), .ZN(n3726) );
  TPOAI21D8BWP12T U4527 ( .A1(n4305), .A2(n4260), .B(n3729), .ZN(result[26])
         );
  TPOAI21D1BWP12T U4528 ( .A1(n3732), .A2(n3731), .B(n3730), .ZN(n3737) );
  CKND0BWP12T U4529 ( .I(n3733), .ZN(n3735) );
  ND2D1BWP12T U4530 ( .A1(n3735), .A2(n3734), .ZN(n3736) );
  XNR2XD4BWP12T U4531 ( .A1(n3737), .A2(n3736), .ZN(n4288) );
  TPND2D0BWP12T U4532 ( .A1(n3738), .A2(n3787), .ZN(n3742) );
  INVD1BWP12T U4533 ( .I(n3739), .ZN(n3786) );
  AOI21D1BWP12T U4534 ( .A1(n3740), .A2(n3787), .B(n3786), .ZN(n3741) );
  OAI21D1BWP12T U4535 ( .A1(n4985), .A2(n3742), .B(n3741), .ZN(n3745) );
  XNR2XD1BWP12T U4536 ( .A1(n3745), .A2(n3789), .ZN(n4979) );
  INVD1BWP12T U4537 ( .I(n4979), .ZN(n3792) );
  XNR2D1BWP12T U4538 ( .A1(n3746), .A2(n3785), .ZN(n4507) );
  INR2XD0BWP12T U4539 ( .A1(n4742), .B1(n4518), .ZN(n3747) );
  INVD1BWP12T U4540 ( .I(n3747), .ZN(n3751) );
  NR2D1BWP12T U4541 ( .A1(n4517), .A2(n3748), .ZN(n3749) );
  INR2D1BWP12T U4542 ( .A1(n4685), .B1(n3749), .ZN(n3750) );
  ND2D1BWP12T U4543 ( .A1(n3751), .A2(n3750), .ZN(n3769) );
  AOI22D1BWP12T U4544 ( .A1(n3755), .A2(n3754), .B1(n3753), .B2(n4801), .ZN(
        n3757) );
  OAI211D1BWP12T U4545 ( .A1(n3758), .A2(n4093), .B(n3757), .C(n3756), .ZN(
        n4808) );
  INVD1BWP12T U4546 ( .I(n4808), .ZN(n3765) );
  TPND3D0BWP12T U4547 ( .A1(n4573), .A2(n3902), .A3(n4583), .ZN(n3759) );
  AO222D1BWP12T U4548 ( .A1(n3762), .A2(n3761), .B1(n3760), .B2(n4158), .C1(
        n3759), .C2(n4890), .Z(n4618) );
  NR2D1BWP12T U4549 ( .A1(n4618), .A2(n5042), .ZN(n3764) );
  AOI211D1BWP12T U4550 ( .A1(n3765), .A2(n5094), .B(n3764), .C(n3763), .ZN(
        n3779) );
  AOI22D1BWP12T U4551 ( .A1(n3767), .A2(n4569), .B1(n3766), .B2(n4624), .ZN(
        n3768) );
  ND2D1BWP12T U4552 ( .A1(n3769), .A2(n3768), .ZN(n4858) );
  OAI21D1BWP12T U4553 ( .A1(n4924), .A2(n5083), .B(n5081), .ZN(n3772) );
  AOI22D1BWP12T U4554 ( .A1(n4427), .A2(n5078), .B1(n336), .B2(n3772), .ZN(
        n3776) );
  MUX2ND0BWP12T U4555 ( .I0(n5045), .I1(n5044), .S(n336), .ZN(n3773) );
  TPND2D0BWP12T U4556 ( .A1(n3773), .A2(n5081), .ZN(n3774) );
  MUX2NXD0BWP12T U4557 ( .I0(n3774), .I1(n5048), .S(n1342), .ZN(n3775) );
  OA211D1BWP12T U4558 ( .A1(n4858), .A2(n3777), .B(n3776), .C(n3775), .Z(n3778) );
  OAI211D1BWP12T U4559 ( .A1(n3899), .A2(n4824), .B(n3779), .C(n3778), .ZN(
        n3780) );
  AOI21D1BWP12T U4560 ( .A1(n4103), .A2(n4507), .B(n3780), .ZN(n3791) );
  AOI22D1BWP12T U4561 ( .A1(n5088), .A2(n4410), .B1(n4330), .B2(n5090), .ZN(
        n3790) );
  OAI211D1BWP12T U4562 ( .A1(n4954), .A2(n3792), .B(n3791), .C(n3790), .ZN(
        n3793) );
  AO21D4BWP12T U4563 ( .A1(n4288), .A2(n5085), .B(n3793), .Z(result[19]) );
  TPAOI21D1BWP12T U4564 ( .A1(n291), .A2(n3795), .B(n302), .ZN(n3800) );
  IND2D1BWP12T U4565 ( .A1(n3798), .B1(n3797), .ZN(n3799) );
  XNR2XD4BWP12T U4566 ( .A1(n3800), .A2(n3799), .ZN(n4304) );
  ND2XD0BWP12T U4567 ( .A1(n3930), .A2(n3802), .ZN(n3804) );
  AOI21D1BWP12T U4568 ( .A1(n3933), .A2(n3802), .B(n3801), .ZN(n3803) );
  OAI21D1BWP12T U4569 ( .A1(n4353), .A2(n3804), .B(n3803), .ZN(n3807) );
  CKND2D1BWP12T U4570 ( .A1(n3806), .A2(n3805), .ZN(n3808) );
  XOR2XD1BWP12T U4571 ( .A1(n3991), .A2(n3808), .Z(n4948) );
  CKND2D1BWP12T U4572 ( .A1(n3809), .A2(n4045), .ZN(n3827) );
  INVD1BWP12T U4573 ( .I(n3810), .ZN(n3836) );
  TPNR2D0BWP12T U4574 ( .A1(n3945), .A2(n3836), .ZN(n3815) );
  CKND1BWP12T U4575 ( .I(n3811), .ZN(n3837) );
  OAI22D0BWP12T U4576 ( .A1(n3813), .A2(n3837), .B1(n3812), .B2(n3835), .ZN(
        n3814) );
  AOI211D1BWP12T U4577 ( .A1(n3941), .A2(n3816), .B(n3815), .C(n3814), .ZN(
        n3819) );
  OAI21D0BWP12T U4578 ( .A1(n3819), .A2(n3818), .B(n3817), .ZN(n3820) );
  AOI31D1BWP12T U4579 ( .A1(n4799), .A2(n3822), .A3(n3821), .B(n3820), .ZN(
        n3826) );
  MUX2ND0BWP12T U4580 ( .I0(n3824), .I1(n3823), .S(n4742), .ZN(n3825) );
  AOI22D1BWP12T U4581 ( .A1(n3827), .A2(n3826), .B1(n4158), .B2(n3825), .ZN(
        n4815) );
  AOI22D1BWP12T U4582 ( .A1(n4509), .A2(n4103), .B1(n4408), .B2(n5088), .ZN(
        n3859) );
  INVD0BWP12T U4583 ( .I(n3833), .ZN(n3841) );
  OAI22D0BWP12T U4584 ( .A1(n3835), .A2(n3961), .B1(n3834), .B2(n3957), .ZN(
        n3839) );
  OAI22D0BWP12T U4585 ( .A1(n3837), .A2(n3959), .B1(n3836), .B2(n3963), .ZN(
        n3838) );
  OAI21D1BWP12T U4586 ( .A1(n3839), .A2(n3838), .B(n4158), .ZN(n3840) );
  OAI211D1BWP12T U4587 ( .A1(n3841), .A2(n3968), .B(n4573), .C(n3840), .ZN(
        n3842) );
  AOI21D1BWP12T U4588 ( .A1(n4843), .A2(n4581), .B(n3842), .ZN(n4619) );
  RCAOI21D0BWP12T U4589 ( .A1(n4685), .A2(n3844), .B(n3843), .ZN(n4876) );
  NR2D1BWP12T U4590 ( .A1(n4876), .A2(n3845), .ZN(n3857) );
  XNR2D1BWP12T U4591 ( .A1(n3848), .A2(n3847), .ZN(n4441) );
  INVD1BWP12T U4592 ( .I(n4441), .ZN(n3855) );
  TPND2D0BWP12T U4593 ( .A1(n3849), .A2(n4532), .ZN(n3854) );
  OAI21D1BWP12T U4594 ( .A1(n4699), .A2(n5083), .B(n5081), .ZN(n3852) );
  AOI21D1BWP12T U4595 ( .A1(n4739), .A2(n3852), .B(n3851), .ZN(n3853) );
  OAI211D1BWP12T U4596 ( .A1(n3855), .A2(n4420), .B(n3854), .C(n3853), .ZN(
        n3856) );
  AOI211D1BWP12T U4597 ( .A1(n4619), .A2(n4167), .B(n3857), .C(n3856), .ZN(
        n3858) );
  OAI211D1BWP12T U4598 ( .A1(n4815), .A2(n5040), .B(n3859), .C(n3858), .ZN(
        n3860) );
  IOA21D2BWP12T U4599 ( .A1(n5090), .A2(n4312), .B(n3861), .ZN(n3862) );
  INVD1P75BWP12T U4600 ( .I(n3862), .ZN(n3863) );
  RCOAI21D4BWP12T U4601 ( .A1(n4304), .A2(n4260), .B(n3863), .ZN(result[25])
         );
  INVD1BWP12T U4602 ( .I(n3867), .ZN(n3869) );
  AN2XD2BWP12T U4603 ( .A1(n3869), .A2(n3868), .Z(n3870) );
  XNR2D2BWP12T U4604 ( .A1(n3871), .A2(n3870), .ZN(n4295) );
  ND2D1BWP12T U4605 ( .A1(n3875), .A2(n3874), .ZN(n3882) );
  ND2D1BWP12T U4606 ( .A1(n4358), .A2(n5090), .ZN(n3918) );
  ND2XD0BWP12T U4607 ( .A1(n3876), .A2(n3878), .ZN(n3881) );
  AOI21D1BWP12T U4608 ( .A1(n3879), .A2(n3878), .B(n3877), .ZN(n3880) );
  OAI21D1BWP12T U4609 ( .A1(n4985), .A2(n3881), .B(n3880), .ZN(n3883) );
  ND2D1BWP12T U4610 ( .A1(n4989), .A2(n5093), .ZN(n3917) );
  INVD1BWP12T U4611 ( .I(n3884), .ZN(n3885) );
  AOI21D1BWP12T U4612 ( .A1(n3887), .A2(n3886), .B(n3885), .ZN(n3890) );
  TPND2D0BWP12T U4613 ( .A1(n3889), .A2(n3888), .ZN(n3913) );
  XOR2XD1BWP12T U4614 ( .A1(n3890), .A2(n3913), .Z(n4501) );
  MUX2ND0BWP12T U4615 ( .I0(n5077), .I1(n5076), .S(n4729), .ZN(n3893) );
  NR2D0BWP12T U4616 ( .A1(n3893), .A2(n905), .ZN(n3894) );
  MUX2ND0BWP12T U4617 ( .I0(n3894), .I1(n5080), .S(n4651), .ZN(n3897) );
  NR2D0BWP12T U4618 ( .A1(n4915), .A2(n5083), .ZN(n3895) );
  OA21XD0BWP12T U4619 ( .A1(n905), .A2(n3895), .B(n4729), .Z(n3896) );
  AOI211D1BWP12T U4620 ( .A1(n4445), .A2(n5078), .B(n3897), .C(n3896), .ZN(
        n3898) );
  OAI211D1BWP12T U4621 ( .A1(n4538), .A2(n3899), .B(n4165), .C(n3898), .ZN(
        n3906) );
  AOI222D1BWP12T U4622 ( .A1(n3900), .A2(n4801), .B1(n4034), .B2(n4797), .C1(
        n4033), .C2(n4799), .ZN(n4805) );
  AOI22D1BWP12T U4623 ( .A1(n3903), .A2(n4863), .B1(n4601), .B2(n4167), .ZN(
        n3904) );
  OAI21D1BWP12T U4624 ( .A1(n4805), .A2(n5040), .B(n3904), .ZN(n3905) );
  AOI211D1BWP12T U4625 ( .A1(n4501), .A2(n4103), .B(n3906), .C(n3905), .ZN(
        n3916) );
  CKND2D1BWP12T U4626 ( .A1(n3907), .A2(n3909), .ZN(n3912) );
  AOI21D1BWP12T U4627 ( .A1(n3910), .A2(n3909), .B(n3908), .ZN(n3911) );
  CKND2D1BWP12T U4628 ( .A1(n4372), .A2(n5088), .ZN(n3915) );
  AN4XD1BWP12T U4629 ( .A1(n3918), .A2(n3917), .A3(n3916), .A4(n3915), .Z(
        n3919) );
  TPOAI21D2BWP12T U4630 ( .A1(n3920), .A2(n4260), .B(n3919), .ZN(result[22])
         );
  TPOAI21D1BWP12T U4631 ( .A1(n3923), .A2(n3922), .B(n3921), .ZN(n3927) );
  INVD1BWP12T U4632 ( .I(n3924), .ZN(n3926) );
  XNR2XD4BWP12T U4633 ( .A1(n3927), .A2(n353), .ZN(n4303) );
  ND2D1BWP12T U4634 ( .A1(n3935), .A2(n3934), .ZN(n3992) );
  ND2D1BWP12T U4635 ( .A1(n4314), .A2(n5090), .ZN(n4003) );
  INVD1BWP12T U4636 ( .I(n3938), .ZN(n4800) );
  AOI22D0BWP12T U4637 ( .A1(n4799), .A2(n4802), .B1(n4800), .B2(n4797), .ZN(
        n3950) );
  AOI22D0BWP12T U4638 ( .A1(n3960), .A2(n3940), .B1(n3939), .B2(n3962), .ZN(
        n3943) );
  TPND2D0BWP12T U4639 ( .A1(n3941), .A2(n3958), .ZN(n3942) );
  OAI211D0BWP12T U4640 ( .A1(n3945), .A2(n3944), .B(n3943), .C(n3942), .ZN(
        n3948) );
  INVD1BWP12T U4641 ( .I(n3946), .ZN(n4798) );
  AOI22D0BWP12T U4642 ( .A1(n3948), .A2(n4801), .B1(n3947), .B2(n4798), .ZN(
        n3949) );
  CKND2D1BWP12T U4643 ( .A1(n3950), .A2(n3949), .ZN(n4839) );
  INVD1BWP12T U4644 ( .I(n4839), .ZN(n3981) );
  OAI22D1BWP12T U4645 ( .A1(n3952), .A2(n3961), .B1(n3951), .B2(n3957), .ZN(
        n3956) );
  OAI22D1BWP12T U4646 ( .A1(n3954), .A2(n3959), .B1(n3953), .B2(n3963), .ZN(
        n3955) );
  NR2D1BWP12T U4647 ( .A1(n3956), .A2(n3955), .ZN(n4612) );
  OAI22D1BWP12T U4648 ( .A1(n3960), .A2(n3959), .B1(n3958), .B2(n3957), .ZN(
        n3966) );
  OAI22D1BWP12T U4649 ( .A1(n3964), .A2(n3963), .B1(n3962), .B2(n3961), .ZN(
        n3965) );
  TPOAI21D0BWP12T U4650 ( .A1(n3966), .A2(n3965), .B(n4158), .ZN(n3967) );
  OAI211D1BWP12T U4651 ( .A1(n4612), .A2(n3968), .B(n4573), .C(n3967), .ZN(
        n3971) );
  INVD1BWP12T U4652 ( .I(n4607), .ZN(n4584) );
  NR2XD0BWP12T U4653 ( .A1(n4584), .A2(n3969), .ZN(n3970) );
  AOI211D1BWP12T U4654 ( .A1(n3972), .A2(n4608), .B(n3971), .C(n3970), .ZN(
        n4590) );
  ND2D1BWP12T U4655 ( .A1(n4590), .A2(n4167), .ZN(n3980) );
  HICIND1BWP12T U4656 ( .A(n4665), .CIN(n3973), .CO(n3584), .S(n4452) );
  MUX2ND0BWP12T U4657 ( .I0(n5077), .I1(n5076), .S(n4733), .ZN(n3974) );
  NR2XD0BWP12T U4658 ( .A1(n3974), .A2(n905), .ZN(n3975) );
  MUX2ND0BWP12T U4659 ( .I0(n3975), .I1(n5080), .S(n4665), .ZN(n3978) );
  TPNR2D0BWP12T U4660 ( .A1(n4459), .A2(n5083), .ZN(n3976) );
  OA21D0BWP12T U4661 ( .A1(n905), .A2(n3976), .B(n4733), .Z(n3977) );
  AOI211D1BWP12T U4662 ( .A1(n4452), .A2(n5078), .B(n3978), .C(n3977), .ZN(
        n3979) );
  OAI211D1BWP12T U4663 ( .A1(n3981), .A2(n5040), .B(n3980), .C(n3979), .ZN(
        n3986) );
  OAI21D1BWP12T U4664 ( .A1(n3983), .A2(n3982), .B(n4874), .ZN(n4871) );
  OAI22D0BWP12T U4665 ( .A1(n3984), .A2(n4173), .B1(n5063), .B2(n4871), .ZN(
        n3985) );
  AOI211XD0BWP12T U4666 ( .A1(n4500), .A2(n4103), .B(n3986), .C(n3985), .ZN(
        n4002) );
  ND2D1BWP12T U4667 ( .A1(n4992), .A2(n5093), .ZN(n4001) );
  ND2D1BWP12T U4668 ( .A1(n4376), .A2(n5088), .ZN(n4000) );
  AN4D2BWP12T U4669 ( .A1(n4003), .A2(n4002), .A3(n4001), .A4(n4000), .Z(n4004) );
  RCOAI21D4BWP12T U4670 ( .A1(n4303), .A2(n4260), .B(n4004), .ZN(result[28])
         );
  TPOAI21D1BWP12T U4671 ( .A1(n4008), .A2(n4007), .B(n4006), .ZN(n4013) );
  INVD0BWP12T U4672 ( .I(n4009), .ZN(n4010) );
  OR2XD1BWP12T U4673 ( .A1(n4011), .A2(n4010), .Z(n4012) );
  XNR2XD4BWP12T U4674 ( .A1(n4013), .A2(n4012), .ZN(n4277) );
  TPND2D2BWP12T U4675 ( .A1(n4277), .A2(n5085), .ZN(n4083) );
  NR2XD0BWP12T U4676 ( .A1(n4014), .A2(n4016), .ZN(n4019) );
  TPOAI21D0BWP12T U4677 ( .A1(n4017), .A2(n4016), .B(n4015), .ZN(n4018) );
  AOI21D1BWP12T U4678 ( .A1(n4971), .A2(n4019), .B(n4018), .ZN(n4022) );
  CKND2D1BWP12T U4679 ( .A1(n4021), .A2(n4020), .ZN(n4076) );
  XOR2XD1BWP12T U4680 ( .A1(n4022), .A2(n4076), .Z(n4950) );
  CKND2D0BWP12T U4681 ( .A1(n4023), .A2(n4025), .ZN(n4028) );
  TPAOI21D0BWP12T U4682 ( .A1(n4026), .A2(n4025), .B(n4024), .ZN(n4027) );
  OAI21D1BWP12T U4683 ( .A1(n4493), .A2(n4028), .B(n4027), .ZN(n4031) );
  ND2D0BWP12T U4684 ( .A1(n4030), .A2(n4029), .ZN(n4055) );
  XNR2XD1BWP12T U4685 ( .A1(n4031), .A2(n4055), .ZN(n4479) );
  AOI22D1BWP12T U4686 ( .A1(n4950), .A2(n5093), .B1(n4103), .B2(n4479), .ZN(
        n4081) );
  MUX2NXD0BWP12T U4687 ( .I0(n4034), .I1(n4033), .S(n4032), .ZN(n4044) );
  CKND0BWP12T U4688 ( .I(n4035), .ZN(n4533) );
  ND2XD0BWP12T U4689 ( .A1(n4533), .A2(n4039), .ZN(n4043) );
  MUX2ND0BWP12T U4690 ( .I0(n4037), .I1(n4036), .S(n4742), .ZN(n4038) );
  CKND2D0BWP12T U4691 ( .A1(n4038), .A2(n4707), .ZN(n4042) );
  AOI222D1BWP12T U4692 ( .A1(n4042), .A2(n4611), .B1(n4041), .B2(n4556), .C1(
        n4040), .C2(n4039), .ZN(n4047) );
  AO21D1BWP12T U4693 ( .A1(n4843), .A2(n4043), .B(n4047), .Z(n4531) );
  OAI21D1BWP12T U4694 ( .A1(n4045), .A2(n4044), .B(n4531), .ZN(n4838) );
  INR2D0BWP12T U4695 ( .A1(n4843), .B1(n4864), .ZN(n4048) );
  TPOAI31D0BWP12T U4696 ( .A1(n4891), .A2(n4048), .A3(n4047), .B(n4046), .ZN(
        n4855) );
  AOI22D1BWP12T U4697 ( .A1(n4838), .A2(n5094), .B1(n5099), .B2(n4855), .ZN(
        n4080) );
  NR2D0BWP12T U4698 ( .A1(n4049), .A2(n4051), .ZN(n4054) );
  OAI21D0BWP12T U4699 ( .A1(n4052), .A2(n4051), .B(n4050), .ZN(n4053) );
  TPAOI21D0BWP12T U4700 ( .A1(n4384), .A2(n4054), .B(n4053), .ZN(n4056) );
  XOR2XD1BWP12T U4701 ( .A1(n4056), .A2(n4055), .Z(n4407) );
  NR2D0BWP12T U4702 ( .A1(n4932), .A2(n5083), .ZN(n4059) );
  OA21XD0BWP12T U4703 ( .A1(n905), .A2(n4059), .B(n4752), .Z(n4063) );
  MUX2ND0BWP12T U4704 ( .I0(n5077), .I1(n5076), .S(n4752), .ZN(n4060) );
  NR2D0BWP12T U4705 ( .A1(n4060), .A2(n905), .ZN(n4061) );
  MUX2NXD0BWP12T U4706 ( .I0(n4061), .I1(n5080), .S(n4680), .ZN(n4062) );
  AOI211D1BWP12T U4707 ( .A1(n4440), .A2(n5078), .B(n4063), .C(n4062), .ZN(
        n4067) );
  MUX2NXD0BWP12T U4708 ( .I0(n4064), .I1(n4586), .S(n4743), .ZN(n4065) );
  NR2XD0BWP12T U4709 ( .A1(n4065), .A2(n4890), .ZN(n4598) );
  CKND2D1BWP12T U4710 ( .A1(n4598), .A2(n4167), .ZN(n4066) );
  OAI211D1BWP12T U4711 ( .A1(n4068), .A2(n4531), .B(n4067), .C(n4066), .ZN(
        n4069) );
  AOI21D1BWP12T U4712 ( .A1(n5088), .A2(n4407), .B(n4069), .ZN(n4079) );
  NR2D0BWP12T U4713 ( .A1(n4070), .A2(n4072), .ZN(n4075) );
  TPOAI21D0BWP12T U4714 ( .A1(n4073), .A2(n4072), .B(n4071), .ZN(n4074) );
  AOI21D1BWP12T U4715 ( .A1(n4333), .A2(n4075), .B(n4074), .ZN(n4077) );
  XOR2XD1BWP12T U4716 ( .A1(n4077), .A2(n4076), .Z(n4344) );
  CKND2D1BWP12T U4717 ( .A1(n4344), .A2(n5090), .ZN(n4078) );
  AN4XD1BWP12T U4718 ( .A1(n4081), .A2(n4080), .A3(n4079), .A4(n4078), .Z(
        n4082) );
  AOI22D0BWP12T U4719 ( .A1(n4200), .A2(n289), .B1(n4561), .B2(n4931), .ZN(
        n4086) );
  AOI22D1BWP12T U4720 ( .A1(n4559), .A2(n4921), .B1(n4562), .B2(n2746), .ZN(
        n4085) );
  TPAOI21D0BWP12T U4721 ( .A1(n4086), .A2(n4085), .B(n4743), .ZN(n4087) );
  AOI211D1BWP12T U4722 ( .A1(n4556), .A2(n4088), .B(n4087), .C(n4843), .ZN(
        n4091) );
  MAOI22D0BWP12T U4723 ( .A1(n4089), .A2(n4569), .B1(n4522), .B2(n4554), .ZN(
        n4090) );
  ND2D1BWP12T U4724 ( .A1(n4091), .A2(n4090), .ZN(n4139) );
  INVD0BWP12T U4725 ( .I(n4139), .ZN(n4092) );
  AOI21D1BWP12T U4726 ( .A1(n4824), .A2(n4843), .B(n4092), .ZN(n4529) );
  INVD1BWP12T U4727 ( .I(n4093), .ZN(n4780) );
  CKND0BWP12T U4728 ( .I(n4094), .ZN(n4107) );
  INVD1BWP12T U4729 ( .I(n4095), .ZN(n4097) );
  ND2D1BWP12T U4730 ( .A1(n4097), .A2(n4096), .ZN(n4099) );
  XNR2D1BWP12T U4731 ( .A1(n4099), .A2(n4098), .ZN(n4263) );
  ND2D1BWP12T U4732 ( .A1(n4263), .A2(n5085), .ZN(n4106) );
  CKND2D1BWP12T U4733 ( .A1(n4101), .A2(n4100), .ZN(n4120) );
  XOR2XD1BWP12T U4734 ( .A1(n4102), .A2(n4120), .Z(n4495) );
  INVD1BWP12T U4735 ( .I(n4104), .ZN(n4105) );
  OAI211D1BWP12T U4736 ( .A1(n4780), .A2(n4107), .B(n4106), .C(n4105), .ZN(
        n4138) );
  OR2D0BWP12T U4737 ( .A1(n4113), .A2(n4114), .Z(n4119) );
  INR2D1BWP12T U4738 ( .A1(n4115), .B1(n4114), .ZN(n4117) );
  NR2D1BWP12T U4739 ( .A1(n4117), .A2(n4116), .ZN(n4118) );
  OAI21D1BWP12T U4740 ( .A1(n5082), .A2(n4119), .B(n4118), .ZN(n4121) );
  XNR2D1BWP12T U4741 ( .A1(n4121), .A2(n4120), .ZN(n4400) );
  MUX2ND0BWP12T U4742 ( .I0(n5045), .I1(n5044), .S(n4743), .ZN(n4122) );
  ND2XD0BWP12T U4743 ( .A1(n4122), .A2(n5081), .ZN(n4123) );
  MUX2ND0BWP12T U4744 ( .I0(n4123), .I1(n5048), .S(n4626), .ZN(n4128) );
  OAI21D1BWP12T U4745 ( .A1(n289), .A2(n5083), .B(n5081), .ZN(n4126) );
  AOI22D1BWP12T U4746 ( .A1(n4419), .A2(n5078), .B1(n4743), .B2(n4126), .ZN(
        n4127) );
  CKND2D1BWP12T U4747 ( .A1(n4128), .A2(n4127), .ZN(n4129) );
  TPAOI21D0BWP12T U4748 ( .A1(n4400), .A2(n5088), .B(n4129), .ZN(n4130) );
  IOA21D1BWP12T U4749 ( .A1(n4957), .A2(n5093), .B(n4130), .ZN(n4136) );
  AOI22D1BWP12T U4750 ( .A1(n4323), .A2(n5090), .B1(n4249), .B2(n4583), .ZN(
        n4135) );
  AOI211D1BWP12T U4751 ( .A1(n5026), .A2(n4529), .B(n4138), .C(n4137), .ZN(
        n4143) );
  TPOAI21D0BWP12T U4752 ( .A1(n4858), .A2(n4891), .B(n4890), .ZN(n4140) );
  INR2D2BWP12T U4753 ( .A1(n5099), .B1(n4880), .ZN(n4141) );
  INVD1P75BWP12T U4754 ( .I(n4141), .ZN(n4142) );
  TPND2D2BWP12T U4755 ( .A1(n4143), .A2(n4142), .ZN(result[3]) );
  INVD1BWP12T U4756 ( .I(n4144), .ZN(n4145) );
  ND2D1BWP12T U4757 ( .A1(n4146), .A2(n4145), .ZN(n4147) );
  XNR2XD2BWP12T U4758 ( .A1(n4148), .A2(n4147), .ZN(n4281) );
  XOR2XD1BWP12T U4759 ( .A1(n4367), .A2(n4187), .Z(n4404) );
  AOI222D1BWP12T U4760 ( .A1(n4152), .A2(n4801), .B1(n4153), .B2(n4797), .C1(
        n4151), .C2(n4799), .ZN(n4169) );
  OAI22D1BWP12T U4761 ( .A1(n4154), .A2(n4685), .B1(n4153), .B2(n4707), .ZN(
        n4155) );
  AOI211D1BWP12T U4762 ( .A1(n4158), .A2(n4157), .B(n4156), .C(n4155), .ZN(
        n4604) );
  XNR2XD1BWP12T U4763 ( .A1(n4426), .A2(n4927), .ZN(n4436) );
  NR2D0BWP12T U4764 ( .A1(n4927), .A2(n5083), .ZN(n4159) );
  OA21D1BWP12T U4765 ( .A1(n905), .A2(n4159), .B(n4761), .Z(n4160) );
  AOI21D1BWP12T U4766 ( .A1(n4436), .A2(n5078), .B(n4160), .ZN(n4164) );
  MUX2ND0BWP12T U4767 ( .I0(n5045), .I1(n5044), .S(n4761), .ZN(n4161) );
  TPND2D0BWP12T U4768 ( .A1(n4161), .A2(n5081), .ZN(n4162) );
  MUX2NXD0BWP12T U4769 ( .I0(n4162), .I1(n5048), .S(n4638), .ZN(n4163) );
  ND3D1BWP12T U4770 ( .A1(n4165), .A2(n4164), .A3(n4163), .ZN(n4166) );
  AOI21D1BWP12T U4771 ( .A1(n4604), .A2(n4167), .B(n4166), .ZN(n4168) );
  OAI21D1BWP12T U4772 ( .A1(n4169), .A2(n5040), .B(n4168), .ZN(n4178) );
  OAI22D1BWP12T U4773 ( .A1(n4171), .A2(n4206), .B1(n4170), .B2(n4521), .ZN(
        n4175) );
  OAI22D1BWP12T U4774 ( .A1(n4173), .A2(n4554), .B1(n4172), .B2(n4566), .ZN(
        n4174) );
  IOA21D1BWP12T U4775 ( .A1(n4404), .A2(n5088), .B(n4179), .ZN(n4180) );
  CKND2D1BWP12T U4776 ( .A1(n4181), .A2(n4183), .ZN(n4186) );
  AOI21D1BWP12T U4777 ( .A1(n4184), .A2(n4183), .B(n4182), .ZN(n4185) );
  OAI21D1BWP12T U4778 ( .A1(n4493), .A2(n4186), .B(n4185), .ZN(n4188) );
  ND2D1BWP12T U4779 ( .A1(n4506), .A2(n4103), .ZN(n4195) );
  XOR2XD1BWP12T U4780 ( .A1(n4985), .A2(n4193), .Z(n4960) );
  INR2D2BWP12T U4781 ( .A1(n4195), .B1(n4194), .ZN(n4196) );
  TPND2D2BWP12T U4782 ( .A1(n4197), .A2(n4196), .ZN(n4198) );
  NR2XD0BWP12T U4783 ( .A1(n4199), .A2(n4521), .ZN(n4205) );
  CKND2D1BWP12T U4784 ( .A1(n4559), .A2(n4912), .ZN(n4202) );
  CKND2D0BWP12T U4785 ( .A1(n4200), .A2(n4911), .ZN(n4201) );
  OAI22D1BWP12T U4786 ( .A1(n4208), .A2(n4554), .B1(n4207), .B2(n4206), .ZN(
        n4817) );
  OR2XD1BWP12T U4787 ( .A1(n4209), .A2(n5099), .Z(n4210) );
  ND2D1BWP12T U4788 ( .A1(n4573), .A2(n4210), .ZN(n4211) );
  NR2D0BWP12T U4789 ( .A1(n4545), .A2(n4211), .ZN(n4213) );
  TPND2D1BWP12T U4790 ( .A1(n4213), .A2(n4212), .ZN(n4256) );
  XNR2D1BWP12T U4791 ( .A1(n4214), .A2(n5079), .ZN(n4421) );
  OAI21D0BWP12T U4792 ( .A1(n4911), .A2(n5083), .B(n5081), .ZN(n4215) );
  AOI22D0BWP12T U4793 ( .A1(n4421), .A2(n5078), .B1(n4645), .B2(n4215), .ZN(
        n4219) );
  MUX2ND0BWP12T U4794 ( .I0(n5045), .I1(n5044), .S(n4738), .ZN(n4216) );
  CKND2D0BWP12T U4795 ( .A1(n4216), .A2(n5081), .ZN(n4217) );
  MUX2ND0BWP12T U4796 ( .I0(n4217), .I1(n5048), .S(n4644), .ZN(n4218) );
  AN2XD1BWP12T U4797 ( .A1(n4219), .A2(n4218), .Z(n4236) );
  INVD0BWP12T U4798 ( .I(n4394), .ZN(n4220) );
  AOI21D1BWP12T U4799 ( .A1(n5075), .A2(n4952), .B(n4220), .ZN(n4223) );
  CKND2D1BWP12T U4800 ( .A1(n4230), .A2(n4221), .ZN(n4222) );
  XOR2XD1BWP12T U4801 ( .A1(n4223), .A2(n4222), .Z(n4397) );
  INR2D1BWP12T U4802 ( .A1(n4397), .B1(n4396), .ZN(n4235) );
  INVD1BWP12T U4803 ( .I(n4224), .ZN(n4952) );
  AOI21D1BWP12T U4804 ( .A1(n4225), .A2(n4952), .B(n4220), .ZN(n4228) );
  XOR2XD1BWP12T U4805 ( .A1(n4228), .A2(n4243), .Z(n4955) );
  CKND2D1BWP12T U4806 ( .A1(n4230), .A2(n4229), .ZN(n4231) );
  XOR2XD1BWP12T U4807 ( .A1(n4231), .A2(n4487), .Z(n4490) );
  INVD1BWP12T U4808 ( .I(n4490), .ZN(n4232) );
  INR3XD1BWP12T U4809 ( .A1(n4236), .B1(n4235), .B2(n4234), .ZN(n4241) );
  ND2D0BWP12T U4810 ( .A1(n4259), .A2(n5085), .ZN(n4240) );
  ND2D1BWP12T U4811 ( .A1(n4241), .A2(n4240), .ZN(n4242) );
  AOI21D1BWP12T U4812 ( .A1(n5100), .A2(n5099), .B(n4242), .ZN(n4250) );
  CKXOR2D1BWP12T U4813 ( .A1(n4244), .A2(n4243), .Z(n4319) );
  TPND2D0BWP12T U4814 ( .A1(n4319), .A2(n5090), .ZN(n4245) );
  TPND2D0BWP12T U4815 ( .A1(n4818), .A2(n4245), .ZN(n4247) );
  CKND2D1BWP12T U4816 ( .A1(n4245), .A2(n5098), .ZN(n4246) );
  INVD1BWP12T U4817 ( .I(n4248), .ZN(n4582) );
  OR2D0BWP12T U4818 ( .A1(n4707), .A2(n5040), .Z(n4252) );
  OAI22D1BWP12T U4819 ( .A1(n4787), .A2(n5040), .B1(n4788), .B2(n4252), .ZN(
        n4253) );
  TPNR2D1BWP12T U4820 ( .A1(n4254), .A2(n4253), .ZN(n4255) );
  TPND2D2BWP12T U4821 ( .A1(n4256), .A2(n4255), .ZN(result[1]) );
  INR2D1BWP12T U4822 ( .A1(n4258), .B1(n4257), .ZN(n5086) );
  OR3D0BWP12T U4823 ( .A1(n5086), .A2(n4260), .A3(n4259), .Z(n4261) );
  IND2D1BWP12T U4824 ( .A1(n4272), .B1(n4271), .ZN(n4273) );
  XNR2XD4BWP12T U4825 ( .A1(n4274), .A2(n4273), .ZN(n5036) );
  CKND0BWP12T U4826 ( .I(n4277), .ZN(n4279) );
  IND4D1BWP12T U4827 ( .A1(n4281), .B1(n4280), .B2(n4279), .B3(n4278), .ZN(
        n4287) );
  ND2D1BWP12T U4828 ( .A1(n311), .A2(n4290), .ZN(n4292) );
  NR4D0BWP12T U4829 ( .A1(n4296), .A2(n5073), .A3(n4295), .A4(n4294), .ZN(
        n4297) );
  TPND2D1BWP12T U4830 ( .A1(n4298), .A2(n4297), .ZN(n5008) );
  CKND3BWP12T U4831 ( .I(n4301), .ZN(n4302) );
  NR2XD2BWP12T U4832 ( .A1(n4308), .A2(n4307), .ZN(n4309) );
  TPND2D2BWP12T U4833 ( .A1(n4310), .A2(n4309), .ZN(n5007) );
  OR4D1BWP12T U4834 ( .A1(n4319), .A2(n5091), .A3(n4318), .A4(n4317), .Z(n4320) );
  OR4D1BWP12T U4835 ( .A1(n4323), .A2(n4322), .A3(n4321), .A4(n4320), .Z(n4326) );
  NR4D0BWP12T U4836 ( .A1(n4327), .A2(n4326), .A3(n4325), .A4(n4324), .ZN(
        n4348) );
  TPNR3D0BWP12T U4837 ( .A1(n4330), .A2(n4329), .A3(n4328), .ZN(n4347) );
  TPAOI21D1BWP12T U4838 ( .A1(n4333), .A2(n4332), .B(n4331), .ZN(n4337) );
  INVD0BWP12T U4839 ( .I(n4334), .ZN(n4335) );
  CKND2D1BWP12T U4840 ( .A1(n4335), .A2(n4972), .ZN(n4336) );
  XOR2XD1BWP12T U4841 ( .A1(n4337), .A2(n4336), .Z(n5011) );
  NR4D0BWP12T U4842 ( .A1(n4340), .A2(n5011), .A3(n4339), .A4(n4338), .ZN(
        n4346) );
  NR4D0BWP12T U4843 ( .A1(n4344), .A2(n4343), .A3(n4342), .A4(n4341), .ZN(
        n4345) );
  ND4D1BWP12T U4844 ( .A1(n4348), .A2(n4347), .A3(n4346), .A4(n4345), .ZN(
        n4361) );
  INVD0BWP12T U4845 ( .I(n4349), .ZN(n4352) );
  INVD1BWP12T U4846 ( .I(n4350), .ZN(n4351) );
  OAI21D1BWP12T U4847 ( .A1(n4353), .A2(n4352), .B(n4351), .ZN(n4356) );
  ND2D1BWP12T U4848 ( .A1(n4355), .A2(n4354), .ZN(n4986) );
  OR4D1BWP12T U4849 ( .A1(n5071), .A2(n4359), .A3(n4358), .A4(n4357), .Z(n4360) );
  NR4D0BWP12T U4850 ( .A1(n4363), .A2(n4362), .A3(n4361), .A4(n4360), .ZN(
        n5004) );
  CKND0BWP12T U4851 ( .I(n4364), .ZN(n5003) );
  OAI21D1BWP12T U4852 ( .A1(n4367), .A2(n4366), .B(n4365), .ZN(n4370) );
  CKND2D1BWP12T U4853 ( .A1(n4369), .A2(n4368), .ZN(n4477) );
  XNR2D1BWP12T U4854 ( .A1(n4370), .A2(n4477), .ZN(n5061) );
  OR4XD1BWP12T U4855 ( .A1(n5061), .A2(n4373), .A3(n4372), .A4(n4371), .Z(
        n4375) );
  NR2D0BWP12T U4856 ( .A1(n4378), .A2(n4380), .ZN(n4383) );
  TPOAI21D0BWP12T U4857 ( .A1(n4381), .A2(n4380), .B(n4379), .ZN(n4382) );
  AOI21D1BWP12T U4858 ( .A1(n4384), .A2(n4383), .B(n4382), .ZN(n4386) );
  CKND2D1BWP12T U4859 ( .A1(n4492), .A2(n4491), .ZN(n4385) );
  XOR2XD1BWP12T U4860 ( .A1(n4386), .A2(n4385), .Z(n5029) );
  OR4D1BWP12T U4861 ( .A1(n4390), .A2(n4389), .A3(n4388), .A4(n4387), .Z(n4391) );
  OR4D1BWP12T U4862 ( .A1(n5029), .A2(n4393), .A3(n4392), .A4(n4391), .Z(n4405) );
  OR4D1BWP12T U4863 ( .A1(n4397), .A2(n5087), .A3(n4396), .A4(n4395), .Z(n4399) );
  OR4D1BWP12T U4864 ( .A1(n4401), .A2(n4400), .A3(n4399), .A4(n4398), .Z(n4402) );
  TPNR2D0BWP12T U4865 ( .A1(n4411), .A2(n4410), .ZN(n4415) );
  NR2D1BWP12T U4866 ( .A1(n4413), .A2(n4412), .ZN(n4414) );
  ND2D1BWP12T U4867 ( .A1(n4415), .A2(n4414), .ZN(n4417) );
  OR4D1BWP12T U4868 ( .A1(n4421), .A2(n4420), .A3(n4419), .A4(n4418), .Z(n4423) );
  NR4D0BWP12T U4869 ( .A1(n4438), .A2(n4437), .A3(n4436), .A4(n4435), .ZN(
        n4456) );
  TPNR3D0BWP12T U4870 ( .A1(n4441), .A2(n4440), .A3(n4439), .ZN(n4455) );
  NR2D1BWP12T U4871 ( .A1(n4446), .A2(n4904), .ZN(n4447) );
  TPND2D0BWP12T U4872 ( .A1(n4448), .A2(n4447), .ZN(n4450) );
  XOR2XD1BWP12T U4873 ( .A1(n4450), .A2(n4449), .Z(n5019) );
  NR4D0BWP12T U4874 ( .A1(n5019), .A2(n4453), .A3(n4452), .A4(n4451), .ZN(
        n4454) );
  NR4D0BWP12T U4875 ( .A1(n848), .A2(n4922), .A3(a[27]), .A4(n4907), .ZN(n4463) );
  NR4D0BWP12T U4876 ( .A1(n4909), .A2(n4459), .A3(n2818), .A4(n4904), .ZN(
        n4462) );
  NR4D0BWP12T U4877 ( .A1(n4932), .A2(n5014), .A3(n4905), .A4(n4906), .ZN(
        n4461) );
  NR4D0BWP12T U4878 ( .A1(n4923), .A2(n2666), .A3(n4926), .A4(n4925), .ZN(
        n4460) );
  ND4D1BWP12T U4879 ( .A1(n4463), .A2(n4462), .A3(n4461), .A4(n4460), .ZN(
        n4469) );
  ND4D0BWP12T U4880 ( .A1(n4651), .A2(n5047), .A3(n4625), .A4(n4631), .ZN(
        n4468) );
  NR4D0BWP12T U4881 ( .A1(n2746), .A2(n4921), .A3(n4560), .A4(n4911), .ZN(
        n4464) );
  ND4D0BWP12T U4882 ( .A1(n4465), .A2(n905), .A3(n4464), .A4(n1810), .ZN(n4467) );
  ND4D0BWP12T U4883 ( .A1(n4638), .A2(n373), .A3(n1342), .A4(n4679), .ZN(n4466) );
  OAI21D1BWP12T U4884 ( .A1(n4473), .A2(n4472), .B(n4471), .ZN(n5001) );
  OAI21D1BWP12T U4885 ( .A1(n4476), .A2(n4475), .B(n4474), .ZN(n4478) );
  OR4D1BWP12T U4886 ( .A1(n5089), .A2(n4490), .A3(n4489), .A4(n4488), .Z(n4494) );
  OR4D1BWP12T U4887 ( .A1(n4496), .A2(n4495), .A3(n4494), .A4(n5030), .Z(n4499) );
  NR4D0BWP12T U4888 ( .A1(n4504), .A2(n4503), .A3(n4502), .A4(n4501), .ZN(
        n4513) );
  INVD0BWP12T U4889 ( .I(n4517), .ZN(n4519) );
  MAOI22D0BWP12T U4890 ( .A1(n4519), .A2(n4569), .B1(n4518), .B2(n4554), .ZN(
        n4526) );
  OAI21D0BWP12T U4891 ( .A1(n4520), .A2(n4566), .B(n4707), .ZN(n4524) );
  NR2D0BWP12T U4892 ( .A1(n4522), .A2(n4521), .ZN(n4523) );
  NR2D1BWP12T U4893 ( .A1(n4524), .A2(n4523), .ZN(n4525) );
  ND2D1BWP12T U4894 ( .A1(n4526), .A2(n4525), .ZN(n4893) );
  INVD1BWP12T U4895 ( .I(n4893), .ZN(n4527) );
  AOI21D1BWP12T U4896 ( .A1(n4821), .A2(n4843), .B(n4527), .ZN(n5027) );
  TPNR3D0BWP12T U4897 ( .A1(n4529), .A2(n5027), .A3(n4528), .ZN(n4827) );
  AOI31D0BWP12T U4898 ( .A1(n4531), .A2(n4827), .A3(n4530), .B(n4891), .ZN(
        n4777) );
  NR4D0BWP12T U4899 ( .A1(n4536), .A2(n4535), .A3(n4534), .A4(n4533), .ZN(
        n4537) );
  ND4D1BWP12T U4900 ( .A1(n4540), .A2(n4539), .A3(n4538), .A4(n4537), .ZN(
        n4784) );
  INVD1BWP12T U4901 ( .I(n4541), .ZN(n5037) );
  TPNR2D0BWP12T U4902 ( .A1(n5037), .A2(n4542), .ZN(n4825) );
  OAI21D0BWP12T U4903 ( .A1(n4552), .A2(n4551), .B(n4573), .ZN(n4579) );
  INVD0BWP12T U4904 ( .I(n4553), .ZN(n4557) );
  INVD1BWP12T U4905 ( .I(n4558), .ZN(n4570) );
  ND2D0BWP12T U4906 ( .A1(n4559), .A2(n4911), .ZN(n4565) );
  CKND2D0BWP12T U4907 ( .A1(n4561), .A2(n4560), .ZN(n4564) );
  CKND2D0BWP12T U4908 ( .A1(n4562), .A2(n4912), .ZN(n4563) );
  TPAOI31D0BWP12T U4909 ( .A1(n4565), .A2(n4564), .A3(n4563), .B(n4743), .ZN(
        n4568) );
  NR2D1BWP12T U4910 ( .A1(n4567), .A2(n4566), .ZN(n5096) );
  AOI211XD0BWP12T U4911 ( .A1(n4570), .A2(n4569), .B(n4568), .C(n5096), .ZN(
        n4571) );
  ND2D1BWP12T U4912 ( .A1(n4572), .A2(n4571), .ZN(n5074) );
  AOI22D1BWP12T U4913 ( .A1(n4605), .A2(n5074), .B1(n5095), .B2(n4573), .ZN(
        n5103) );
  INVD1BWP12T U4914 ( .I(n5103), .ZN(n5101) );
  NR4D0BWP12T U4915 ( .A1(n5101), .A2(n4575), .A3(n4574), .A4(n5102), .ZN(
        n4578) );
  ND4D0BWP12T U4916 ( .A1(n4579), .A2(n4578), .A3(n4577), .A4(n4576), .ZN(
        n4775) );
  NR3D1BWP12T U4917 ( .A1(n4586), .A2(n4585), .A3(n4584), .ZN(n4587) );
  ND4D1BWP12T U4918 ( .A1(n4595), .A2(n4594), .A3(n4593), .A4(n4592), .ZN(
        n4596) );
  NR4D0BWP12T U4919 ( .A1(n4599), .A2(n4598), .A3(n4597), .A4(n4596), .ZN(
        n4773) );
  NR4D0BWP12T U4920 ( .A1(n4603), .A2(n4602), .A3(n4601), .A4(n4600), .ZN(
        n4615) );
  AOI211D1BWP12T U4921 ( .A1(n4606), .A2(n4605), .B(n4604), .C(n5042), .ZN(
        n4614) );
  AOI22D1BWP12T U4922 ( .A1(n4743), .A2(n4608), .B1(n4607), .B2(n4843), .ZN(
        n4609) );
  OAI211D1BWP12T U4923 ( .A1(n4612), .A2(n4611), .B(n4610), .C(n4609), .ZN(
        n5043) );
  ND4D0BWP12T U4924 ( .A1(n4615), .A2(n4614), .A3(n5043), .A4(n4613), .ZN(
        n4622) );
  ND3D0BWP12T U4925 ( .A1(n4618), .A2(n4617), .A3(n4616), .ZN(n4621) );
  NR4D0BWP12T U4926 ( .A1(n4622), .A2(n4621), .A3(n4620), .A4(n4619), .ZN(
        n4772) );
  OAI21D1BWP12T U4927 ( .A1(n4751), .A2(n4624), .B(n4623), .ZN(n4725) );
  AOI22D1BWP12T U4928 ( .A1(n4726), .A2(n4625), .B1(n5053), .B2(n5047), .ZN(
        n4642) );
  AOI22D0BWP12T U4929 ( .A1(n4743), .A2(n4626), .B1(n4742), .B2(n373), .ZN(
        n4630) );
  ND2D1BWP12T U4930 ( .A1(n4628), .A2(n4627), .ZN(n4629) );
  OAI211D0BWP12T U4931 ( .A1(n4921), .A2(n4707), .B(n4630), .C(n4629), .ZN(
        n4635) );
  CKND2D0BWP12T U4932 ( .A1(n4748), .A2(n4631), .ZN(n4632) );
  OAI211D0BWP12T U4933 ( .A1(n4906), .A2(n4704), .B(n4633), .C(n4632), .ZN(
        n4634) );
  AOI211D1BWP12T U4934 ( .A1(n4727), .A2(n4636), .B(n4635), .C(n4634), .ZN(
        n4641) );
  AOI22D0BWP12T U4935 ( .A1(n4762), .A2(n4637), .B1(n1342), .B2(n4764), .ZN(
        n4640) );
  AOI22D0BWP12T U4936 ( .A1(n4761), .A2(n4638), .B1(n279), .B2(n1810), .ZN(
        n4639) );
  ND4D1BWP12T U4937 ( .A1(n4642), .A2(n4641), .A3(n4640), .A4(n4639), .ZN(
        n4663) );
  CKND0BWP12T U4938 ( .I(n5084), .ZN(n4643) );
  AOI21D0BWP12T U4939 ( .A1(n4759), .A2(n4930), .B(n4643), .ZN(n4647) );
  AOI22D0BWP12T U4940 ( .A1(n4750), .A2(n4679), .B1(n4645), .B2(n4644), .ZN(
        n4646) );
  OAI211D0BWP12T U4941 ( .A1(n4648), .A2(n4688), .B(n4647), .C(n4646), .ZN(
        n4662) );
  AO22XD0BWP12T U4942 ( .A1(n4740), .A2(n4650), .B1(n4739), .B2(n4649), .Z(
        n4661) );
  CKND2D0BWP12T U4943 ( .A1(n4729), .A2(n4651), .ZN(n4659) );
  AOI22D0BWP12T U4944 ( .A1(n4760), .A2(n4652), .B1(n4752), .B2(n4680), .ZN(
        n4658) );
  AOI22D0BWP12T U4945 ( .A1(n342), .A2(n4654), .B1(n295), .B2(n4653), .ZN(
        n4657) );
  AOI22D0BWP12T U4946 ( .A1(n4749), .A2(n4655), .B1(n5015), .B2(n777), .ZN(
        n4656) );
  ND4D1BWP12T U4947 ( .A1(n4659), .A2(n4658), .A3(n4657), .A4(n4656), .ZN(
        n4660) );
  NR4D0BWP12T U4948 ( .A1(n4663), .A2(n4662), .A3(n4661), .A4(n4660), .ZN(
        n4672) );
  AOI22D0BWP12T U4949 ( .A1(n4733), .A2(n4665), .B1(n4730), .B2(n4664), .ZN(
        n4671) );
  AOI22D0BWP12T U4950 ( .A1(n4731), .A2(n4667), .B1(b[26]), .B2(n4666), .ZN(
        n4670) );
  CKND0BWP12T U4951 ( .I(n4668), .ZN(n4669) );
  ND4D1BWP12T U4952 ( .A1(n4672), .A2(n4671), .A3(n4670), .A4(n4669), .ZN(
        n4724) );
  AOI22D1BWP12T U4953 ( .A1(n4925), .A2(n4674), .B1(n4673), .B2(n4926), .ZN(
        n4678) );
  AOI22D0BWP12T U4954 ( .A1(n4904), .A2(n4676), .B1(n4675), .B2(n5014), .ZN(
        n4677) );
  CKND2D1BWP12T U4955 ( .A1(n4678), .A2(n4677), .ZN(n4682) );
  OAI22D0BWP12T U4956 ( .A1(n4752), .A2(n4680), .B1(n4750), .B2(n4679), .ZN(
        n4681) );
  AOI211D1BWP12T U4957 ( .A1(n4728), .A2(n4683), .B(n4682), .C(n4681), .ZN(
        n4692) );
  AOI22D0BWP12T U4958 ( .A1(n2746), .A2(n4684), .B1(n4848), .B2(n4912), .ZN(
        n4691) );
  AOI22D0BWP12T U4959 ( .A1(n4911), .A2(n4686), .B1(n4685), .B2(n289), .ZN(
        n4690) );
  AOI22D1BWP12T U4960 ( .A1(n4916), .A2(n4688), .B1(n4687), .B2(n2666), .ZN(
        n4689) );
  AN4XD1BWP12T U4961 ( .A1(n4692), .A2(n4691), .A3(n4690), .A4(n4689), .Z(
        n4703) );
  AOI22D1BWP12T U4962 ( .A1(n4908), .A2(n4694), .B1(n4693), .B2(n4909), .ZN(
        n4702) );
  AOI22D1BWP12T U4963 ( .A1(a[27]), .A2(n4696), .B1(n4695), .B2(n4922), .ZN(
        n4701) );
  AOI22D1BWP12T U4964 ( .A1(n4699), .A2(n4698), .B1(n4697), .B2(n4907), .ZN(
        n4700) );
  ND4D1BWP12T U4965 ( .A1(n4703), .A2(n4702), .A3(n4701), .A4(n4700), .ZN(
        n4723) );
  AOI22D0BWP12T U4966 ( .A1(n4905), .A2(n4705), .B1(n4704), .B2(n4906), .ZN(
        n4709) );
  AOI22D0BWP12T U4967 ( .A1(n4707), .A2(n4921), .B1(n4706), .B2(n4931), .ZN(
        n4708) );
  OAI211D0BWP12T U4968 ( .A1(n5075), .A2(n5079), .B(n4709), .C(n4708), .ZN(
        n4710) );
  AOI21D0BWP12T U4969 ( .A1(n4933), .A2(n4711), .B(n4710), .ZN(n4721) );
  AOI22D1BWP12T U4970 ( .A1(n5051), .A2(n4713), .B1(n4712), .B2(n4914), .ZN(
        n4720) );
  AOI22D1BWP12T U4971 ( .A1(n4924), .A2(n4715), .B1(n4714), .B2(n4923), .ZN(
        n4719) );
  AOI22D0BWP12T U4972 ( .A1(n2688), .A2(n4717), .B1(n4716), .B2(n4927), .ZN(
        n4718) );
  ND4D1BWP12T U4973 ( .A1(n4721), .A2(n4720), .A3(n4719), .A4(n4718), .ZN(
        n4722) );
  AOI211D1BWP12T U4974 ( .A1(n4725), .A2(n4724), .B(n4723), .C(n4722), .ZN(
        n4771) );
  AOI22D1BWP12T U4975 ( .A1(n4726), .A2(n4914), .B1(n5053), .B2(n5051), .ZN(
        n4737) );
  AOI22D1BWP12T U4976 ( .A1(n4729), .A2(n4728), .B1(n4727), .B2(n4933), .ZN(
        n4736) );
  AOI22D1BWP12T U4977 ( .A1(n4731), .A2(a[27]), .B1(n4730), .B2(n4909), .ZN(
        n4735) );
  AOI22D0BWP12T U4978 ( .A1(n4733), .A2(n4908), .B1(n4732), .B2(n4916), .ZN(
        n4734) );
  ND4D1BWP12T U4979 ( .A1(n4737), .A2(n4736), .A3(n4735), .A4(n4734), .ZN(
        n4769) );
  AOI22D1BWP12T U4980 ( .A1(b[26]), .A2(n4922), .B1(n4738), .B2(n4911), .ZN(
        n4747) );
  AOI22D1BWP12T U4981 ( .A1(n4740), .A2(n4907), .B1(n4739), .B2(n2818), .ZN(
        n4746) );
  AOI22D0BWP12T U4982 ( .A1(n4741), .A2(n2746), .B1(n4843), .B2(n4921), .ZN(
        n4745) );
  AOI22D0BWP12T U4983 ( .A1(n4743), .A2(n289), .B1(n4742), .B2(n4912), .ZN(
        n4744) );
  ND4D1BWP12T U4984 ( .A1(n4747), .A2(n4746), .A3(n4745), .A4(n4744), .ZN(
        n4768) );
  AOI22D1BWP12T U4985 ( .A1(n4749), .A2(n4905), .B1(n4748), .B2(n4931), .ZN(
        n4758) );
  AOI22D0BWP12T U4986 ( .A1(n848), .A2(n4751), .B1(n4750), .B2(n288), .ZN(
        n4757) );
  AOI22D1BWP12T U4987 ( .A1(n295), .A2(n4926), .B1(n4752), .B2(n4932), .ZN(
        n4756) );
  AOI22D0BWP12T U4988 ( .A1(n5015), .A2(n5014), .B1(n342), .B2(n4904), .ZN(
        n4755) );
  ND4D1BWP12T U4989 ( .A1(n4758), .A2(n4757), .A3(n4756), .A4(n4755), .ZN(
        n4767) );
  NR4D0BWP12T U4990 ( .A1(n4769), .A2(n4768), .A3(n4767), .A4(n4766), .ZN(
        n4770) );
  RCAOI211D1BWP12T U4991 ( .A1(n4773), .A2(n4772), .B(n4771), .C(n4770), .ZN(
        n4774) );
  TPOAI31D0BWP12T U4992 ( .A1(n4777), .A2(n4776), .A3(n4775), .B(n4774), .ZN(
        n4942) );
  TPNR2D0BWP12T U4993 ( .A1(n4779), .A2(n4778), .ZN(n4782) );
  ND4D1BWP12T U4994 ( .A1(n4782), .A2(n4781), .A3(n5094), .A4(n4780), .ZN(
        n4783) );
  AOI211D1BWP12T U4995 ( .A1(n4786), .A2(n4785), .B(n4784), .C(n4783), .ZN(
        n4792) );
  CKND2D0BWP12T U4996 ( .A1(n4788), .A2(n4787), .ZN(n4790) );
  NR4D0BWP12T U4997 ( .A1(n4790), .A2(n5095), .A3(n4789), .A4(n5074), .ZN(
        n4791) );
  CKND2D1BWP12T U4998 ( .A1(n4792), .A2(n4791), .ZN(n4812) );
  ND4D0BWP12T U4999 ( .A1(n4796), .A2(n4795), .A3(n4794), .A4(n4793), .ZN(
        n4811) );
  AOI222D1BWP12T U5000 ( .A1(n4802), .A2(n4801), .B1(n4800), .B2(n4799), .C1(
        n4798), .C2(n4797), .ZN(n5041) );
  ND4D1BWP12T U5001 ( .A1(n4805), .A2(n4804), .A3(n5041), .A4(n4803), .ZN(
        n4810) );
  ND4D0BWP12T U5002 ( .A1(n4808), .A2(n4807), .A3(n5023), .A4(n4806), .ZN(
        n4809) );
  NR4D0BWP12T U5003 ( .A1(n4812), .A2(n4811), .A3(n4810), .A4(n4809), .ZN(
        n4816) );
  ND4D1BWP12T U5004 ( .A1(n4816), .A2(n4815), .A3(n4814), .A4(n4813), .ZN(
        n4845) );
  INR2D0BWP12T U5005 ( .A1(n4818), .B1(n4817), .ZN(n4820) );
  CKND2D0BWP12T U5006 ( .A1(n4830), .A2(n4829), .ZN(n4831) );
  NR2D0BWP12T U5007 ( .A1(n4832), .A2(n4831), .ZN(n4834) );
  NR2D1BWP12T U5008 ( .A1(n4845), .A2(n4844), .ZN(n4941) );
  TPAOI21D0BWP12T U5009 ( .A1(n4848), .A2(n4847), .B(n4846), .ZN(n4849) );
  OAI21D1BWP12T U5010 ( .A1(n4849), .A2(n5037), .B(n4874), .ZN(n5064) );
  ND4D0BWP12T U5011 ( .A1(n5064), .A2(n4852), .A3(n4851), .A4(n4850), .ZN(
        n4857) );
  NR2D0BWP12T U5012 ( .A1(n4854), .A2(n4853), .ZN(n4856) );
  NR3XD0BWP12T U5013 ( .A1(n4857), .A2(n4856), .A3(n4855), .ZN(n4903) );
  ND4D1BWP12T U5014 ( .A1(n4861), .A2(n4860), .A3(n4859), .A4(n4858), .ZN(
        n4862) );
  TPOAI31D0BWP12T U5015 ( .A1(n4864), .A2(n4863), .A3(n4862), .B(n4889), .ZN(
        n4870) );
  CKND2D0BWP12T U5016 ( .A1(n4866), .A2(n4865), .ZN(n4869) );
  ND4D0BWP12T U5017 ( .A1(n4870), .A2(n4869), .A3(n4868), .A4(n4867), .ZN(
        n4884) );
  ND4D0BWP12T U5018 ( .A1(n4873), .A2(n5103), .A3(n4872), .A4(n4871), .ZN(
        n4883) );
  CKND0BWP12T U5019 ( .I(n4874), .ZN(n4875) );
  AOI21D0BWP12T U5020 ( .A1(n4877), .A2(n4876), .B(n4875), .ZN(n4882) );
  ND3D0BWP12T U5021 ( .A1(n4880), .A2(n4879), .A3(n4878), .ZN(n4881) );
  NR4D0BWP12T U5022 ( .A1(n4884), .A2(n4883), .A3(n4882), .A4(n4881), .ZN(
        n4902) );
  CKND2D0BWP12T U5023 ( .A1(n4886), .A2(n4885), .ZN(n4901) );
  AOI211D0BWP12T U5024 ( .A1(n4889), .A2(n4888), .B(n4887), .C(n5063), .ZN(
        n4895) );
  OAI21D0BWP12T U5025 ( .A1(n4892), .A2(n4891), .B(n4890), .ZN(n4894) );
  AOI21D1BWP12T U5026 ( .A1(n4894), .A2(n4893), .B(n5100), .ZN(n5028) );
  CKND2D0BWP12T U5027 ( .A1(n4895), .A2(n5028), .ZN(n4897) );
  NR4D0BWP12T U5028 ( .A1(n4899), .A2(n4898), .A3(n4897), .A4(n4896), .ZN(
        n4900) );
  ND4D1BWP12T U5029 ( .A1(n4903), .A2(n4902), .A3(n4901), .A4(n4900), .ZN(
        n4939) );
  ND4D0BWP12T U5030 ( .A1(n4906), .A2(n4905), .A3(n4904), .A4(n5014), .ZN(
        n4920) );
  ND4D1BWP12T U5031 ( .A1(n4909), .A2(n4908), .A3(n2818), .A4(n4907), .ZN(
        n4919) );
  ND4D0BWP12T U5032 ( .A1(n289), .A2(n4912), .A3(n4911), .A4(n4910), .ZN(n4918) );
  ND4D1BWP12T U5033 ( .A1(n4916), .A2(n4915), .A3(n4914), .A4(n5051), .ZN(
        n4917) );
  NR4D0BWP12T U5034 ( .A1(n4920), .A2(n4919), .A3(n4918), .A4(n4917), .ZN(
        n4937) );
  AN4XD1BWP12T U5035 ( .A1(a[27]), .A2(n4922), .A3(n4921), .A4(n2746), .Z(
        n4936) );
  ND2D1BWP12T U5036 ( .A1(n4924), .A2(n4923), .ZN(n4929) );
  ND4D0BWP12T U5037 ( .A1(n2688), .A2(n4927), .A3(n4926), .A4(n4925), .ZN(
        n4928) );
  NR4D0BWP12T U5038 ( .A1(n4930), .A2(n4929), .A3(n4928), .A4(n5080), .ZN(
        n4935) );
  AN4D0BWP12T U5039 ( .A1(n4933), .A2(n4932), .A3(n4931), .A4(n288), .Z(n4934)
         );
  ND4D1BWP12T U5040 ( .A1(n4937), .A2(n4936), .A3(n4935), .A4(n4934), .ZN(
        n4938) );
  MUX2ND0BWP12T U5041 ( .I0(n4939), .I1(n4938), .S(n848), .ZN(n4940) );
  OR3D2BWP12T U5042 ( .A1(n4942), .A2(n4941), .A3(n4940), .Z(n4943) );
  NR2D1BWP12T U5043 ( .A1(n4944), .A2(n4943), .ZN(n5000) );
  NR2D0BWP12T U5044 ( .A1(n4946), .A2(n4945), .ZN(n4997) );
  OR4D1BWP12T U5045 ( .A1(n4950), .A2(n4949), .A3(n4948), .A4(n4947), .Z(n4982) );
  NR2D0BWP12T U5046 ( .A1(n4965), .A2(n4967), .ZN(n4970) );
  TPOAI21D0BWP12T U5047 ( .A1(n4968), .A2(n4967), .B(n4966), .ZN(n4969) );
  AOI21D1BWP12T U5048 ( .A1(n4971), .A2(n4970), .B(n4969), .ZN(n4975) );
  CKND2D1BWP12T U5049 ( .A1(n4973), .A2(n4972), .ZN(n4974) );
  XOR2XD1BWP12T U5050 ( .A1(n4975), .A2(n4974), .Z(n5010) );
  NR4D0BWP12T U5051 ( .A1(n4982), .A2(n4981), .A3(n4980), .A4(n4979), .ZN(
        n4996) );
  OAI21D1BWP12T U5052 ( .A1(n4985), .A2(n4984), .B(n4983), .ZN(n4987) );
  XNR2XD1BWP12T U5053 ( .A1(n4987), .A2(n4986), .ZN(n5065) );
  OR4XD1BWP12T U5054 ( .A1(n5065), .A2(n4990), .A3(n4989), .A4(n4988), .Z(
        n4991) );
  NR4D0BWP12T U5055 ( .A1(n4994), .A2(n4993), .A3(n4992), .A4(n4991), .ZN(
        n4995) );
  IND4D1BWP12T U5056 ( .A1(n4998), .B1(n4997), .B2(n4996), .B3(n4995), .ZN(
        n4999) );
  IND3D1BWP12T U5057 ( .A1(n5001), .B1(n5000), .B2(n4999), .ZN(n5002) );
  TPAOI31D1BWP12T U5058 ( .A1(n5005), .A2(n5004), .A3(n5003), .B(n5002), .ZN(
        n5006) );
  MUX2ND0BWP12T U5059 ( .I0(n5077), .I1(n5076), .S(n5015), .ZN(n5012) );
  NR2D0BWP12T U5060 ( .A1(n5012), .A2(n905), .ZN(n5013) );
  MUX2NXD0BWP12T U5061 ( .I0(n5013), .I1(n5080), .S(n777), .ZN(n5018) );
  NR2D0BWP12T U5062 ( .A1(n5014), .A2(n5083), .ZN(n5016) );
  OA21XD0BWP12T U5063 ( .A1(n905), .A2(n5016), .B(n5015), .Z(n5017) );
  AOI211D1BWP12T U5064 ( .A1(n5019), .A2(n5078), .B(n5018), .C(n5017), .ZN(
        n5022) );
  CKND2D1BWP12T U5065 ( .A1(n5020), .A2(n5097), .ZN(n5021) );
  OAI211D1BWP12T U5066 ( .A1(n5024), .A2(n5023), .B(n5022), .C(n5021), .ZN(
        n5025) );
  AOI21D1BWP12T U5067 ( .A1(n5027), .A2(n5026), .B(n5025), .ZN(n5033) );
  MAOI22D0BWP12T U5068 ( .A1(n5029), .A2(n5088), .B1(n5028), .B2(n5063), .ZN(
        n5032) );
  CKND2D1BWP12T U5069 ( .A1(n5030), .A2(n4103), .ZN(n5031) );
  AO21D4BWP12T U5070 ( .A1(n5036), .A2(n5085), .B(n5035), .Z(result[11]) );
  ND2D1BWP12T U5071 ( .A1(n5038), .A2(n5037), .ZN(n5039) );
  OAI21D1BWP12T U5072 ( .A1(n5041), .A2(n5040), .B(n5039), .ZN(n5059) );
  NR2D1BWP12T U5073 ( .A1(n5043), .A2(n5042), .ZN(n5058) );
  MUX2ND0BWP12T U5074 ( .I0(n5045), .I1(n5044), .S(n5053), .ZN(n5046) );
  TPND2D0BWP12T U5075 ( .A1(n5046), .A2(n5081), .ZN(n5049) );
  MUX2NXD0BWP12T U5076 ( .I0(n5049), .I1(n5048), .S(n5047), .ZN(n5056) );
  ND2D1BWP12T U5077 ( .A1(n5050), .A2(n5078), .ZN(n5055) );
  OAI21D1BWP12T U5078 ( .A1(n5051), .A2(n5083), .B(n5081), .ZN(n5052) );
  ND2D1BWP12T U5079 ( .A1(n5053), .A2(n5052), .ZN(n5054) );
  ND3D1BWP12T U5080 ( .A1(n5056), .A2(n5055), .A3(n5054), .ZN(n5057) );
  NR3D1BWP12T U5081 ( .A1(n5059), .A2(n5058), .A3(n5057), .ZN(n5060) );
  IOA21D1BWP12T U5082 ( .A1(n5061), .A2(n5088), .B(n5060), .ZN(n5069) );
  ND2D1BWP12T U5083 ( .A1(n5062), .A2(n4103), .ZN(n5067) );
  ND2D1BWP12T U5084 ( .A1(n5067), .A2(n5066), .ZN(n5068) );
  TPNR2D1BWP12T U5085 ( .A1(n5069), .A2(n5068), .ZN(n5070) );
  IOA21D2BWP12T U5086 ( .A1(n5071), .A2(n5090), .B(n5070), .ZN(n5072) );
  AO21D4BWP12T U5087 ( .A1(n5073), .A2(n5085), .B(n5072), .Z(result[20]) );
endmodule


module memory_interface_simple ( clock, reset, interface_cpu_sign_extend, 
        interface_cpu_word_type, interface_cpu_load_request, 
        interface_cpu_address_in, interface_cpu_data_in, from_mem_data_out, 
        interface_cpu_read_finished, interface_cpu_write_finished, 
        interface_cpu_data_out, to_mem_address, to_mem_data_in, 
        to_mem_read_enable, to_mem_write_enable, to_mem_enable, 
        interface_cpu_store_request_BAR );
  input [1:0] interface_cpu_word_type;
  input [12:0] interface_cpu_address_in;
  input [31:0] interface_cpu_data_in;
  input [15:0] from_mem_data_out;
  output [31:0] interface_cpu_data_out;
  output [11:0] to_mem_address;
  output [15:0] to_mem_data_in;
  input clock, reset, interface_cpu_sign_extend, interface_cpu_load_request,
         interface_cpu_store_request_BAR;
  output interface_cpu_read_finished, interface_cpu_write_finished,
         to_mem_read_enable, to_mem_write_enable, to_mem_enable;
  wire   sign_extend, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76,
         N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90,
         N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N183, N184, N185, N186, N187, N188, N189, N190, N191,
         N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202,
         N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, n346,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n347, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453;
  wire   [5:0] state;
  wire   [15:0] tmp_value_1;
  wire   [15:0] tmp_value_2;
  wire   [31:0] cpu_data_in;
  wire   [12:1] cpu_address_in;

  DFQD1BWP12T state_reg_0_ ( .D(N66), .CP(clock), .Q(state[0]) );
  DFQD1BWP12T state_reg_5_ ( .D(N71), .CP(clock), .Q(state[5]) );
  DFQD1BWP12T state_reg_1_ ( .D(N67), .CP(clock), .Q(state[1]) );
  DFQD1BWP12T state_reg_4_ ( .D(N70), .CP(clock), .Q(state[4]) );
  DFQD1BWP12T state_reg_2_ ( .D(N68), .CP(clock), .Q(state[2]) );
  DFQD1BWP12T state_reg_3_ ( .D(N69), .CP(clock), .Q(state[3]) );
  DFQD1BWP12T to_mem_write_enable_reg ( .D(N212), .CP(clock), .Q(
        to_mem_write_enable) );
  DFQD1BWP12T interface_cpu_read_finished_reg ( .D(N72), .CP(clock), .Q(
        interface_cpu_read_finished) );
  DFQD1BWP12T interface_cpu_write_finished_reg ( .D(N73), .CP(clock), .Q(
        interface_cpu_write_finished) );
  DFQD1BWP12T tmp_value_1_reg_15_ ( .D(n423), .CP(clock), .Q(tmp_value_1[15])
         );
  DFQD1BWP12T tmp_value_1_reg_14_ ( .D(n422), .CP(clock), .Q(tmp_value_1[14])
         );
  DFQD1BWP12T tmp_value_1_reg_13_ ( .D(n421), .CP(clock), .Q(tmp_value_1[13])
         );
  DFQD1BWP12T tmp_value_1_reg_12_ ( .D(n420), .CP(clock), .Q(tmp_value_1[12])
         );
  DFQD1BWP12T tmp_value_1_reg_11_ ( .D(n419), .CP(clock), .Q(tmp_value_1[11])
         );
  DFQD1BWP12T tmp_value_1_reg_10_ ( .D(n418), .CP(clock), .Q(tmp_value_1[10])
         );
  DFQD1BWP12T tmp_value_1_reg_9_ ( .D(n417), .CP(clock), .Q(tmp_value_1[9]) );
  DFQD1BWP12T tmp_value_1_reg_8_ ( .D(n416), .CP(clock), .Q(tmp_value_1[8]) );
  DFQD1BWP12T tmp_value_1_reg_7_ ( .D(n415), .CP(clock), .Q(tmp_value_1[7]) );
  DFQD1BWP12T interface_cpu_data_out_reg_7_ ( .D(N81), .CP(clock), .Q(
        interface_cpu_data_out[7]) );
  DFQD1BWP12T tmp_value_1_reg_6_ ( .D(n414), .CP(clock), .Q(tmp_value_1[6]) );
  DFQD1BWP12T interface_cpu_data_out_reg_6_ ( .D(N80), .CP(clock), .Q(
        interface_cpu_data_out[6]) );
  DFQD1BWP12T tmp_value_1_reg_5_ ( .D(n413), .CP(clock), .Q(tmp_value_1[5]) );
  DFQD1BWP12T interface_cpu_data_out_reg_5_ ( .D(N79), .CP(clock), .Q(
        interface_cpu_data_out[5]) );
  DFQD1BWP12T tmp_value_1_reg_4_ ( .D(n412), .CP(clock), .Q(tmp_value_1[4]) );
  DFQD1BWP12T interface_cpu_data_out_reg_4_ ( .D(N78), .CP(clock), .Q(
        interface_cpu_data_out[4]) );
  DFQD1BWP12T tmp_value_1_reg_3_ ( .D(n411), .CP(clock), .Q(tmp_value_1[3]) );
  DFQD1BWP12T interface_cpu_data_out_reg_3_ ( .D(N77), .CP(clock), .Q(
        interface_cpu_data_out[3]) );
  DFQD1BWP12T tmp_value_1_reg_2_ ( .D(n410), .CP(clock), .Q(tmp_value_1[2]) );
  DFQD1BWP12T interface_cpu_data_out_reg_2_ ( .D(N76), .CP(clock), .Q(
        interface_cpu_data_out[2]) );
  DFQD1BWP12T tmp_value_1_reg_1_ ( .D(n409), .CP(clock), .Q(tmp_value_1[1]) );
  DFQD1BWP12T interface_cpu_data_out_reg_1_ ( .D(N75), .CP(clock), .Q(
        interface_cpu_data_out[1]) );
  DFQD1BWP12T tmp_value_1_reg_0_ ( .D(n408), .CP(clock), .Q(tmp_value_1[0]) );
  DFQD1BWP12T interface_cpu_data_out_reg_0_ ( .D(N74), .CP(clock), .Q(
        interface_cpu_data_out[0]) );
  DFQD1BWP12T tmp_value_2_reg_15_ ( .D(n407), .CP(clock), .Q(tmp_value_2[15])
         );
  DFQD1BWP12T tmp_value_2_reg_14_ ( .D(n406), .CP(clock), .Q(tmp_value_2[14])
         );
  DFQD1BWP12T tmp_value_2_reg_13_ ( .D(n405), .CP(clock), .Q(tmp_value_2[13])
         );
  DFQD1BWP12T tmp_value_2_reg_12_ ( .D(n404), .CP(clock), .Q(tmp_value_2[12])
         );
  DFQD1BWP12T tmp_value_2_reg_11_ ( .D(n403), .CP(clock), .Q(tmp_value_2[11])
         );
  DFQD1BWP12T tmp_value_2_reg_10_ ( .D(n402), .CP(clock), .Q(tmp_value_2[10])
         );
  DFQD1BWP12T tmp_value_2_reg_9_ ( .D(n401), .CP(clock), .Q(tmp_value_2[9]) );
  DFQD1BWP12T tmp_value_2_reg_8_ ( .D(n400), .CP(clock), .Q(tmp_value_2[8]) );
  DFQD1BWP12T tmp_value_2_reg_7_ ( .D(n399), .CP(clock), .Q(tmp_value_2[7]) );
  DFQD1BWP12T tmp_value_2_reg_6_ ( .D(n398), .CP(clock), .Q(tmp_value_2[6]) );
  DFQD1BWP12T tmp_value_2_reg_5_ ( .D(n397), .CP(clock), .Q(tmp_value_2[5]) );
  DFQD1BWP12T tmp_value_2_reg_4_ ( .D(n396), .CP(clock), .Q(tmp_value_2[4]) );
  DFQD1BWP12T tmp_value_2_reg_3_ ( .D(n395), .CP(clock), .Q(tmp_value_2[3]) );
  DFQD1BWP12T tmp_value_2_reg_2_ ( .D(n394), .CP(clock), .Q(tmp_value_2[2]) );
  DFQD1BWP12T tmp_value_2_reg_1_ ( .D(n393), .CP(clock), .Q(tmp_value_2[1]) );
  DFQD1BWP12T tmp_value_2_reg_0_ ( .D(n392), .CP(clock), .Q(tmp_value_2[0]) );
  DFQD1BWP12T cpu_data_in_reg_31_ ( .D(n391), .CP(clock), .Q(cpu_data_in[31])
         );
  DFQD1BWP12T cpu_data_in_reg_30_ ( .D(n390), .CP(clock), .Q(cpu_data_in[30])
         );
  DFQD1BWP12T cpu_data_in_reg_29_ ( .D(n389), .CP(clock), .Q(cpu_data_in[29])
         );
  DFQD1BWP12T cpu_data_in_reg_28_ ( .D(n388), .CP(clock), .Q(cpu_data_in[28])
         );
  DFQD1BWP12T cpu_data_in_reg_27_ ( .D(n387), .CP(clock), .Q(cpu_data_in[27])
         );
  DFQD1BWP12T cpu_data_in_reg_26_ ( .D(n386), .CP(clock), .Q(cpu_data_in[26])
         );
  DFQD1BWP12T cpu_data_in_reg_25_ ( .D(n385), .CP(clock), .Q(cpu_data_in[25])
         );
  DFQD1BWP12T cpu_data_in_reg_24_ ( .D(n384), .CP(clock), .Q(cpu_data_in[24])
         );
  DFQD1BWP12T cpu_data_in_reg_23_ ( .D(n383), .CP(clock), .Q(cpu_data_in[23])
         );
  DFQD1BWP12T cpu_data_in_reg_22_ ( .D(n382), .CP(clock), .Q(cpu_data_in[22])
         );
  DFQD1BWP12T cpu_data_in_reg_21_ ( .D(n381), .CP(clock), .Q(cpu_data_in[21])
         );
  DFQD1BWP12T cpu_data_in_reg_20_ ( .D(n380), .CP(clock), .Q(cpu_data_in[20])
         );
  DFQD1BWP12T cpu_data_in_reg_19_ ( .D(n379), .CP(clock), .Q(cpu_data_in[19])
         );
  DFQD1BWP12T cpu_data_in_reg_18_ ( .D(n378), .CP(clock), .Q(cpu_data_in[18])
         );
  DFQD1BWP12T cpu_data_in_reg_17_ ( .D(n377), .CP(clock), .Q(cpu_data_in[17])
         );
  DFQD1BWP12T cpu_data_in_reg_16_ ( .D(n376), .CP(clock), .Q(cpu_data_in[16])
         );
  DFQD1BWP12T cpu_data_in_reg_15_ ( .D(n375), .CP(clock), .Q(cpu_data_in[15])
         );
  DFQD1BWP12T cpu_data_in_reg_14_ ( .D(n374), .CP(clock), .Q(cpu_data_in[14])
         );
  DFQD1BWP12T cpu_data_in_reg_13_ ( .D(n373), .CP(clock), .Q(cpu_data_in[13])
         );
  DFQD1BWP12T cpu_data_in_reg_12_ ( .D(n372), .CP(clock), .Q(cpu_data_in[12])
         );
  DFQD1BWP12T cpu_data_in_reg_11_ ( .D(n371), .CP(clock), .Q(cpu_data_in[11])
         );
  DFQD1BWP12T cpu_data_in_reg_10_ ( .D(n370), .CP(clock), .Q(cpu_data_in[10])
         );
  DFQD1BWP12T cpu_data_in_reg_9_ ( .D(n369), .CP(clock), .Q(cpu_data_in[9]) );
  DFQD1BWP12T cpu_data_in_reg_8_ ( .D(n368), .CP(clock), .Q(cpu_data_in[8]) );
  DFQD1BWP12T cpu_data_in_reg_7_ ( .D(n367), .CP(clock), .Q(cpu_data_in[7]) );
  DFQD1BWP12T cpu_data_in_reg_6_ ( .D(n366), .CP(clock), .Q(cpu_data_in[6]) );
  DFQD1BWP12T cpu_data_in_reg_5_ ( .D(n365), .CP(clock), .Q(cpu_data_in[5]) );
  DFQD1BWP12T cpu_data_in_reg_4_ ( .D(n364), .CP(clock), .Q(cpu_data_in[4]) );
  DFQD1BWP12T cpu_data_in_reg_3_ ( .D(n363), .CP(clock), .Q(cpu_data_in[3]) );
  DFQD1BWP12T cpu_data_in_reg_2_ ( .D(n362), .CP(clock), .Q(cpu_data_in[2]) );
  DFQD1BWP12T cpu_data_in_reg_1_ ( .D(n361), .CP(clock), .Q(cpu_data_in[1]) );
  DFQD1BWP12T cpu_data_in_reg_0_ ( .D(n360), .CP(clock), .Q(cpu_data_in[0]) );
  DFQD1BWP12T cpu_address_in_reg_12_ ( .D(n359), .CP(clock), .Q(
        cpu_address_in[12]) );
  DFQD1BWP12T cpu_address_in_reg_11_ ( .D(n358), .CP(clock), .Q(
        cpu_address_in[11]) );
  DFQD1BWP12T cpu_address_in_reg_10_ ( .D(n357), .CP(clock), .Q(
        cpu_address_in[10]) );
  DFQD1BWP12T cpu_address_in_reg_9_ ( .D(n356), .CP(clock), .Q(
        cpu_address_in[9]) );
  DFQD1BWP12T cpu_address_in_reg_8_ ( .D(n355), .CP(clock), .Q(
        cpu_address_in[8]) );
  DFQD1BWP12T cpu_address_in_reg_7_ ( .D(n354), .CP(clock), .Q(
        cpu_address_in[7]) );
  DFQD1BWP12T cpu_address_in_reg_6_ ( .D(n353), .CP(clock), .Q(
        cpu_address_in[6]) );
  DFQD1BWP12T cpu_address_in_reg_5_ ( .D(n352), .CP(clock), .Q(
        cpu_address_in[5]) );
  DFQD1BWP12T cpu_address_in_reg_4_ ( .D(n351), .CP(clock), .Q(
        cpu_address_in[4]) );
  DFQD1BWP12T cpu_address_in_reg_3_ ( .D(n350), .CP(clock), .Q(
        cpu_address_in[3]) );
  DFQD1BWP12T cpu_address_in_reg_2_ ( .D(n349), .CP(clock), .Q(
        cpu_address_in[2]) );
  DFQD1BWP12T cpu_address_in_reg_1_ ( .D(n348), .CP(clock), .Q(
        cpu_address_in[1]) );
  DFQD1BWP12T sign_extend_reg ( .D(n346), .CP(clock), .Q(sign_extend) );
  DFQD1BWP12T interface_cpu_data_out_reg_8_ ( .D(N82), .CP(clock), .Q(
        interface_cpu_data_out[8]) );
  DFQD1BWP12T interface_cpu_data_out_reg_9_ ( .D(N83), .CP(clock), .Q(
        interface_cpu_data_out[9]) );
  DFQD1BWP12T interface_cpu_data_out_reg_10_ ( .D(N84), .CP(clock), .Q(
        interface_cpu_data_out[10]) );
  DFQD1BWP12T interface_cpu_data_out_reg_11_ ( .D(N85), .CP(clock), .Q(
        interface_cpu_data_out[11]) );
  DFQD1BWP12T interface_cpu_data_out_reg_12_ ( .D(N86), .CP(clock), .Q(
        interface_cpu_data_out[12]) );
  DFQD1BWP12T interface_cpu_data_out_reg_13_ ( .D(N87), .CP(clock), .Q(
        interface_cpu_data_out[13]) );
  DFQD1BWP12T interface_cpu_data_out_reg_14_ ( .D(N88), .CP(clock), .Q(
        interface_cpu_data_out[14]) );
  DFQD1BWP12T interface_cpu_data_out_reg_15_ ( .D(N89), .CP(clock), .Q(
        interface_cpu_data_out[15]) );
  DFQD1BWP12T interface_cpu_data_out_reg_16_ ( .D(N90), .CP(clock), .Q(
        interface_cpu_data_out[16]) );
  DFQD1BWP12T interface_cpu_data_out_reg_17_ ( .D(N91), .CP(clock), .Q(
        interface_cpu_data_out[17]) );
  DFQD1BWP12T interface_cpu_data_out_reg_18_ ( .D(N92), .CP(clock), .Q(
        interface_cpu_data_out[18]) );
  DFQD1BWP12T interface_cpu_data_out_reg_19_ ( .D(N93), .CP(clock), .Q(
        interface_cpu_data_out[19]) );
  DFQD1BWP12T interface_cpu_data_out_reg_20_ ( .D(N94), .CP(clock), .Q(
        interface_cpu_data_out[20]) );
  DFQD1BWP12T interface_cpu_data_out_reg_21_ ( .D(N95), .CP(clock), .Q(
        interface_cpu_data_out[21]) );
  DFQD1BWP12T interface_cpu_data_out_reg_22_ ( .D(N96), .CP(clock), .Q(
        interface_cpu_data_out[22]) );
  DFQD1BWP12T interface_cpu_data_out_reg_23_ ( .D(N97), .CP(clock), .Q(
        interface_cpu_data_out[23]) );
  DFQD1BWP12T interface_cpu_data_out_reg_24_ ( .D(N98), .CP(clock), .Q(
        interface_cpu_data_out[24]) );
  DFQD1BWP12T interface_cpu_data_out_reg_25_ ( .D(N99), .CP(clock), .Q(
        interface_cpu_data_out[25]) );
  DFQD1BWP12T interface_cpu_data_out_reg_26_ ( .D(N100), .CP(clock), .Q(
        interface_cpu_data_out[26]) );
  DFQD1BWP12T interface_cpu_data_out_reg_27_ ( .D(N101), .CP(clock), .Q(
        interface_cpu_data_out[27]) );
  DFQD1BWP12T interface_cpu_data_out_reg_28_ ( .D(N102), .CP(clock), .Q(
        interface_cpu_data_out[28]) );
  DFQD1BWP12T interface_cpu_data_out_reg_29_ ( .D(N103), .CP(clock), .Q(
        interface_cpu_data_out[29]) );
  DFQD1BWP12T interface_cpu_data_out_reg_30_ ( .D(N104), .CP(clock), .Q(
        interface_cpu_data_out[30]) );
  DFQD1BWP12T interface_cpu_data_out_reg_31_ ( .D(N105), .CP(clock), .Q(
        interface_cpu_data_out[31]) );
  DFQD1BWP12T to_mem_address_reg_11_ ( .D(N194), .CP(clock), .Q(
        to_mem_address[11]) );
  DFQD1BWP12T to_mem_address_reg_10_ ( .D(N193), .CP(clock), .Q(
        to_mem_address[10]) );
  DFQD1BWP12T to_mem_address_reg_9_ ( .D(N192), .CP(clock), .Q(
        to_mem_address[9]) );
  DFQD1BWP12T to_mem_address_reg_8_ ( .D(N191), .CP(clock), .Q(
        to_mem_address[8]) );
  DFQD1BWP12T to_mem_address_reg_7_ ( .D(N190), .CP(clock), .Q(
        to_mem_address[7]) );
  DFQD1BWP12T to_mem_address_reg_6_ ( .D(N189), .CP(clock), .Q(
        to_mem_address[6]) );
  DFQD1BWP12T to_mem_address_reg_5_ ( .D(N188), .CP(clock), .Q(
        to_mem_address[5]) );
  DFQD1BWP12T to_mem_address_reg_4_ ( .D(N187), .CP(clock), .Q(
        to_mem_address[4]) );
  DFQD1BWP12T to_mem_address_reg_3_ ( .D(N186), .CP(clock), .Q(
        to_mem_address[3]) );
  DFQD1BWP12T to_mem_address_reg_2_ ( .D(N185), .CP(clock), .Q(
        to_mem_address[2]) );
  DFQD1BWP12T to_mem_address_reg_1_ ( .D(N184), .CP(clock), .Q(
        to_mem_address[1]) );
  DFQD1BWP12T to_mem_address_reg_0_ ( .D(N183), .CP(clock), .Q(
        to_mem_address[0]) );
  DFQD1BWP12T to_mem_data_in_reg_15_ ( .D(N210), .CP(clock), .Q(
        to_mem_data_in[15]) );
  DFQD1BWP12T to_mem_data_in_reg_14_ ( .D(N209), .CP(clock), .Q(
        to_mem_data_in[14]) );
  DFQD1BWP12T to_mem_data_in_reg_13_ ( .D(N208), .CP(clock), .Q(
        to_mem_data_in[13]) );
  DFQD1BWP12T to_mem_data_in_reg_12_ ( .D(N207), .CP(clock), .Q(
        to_mem_data_in[12]) );
  DFQD1BWP12T to_mem_data_in_reg_11_ ( .D(N206), .CP(clock), .Q(
        to_mem_data_in[11]) );
  DFQD1BWP12T to_mem_data_in_reg_10_ ( .D(N205), .CP(clock), .Q(
        to_mem_data_in[10]) );
  DFQD1BWP12T to_mem_data_in_reg_9_ ( .D(N204), .CP(clock), .Q(
        to_mem_data_in[9]) );
  DFQD1BWP12T to_mem_data_in_reg_8_ ( .D(N203), .CP(clock), .Q(
        to_mem_data_in[8]) );
  DFQD1BWP12T to_mem_data_in_reg_7_ ( .D(N202), .CP(clock), .Q(
        to_mem_data_in[7]) );
  DFQD1BWP12T to_mem_data_in_reg_6_ ( .D(N201), .CP(clock), .Q(
        to_mem_data_in[6]) );
  DFQD1BWP12T to_mem_data_in_reg_5_ ( .D(N200), .CP(clock), .Q(
        to_mem_data_in[5]) );
  DFQD1BWP12T to_mem_data_in_reg_4_ ( .D(N199), .CP(clock), .Q(
        to_mem_data_in[4]) );
  DFQD1BWP12T to_mem_data_in_reg_3_ ( .D(N198), .CP(clock), .Q(
        to_mem_data_in[3]) );
  DFQD1BWP12T to_mem_data_in_reg_2_ ( .D(N197), .CP(clock), .Q(
        to_mem_data_in[2]) );
  DFQD1BWP12T to_mem_data_in_reg_1_ ( .D(N196), .CP(clock), .Q(
        to_mem_data_in[1]) );
  DFQD1BWP12T to_mem_data_in_reg_0_ ( .D(N195), .CP(clock), .Q(
        to_mem_data_in[0]) );
  DFQD1BWP12T to_mem_read_enable_reg ( .D(N211), .CP(clock), .Q(
        to_mem_read_enable) );
  INVD1BWP12T U3 ( .I(n314), .ZN(n60) );
  INR2D1BWP12T U4 ( .A1(n226), .B1(n34), .ZN(n41) );
  IND2D1BWP12T U5 ( .A1(state[4]), .B1(state[5]), .ZN(n33) );
  ND2D1BWP12T U6 ( .A1(n20), .A2(n30), .ZN(n34) );
  NR2D1BWP12T U7 ( .A1(state[2]), .A2(state[3]), .ZN(n226) );
  INVD1BWP12T U8 ( .I(n29), .ZN(n24) );
  INR2D1BWP12T U9 ( .A1(n22), .B1(n33), .ZN(n68) );
  INR2D1BWP12T U10 ( .A1(state[3]), .B1(n92), .ZN(n31) );
  INVD1BWP12T U11 ( .I(n126), .ZN(n288) );
  NR4D0BWP12T U12 ( .A1(n40), .A2(n39), .A3(n38), .A4(n271), .ZN(n321) );
  INVD1BWP12T U13 ( .I(state[0]), .ZN(n20) );
  NR2D1BWP12T U14 ( .A1(n34), .A2(n33), .ZN(n251) );
  ND2D1BWP12T U15 ( .A1(n105), .A2(n31), .ZN(n170) );
  ND2D1BWP12T U16 ( .A1(n222), .A2(n31), .ZN(n203) );
  HA1D0BWP12T U17 ( .A(n241), .B(cpu_address_in[3]), .CO(n277), .S(n242) );
  HA1D0BWP12T U18 ( .A(n277), .B(cpu_address_in[4]), .CO(n279), .S(n278) );
  HA1D0BWP12T U19 ( .A(n279), .B(cpu_address_in[5]), .CO(n281), .S(n280) );
  HA1D0BWP12T U20 ( .A(n281), .B(cpu_address_in[6]), .CO(n283), .S(n282) );
  HA1D0BWP12T U21 ( .A(n283), .B(cpu_address_in[7]), .CO(n285), .S(n284) );
  HA1D0BWP12T U22 ( .A(n285), .B(cpu_address_in[8]), .CO(n287), .S(n286) );
  HA1D0BWP12T U23 ( .A(n287), .B(cpu_address_in[9]), .CO(n124), .S(n290) );
  HA1D0BWP12T U24 ( .A(n124), .B(cpu_address_in[10]), .CO(n121), .S(n125) );
  OAI31D1BWP12T U25 ( .A1(n297), .A2(n49), .A3(n48), .B(n256), .ZN(n126) );
  HA1D0BWP12T U26 ( .A(n121), .B(cpu_address_in[11]), .CO(n119), .S(n122) );
  ND2D1BWP12T U27 ( .A1(n256), .A2(n130), .ZN(n169) );
  NR2D1BWP12T U28 ( .A1(n61), .A2(n60), .ZN(n273) );
  NR2D1BWP12T U29 ( .A1(reset), .A2(n127), .ZN(n272) );
  INR2D1BWP12T U30 ( .A1(n105), .B1(n95), .ZN(n270) );
  INVD1BWP12T U31 ( .I(n321), .ZN(n94) );
  AOI21D1BWP12T U32 ( .A1(n308), .A2(n44), .B(reset), .ZN(n451) );
  INVD1BWP12T U33 ( .I(n324), .ZN(n340) );
  ND2D1BWP12T U34 ( .A1(n68), .A2(n37), .ZN(n248) );
  ND4D1BWP12T U35 ( .A1(n324), .A2(n248), .A3(n247), .A4(n342), .ZN(n322) );
  INVD1BWP12T U36 ( .I(n322), .ZN(n265) );
  ND2D1BWP12T U37 ( .A1(n256), .A2(n295), .ZN(n323) );
  INVD1BWP12T U38 ( .I(n248), .ZN(n271) );
  NR2D1BWP12T U39 ( .A1(state[4]), .A2(state[5]), .ZN(n107) );
  NR2D1BWP12T U40 ( .A1(n106), .A2(n33), .ZN(n105) );
  INVD1BWP12T U41 ( .I(reset), .ZN(n256) );
  INR2D1BWP12T U42 ( .A1(state[3]), .B1(state[2]), .ZN(n312) );
  INR2D1BWP12T U43 ( .A1(state[2]), .B1(state[3]), .ZN(n314) );
  OAI21D1BWP12T U44 ( .A1(n246), .A2(n245), .B(n256), .ZN(n342) );
  INR2D1BWP12T U45 ( .A1(n312), .B1(n51), .ZN(n245) );
  ND2D1BWP12T U46 ( .A1(n41), .A2(n107), .ZN(n308) );
  INR2D1BWP12T U47 ( .A1(n170), .B1(n50), .ZN(n293) );
  ND3D1BWP12T U48 ( .A1(n251), .A2(n312), .A3(n256), .ZN(n302) );
  MOAI22D0BWP12T U49 ( .A1(n320), .A2(n126), .B1(n125), .B2(n289), .ZN(N192)
         );
  MOAI22D0BWP12T U50 ( .A1(n123), .A2(n126), .B1(n122), .B2(n289), .ZN(N193)
         );
  MOAI22D0BWP12T U51 ( .A1(n321), .A2(n120), .B1(interface_cpu_address_in[12]), 
        .B2(n451), .ZN(n359) );
  AO22D0BWP12T U52 ( .A1(n94), .A2(cpu_address_in[1]), .B1(n451), .B2(
        interface_cpu_address_in[1]), .Z(n348) );
  MOAI22D0BWP12T U53 ( .A1(n453), .A2(n431), .B1(n451), .B2(
        interface_cpu_data_in[20]), .ZN(n380) );
  AO22D0BWP12T U54 ( .A1(n94), .A2(cpu_address_in[2]), .B1(n451), .B2(
        interface_cpu_address_in[2]), .Z(n349) );
  AO22D0BWP12T U55 ( .A1(n94), .A2(cpu_address_in[3]), .B1(n451), .B2(
        interface_cpu_address_in[3]), .Z(n350) );
  AO22D0BWP12T U56 ( .A1(n94), .A2(cpu_address_in[4]), .B1(n451), .B2(
        interface_cpu_address_in[4]), .Z(n351) );
  AO22D0BWP12T U57 ( .A1(n94), .A2(cpu_address_in[5]), .B1(n451), .B2(
        interface_cpu_address_in[5]), .Z(n352) );
  AO22D0BWP12T U58 ( .A1(n94), .A2(cpu_address_in[6]), .B1(n451), .B2(
        interface_cpu_address_in[6]), .Z(n353) );
  CKND2D0BWP12T U59 ( .A1(n312), .A2(n68), .ZN(n1) );
  OAI211D0BWP12T U60 ( .A1(n51), .A2(n60), .B(n244), .C(n1), .ZN(n71) );
  MAOI22D0BWP12T U61 ( .A1(cpu_address_in[12]), .A2(n119), .B1(
        cpu_address_in[12]), .B2(n119), .ZN(n2) );
  MOAI22D0BWP12T U62 ( .A1(n120), .A2(n126), .B1(n289), .B2(n2), .ZN(N194) );
  AO22D0BWP12T U63 ( .A1(n94), .A2(cpu_address_in[7]), .B1(n451), .B2(
        interface_cpu_address_in[7]), .Z(n354) );
  ND4D0BWP12T U64 ( .A1(n182), .A2(n73), .A3(n103), .A4(n230), .ZN(n3) );
  ND2D1BWP12T U65 ( .A1(n181), .A2(n303), .ZN(n4) );
  AOI211D1BWP12T U66 ( .A1(n256), .A2(n3), .B(N212), .C(n4), .ZN(n453) );
  AO22D0BWP12T U67 ( .A1(n94), .A2(cpu_address_in[8]), .B1(n451), .B2(
        interface_cpu_address_in[8]), .Z(n355) );
  OAI22D0BWP12T U68 ( .A1(n100), .A2(state[5]), .B1(n254), .B2(n101), .ZN(n5)
         );
  INR3D0BWP12T U69 ( .A1(n171), .B1(n102), .B2(n5), .ZN(n6) );
  OAI211D0BWP12T U70 ( .A1(n305), .A2(n104), .B(n103), .C(n6), .ZN(n319) );
  AO22D0BWP12T U71 ( .A1(n94), .A2(cpu_address_in[9]), .B1(n451), .B2(
        interface_cpu_address_in[9]), .Z(n356) );
  IND2D0BWP12T U72 ( .A1(state[4]), .B1(n23), .ZN(n108) );
  MOAI22D0BWP12T U73 ( .A1(n321), .A2(n320), .B1(n451), .B2(
        interface_cpu_address_in[10]), .ZN(n357) );
  OA21D0BWP12T U74 ( .A1(n316), .A2(n315), .B(n314), .Z(n7) );
  AOI21D0BWP12T U75 ( .A1(n312), .A2(n313), .B(n311), .ZN(n8) );
  OAI211D0BWP12T U76 ( .A1(n310), .A2(state[1]), .B(n317), .C(n8), .ZN(n9) );
  NR4D0BWP12T U77 ( .A1(n319), .A2(n318), .A3(n7), .A4(n9), .ZN(n10) );
  NR3D0BWP12T U78 ( .A1(interface_cpu_word_type[0]), .A2(n309), .A3(n308), 
        .ZN(n11) );
  NR2D0BWP12T U79 ( .A1(n305), .A2(n306), .ZN(n12) );
  AOI22D0BWP12T U80 ( .A1(interface_cpu_address_in[0]), .A2(n11), .B1(n307), 
        .B2(n12), .ZN(n13) );
  AOI32D0BWP12T U81 ( .A1(n10), .A2(n342), .A3(n13), .B1(reset), .B2(n342), 
        .ZN(N68) );
  AO21D0BWP12T U82 ( .A1(n222), .A2(state[3]), .B(n318), .Z(n118) );
  OAI21D0BWP12T U83 ( .A1(interface_cpu_word_type[1]), .A2(
        interface_cpu_address_in[0]), .B(n292), .ZN(n14) );
  OR4D0BWP12T U84 ( .A1(n109), .A2(n246), .A3(n227), .A4(n102), .Z(n15) );
  AOI211D0BWP12T U85 ( .A1(n114), .A2(n14), .B(n294), .C(n15), .ZN(n16) );
  OAI32D0BWP12T U86 ( .A1(reset), .A2(n104), .A3(n308), .B1(n16), .B2(reset), 
        .ZN(N67) );
  CKND0BWP12T U87 ( .I(n224), .ZN(n17) );
  AOI22D0BWP12T U88 ( .A1(n89), .A2(n314), .B1(n226), .B2(n17), .ZN(n212) );
  AOI21D0BWP12T U89 ( .A1(n243), .A2(n244), .B(reset), .ZN(n18) );
  NR2D0BWP12T U90 ( .A1(n270), .A2(n18), .ZN(n324) );
  AN2D0BWP12T U91 ( .A1(n107), .A2(n22), .Z(n227) );
  MOAI22D0BWP12T U92 ( .A1(n321), .A2(n123), .B1(n451), .B2(
        interface_cpu_address_in[11]), .ZN(n358) );
  IND2D0BWP12T U93 ( .A1(n50), .B1(n203), .ZN(n176) );
  IND2D0BWP12T U94 ( .A1(n315), .B1(n83), .ZN(n299) );
  OA21D0BWP12T U95 ( .A1(n231), .A2(n118), .B(n256), .Z(n289) );
  AOI211D0BWP12T U96 ( .A1(n80), .A2(n79), .B(n81), .C(n82), .ZN(n19) );
  AOI21D0BWP12T U97 ( .A1(n19), .A2(n83), .B(reset), .ZN(N71) );
  INVD1BWP12T U98 ( .I(state[5]), .ZN(n27) );
  INR2D1BWP12T U99 ( .A1(state[1]), .B1(n20), .ZN(n23) );
  INR2D1BWP12T U100 ( .A1(n27), .B1(n108), .ZN(n313) );
  ND2D1BWP12T U101 ( .A1(n20), .A2(state[1]), .ZN(n106) );
  INVD1BWP12T U102 ( .I(state[1]), .ZN(n30) );
  IND2D1BWP12T U103 ( .A1(state[5]), .B1(state[4]), .ZN(n29) );
  NR2XD0BWP12T U104 ( .A1(n34), .A2(n29), .ZN(n315) );
  OA31D0BWP12T U105 ( .A1(n105), .A2(n313), .A3(n315), .B(n312), .Z(n21) );
  RCAOI21D0BWP12T U106 ( .A1(n314), .A2(n313), .B(n21), .ZN(n230) );
  INR2D1BWP12T U107 ( .A1(state[5]), .B1(n108), .ZN(n222) );
  INVD1BWP12T U108 ( .I(n34), .ZN(n26) );
  INVD1BWP12T U109 ( .I(state[2]), .ZN(n92) );
  ND2D1BWP12T U110 ( .A1(n26), .A2(n31), .ZN(n100) );
  NR2D1BWP12T U111 ( .A1(n100), .A2(n33), .ZN(n249) );
  AOI21D0BWP12T U112 ( .A1(n312), .A2(n222), .B(n249), .ZN(n103) );
  INR2D1BWP12T U113 ( .A1(state[0]), .B1(state[1]), .ZN(n22) );
  ND2D1BWP12T U114 ( .A1(n24), .A2(n22), .ZN(n224) );
  INVD1BWP12T U115 ( .I(n224), .ZN(n52) );
  NR2D1BWP12T U116 ( .A1(n106), .A2(n29), .ZN(n316) );
  TPOAI21D0BWP12T U117 ( .A1(n52), .A2(n316), .B(n312), .ZN(n73) );
  INR2XD0BWP12T U118 ( .A1(n107), .B1(n106), .ZN(n89) );
  CKND2D0BWP12T U119 ( .A1(n89), .A2(state[3]), .ZN(n182) );
  OAI21D1BWP12T U120 ( .A1(n316), .A2(n222), .B(n314), .ZN(n172) );
  ND2D1BWP12T U121 ( .A1(n227), .A2(n31), .ZN(n171) );
  ND2D1BWP12T U122 ( .A1(n172), .A2(n171), .ZN(n206) );
  ND2D1BWP12T U123 ( .A1(n24), .A2(n23), .ZN(n51) );
  AOI21D1BWP12T U124 ( .A1(n68), .A2(n31), .B(n245), .ZN(n202) );
  ND2D1BWP12T U125 ( .A1(n227), .A2(n312), .ZN(n201) );
  ND2D1BWP12T U126 ( .A1(n202), .A2(n201), .ZN(n145) );
  NR2D1BWP12T U127 ( .A1(n206), .A2(n145), .ZN(n47) );
  INVD1BWP12T U128 ( .I(n170), .ZN(n102) );
  INR2D1BWP12T U129 ( .A1(n24), .B1(n100), .ZN(n50) );
  NR2D1BWP12T U130 ( .A1(n102), .A2(n176), .ZN(n243) );
  IOA21D1BWP12T U131 ( .A1(n47), .A2(n243), .B(n256), .ZN(n25) );
  ND2D1BWP12T U132 ( .A1(n25), .A2(n302), .ZN(N212) );
  ND4D1BWP12T U133 ( .A1(n26), .A2(n107), .A3(state[3]), .A4(n256), .ZN(n303)
         );
  INR2D1BWP12T U134 ( .A1(state[4]), .B1(n27), .ZN(n42) );
  AOI22D1BWP12T U135 ( .A1(n41), .A2(n42), .B1(n52), .B2(n31), .ZN(n244) );
  ND2D1BWP12T U136 ( .A1(n256), .A2(n71), .ZN(n181) );
  INVD1BWP12T U137 ( .I(n453), .ZN(n40) );
  INR2D1BWP12T U138 ( .A1(n256), .B1(n224), .ZN(n59) );
  ND2D1BWP12T U139 ( .A1(n59), .A2(n226), .ZN(n276) );
  INVD1BWP12T U140 ( .I(n276), .ZN(n39) );
  INR2D1BWP12T U141 ( .A1(n251), .B1(n60), .ZN(n318) );
  INR2XD0BWP12T U142 ( .A1(n31), .B1(n51), .ZN(n82) );
  INVD1BWP12T U143 ( .I(n82), .ZN(n28) );
  ND2XD0BWP12T U144 ( .A1(n222), .A2(n226), .ZN(n317) );
  ND2D1BWP12T U145 ( .A1(n28), .A2(n317), .ZN(n55) );
  CKND0BWP12T U146 ( .I(n226), .ZN(n69) );
  ND2XD0BWP12T U147 ( .A1(n313), .A2(n31), .ZN(n46) );
  OAI31D0BWP12T U148 ( .A1(n30), .A2(n69), .A3(n29), .B(n46), .ZN(n62) );
  INVD0BWP12T U149 ( .I(n105), .ZN(n87) );
  INVD1BWP12T U150 ( .I(n316), .ZN(n254) );
  INVD0BWP12T U151 ( .I(n31), .ZN(n101) );
  OAI22D0BWP12T U152 ( .A1(n69), .A2(n87), .B1(n254), .B2(n101), .ZN(n32) );
  NR4D0BWP12T U153 ( .A1(n318), .A2(n55), .A3(n62), .A4(n32), .ZN(n229) );
  CKND0BWP12T U154 ( .I(n33), .ZN(n81) );
  CKND2D1BWP12T U155 ( .A1(n314), .A2(n107), .ZN(n310) );
  NR2D1BWP12T U156 ( .A1(n310), .A2(n34), .ZN(n297) );
  CKND0BWP12T U157 ( .I(state[3]), .ZN(n250) );
  OAI31D0BWP12T U158 ( .A1(n89), .A2(n315), .A3(n227), .B(n250), .ZN(n35) );
  ND2D1BWP12T U159 ( .A1(n313), .A2(n226), .ZN(n96) );
  IND3D0BWP12T U160 ( .A1(n297), .B1(n35), .B2(n96), .ZN(n63) );
  AOI21D1BWP12T U161 ( .A1(n87), .A2(n224), .B(n60), .ZN(n219) );
  RCAOI211D0BWP12T U162 ( .A1(n81), .A2(n41), .B(n63), .C(n219), .ZN(n36) );
  AOI21D1BWP12T U163 ( .A1(n229), .A2(n36), .B(reset), .ZN(n38) );
  INR2D1BWP12T U164 ( .A1(n226), .B1(reset), .ZN(n37) );
  INVD1BWP12T U165 ( .I(cpu_address_in[12]), .ZN(n120) );
  INVD1BWP12T U166 ( .I(n41), .ZN(n43) );
  ND2D1BWP12T U167 ( .A1(n43), .A2(n42), .ZN(n44) );
  INVD1BWP12T U168 ( .I(cpu_address_in[11]), .ZN(n123) );
  AOI21D1BWP12T U169 ( .A1(n69), .A2(n101), .B(n254), .ZN(n49) );
  OAI21D0BWP12T U170 ( .A1(n227), .A2(n105), .B(n226), .ZN(n45) );
  ND4D1BWP12T U171 ( .A1(n230), .A2(n47), .A3(n46), .A4(n45), .ZN(n48) );
  INR2XD0BWP12T U172 ( .A1(n226), .B1(n51), .ZN(n311) );
  INVD1BWP12T U173 ( .I(n311), .ZN(n54) );
  OAI21D0BWP12T U174 ( .A1(n52), .A2(n251), .B(n312), .ZN(n53) );
  AN3XD1BWP12T U175 ( .A1(n293), .A2(n54), .A3(n53), .Z(n57) );
  INVD1BWP12T U176 ( .I(n55), .ZN(n56) );
  ND2D1BWP12T U177 ( .A1(n57), .A2(n56), .ZN(n231) );
  AO22XD1BWP12T U178 ( .A1(n288), .A2(cpu_address_in[2]), .B1(n58), .B2(n289), 
        .Z(N184) );
  INVD1BWP12T U179 ( .I(n59), .ZN(n61) );
  INVD1BWP12T U180 ( .I(n273), .ZN(n247) );
  OAI21D0BWP12T U181 ( .A1(n63), .A2(n62), .B(n256), .ZN(n64) );
  ND4D0BWP12T U182 ( .A1(n276), .A2(n303), .A3(n247), .A4(n64), .ZN(n65) );
  AO22XD1BWP12T U183 ( .A1(n451), .A2(interface_cpu_sign_extend), .B1(
        sign_extend), .B2(n65), .Z(n346) );
  INVD1BWP12T U184 ( .I(n96), .ZN(n218) );
  NR2D0BWP12T U185 ( .A1(n218), .A2(n219), .ZN(n66) );
  CKND2D1BWP12T U186 ( .A1(n212), .A2(n66), .ZN(n72) );
  AO21D0BWP12T U187 ( .A1(n72), .A2(n256), .B(n271), .Z(N72) );
  CKND0BWP12T U188 ( .I(interface_cpu_word_type[1]), .ZN(n84) );
  INVD1BWP12T U189 ( .I(n308), .ZN(n67) );
  NR2D1BWP12T U190 ( .A1(interface_cpu_load_request), .A2(
        interface_cpu_store_request_BAR), .ZN(n291) );
  ND2D1BWP12T U191 ( .A1(n67), .A2(n291), .ZN(n91) );
  INVD1BWP12T U192 ( .I(n91), .ZN(n114) );
  AO31D1BWP12T U193 ( .A1(interface_cpu_address_in[0]), .A2(
        interface_cpu_load_request), .A3(n67), .B(n114), .Z(n80) );
  IND2XD1BWP12T U194 ( .A1(interface_cpu_word_type[0]), .B1(
        interface_cpu_word_type[1]), .ZN(n292) );
  INVD1BWP12T U195 ( .I(n292), .ZN(n79) );
  CKND2D1BWP12T U196 ( .A1(n79), .A2(interface_cpu_load_request), .ZN(n85) );
  NR2D1BWP12T U197 ( .A1(interface_cpu_address_in[0]), .A2(n308), .ZN(n301) );
  INVD1BWP12T U198 ( .I(n301), .ZN(n305) );
  INVD1BWP12T U199 ( .I(n68), .ZN(n93) );
  OAI21D0BWP12T U200 ( .A1(n93), .A2(n69), .B(n182), .ZN(n70) );
  NR3XD0BWP12T U201 ( .A1(n72), .A2(n71), .A3(n70), .ZN(n83) );
  INVD1BWP12T U202 ( .I(n299), .ZN(n76) );
  INVD1BWP12T U203 ( .I(n73), .ZN(n109) );
  OAI21D0BWP12T U204 ( .A1(n108), .A2(n101), .B(n254), .ZN(n74) );
  NR4D0BWP12T U205 ( .A1(n109), .A2(n245), .A3(n311), .A4(n74), .ZN(n75) );
  OAI211D1BWP12T U206 ( .A1(n85), .A2(n305), .B(n76), .C(n75), .ZN(n77) );
  AOI31D1BWP12T U207 ( .A1(interface_cpu_word_type[0]), .A2(n84), .A3(n80), 
        .B(n77), .ZN(n78) );
  NR2D1BWP12T U208 ( .A1(n78), .A2(reset), .ZN(N70) );
  CKND0BWP12T U209 ( .I(interface_cpu_word_type[0]), .ZN(n86) );
  CKND2D1BWP12T U210 ( .A1(n84), .A2(interface_cpu_load_request), .ZN(n309) );
  OA21D1BWP12T U211 ( .A1(n86), .A2(n309), .B(n85), .Z(n104) );
  NR2D0BWP12T U212 ( .A1(n87), .A2(state[2]), .ZN(n88) );
  AOI211D0BWP12T U213 ( .A1(n226), .A2(n89), .B(n88), .C(n316), .ZN(n90) );
  TPOAI31D0BWP12T U214 ( .A1(interface_cpu_word_type[1]), .A2(
        interface_cpu_word_type[0]), .A3(n91), .B(n90), .ZN(n294) );
  NR2D1BWP12T U215 ( .A1(n93), .A2(n92), .ZN(n246) );
  INVD1BWP12T U216 ( .I(from_mem_data_out[7]), .ZN(n333) );
  ND2D1BWP12T U217 ( .A1(n314), .A2(n256), .ZN(n95) );
  AOI22D0BWP12T U218 ( .A1(n271), .A2(tmp_value_1[7]), .B1(n270), .B2(
        tmp_value_2[15]), .ZN(n99) );
  TPNR2D0BWP12T U219 ( .A1(n106), .A2(n310), .ZN(n97) );
  NR2D1BWP12T U220 ( .A1(n96), .A2(n333), .ZN(n214) );
  AOI32D1BWP12T U221 ( .A1(from_mem_data_out[15]), .A2(sign_extend), .A3(n97), 
        .B1(n214), .B2(sign_extend), .ZN(n127) );
  AOI21D0BWP12T U222 ( .A1(n273), .A2(from_mem_data_out[15]), .B(n272), .ZN(
        n98) );
  OAI211D0BWP12T U223 ( .A1(n276), .A2(n333), .B(n99), .C(n98), .ZN(N89) );
  CKND2D0BWP12T U224 ( .A1(interface_cpu_word_type[0]), .A2(
        interface_cpu_word_type[1]), .ZN(n307) );
  AOI211D0BWP12T U225 ( .A1(n107), .A2(n106), .B(n105), .C(n315), .ZN(n112) );
  INVD0BWP12T U226 ( .I(n312), .ZN(n255) );
  CKND0BWP12T U227 ( .I(n108), .ZN(n110) );
  AOI21D0BWP12T U228 ( .A1(n110), .A2(n314), .B(n109), .ZN(n111) );
  OAI211D1BWP12T U229 ( .A1(n112), .A2(n255), .B(n111), .C(n202), .ZN(n113) );
  AO31D1BWP12T U230 ( .A1(interface_cpu_address_in[0]), .A2(n114), .A3(n307), 
        .B(n113), .Z(n115) );
  OAI21D1BWP12T U231 ( .A1(n319), .A2(n115), .B(n256), .ZN(n116) );
  CKND2D1BWP12T U232 ( .A1(n116), .A2(n302), .ZN(N69) );
  FA1D0BWP12T U233 ( .A(cpu_address_in[2]), .B(n118), .CI(n117), .CO(n241), 
        .S(n58) );
  INVD1BWP12T U234 ( .I(cpu_address_in[10]), .ZN(n320) );
  INVD1BWP12T U235 ( .I(from_mem_data_out[14]), .ZN(n326) );
  AOI22D0BWP12T U236 ( .A1(n226), .A2(from_mem_data_out[7]), .B1(n314), .B2(
        from_mem_data_out[15]), .ZN(n129) );
  CKND0BWP12T U237 ( .I(sign_extend), .ZN(n128) );
  OAI31D1BWP12T U238 ( .A1(n129), .A2(n128), .A3(n224), .B(n127), .ZN(n130) );
  TPND2D0BWP12T U239 ( .A1(n270), .A2(tmp_value_2[6]), .ZN(n131) );
  OAI211D0BWP12T U240 ( .A1(n326), .A2(n248), .B(n169), .C(n131), .ZN(N96) );
  INVD1BWP12T U241 ( .I(from_mem_data_out[0]), .ZN(n341) );
  TPND2D0BWP12T U242 ( .A1(n270), .A2(from_mem_data_out[8]), .ZN(n132) );
  OAI211D0BWP12T U243 ( .A1(n341), .A2(n248), .B(n169), .C(n132), .ZN(N98) );
  INVD1BWP12T U244 ( .I(from_mem_data_out[15]), .ZN(n325) );
  TPND2D0BWP12T U245 ( .A1(n270), .A2(tmp_value_2[7]), .ZN(n133) );
  OAI211D0BWP12T U246 ( .A1(n325), .A2(n248), .B(n169), .C(n133), .ZN(N97) );
  INVD1BWP12T U247 ( .I(from_mem_data_out[4]), .ZN(n336) );
  TPND2D0BWP12T U248 ( .A1(n270), .A2(from_mem_data_out[12]), .ZN(n134) );
  OAI211D0BWP12T U249 ( .A1(n336), .A2(n248), .B(n169), .C(n134), .ZN(N102) );
  INVD1BWP12T U250 ( .I(from_mem_data_out[5]), .ZN(n335) );
  TPND2D0BWP12T U251 ( .A1(n270), .A2(from_mem_data_out[13]), .ZN(n135) );
  OAI211D0BWP12T U252 ( .A1(n335), .A2(n248), .B(n169), .C(n135), .ZN(N103) );
  INVD1BWP12T U253 ( .I(from_mem_data_out[1]), .ZN(n339) );
  TPND2D0BWP12T U254 ( .A1(n270), .A2(from_mem_data_out[9]), .ZN(n136) );
  OAI211D0BWP12T U255 ( .A1(n339), .A2(n248), .B(n169), .C(n136), .ZN(N99) );
  INVD1BWP12T U256 ( .I(from_mem_data_out[13]), .ZN(n327) );
  TPND2D0BWP12T U257 ( .A1(n270), .A2(tmp_value_2[5]), .ZN(n137) );
  OAI211D0BWP12T U258 ( .A1(n327), .A2(n248), .B(n169), .C(n137), .ZN(N95) );
  INVD1BWP12T U259 ( .I(from_mem_data_out[12]), .ZN(n328) );
  TPND2D0BWP12T U260 ( .A1(n270), .A2(tmp_value_2[4]), .ZN(n138) );
  OAI211D0BWP12T U261 ( .A1(n328), .A2(n248), .B(n169), .C(n138), .ZN(N94) );
  INVD1BWP12T U262 ( .I(from_mem_data_out[11]), .ZN(n329) );
  TPND2D0BWP12T U263 ( .A1(n270), .A2(tmp_value_2[3]), .ZN(n139) );
  OAI211D0BWP12T U264 ( .A1(n329), .A2(n248), .B(n169), .C(n139), .ZN(N93) );
  INVD1BWP12T U265 ( .I(from_mem_data_out[10]), .ZN(n330) );
  TPND2D0BWP12T U266 ( .A1(n270), .A2(tmp_value_2[2]), .ZN(n140) );
  OAI211D0BWP12T U267 ( .A1(n330), .A2(n248), .B(n169), .C(n140), .ZN(N92) );
  INVD1BWP12T U268 ( .I(from_mem_data_out[9]), .ZN(n331) );
  TPND2D0BWP12T U269 ( .A1(n270), .A2(tmp_value_2[1]), .ZN(n141) );
  OAI211D0BWP12T U270 ( .A1(n331), .A2(n248), .B(n169), .C(n141), .ZN(N91) );
  INVD1BWP12T U271 ( .I(from_mem_data_out[2]), .ZN(n338) );
  TPND2D0BWP12T U272 ( .A1(n270), .A2(from_mem_data_out[10]), .ZN(n142) );
  OAI211D0BWP12T U273 ( .A1(n338), .A2(n248), .B(n169), .C(n142), .ZN(N100) );
  INVD1BWP12T U274 ( .I(from_mem_data_out[8]), .ZN(n332) );
  TPND2D0BWP12T U275 ( .A1(n270), .A2(tmp_value_2[0]), .ZN(n143) );
  OAI211D0BWP12T U276 ( .A1(n332), .A2(n248), .B(n169), .C(n143), .ZN(N90) );
  INVD1BWP12T U277 ( .I(from_mem_data_out[3]), .ZN(n337) );
  TPND2D0BWP12T U278 ( .A1(n270), .A2(from_mem_data_out[11]), .ZN(n144) );
  OAI211D0BWP12T U279 ( .A1(n337), .A2(n248), .B(n169), .C(n144), .ZN(N101) );
  INVD1BWP12T U280 ( .I(cpu_data_in[23]), .ZN(n428) );
  OAI22D0BWP12T U281 ( .A1(n171), .A2(n333), .B1(n170), .B2(n428), .ZN(n147)
         );
  INVD1BWP12T U282 ( .I(n145), .ZN(n173) );
  INVD1BWP12T U283 ( .I(cpu_data_in[7]), .ZN(n444) );
  INVD1BWP12T U284 ( .I(cpu_data_in[15]), .ZN(n436) );
  OAI22D0BWP12T U285 ( .A1(n173), .A2(n444), .B1(n172), .B2(n436), .ZN(n146)
         );
  AOI211D0BWP12T U286 ( .A1(tmp_value_2[7]), .A2(n176), .B(n147), .C(n146), 
        .ZN(n148) );
  INVD1BWP12T U287 ( .I(cpu_data_in[31]), .ZN(n343) );
  OAI22D0BWP12T U288 ( .A1(reset), .A2(n148), .B1(n343), .B2(n302), .ZN(N202)
         );
  INVD1BWP12T U289 ( .I(from_mem_data_out[6]), .ZN(n334) );
  INVD1BWP12T U290 ( .I(cpu_data_in[22]), .ZN(n429) );
  OAI22D0BWP12T U291 ( .A1(n171), .A2(n334), .B1(n170), .B2(n429), .ZN(n150)
         );
  INVD1BWP12T U292 ( .I(cpu_data_in[6]), .ZN(n445) );
  INVD1BWP12T U293 ( .I(cpu_data_in[14]), .ZN(n437) );
  OAI22D0BWP12T U294 ( .A1(n173), .A2(n445), .B1(n172), .B2(n437), .ZN(n149)
         );
  AOI211D0BWP12T U295 ( .A1(tmp_value_2[6]), .A2(n176), .B(n150), .C(n149), 
        .ZN(n151) );
  INVD1BWP12T U296 ( .I(cpu_data_in[30]), .ZN(n344) );
  OAI22D0BWP12T U297 ( .A1(reset), .A2(n151), .B1(n344), .B2(n302), .ZN(N201)
         );
  INVD1BWP12T U298 ( .I(cpu_data_in[21]), .ZN(n430) );
  OAI22D0BWP12T U299 ( .A1(n171), .A2(n335), .B1(n170), .B2(n430), .ZN(n153)
         );
  INVD1BWP12T U300 ( .I(cpu_data_in[5]), .ZN(n446) );
  INVD1BWP12T U301 ( .I(cpu_data_in[13]), .ZN(n438) );
  OAI22D0BWP12T U302 ( .A1(n173), .A2(n446), .B1(n172), .B2(n438), .ZN(n152)
         );
  AOI211D0BWP12T U303 ( .A1(tmp_value_2[5]), .A2(n176), .B(n153), .C(n152), 
        .ZN(n154) );
  INVD1BWP12T U304 ( .I(cpu_data_in[29]), .ZN(n345) );
  OAI22D0BWP12T U305 ( .A1(reset), .A2(n154), .B1(n345), .B2(n302), .ZN(N200)
         );
  INVD1BWP12T U306 ( .I(cpu_data_in[20]), .ZN(n431) );
  OAI22D0BWP12T U307 ( .A1(n171), .A2(n336), .B1(n170), .B2(n431), .ZN(n156)
         );
  INVD1BWP12T U308 ( .I(cpu_data_in[4]), .ZN(n447) );
  INVD1BWP12T U309 ( .I(cpu_data_in[12]), .ZN(n439) );
  OAI22D0BWP12T U310 ( .A1(n173), .A2(n447), .B1(n172), .B2(n439), .ZN(n155)
         );
  AOI211D0BWP12T U311 ( .A1(tmp_value_2[4]), .A2(n176), .B(n156), .C(n155), 
        .ZN(n157) );
  INVD1BWP12T U312 ( .I(cpu_data_in[28]), .ZN(n347) );
  OAI22D0BWP12T U313 ( .A1(reset), .A2(n157), .B1(n347), .B2(n302), .ZN(N199)
         );
  INVD1BWP12T U314 ( .I(cpu_data_in[19]), .ZN(n432) );
  OAI22D0BWP12T U315 ( .A1(n171), .A2(n337), .B1(n170), .B2(n432), .ZN(n159)
         );
  INVD1BWP12T U316 ( .I(cpu_data_in[3]), .ZN(n448) );
  INVD1BWP12T U317 ( .I(cpu_data_in[11]), .ZN(n440) );
  OAI22D0BWP12T U318 ( .A1(n173), .A2(n448), .B1(n172), .B2(n440), .ZN(n158)
         );
  AOI211D0BWP12T U319 ( .A1(tmp_value_2[3]), .A2(n176), .B(n159), .C(n158), 
        .ZN(n160) );
  INVD1BWP12T U320 ( .I(cpu_data_in[27]), .ZN(n424) );
  OAI22D0BWP12T U321 ( .A1(reset), .A2(n160), .B1(n424), .B2(n302), .ZN(N198)
         );
  INVD1BWP12T U322 ( .I(cpu_data_in[18]), .ZN(n433) );
  OAI22D0BWP12T U323 ( .A1(n171), .A2(n338), .B1(n170), .B2(n433), .ZN(n162)
         );
  INVD1BWP12T U324 ( .I(cpu_data_in[2]), .ZN(n449) );
  INVD1BWP12T U325 ( .I(cpu_data_in[10]), .ZN(n441) );
  OAI22D0BWP12T U326 ( .A1(n173), .A2(n449), .B1(n172), .B2(n441), .ZN(n161)
         );
  AOI211D0BWP12T U327 ( .A1(tmp_value_2[2]), .A2(n176), .B(n162), .C(n161), 
        .ZN(n163) );
  INVD1BWP12T U328 ( .I(cpu_data_in[26]), .ZN(n425) );
  OAI22D0BWP12T U329 ( .A1(reset), .A2(n163), .B1(n425), .B2(n302), .ZN(N197)
         );
  TPND2D0BWP12T U330 ( .A1(n270), .A2(from_mem_data_out[14]), .ZN(n164) );
  OAI211D0BWP12T U331 ( .A1(n334), .A2(n248), .B(n169), .C(n164), .ZN(N104) );
  INVD1BWP12T U332 ( .I(cpu_data_in[17]), .ZN(n434) );
  OAI22D0BWP12T U333 ( .A1(n171), .A2(n339), .B1(n170), .B2(n434), .ZN(n166)
         );
  INVD1BWP12T U334 ( .I(cpu_data_in[1]), .ZN(n450) );
  INVD1BWP12T U335 ( .I(cpu_data_in[9]), .ZN(n442) );
  OAI22D0BWP12T U336 ( .A1(n173), .A2(n450), .B1(n172), .B2(n442), .ZN(n165)
         );
  AOI211D0BWP12T U337 ( .A1(tmp_value_2[1]), .A2(n176), .B(n166), .C(n165), 
        .ZN(n167) );
  INVD1BWP12T U338 ( .I(cpu_data_in[25]), .ZN(n426) );
  OAI22D0BWP12T U339 ( .A1(reset), .A2(n167), .B1(n426), .B2(n302), .ZN(N196)
         );
  CKND2D0BWP12T U340 ( .A1(from_mem_data_out[15]), .A2(n270), .ZN(n168) );
  OAI211D0BWP12T U341 ( .A1(n333), .A2(n248), .B(n169), .C(n168), .ZN(N105) );
  INVD1BWP12T U342 ( .I(cpu_data_in[16]), .ZN(n435) );
  OAI22D0BWP12T U343 ( .A1(n171), .A2(n341), .B1(n170), .B2(n435), .ZN(n175)
         );
  INVD1BWP12T U344 ( .I(cpu_data_in[0]), .ZN(n452) );
  INVD1BWP12T U345 ( .I(cpu_data_in[8]), .ZN(n443) );
  OAI22D0BWP12T U346 ( .A1(n173), .A2(n452), .B1(n172), .B2(n443), .ZN(n174)
         );
  AOI211D0BWP12T U347 ( .A1(tmp_value_2[0]), .A2(n176), .B(n175), .C(n174), 
        .ZN(n177) );
  INVD1BWP12T U348 ( .I(cpu_data_in[24]), .ZN(n427) );
  OAI22D0BWP12T U349 ( .A1(reset), .A2(n177), .B1(n427), .B2(n302), .ZN(N195)
         );
  INVD1BWP12T U350 ( .I(tmp_value_1[15]), .ZN(n264) );
  OAI22D0BWP12T U351 ( .A1(n202), .A2(n264), .B1(n201), .B2(n325), .ZN(n179)
         );
  OAI22D0BWP12T U352 ( .A1(n293), .A2(n436), .B1(n203), .B2(n343), .ZN(n178)
         );
  AOI211D0BWP12T U353 ( .A1(cpu_data_in[7]), .A2(n206), .B(n179), .C(n178), 
        .ZN(n180) );
  OAI22D0BWP12T U354 ( .A1(reset), .A2(n180), .B1(n428), .B2(n302), .ZN(N210)
         );
  OAI21D0BWP12T U355 ( .A1(reset), .A2(n182), .B(n181), .ZN(N73) );
  INVD1BWP12T U356 ( .I(tmp_value_1[14]), .ZN(n262) );
  OAI22D0BWP12T U357 ( .A1(n202), .A2(n262), .B1(n201), .B2(n326), .ZN(n184)
         );
  OAI22D0BWP12T U358 ( .A1(n293), .A2(n437), .B1(n203), .B2(n344), .ZN(n183)
         );
  AOI211D0BWP12T U359 ( .A1(cpu_data_in[6]), .A2(n206), .B(n184), .C(n183), 
        .ZN(n185) );
  OAI22D0BWP12T U360 ( .A1(reset), .A2(n185), .B1(n429), .B2(n302), .ZN(N209)
         );
  INVD1BWP12T U361 ( .I(tmp_value_1[13]), .ZN(n263) );
  OAI22D0BWP12T U362 ( .A1(n202), .A2(n263), .B1(n201), .B2(n327), .ZN(n187)
         );
  OAI22D0BWP12T U363 ( .A1(n293), .A2(n438), .B1(n203), .B2(n345), .ZN(n186)
         );
  AOI211D0BWP12T U364 ( .A1(cpu_data_in[5]), .A2(n206), .B(n187), .C(n186), 
        .ZN(n188) );
  OAI22D0BWP12T U365 ( .A1(reset), .A2(n188), .B1(n430), .B2(n302), .ZN(N208)
         );
  INVD1BWP12T U366 ( .I(tmp_value_1[12]), .ZN(n260) );
  OAI22D0BWP12T U367 ( .A1(n202), .A2(n260), .B1(n201), .B2(n328), .ZN(n190)
         );
  OAI22D0BWP12T U368 ( .A1(n293), .A2(n439), .B1(n203), .B2(n347), .ZN(n189)
         );
  AOI211D0BWP12T U369 ( .A1(cpu_data_in[4]), .A2(n206), .B(n190), .C(n189), 
        .ZN(n191) );
  OAI22D0BWP12T U370 ( .A1(reset), .A2(n191), .B1(n431), .B2(n302), .ZN(N207)
         );
  INVD1BWP12T U371 ( .I(tmp_value_1[11]), .ZN(n261) );
  OAI22D0BWP12T U372 ( .A1(n202), .A2(n261), .B1(n201), .B2(n329), .ZN(n193)
         );
  OAI22D0BWP12T U373 ( .A1(n293), .A2(n440), .B1(n203), .B2(n424), .ZN(n192)
         );
  AOI211D0BWP12T U374 ( .A1(cpu_data_in[3]), .A2(n206), .B(n193), .C(n192), 
        .ZN(n194) );
  OAI22D0BWP12T U375 ( .A1(reset), .A2(n194), .B1(n432), .B2(n302), .ZN(N206)
         );
  INVD1BWP12T U376 ( .I(tmp_value_1[10]), .ZN(n258) );
  OAI22D0BWP12T U377 ( .A1(n202), .A2(n258), .B1(n201), .B2(n330), .ZN(n196)
         );
  OAI22D0BWP12T U378 ( .A1(n293), .A2(n441), .B1(n203), .B2(n425), .ZN(n195)
         );
  AOI211D0BWP12T U379 ( .A1(cpu_data_in[2]), .A2(n206), .B(n196), .C(n195), 
        .ZN(n197) );
  OAI22D0BWP12T U380 ( .A1(reset), .A2(n197), .B1(n433), .B2(n302), .ZN(N205)
         );
  INVD1BWP12T U381 ( .I(tmp_value_1[9]), .ZN(n259) );
  OAI22D0BWP12T U382 ( .A1(n202), .A2(n259), .B1(n201), .B2(n331), .ZN(n199)
         );
  OAI22D0BWP12T U383 ( .A1(n293), .A2(n442), .B1(n203), .B2(n426), .ZN(n198)
         );
  AOI211D0BWP12T U384 ( .A1(cpu_data_in[1]), .A2(n206), .B(n199), .C(n198), 
        .ZN(n200) );
  OAI22D0BWP12T U385 ( .A1(reset), .A2(n200), .B1(n434), .B2(n302), .ZN(N204)
         );
  INVD1BWP12T U386 ( .I(tmp_value_1[8]), .ZN(n257) );
  OAI22D0BWP12T U387 ( .A1(n202), .A2(n257), .B1(n201), .B2(n332), .ZN(n205)
         );
  OAI22D0BWP12T U388 ( .A1(n293), .A2(n443), .B1(n203), .B2(n427), .ZN(n204)
         );
  AOI211D0BWP12T U389 ( .A1(cpu_data_in[0]), .A2(n206), .B(n205), .C(n204), 
        .ZN(n207) );
  OAI22D0BWP12T U390 ( .A1(reset), .A2(n207), .B1(n435), .B2(n302), .ZN(N203)
         );
  INVD1BWP12T U391 ( .I(n212), .ZN(n220) );
  AOI222D0BWP12T U392 ( .A1(n220), .A2(from_mem_data_out[12]), .B1(n219), .B2(
        tmp_value_1[4]), .C1(n218), .C2(from_mem_data_out[4]), .ZN(n208) );
  OAI22D0BWP12T U393 ( .A1(n208), .A2(reset), .B1(n260), .B2(n248), .ZN(N78)
         );
  AOI222D0BWP12T U394 ( .A1(n220), .A2(from_mem_data_out[10]), .B1(n219), .B2(
        tmp_value_1[2]), .C1(n218), .C2(from_mem_data_out[2]), .ZN(n209) );
  OAI22D0BWP12T U395 ( .A1(n209), .A2(reset), .B1(n258), .B2(n248), .ZN(N76)
         );
  AOI222D0BWP12T U396 ( .A1(n220), .A2(from_mem_data_out[9]), .B1(n219), .B2(
        tmp_value_1[1]), .C1(n218), .C2(from_mem_data_out[1]), .ZN(n210) );
  OAI22D0BWP12T U397 ( .A1(n210), .A2(reset), .B1(n259), .B2(n248), .ZN(N75)
         );
  AOI222D0BWP12T U398 ( .A1(n220), .A2(from_mem_data_out[8]), .B1(n219), .B2(
        tmp_value_1[0]), .C1(n218), .C2(from_mem_data_out[0]), .ZN(n211) );
  OAI22D0BWP12T U399 ( .A1(n211), .A2(reset), .B1(n257), .B2(n248), .ZN(N74)
         );
  TPNR2D0BWP12T U400 ( .A1(n212), .A2(n325), .ZN(n213) );
  AOI211D0BWP12T U401 ( .A1(n219), .A2(tmp_value_1[7]), .B(n214), .C(n213), 
        .ZN(n215) );
  OAI22D0BWP12T U402 ( .A1(n215), .A2(reset), .B1(n264), .B2(n248), .ZN(N81)
         );
  AOI222D0BWP12T U403 ( .A1(n220), .A2(from_mem_data_out[14]), .B1(n219), .B2(
        tmp_value_1[6]), .C1(n218), .C2(from_mem_data_out[6]), .ZN(n216) );
  OAI22D0BWP12T U404 ( .A1(n216), .A2(reset), .B1(n262), .B2(n248), .ZN(N80)
         );
  AOI222D0BWP12T U405 ( .A1(n220), .A2(from_mem_data_out[13]), .B1(n219), .B2(
        tmp_value_1[5]), .C1(n218), .C2(from_mem_data_out[5]), .ZN(n217) );
  OAI22D0BWP12T U406 ( .A1(n217), .A2(reset), .B1(n263), .B2(n248), .ZN(N79)
         );
  AOI222D0BWP12T U407 ( .A1(n220), .A2(from_mem_data_out[11]), .B1(n219), .B2(
        tmp_value_1[3]), .C1(n218), .C2(from_mem_data_out[3]), .ZN(n221) );
  OAI22D0BWP12T U408 ( .A1(n221), .A2(reset), .B1(n261), .B2(n248), .ZN(N77)
         );
  CKND0BWP12T U409 ( .I(n222), .ZN(n223) );
  AOI21D0BWP12T U410 ( .A1(n224), .A2(n223), .B(n255), .ZN(n225) );
  AOI211D0BWP12T U411 ( .A1(n227), .A2(n226), .B(n297), .C(n225), .ZN(n228) );
  TPAOI31D0BWP12T U412 ( .A1(n230), .A2(n229), .A3(n228), .B(reset), .ZN(N211)
         );
  HA1D0BWP12T U413 ( .A(cpu_address_in[1]), .B(n231), .CO(n117), .S(n232) );
  AO22D1BWP12T U414 ( .A1(n288), .A2(cpu_address_in[1]), .B1(n289), .B2(n232), 
        .Z(N183) );
  AOI22D0BWP12T U415 ( .A1(n271), .A2(tmp_value_1[3]), .B1(n270), .B2(
        tmp_value_2[11]), .ZN(n233) );
  OAI21D0BWP12T U416 ( .A1(n276), .A2(n337), .B(n233), .ZN(n234) );
  AO211D1BWP12T U417 ( .A1(n273), .A2(from_mem_data_out[11]), .B(n272), .C(
        n234), .Z(N85) );
  AOI22D0BWP12T U418 ( .A1(n271), .A2(tmp_value_1[1]), .B1(n270), .B2(
        tmp_value_2[9]), .ZN(n235) );
  OAI21D0BWP12T U419 ( .A1(n276), .A2(n339), .B(n235), .ZN(n236) );
  AO211D1BWP12T U420 ( .A1(from_mem_data_out[9]), .A2(n273), .B(n272), .C(n236), .Z(N83) );
  AOI22D0BWP12T U421 ( .A1(n271), .A2(tmp_value_1[2]), .B1(n270), .B2(
        tmp_value_2[10]), .ZN(n237) );
  OAI21D0BWP12T U422 ( .A1(n276), .A2(n338), .B(n237), .ZN(n238) );
  AO211D1BWP12T U423 ( .A1(n273), .A2(from_mem_data_out[10]), .B(n272), .C(
        n238), .Z(N84) );
  AOI22D0BWP12T U424 ( .A1(n271), .A2(tmp_value_1[0]), .B1(n270), .B2(
        tmp_value_2[8]), .ZN(n239) );
  OAI21D0BWP12T U425 ( .A1(n276), .A2(n341), .B(n239), .ZN(n240) );
  AO211D1BWP12T U426 ( .A1(n273), .A2(from_mem_data_out[8]), .B(n272), .C(n240), .Z(N82) );
  AO22D1BWP12T U427 ( .A1(n242), .A2(n289), .B1(cpu_address_in[3]), .B2(n288), 
        .Z(N185) );
  INVD1BWP12T U428 ( .I(n249), .ZN(n253) );
  AOI22D0BWP12T U429 ( .A1(n314), .A2(n315), .B1(n251), .B2(n250), .ZN(n252)
         );
  OAI211D1BWP12T U430 ( .A1(n255), .A2(n254), .B(n253), .C(n252), .ZN(n295) );
  OAI22D1BWP12T U431 ( .A1(n265), .A2(n257), .B1(n323), .B2(n332), .ZN(n416)
         );
  OAI22D1BWP12T U432 ( .A1(n265), .A2(n258), .B1(n323), .B2(n330), .ZN(n418)
         );
  OAI22D1BWP12T U433 ( .A1(n265), .A2(n259), .B1(n323), .B2(n331), .ZN(n417)
         );
  OAI22D1BWP12T U434 ( .A1(n265), .A2(n260), .B1(n323), .B2(n328), .ZN(n420)
         );
  OAI22D1BWP12T U435 ( .A1(n265), .A2(n261), .B1(n323), .B2(n329), .ZN(n419)
         );
  OAI22D1BWP12T U436 ( .A1(n265), .A2(n262), .B1(n323), .B2(n326), .ZN(n422)
         );
  OAI22D1BWP12T U437 ( .A1(n265), .A2(n263), .B1(n323), .B2(n327), .ZN(n421)
         );
  OAI22D1BWP12T U438 ( .A1(n265), .A2(n264), .B1(n323), .B2(n325), .ZN(n423)
         );
  AOI22D0BWP12T U439 ( .A1(n271), .A2(tmp_value_1[6]), .B1(n270), .B2(
        tmp_value_2[14]), .ZN(n267) );
  AOI21D0BWP12T U440 ( .A1(from_mem_data_out[14]), .A2(n273), .B(n272), .ZN(
        n266) );
  OAI211D1BWP12T U441 ( .A1(n276), .A2(n334), .B(n267), .C(n266), .ZN(N88) );
  AOI22D0BWP12T U442 ( .A1(n271), .A2(tmp_value_1[4]), .B1(n270), .B2(
        tmp_value_2[12]), .ZN(n269) );
  AOI21D0BWP12T U443 ( .A1(from_mem_data_out[12]), .A2(n273), .B(n272), .ZN(
        n268) );
  OAI211D1BWP12T U444 ( .A1(n276), .A2(n336), .B(n269), .C(n268), .ZN(N86) );
  AOI22D0BWP12T U445 ( .A1(n271), .A2(tmp_value_1[5]), .B1(n270), .B2(
        tmp_value_2[13]), .ZN(n275) );
  AOI21D0BWP12T U446 ( .A1(from_mem_data_out[13]), .A2(n273), .B(n272), .ZN(
        n274) );
  OAI211D1BWP12T U447 ( .A1(n276), .A2(n335), .B(n275), .C(n274), .ZN(N87) );
  AO22D1BWP12T U448 ( .A1(n278), .A2(n289), .B1(cpu_address_in[4]), .B2(n288), 
        .Z(N186) );
  AO22D1BWP12T U449 ( .A1(n280), .A2(n289), .B1(cpu_address_in[5]), .B2(n288), 
        .Z(N187) );
  AO22D1BWP12T U450 ( .A1(n282), .A2(n289), .B1(cpu_address_in[6]), .B2(n288), 
        .Z(N188) );
  AO22D1BWP12T U451 ( .A1(n284), .A2(n289), .B1(cpu_address_in[7]), .B2(n288), 
        .Z(N189) );
  AO22D1BWP12T U452 ( .A1(n286), .A2(n289), .B1(cpu_address_in[8]), .B2(n288), 
        .Z(N190) );
  AO22D1BWP12T U453 ( .A1(n290), .A2(n289), .B1(cpu_address_in[9]), .B2(n288), 
        .Z(N191) );
  CKND0BWP12T U454 ( .I(n291), .ZN(n306) );
  OAI21D0BWP12T U455 ( .A1(n292), .A2(n306), .B(n309), .ZN(n300) );
  INVD0BWP12T U456 ( .I(n293), .ZN(n296) );
  OR4D0BWP12T U457 ( .A1(n297), .A2(n296), .A3(n295), .A4(n294), .Z(n298) );
  AOI211D1BWP12T U458 ( .A1(n301), .A2(n300), .B(n299), .C(n298), .ZN(n304) );
  OAI211D1BWP12T U459 ( .A1(reset), .A2(n304), .B(n303), .C(n302), .ZN(N66) );
  MOAI22D0BWP12T U460 ( .A1(n323), .A2(n333), .B1(tmp_value_1[7]), .B2(n322), 
        .ZN(n415) );
  MOAI22D0BWP12T U461 ( .A1(n323), .A2(n334), .B1(tmp_value_1[6]), .B2(n322), 
        .ZN(n414) );
  MOAI22D0BWP12T U462 ( .A1(n323), .A2(n335), .B1(tmp_value_1[5]), .B2(n322), 
        .ZN(n413) );
  MOAI22D0BWP12T U463 ( .A1(n323), .A2(n336), .B1(tmp_value_1[4]), .B2(n322), 
        .ZN(n412) );
  MOAI22D0BWP12T U464 ( .A1(n323), .A2(n337), .B1(tmp_value_1[3]), .B2(n322), 
        .ZN(n411) );
  MOAI22D0BWP12T U465 ( .A1(n323), .A2(n338), .B1(tmp_value_1[2]), .B2(n322), 
        .ZN(n410) );
  MOAI22D0BWP12T U466 ( .A1(n323), .A2(n339), .B1(tmp_value_1[1]), .B2(n322), 
        .ZN(n409) );
  MOAI22D0BWP12T U467 ( .A1(n323), .A2(n341), .B1(tmp_value_1[0]), .B2(n322), 
        .ZN(n408) );
  MOAI22D0BWP12T U468 ( .A1(n325), .A2(n342), .B1(tmp_value_2[15]), .B2(n340), 
        .ZN(n407) );
  MOAI22D0BWP12T U469 ( .A1(n342), .A2(n326), .B1(tmp_value_2[14]), .B2(n340), 
        .ZN(n406) );
  MOAI22D0BWP12T U470 ( .A1(n342), .A2(n327), .B1(tmp_value_2[13]), .B2(n340), 
        .ZN(n405) );
  MOAI22D0BWP12T U471 ( .A1(n342), .A2(n328), .B1(tmp_value_2[12]), .B2(n340), 
        .ZN(n404) );
  MOAI22D0BWP12T U472 ( .A1(n342), .A2(n329), .B1(tmp_value_2[11]), .B2(n340), 
        .ZN(n403) );
  MOAI22D0BWP12T U473 ( .A1(n342), .A2(n330), .B1(tmp_value_2[10]), .B2(n340), 
        .ZN(n402) );
  MOAI22D0BWP12T U474 ( .A1(n342), .A2(n331), .B1(tmp_value_2[9]), .B2(n340), 
        .ZN(n401) );
  MOAI22D0BWP12T U475 ( .A1(n342), .A2(n332), .B1(tmp_value_2[8]), .B2(n340), 
        .ZN(n400) );
  MOAI22D0BWP12T U476 ( .A1(n342), .A2(n333), .B1(tmp_value_2[7]), .B2(n340), 
        .ZN(n399) );
  MOAI22D0BWP12T U477 ( .A1(n342), .A2(n334), .B1(tmp_value_2[6]), .B2(n340), 
        .ZN(n398) );
  MOAI22D0BWP12T U478 ( .A1(n342), .A2(n335), .B1(tmp_value_2[5]), .B2(n340), 
        .ZN(n397) );
  MOAI22D0BWP12T U479 ( .A1(n342), .A2(n336), .B1(tmp_value_2[4]), .B2(n340), 
        .ZN(n396) );
  MOAI22D0BWP12T U480 ( .A1(n342), .A2(n337), .B1(tmp_value_2[3]), .B2(n340), 
        .ZN(n395) );
  MOAI22D0BWP12T U481 ( .A1(n342), .A2(n338), .B1(tmp_value_2[2]), .B2(n340), 
        .ZN(n394) );
  MOAI22D0BWP12T U482 ( .A1(n342), .A2(n339), .B1(tmp_value_2[1]), .B2(n340), 
        .ZN(n393) );
  MOAI22D0BWP12T U483 ( .A1(n342), .A2(n341), .B1(tmp_value_2[0]), .B2(n340), 
        .ZN(n392) );
  MOAI22D0BWP12T U484 ( .A1(n453), .A2(n343), .B1(n451), .B2(
        interface_cpu_data_in[31]), .ZN(n391) );
  MOAI22D0BWP12T U485 ( .A1(n453), .A2(n344), .B1(n451), .B2(
        interface_cpu_data_in[30]), .ZN(n390) );
  MOAI22D0BWP12T U486 ( .A1(n453), .A2(n345), .B1(n451), .B2(
        interface_cpu_data_in[29]), .ZN(n389) );
  MOAI22D0BWP12T U487 ( .A1(n453), .A2(n347), .B1(n451), .B2(
        interface_cpu_data_in[28]), .ZN(n388) );
  MOAI22D0BWP12T U488 ( .A1(n453), .A2(n424), .B1(n451), .B2(
        interface_cpu_data_in[27]), .ZN(n387) );
  MOAI22D0BWP12T U489 ( .A1(n453), .A2(n425), .B1(n451), .B2(
        interface_cpu_data_in[26]), .ZN(n386) );
  MOAI22D0BWP12T U490 ( .A1(n453), .A2(n426), .B1(n451), .B2(
        interface_cpu_data_in[25]), .ZN(n385) );
  MOAI22D0BWP12T U491 ( .A1(n453), .A2(n427), .B1(n451), .B2(
        interface_cpu_data_in[24]), .ZN(n384) );
  MOAI22D0BWP12T U492 ( .A1(n453), .A2(n428), .B1(n451), .B2(
        interface_cpu_data_in[23]), .ZN(n383) );
  MOAI22D0BWP12T U493 ( .A1(n453), .A2(n429), .B1(n451), .B2(
        interface_cpu_data_in[22]), .ZN(n382) );
  MOAI22D0BWP12T U494 ( .A1(n453), .A2(n430), .B1(n451), .B2(
        interface_cpu_data_in[21]), .ZN(n381) );
  MOAI22D0BWP12T U495 ( .A1(n453), .A2(n432), .B1(n451), .B2(
        interface_cpu_data_in[19]), .ZN(n379) );
  MOAI22D0BWP12T U496 ( .A1(n453), .A2(n433), .B1(n451), .B2(
        interface_cpu_data_in[18]), .ZN(n378) );
  MOAI22D0BWP12T U497 ( .A1(n453), .A2(n434), .B1(n451), .B2(
        interface_cpu_data_in[17]), .ZN(n377) );
  MOAI22D0BWP12T U498 ( .A1(n453), .A2(n435), .B1(n451), .B2(
        interface_cpu_data_in[16]), .ZN(n376) );
  MOAI22D0BWP12T U499 ( .A1(n453), .A2(n436), .B1(n451), .B2(
        interface_cpu_data_in[15]), .ZN(n375) );
  MOAI22D0BWP12T U500 ( .A1(n453), .A2(n437), .B1(n451), .B2(
        interface_cpu_data_in[14]), .ZN(n374) );
  MOAI22D0BWP12T U501 ( .A1(n453), .A2(n438), .B1(n451), .B2(
        interface_cpu_data_in[13]), .ZN(n373) );
  MOAI22D0BWP12T U502 ( .A1(n453), .A2(n439), .B1(n451), .B2(
        interface_cpu_data_in[12]), .ZN(n372) );
  MOAI22D0BWP12T U503 ( .A1(n453), .A2(n440), .B1(n451), .B2(
        interface_cpu_data_in[11]), .ZN(n371) );
  MOAI22D0BWP12T U504 ( .A1(n453), .A2(n441), .B1(n451), .B2(
        interface_cpu_data_in[10]), .ZN(n370) );
  MOAI22D0BWP12T U505 ( .A1(n453), .A2(n442), .B1(n451), .B2(
        interface_cpu_data_in[9]), .ZN(n369) );
  MOAI22D0BWP12T U506 ( .A1(n453), .A2(n443), .B1(n451), .B2(
        interface_cpu_data_in[8]), .ZN(n368) );
  MOAI22D0BWP12T U507 ( .A1(n453), .A2(n444), .B1(n451), .B2(
        interface_cpu_data_in[7]), .ZN(n367) );
  MOAI22D0BWP12T U508 ( .A1(n453), .A2(n445), .B1(n451), .B2(
        interface_cpu_data_in[6]), .ZN(n366) );
  MOAI22D0BWP12T U509 ( .A1(n453), .A2(n446), .B1(n451), .B2(
        interface_cpu_data_in[5]), .ZN(n365) );
  MOAI22D0BWP12T U510 ( .A1(n453), .A2(n447), .B1(n451), .B2(
        interface_cpu_data_in[4]), .ZN(n364) );
  MOAI22D0BWP12T U511 ( .A1(n453), .A2(n448), .B1(n451), .B2(
        interface_cpu_data_in[3]), .ZN(n363) );
  MOAI22D0BWP12T U512 ( .A1(n453), .A2(n449), .B1(n451), .B2(
        interface_cpu_data_in[2]), .ZN(n362) );
  MOAI22D0BWP12T U513 ( .A1(n453), .A2(n450), .B1(n451), .B2(
        interface_cpu_data_in[1]), .ZN(n361) );
  MOAI22D0BWP12T U514 ( .A1(n453), .A2(n452), .B1(n451), .B2(
        interface_cpu_data_in[0]), .ZN(n360) );
endmodule


module cpu ( clock, reset, MEM_MEMCTRL_from_mem_data, 
        MEMCTRL_MEM_to_mem_read_enable, MEMCTRL_MEM_to_mem_write_enable, 
        MEMCTRL_MEM_to_mem_mem_enable, MEMCTRL_MEM_to_mem_address, 
        MEMCTRL_MEM_to_mem_data );
  input [15:0] MEM_MEMCTRL_from_mem_data;
  output [11:0] MEMCTRL_MEM_to_mem_address;
  output [15:0] MEMCTRL_MEM_to_mem_data;
  input clock, reset;
  output MEMCTRL_MEM_to_mem_read_enable, MEMCTRL_MEM_to_mem_write_enable,
         MEMCTRL_MEM_to_mem_mem_enable;
  wire   new_n, ALU_OUT_n, RF_OUT_n, DEC_CPSR_update_flag_c, new_c, ALU_OUT_c,
         RF_OUT_c, DEC_CPSR_update_flag_z, new_z, ALU_OUT_z, RF_OUT_z,
         DEC_CPSR_update_flag_v, new_v, ALU_OUT_v, RF_OUT_v,
         MEMCTRL_write_finished, MEMCTRL_read_finished,
         DEC_MISC_OUT_pc_mask_bit, DEC_RF_alu_write_to_reg_enable,
         DEC_RF_memory_write_to_reg_enable,
         DEC_MISC_OUT_memory_address_source_is_reg,
         DEC_MEMCTRL_memorycontroller_sign_extend,
         DEC_MEMCTRL_memory_load_request, DEC_MEMCTRL_memory_store_request,
         DEC_IF_stall_to_instructionfetch, ALU_IN_c, MEMCTRL_load_in,
         irdecode_inst1_N915, irdecode_inst1_N914, irdecode_inst1_N910,
         irdecode_inst1_N909, irdecode_inst1_N710, irdecode_inst1_N709,
         irdecode_inst1_N708, irdecode_inst1_N707, irdecode_inst1_N706,
         irdecode_inst1_N705, irdecode_inst1_N704, irdecode_inst1_N549,
         irdecode_inst1_N548, irdecode_inst1_N547, irdecode_inst1_N546,
         irdecode_inst1_N545, irdecode_inst1_N544, irdecode_inst1_N543,
         irdecode_inst1_N542, irdecode_inst1_split_instruction,
         irdecode_inst1_next_step_0_, irdecode_inst1_next_step_1_,
         irdecode_inst1_next_step_2_, irdecode_inst1_next_step_3_,
         irdecode_inst1_next_step_4_, irdecode_inst1_next_step_5_,
         irdecode_inst1_next_step_6_, irdecode_inst1_next_step_7_,
         irdecode_inst1_itstate_0_, irdecode_inst1_itstate_1_,
         irdecode_inst1_itstate_2_, irdecode_inst1_itstate_3_,
         irdecode_inst1_itstate_4_, irdecode_inst1_itstate_5_,
         irdecode_inst1_itstate_6_, irdecode_inst1_itstate_7_,
         irdecode_inst1_next_alu_write_to_reg_enable,
         irdecode_inst1_next_update_flag_v, irdecode_inst1_next_update_flag_c,
         irdecode_inst1_next_update_flag_n, Instruction_Fetch_v2_inst1_N98,
         Instruction_Fetch_v2_inst1_N97, Instruction_Fetch_v2_inst1_N96,
         Instruction_Fetch_v2_inst1_N95, Instruction_Fetch_v2_inst1_N93,
         Instruction_Fetch_v2_inst1_N92, Instruction_Fetch_v2_inst1_N91,
         Instruction_Fetch_v2_inst1_N90, Instruction_Fetch_v2_inst1_N89,
         Instruction_Fetch_v2_inst1_N88, Instruction_Fetch_v2_inst1_N87,
         Instruction_Fetch_v2_inst1_N86, Instruction_Fetch_v2_inst1_N85,
         Instruction_Fetch_v2_inst1_N84, Instruction_Fetch_v2_inst1_N83,
         Instruction_Fetch_v2_inst1_N80, Instruction_Fetch_v2_inst1_N79,
         Instruction_Fetch_v2_inst1_first_instruction_fetched,
         Instruction_Fetch_v2_inst1_fetched_instruction_reg_0_,
         Instruction_Fetch_v2_inst1_fetched_instruction_reg_1_,
         Instruction_Fetch_v2_inst1_fetched_instruction_reg_2_,
         Instruction_Fetch_v2_inst1_fetched_instruction_reg_3_,
         Instruction_Fetch_v2_inst1_fetched_instruction_reg_4_,
         Instruction_Fetch_v2_inst1_fetched_instruction_reg_5_,
         Instruction_Fetch_v2_inst1_fetched_instruction_reg_6_,
         Instruction_Fetch_v2_inst1_fetched_instruction_reg_7_,
         Instruction_Fetch_v2_inst1_fetched_instruction_reg_8_,
         Instruction_Fetch_v2_inst1_fetched_instruction_reg_9_,
         Instruction_Fetch_v2_inst1_fetched_instruction_reg_10_,
         Instruction_Fetch_v2_inst1_fetched_instruction_reg_11_,
         Instruction_Fetch_v2_inst1_fetched_instruction_reg_12_,
         Instruction_Fetch_v2_inst1_fetched_instruction_reg_13_,
         Instruction_Fetch_v2_inst1_fetched_instruction_reg_14_,
         Instruction_Fetch_v2_inst1_fetched_instruction_reg_15_,
         Instruction_Fetch_v2_inst1_currentState_0_,
         Instruction_Fetch_v2_inst1_currentState_1_,
         Instruction_Fetch_v2_inst1_current_pc_modified_0_, n770, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51;
  wire   [7:0] IF_DEC_instruction;
  wire   [4:0] DEC_RF_operand_a;
  wire   [4:0] DEC_RF_operand_b;
  wire   [15:0] DEC_RF_offset_a;
  wire   [31:0] DEC_RF_offset_b;
  wire   [4:0] DEC_ALU_alu_opcode;
  wire   [2:0] DEC_MISC_OUT_operator_b_modification;
  wire   [4:0] DEC_RF_alu_write_to_reg;
  wire   [4:0] DEC_RF_memory_write_to_reg;
  wire   [4:0] DEC_RF_memory_store_data_reg;
  wire   [4:0] DEC_RF_memory_store_address_reg;
  wire   [1:0] DEC_MEMCTRL_load_store_width;
  wire   [31:0] ALU_MISC_OUT_result;
  wire   [31:0] MEMCTRL_RF_IF_data_in;
  wire   [31:0] IF_RF_incremented_pc_out;
  wire   [31:0] RF_ALU_operand_a;
  wire   [31:0] RF_ALU_operand_b;
  wire   [31:0] RF_MEMCTRL_data_reg;
  wire   [12:0] RF_MEMCTRL_address_reg;
  wire   [31:1] RF_pc_out;
  wire   [31:0] RF_ALU_operand_b_modified;
  wire   [1:0] MEMCTRL_IN_load_store_width;
  wire   [12:0] MEMCTRL_IN_address;
  wire   [7:0] irdecode_inst1_step;

  register_file_v2 register_file_v2_inst1 ( .readA_sel({DEC_RF_operand_a[4], 
        n1770, DEC_RF_operand_a[2:0]}), .readB_sel({DEC_RF_operand_b[4], n994, 
        DEC_RF_operand_b[2], n999, DEC_RF_operand_b[0]}), .readC_sel(
        DEC_RF_memory_store_data_reg), .readD_sel(
        DEC_RF_memory_store_address_reg), .write1_sel(DEC_RF_alu_write_to_reg), 
        .write2_sel(DEC_RF_memory_write_to_reg), .write1_en(
        DEC_RF_alu_write_to_reg_enable), .write2_en(
        DEC_RF_memory_write_to_reg_enable), .write1_in(ALU_MISC_OUT_result), 
        .write2_in(MEMCTRL_RF_IF_data_in), .immediate1_in({n877, n877, n877, 
        n877, n877, n877, n877, n877, n877, n877, n877, n877, n877, n877, n877, 
        n877, DEC_RF_offset_a}), .immediate2_in(DEC_RF_offset_b), .next_pc_in(
        {IF_RF_incremented_pc_out[31:30], n1779, IF_RF_incremented_pc_out[28], 
        n1775, IF_RF_incremented_pc_out[26], n1778, 
        IF_RF_incremented_pc_out[24], n1774, IF_RF_incremented_pc_out[22], 
        n1773, IF_RF_incremented_pc_out[20], n1777, 
        IF_RF_incremented_pc_out[18], n1776, IF_RF_incremented_pc_out[16:0]}), 
        .next_cpsr_in({new_n, new_c, new_z, new_v}), .next_sp_in({n877, n877, 
        n877, n877, n877, n877, n877, n877, n877, n877, n877, n877, n877, n877, 
        n877, n877, n877, n877, n877, n877, n877, n877, n877, n877, n877, n877, 
        n877, n877, n877, n877, n877, n877}), .clk(clock), .reset(reset), 
        .regA_out(RF_ALU_operand_a), .regB_out(RF_ALU_operand_b), .regC_out(
        RF_MEMCTRL_data_reg), .regD_out({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        RF_MEMCTRL_address_reg}), .pc_out({RF_pc_out, 
        Instruction_Fetch_v2_inst1_current_pc_modified_0_}), .cpsr_out({
        RF_OUT_n, RF_OUT_c, RF_OUT_z, RF_OUT_v}), .sp_out({
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51}), .next_pc_en_BAR(
        n1780) );
  ALU_VARIABLE ALU_VARIABLE_inst1 ( .a({RF_ALU_operand_a[31:28], n1784, 
        RF_ALU_operand_a[26:2], n1772, RF_ALU_operand_a[0]}), .b(
        RF_ALU_operand_b_modified), .op(DEC_ALU_alu_opcode[3:0]), .c_in(
        ALU_IN_c), .result(ALU_MISC_OUT_result), .c_out(ALU_OUT_c), .z(
        ALU_OUT_z), .n(ALU_OUT_n), .v(ALU_OUT_v) );
  memory_interface_simple memory_interface_simple_inst1 ( .clock(clock), 
        .reset(reset), .interface_cpu_sign_extend(
        DEC_MEMCTRL_memorycontroller_sign_extend), .interface_cpu_word_type(
        MEMCTRL_IN_load_store_width), .interface_cpu_load_request(
        MEMCTRL_load_in), .interface_cpu_address_in(MEMCTRL_IN_address), 
        .interface_cpu_data_in(RF_MEMCTRL_data_reg), .from_mem_data_out(
        MEM_MEMCTRL_from_mem_data), .interface_cpu_read_finished(
        MEMCTRL_read_finished), .interface_cpu_write_finished(
        MEMCTRL_write_finished), .interface_cpu_data_out(MEMCTRL_RF_IF_data_in), .to_mem_address(MEMCTRL_MEM_to_mem_address), .to_mem_data_in(
        MEMCTRL_MEM_to_mem_data), .to_mem_read_enable(
        MEMCTRL_MEM_to_mem_read_enable), .to_mem_write_enable(
        MEMCTRL_MEM_to_mem_write_enable), .interface_cpu_store_request_BAR(
        n1554) );
  CKAN2D2BWP12T irdecode_inst1_C5480 ( .A1(irdecode_inst1_next_step_7_), .A2(
        IF_DEC_instruction[7]), .Z(irdecode_inst1_N542) );
  CKAN2D2BWP12T irdecode_inst1_C5481 ( .A1(irdecode_inst1_next_step_6_), .A2(
        IF_DEC_instruction[6]), .Z(irdecode_inst1_N543) );
  CKAN2D2BWP12T irdecode_inst1_C5482 ( .A1(irdecode_inst1_next_step_5_), .A2(
        IF_DEC_instruction[5]), .Z(irdecode_inst1_N544) );
  CKAN2D2BWP12T irdecode_inst1_C5483 ( .A1(irdecode_inst1_next_step_4_), .A2(
        IF_DEC_instruction[4]), .Z(irdecode_inst1_N545) );
  CKAN2D2BWP12T irdecode_inst1_C5484 ( .A1(irdecode_inst1_next_step_3_), .A2(
        IF_DEC_instruction[3]), .Z(irdecode_inst1_N546) );
  CKAN2D2BWP12T irdecode_inst1_C5485 ( .A1(irdecode_inst1_next_step_2_), .A2(
        IF_DEC_instruction[2]), .Z(irdecode_inst1_N547) );
  CKAN2D2BWP12T irdecode_inst1_C5486 ( .A1(irdecode_inst1_next_step_1_), .A2(
        IF_DEC_instruction[1]), .Z(irdecode_inst1_N548) );
  CKAN2D2BWP12T irdecode_inst1_C5487 ( .A1(irdecode_inst1_next_step_0_), .A2(
        IF_DEC_instruction[0]), .Z(irdecode_inst1_N549) );
  CKAN2D2BWP12T irdecode_inst1_C5567 ( .A1(irdecode_inst1_next_step_6_), .A2(
        IF_DEC_instruction[6]), .Z(irdecode_inst1_N704) );
  CKAN2D2BWP12T irdecode_inst1_C5568 ( .A1(irdecode_inst1_next_step_5_), .A2(
        IF_DEC_instruction[5]), .Z(irdecode_inst1_N705) );
  CKAN2D2BWP12T irdecode_inst1_C5569 ( .A1(irdecode_inst1_next_step_4_), .A2(
        IF_DEC_instruction[4]), .Z(irdecode_inst1_N706) );
  CKAN2D2BWP12T irdecode_inst1_C5570 ( .A1(irdecode_inst1_next_step_3_), .A2(
        IF_DEC_instruction[3]), .Z(irdecode_inst1_N707) );
  CKAN2D2BWP12T irdecode_inst1_C5571 ( .A1(irdecode_inst1_next_step_2_), .A2(
        IF_DEC_instruction[2]), .Z(irdecode_inst1_N708) );
  CKAN2D2BWP12T irdecode_inst1_C5572 ( .A1(irdecode_inst1_next_step_1_), .A2(
        IF_DEC_instruction[1]), .Z(irdecode_inst1_N709) );
  CKAN2D2BWP12T irdecode_inst1_C5573 ( .A1(irdecode_inst1_next_step_0_), .A2(
        IF_DEC_instruction[0]), .Z(irdecode_inst1_N710) );
  CKAN2D2BWP12T irdecode_inst1_C2473 ( .A1(irdecode_inst1_next_step_1_), .A2(
        irdecode_inst1_next_step_0_), .Z(irdecode_inst1_N909) );
  CKAN2D2BWP12T irdecode_inst1_C2479 ( .A1(irdecode_inst1_N910), .A2(n1785), 
        .Z(irdecode_inst1_N914) );
  OR2XD4BWP12T irdecode_inst1_C2481 ( .A1(irdecode_inst1_next_step_1_), .A2(
        n1785), .Z(irdecode_inst1_N915) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_fetched_instruction_reg_reg_0_ ( .D(
        Instruction_Fetch_v2_inst1_N83), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_0_) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_fetched_instruction_reg_reg_1_ ( .D(
        Instruction_Fetch_v2_inst1_N84), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_1_) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_fetched_instruction_reg_reg_2_ ( .D(
        Instruction_Fetch_v2_inst1_N85), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_2_) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_fetched_instruction_reg_reg_3_ ( .D(
        Instruction_Fetch_v2_inst1_N86), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_3_) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_fetched_instruction_reg_reg_4_ ( .D(
        Instruction_Fetch_v2_inst1_N87), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_4_) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_fetched_instruction_reg_reg_5_ ( .D(
        Instruction_Fetch_v2_inst1_N88), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_5_) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_fetched_instruction_reg_reg_6_ ( .D(
        Instruction_Fetch_v2_inst1_N89), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_6_) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_fetched_instruction_reg_reg_7_ ( .D(
        Instruction_Fetch_v2_inst1_N90), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_7_) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_fetched_instruction_reg_reg_8_ ( .D(
        Instruction_Fetch_v2_inst1_N91), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_8_) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_fetched_instruction_reg_reg_9_ ( .D(
        Instruction_Fetch_v2_inst1_N92), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_9_) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_fetched_instruction_reg_reg_10_ ( .D(
        Instruction_Fetch_v2_inst1_N93), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_10_) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_fetched_instruction_reg_reg_12_ ( .D(
        Instruction_Fetch_v2_inst1_N95), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_12_) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_fetched_instruction_reg_reg_13_ ( .D(
        Instruction_Fetch_v2_inst1_N96), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_13_) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_fetched_instruction_reg_reg_14_ ( .D(
        Instruction_Fetch_v2_inst1_N97), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_14_) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_fetched_instruction_reg_reg_15_ ( .D(
        Instruction_Fetch_v2_inst1_N98), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_15_) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_first_instruction_fetched_reg ( .D(
        n874), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_first_instruction_fetched) );
  DFQD1BWP12T irdecode_inst1_stall_to_instructionfetch_reg ( .D(n841), .CP(
        clock), .Q(DEC_IF_stall_to_instructionfetch) );
  DFQD1BWP12T Instruction_Fetch_v2_inst1_currentState_reg_0_ ( .D(
        Instruction_Fetch_v2_inst1_N79), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_currentState_0_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_0_ ( .D(n840), .CP(clock), .Q(
        irdecode_inst1_itstate_0_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_1_ ( .D(n839), .CP(clock), .Q(
        irdecode_inst1_itstate_1_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_2_ ( .D(n838), .CP(clock), .Q(
        irdecode_inst1_itstate_2_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_3_ ( .D(n837), .CP(clock), .Q(
        irdecode_inst1_itstate_3_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_4_ ( .D(n836), .CP(clock), .Q(
        irdecode_inst1_itstate_4_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_5_ ( .D(n835), .CP(clock), .Q(
        irdecode_inst1_itstate_5_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_6_ ( .D(n834), .CP(clock), .Q(
        irdecode_inst1_itstate_6_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_7_ ( .D(n833), .CP(clock), .Q(
        irdecode_inst1_itstate_7_) );
  DFQD1BWP12T irdecode_inst1_offset_a_reg_0_ ( .D(n796), .CP(clock), .Q(
        DEC_RF_offset_a[0]) );
  DFQD1BWP12T irdecode_inst1_offset_a_reg_1_ ( .D(n795), .CP(clock), .Q(
        DEC_RF_offset_a[1]) );
  DFQD1BWP12T irdecode_inst1_offset_a_reg_2_ ( .D(n794), .CP(clock), .Q(
        DEC_RF_offset_a[2]) );
  DFQD1BWP12T irdecode_inst1_offset_a_reg_3_ ( .D(n793), .CP(clock), .Q(
        DEC_RF_offset_a[3]) );
  DFQD1BWP12T irdecode_inst1_offset_a_reg_4_ ( .D(n792), .CP(clock), .Q(
        DEC_RF_offset_a[4]) );
  DFQD1BWP12T irdecode_inst1_offset_a_reg_5_ ( .D(n791), .CP(clock), .Q(
        DEC_RF_offset_a[5]) );
  DFQD1BWP12T irdecode_inst1_offset_a_reg_6_ ( .D(n790), .CP(clock), .Q(
        DEC_RF_offset_a[6]) );
  DFQD1BWP12T irdecode_inst1_offset_a_reg_7_ ( .D(n789), .CP(clock), .Q(
        DEC_RF_offset_a[7]) );
  DFQD1BWP12T irdecode_inst1_offset_a_reg_8_ ( .D(n788), .CP(clock), .Q(
        DEC_RF_offset_a[8]) );
  DFQD1BWP12T irdecode_inst1_offset_a_reg_9_ ( .D(n787), .CP(clock), .Q(
        DEC_RF_offset_a[9]) );
  DFQD1BWP12T irdecode_inst1_offset_a_reg_10_ ( .D(n786), .CP(clock), .Q(
        DEC_RF_offset_a[10]) );
  DFQD1BWP12T irdecode_inst1_offset_a_reg_11_ ( .D(n785), .CP(clock), .Q(
        DEC_RF_offset_a[11]) );
  DFQD1BWP12T irdecode_inst1_offset_a_reg_12_ ( .D(n784), .CP(clock), .Q(
        DEC_RF_offset_a[12]) );
  DFQD1BWP12T irdecode_inst1_offset_a_reg_13_ ( .D(n783), .CP(clock), .Q(
        DEC_RF_offset_a[13]) );
  DFQD1BWP12T irdecode_inst1_offset_a_reg_14_ ( .D(n782), .CP(clock), .Q(
        DEC_RF_offset_a[14]) );
  DFQD1BWP12T irdecode_inst1_offset_a_reg_15_ ( .D(n781), .CP(clock), .Q(
        DEC_RF_offset_a[15]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_31_ ( .D(n875), .CP(clock), .Q(
        DEC_RF_offset_b[31]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_30_ ( .D(n873), .CP(clock), .Q(
        DEC_RF_offset_b[30]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_29_ ( .D(n872), .CP(clock), .Q(
        DEC_RF_offset_b[29]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_28_ ( .D(n871), .CP(clock), .Q(
        DEC_RF_offset_b[28]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_27_ ( .D(n870), .CP(clock), .Q(
        DEC_RF_offset_b[27]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_26_ ( .D(n869), .CP(clock), .Q(
        DEC_RF_offset_b[26]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_25_ ( .D(n868), .CP(clock), .Q(
        DEC_RF_offset_b[25]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_24_ ( .D(n867), .CP(clock), .Q(
        DEC_RF_offset_b[24]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_23_ ( .D(n866), .CP(clock), .Q(
        DEC_RF_offset_b[23]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_22_ ( .D(n865), .CP(clock), .Q(
        DEC_RF_offset_b[22]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_21_ ( .D(n864), .CP(clock), .Q(
        DEC_RF_offset_b[21]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_20_ ( .D(n863), .CP(clock), .Q(
        DEC_RF_offset_b[20]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_19_ ( .D(n862), .CP(clock), .Q(
        DEC_RF_offset_b[19]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_18_ ( .D(n861), .CP(clock), .Q(
        DEC_RF_offset_b[18]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_17_ ( .D(n860), .CP(clock), .Q(
        DEC_RF_offset_b[17]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_16_ ( .D(n859), .CP(clock), .Q(
        DEC_RF_offset_b[16]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_15_ ( .D(n858), .CP(clock), .Q(
        DEC_RF_offset_b[15]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_14_ ( .D(n857), .CP(clock), .Q(
        DEC_RF_offset_b[14]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_13_ ( .D(n856), .CP(clock), .Q(
        DEC_RF_offset_b[13]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_12_ ( .D(n855), .CP(clock), .Q(
        DEC_RF_offset_b[12]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_enable_reg ( .D(
        irdecode_inst1_next_alu_write_to_reg_enable), .CP(clock), .Q(
        DEC_RF_alu_write_to_reg_enable) );
  DFQD1BWP12T irdecode_inst1_update_flag_c_reg ( .D(
        irdecode_inst1_next_update_flag_c), .CP(clock), .Q(
        DEC_CPSR_update_flag_c) );
  DFQD1BWP12T irdecode_inst1_update_flag_z_reg ( .D(
        irdecode_inst1_next_update_flag_n), .CP(clock), .Q(
        DEC_CPSR_update_flag_z) );
  DFQD1BWP12T irdecode_inst1_update_flag_v_reg ( .D(
        irdecode_inst1_next_update_flag_v), .CP(clock), .Q(
        DEC_CPSR_update_flag_v) );
  DFQD1BWP12T irdecode_inst1_memorycontroller_sign_extend_reg ( .D(n825), .CP(
        clock), .Q(DEC_MEMCTRL_memorycontroller_sign_extend) );
  DFQD1BWP12T irdecode_inst1_load_store_width_reg_0_ ( .D(n824), .CP(clock), 
        .Q(DEC_MEMCTRL_load_store_width[0]) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_1_ ( .D(n820), .CP(
        clock), .Q(DEC_RF_memory_store_address_reg[1]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_1_ ( .D(n805), .CP(clock), 
        .Q(DEC_RF_alu_write_to_reg[1]) );
  DFQD1BWP12T irdecode_inst1_operator_b_modification_reg_0_ ( .D(n800), .CP(
        clock), .Q(DEC_MISC_OUT_operator_b_modification[0]) );
  DFQD1BWP12T irdecode_inst1_pc_mask_bit_reg ( .D(n797), .CP(clock), .Q(
        DEC_MISC_OUT_pc_mask_bit) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_2_ ( .D(n832), .CP(clock), .Q(
        DEC_ALU_alu_opcode[2]) );
  DFQD1BWP12T irdecode_inst1_load_store_width_reg_1_ ( .D(n823), .CP(clock), 
        .Q(DEC_MEMCTRL_load_store_width[1]) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_4_ ( .D(n817), .CP(
        clock), .Q(DEC_RF_memory_store_address_reg[4]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_2_ ( .D(n804), .CP(clock), 
        .Q(DEC_RF_alu_write_to_reg[2]) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_0_ ( .D(n821), .CP(
        clock), .Q(DEC_RF_memory_store_address_reg[0]) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_2_ ( .D(n819), .CP(
        clock), .Q(DEC_RF_memory_store_address_reg[2]) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_3_ ( .D(n818), .CP(
        clock), .Q(DEC_RF_memory_store_address_reg[3]) );
  DFQD1BWP12T irdecode_inst1_step_reg_6_ ( .D(irdecode_inst1_next_step_6_), 
        .CP(clock), .Q(irdecode_inst1_step[6]) );
  DFQD1BWP12T irdecode_inst1_step_reg_1_ ( .D(irdecode_inst1_next_step_1_), 
        .CP(clock), .Q(irdecode_inst1_step[1]) );
  DFQD1BWP12T irdecode_inst1_step_reg_0_ ( .D(irdecode_inst1_next_step_0_), 
        .CP(clock), .Q(irdecode_inst1_step[0]) );
  DFQD1BWP12T irdecode_inst1_step_reg_2_ ( .D(irdecode_inst1_next_step_2_), 
        .CP(clock), .Q(irdecode_inst1_step[2]) );
  DFQD1BWP12T irdecode_inst1_step_reg_3_ ( .D(irdecode_inst1_next_step_3_), 
        .CP(clock), .Q(irdecode_inst1_step[3]) );
  DFQD1BWP12T irdecode_inst1_step_reg_4_ ( .D(irdecode_inst1_next_step_4_), 
        .CP(clock), .Q(irdecode_inst1_step[4]) );
  DFQD1BWP12T irdecode_inst1_step_reg_5_ ( .D(irdecode_inst1_next_step_5_), 
        .CP(clock), .Q(irdecode_inst1_step[5]) );
  DFQD1BWP12T irdecode_inst1_step_reg_7_ ( .D(irdecode_inst1_next_step_7_), 
        .CP(clock), .Q(irdecode_inst1_step[7]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_1_ ( .D(n815), .CP(
        clock), .Q(DEC_RF_memory_store_data_reg[1]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_1_ ( .D(n809), .CP(clock), 
        .Q(DEC_RF_memory_write_to_reg[1]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_0_ ( .D(n816), .CP(
        clock), .Q(DEC_RF_memory_store_data_reg[0]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_0_ ( .D(n810), .CP(clock), 
        .Q(DEC_RF_memory_write_to_reg[0]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_2_ ( .D(n814), .CP(
        clock), .Q(DEC_RF_memory_store_data_reg[2]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_2_ ( .D(n808), .CP(clock), 
        .Q(DEC_RF_memory_write_to_reg[2]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_9_ ( .D(n844), .CP(clock), .Q(
        DEC_RF_offset_b[9]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_10_ ( .D(n843), .CP(clock), .Q(
        DEC_RF_offset_b[10]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_11_ ( .D(n842), .CP(clock), .Q(
        DEC_RF_offset_b[11]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_3_ ( .D(n850), .CP(clock), .Q(
        DEC_RF_offset_b[3]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_5_ ( .D(n848), .CP(clock), .Q(
        DEC_RF_offset_b[5]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_6_ ( .D(n847), .CP(clock), .Q(
        DEC_RF_offset_b[6]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_8_ ( .D(n845), .CP(clock), .Q(
        DEC_RF_offset_b[8]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_0_ ( .D(n802), .CP(clock), 
        .Q(DEC_RF_alu_write_to_reg[0]) );
  DFQD1BWP12T irdecode_inst1_split_instruction_reg ( .D(n854), .CP(clock), .Q(
        irdecode_inst1_split_instruction) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_4_ ( .D(n801), .CP(clock), 
        .Q(DEC_RF_alu_write_to_reg[4]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_0_ ( .D(n853), .CP(clock), .Q(
        DEC_RF_offset_b[0]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_3_ ( .D(n829), .CP(clock), .Q(
        DEC_ALU_alu_opcode[3]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_3_ ( .D(n813), .CP(
        clock), .Q(DEC_RF_memory_store_data_reg[3]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_3_ ( .D(n807), .CP(clock), 
        .Q(DEC_RF_memory_write_to_reg[3]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_4_ ( .D(n828), .CP(clock), .Q(
        DEC_ALU_alu_opcode[4]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_4_ ( .D(n812), .CP(
        clock), .Q(DEC_RF_memory_store_data_reg[4]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_0_ ( .D(n831), .CP(clock), .Q(
        DEC_ALU_alu_opcode[0]) );
  DFQD1BWP12T irdecode_inst1_memory_load_request_reg ( .D(n826), .CP(clock), 
        .Q(DEC_MEMCTRL_memory_load_request) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_enable_reg ( .D(n811), .CP(
        clock), .Q(DEC_RF_memory_write_to_reg_enable) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_1_ ( .D(n830), .CP(clock), .Q(
        DEC_ALU_alu_opcode[1]) );
  DFQD1BWP12T irdecode_inst1_memory_store_request_reg ( .D(n827), .CP(clock), 
        .Q(DEC_MEMCTRL_memory_store_request) );
  DFQD1BWP12T irdecode_inst1_memory_address_source_is_reg_reg ( .D(n822), .CP(
        clock), .Q(DEC_MISC_OUT_memory_address_source_is_reg) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_4_ ( .D(n806), .CP(clock), 
        .Q(DEC_RF_memory_write_to_reg[4]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_3_ ( .D(n803), .CP(clock), 
        .Q(DEC_RF_alu_write_to_reg[3]) );
  DFQD4BWP12T irdecode_inst1_operator_b_modification_reg_1_ ( .D(n799), .CP(
        clock), .Q(DEC_MISC_OUT_operator_b_modification[1]) );
  DFQD4BWP12T irdecode_inst1_operator_b_modification_reg_2_ ( .D(n798), .CP(
        clock), .Q(DEC_MISC_OUT_operator_b_modification[2]) );
  DFD4BWP12T irdecode_inst1_operand_a_reg_2_ ( .D(n779), .CP(clock), .Q(
        DEC_RF_operand_a[2]) );
  DFD4BWP12T irdecode_inst1_operand_a_reg_4_ ( .D(n776), .CP(clock), .Q(
        DEC_RF_operand_a[4]), .QN(n1781) );
  DFD4BWP12T irdecode_inst1_operand_b_reg_0_ ( .D(n775), .CP(clock), .Q(
        DEC_RF_operand_b[0]), .QN(n1001) );
  DFD4BWP12T irdecode_inst1_operand_a_reg_1_ ( .D(n780), .CP(clock), .Q(
        DEC_RF_operand_a[1]) );
  DFD4BWP12T irdecode_inst1_operand_a_reg_0_ ( .D(n777), .CP(clock), .Q(
        DEC_RF_operand_a[0]) );
  DFD4BWP12T irdecode_inst1_operand_b_reg_2_ ( .D(n773), .CP(clock), .Q(
        DEC_RF_operand_b[2]), .QN(n1771) );
  DFXD1BWP12T irdecode_inst1_offset_b_reg_2_ ( .D(n851), .CP(clock), .Q(
        DEC_RF_offset_b[2]) );
  DFXD1BWP12T irdecode_inst1_offset_b_reg_4_ ( .D(n849), .CP(clock), .Q(
        DEC_RF_offset_b[4]) );
  DFQD4BWP12T Instruction_Fetch_v2_inst1_currentState_reg_1_ ( .D(
        Instruction_Fetch_v2_inst1_N80), .CP(clock), .Q(
        Instruction_Fetch_v2_inst1_currentState_1_) );
  DFKCNXD1BWP12T Instruction_Fetch_v2_inst1_fetched_instruction_reg_reg_11_ ( 
        .CN(n1783), .D(n1782), .CP(clock), .QN(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_11_) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_1_ ( .D(n852), .CP(clock), .Q(
        DEC_RF_offset_b[1]) );
  DFMQD4BWP12T irdecode_inst1_operand_a_reg_3_ ( .DB(n877), .DA(n778), .SA(
        n1769), .CP(clock), .Q(n1770) );
  DFKCNQD4BWP12T irdecode_inst1_operand_b_reg_4_ ( .CN(n770), .D(n1769), .CP(
        clock), .Q(DEC_RF_operand_b[4]) );
  DFMD4BWP12T irdecode_inst1_operand_b_reg_1_ ( .DB(n877), .DA(n774), .SA(
        n1769), .CP(clock), .Q(n999), .QN(n998) );
  DFMD4BWP12T irdecode_inst1_operand_b_reg_3_ ( .DB(n877), .DA(n772), .SA(
        n1769), .CP(clock), .Q(n994), .QN(n995) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_7_ ( .D(n846), .CP(clock), .Q(
        DEC_RF_offset_b[7]) );
  TIELBWP12T U1007 ( .ZN(n877) );
  INVD1BWP12T U1008 ( .I(n877), .ZN(MEMCTRL_MEM_to_mem_mem_enable) );
  NR2D1BWP12T U1009 ( .A1(n1765), .A2(n1764), .ZN(n1768) );
  INVD1BWP12T U1010 ( .I(DEC_MISC_OUT_pc_mask_bit), .ZN(n1422) );
  INVD1BWP12T U1011 ( .I(DEC_MEMCTRL_memory_store_request), .ZN(n1554) );
  INVD1BWP12T U1012 ( .I(DEC_MEMCTRL_memory_load_request), .ZN(n1319) );
  INVD1BWP12T U1013 ( .I(IF_DEC_instruction[7]), .ZN(n1753) );
  INVD1BWP12T U1014 ( .I(IF_DEC_instruction[6]), .ZN(n1747) );
  INR2D1BWP12T U1015 ( .A1(Instruction_Fetch_v2_inst1_currentState_0_), .B1(
        Instruction_Fetch_v2_inst1_currentState_1_), .ZN(n1636) );
  ND2D1BWP12T U1016 ( .A1(RF_ALU_operand_b[26]), .A2(n1763), .ZN(n1389) );
  INR2D1BWP12T U1017 ( .A1(n1682), .B1(n1681), .ZN(n1683) );
  INVD1BWP12T U1018 ( .I(n1459), .ZN(n1391) );
  ND2D1BWP12T U1019 ( .A1(n1195), .A2(n1226), .ZN(n1234) );
  HICIND1BWP12T U1020 ( .A(RF_pc_out[24]), .CIN(n1211), .CO(n1202), .S(n1212)
         );
  INR2D1BWP12T U1021 ( .A1(n1013), .B1(n1638), .ZN(n1084) );
  INVD1BWP12T U1022 ( .I(n1084), .ZN(n1088) );
  INR2D1BWP12T U1023 ( .A1(n1012), .B1(n1011), .ZN(n1087) );
  INVD1BWP12T U1024 ( .I(n1607), .ZN(n1730) );
  INR2D1BWP12T U1025 ( .A1(n1010), .B1(n1638), .ZN(n1086) );
  INVD1BWP12T U1026 ( .I(n1087), .ZN(n1021) );
  INVD1BWP12T U1027 ( .I(n1215), .ZN(n1023) );
  INVD1BWP12T U1028 ( .I(DEC_MISC_OUT_operator_b_modification[1]), .ZN(n1052)
         );
  NR2D1BWP12T U1029 ( .A1(DEC_MISC_OUT_operator_b_modification[0]), .A2(
        DEC_MISC_OUT_operator_b_modification[2]), .ZN(n1050) );
  IOA21D1BWP12T U1030 ( .A1(ALU_MISC_OUT_result[0]), .A2(n1604), .B(n1306), 
        .ZN(MEMCTRL_IN_address[0]) );
  ND2D1BWP12T U1031 ( .A1(n1238), .A2(RF_pc_out[11]), .ZN(n1232) );
  NR2D1BWP12T U1032 ( .A1(n1761), .A2(n1753), .ZN(n1674) );
  ND2D1BWP12T U1033 ( .A1(n1033), .A2(n1783), .ZN(n1369) );
  ND2D1BWP12T U1034 ( .A1(n1365), .A2(n1032), .ZN(n1033) );
  NR2D1BWP12T U1035 ( .A1(n1026), .A2(n1031), .ZN(n1622) );
  INR2D1BWP12T U1036 ( .A1(n1025), .B1(n1634), .ZN(n1026) );
  INVD1BWP12T U1037 ( .I(n1369), .ZN(n1364) );
  INVD1BWP12T U1038 ( .I(n1761), .ZN(n1740) );
  INVD1BWP12T U1039 ( .I(n1674), .ZN(n1649) );
  INR2D1BWP12T U1040 ( .A1(n1005), .B1(n1638), .ZN(n1756) );
  INVD1BWP12T U1041 ( .I(n1756), .ZN(n1745) );
  INR2D1BWP12T U1042 ( .A1(n1004), .B1(n1638), .ZN(n1746) );
  INR2D1BWP12T U1043 ( .A1(n1007), .B1(n1638), .ZN(n1549) );
  ND2D1BWP12T U1044 ( .A1(n1674), .A2(n1381), .ZN(n1640) );
  ND2D1BWP12T U1045 ( .A1(n1414), .A2(n1747), .ZN(n1711) );
  NR2D1BWP12T U1046 ( .A1(n1649), .A2(n1329), .ZN(n1414) );
  ND2D1BWP12T U1047 ( .A1(n1351), .A2(n1622), .ZN(n1761) );
  INR2D1BWP12T U1048 ( .A1(n1783), .B1(n1780), .ZN(n1634) );
  INVD1BWP12T U1049 ( .I(n1586), .ZN(n1627) );
  INR2D1BWP12T U1050 ( .A1(DEC_MISC_OUT_operator_b_modification[0]), .B1(
        DEC_MISC_OUT_operator_b_modification[2]), .ZN(n1684) );
  INVD1BWP12T U1051 ( .I(reset), .ZN(n1783) );
  OAI21D1BWP12T U1052 ( .A1(n1780), .A2(n1688), .B(n1136), .ZN(
        IF_DEC_instruction[0]) );
  OAI21D1BWP12T U1053 ( .A1(n1780), .A2(n1687), .B(n1217), .ZN(
        IF_DEC_instruction[1]) );
  OAI21D1BWP12T U1054 ( .A1(n1780), .A2(n1693), .B(n1062), .ZN(
        IF_DEC_instruction[2]) );
  OAI21D1BWP12T U1055 ( .A1(n1780), .A2(n1695), .B(n1133), .ZN(
        IF_DEC_instruction[6]) );
  OAI21D1BWP12T U1056 ( .A1(n1780), .A2(n1689), .B(n1024), .ZN(
        IF_DEC_instruction[7]) );
  ND2D1BWP12T U1057 ( .A1(RF_ALU_operand_b[22]), .A2(n1040), .ZN(n1466) );
  ND2D1BWP12T U1058 ( .A1(RF_ALU_operand_b[22]), .A2(n1039), .ZN(n1489) );
  ND2D1BWP12T U1059 ( .A1(RF_ALU_operand_b[9]), .A2(n1039), .ZN(n1453) );
  ND3D1BWP12T U1060 ( .A1(n1766), .A2(n1686), .A3(n1685), .ZN(
        RF_ALU_operand_b_modified[31]) );
  AN2D1BWP12T U1061 ( .A1(n1684), .A2(n1052), .Z(n1053) );
  ND2D1BWP12T U1062 ( .A1(RF_ALU_operand_b[7]), .A2(n1446), .ZN(n1447) );
  ND2D1BWP12T U1063 ( .A1(RF_ALU_operand_b[17]), .A2(n1763), .ZN(n1452) );
  ND2D1BWP12T U1064 ( .A1(RF_ALU_operand_b[25]), .A2(n1040), .ZN(n1455) );
  INVD1BWP12T U1065 ( .I(n1496), .ZN(n1485) );
  ND2D1BWP12T U1066 ( .A1(RF_ALU_operand_b[12]), .A2(n1508), .ZN(n1509) );
  NR2D1BWP12T U1067 ( .A1(n1051), .A2(n1391), .ZN(n1054) );
  ND2D1BWP12T U1068 ( .A1(n1058), .A2(n1057), .ZN(n1059) );
  INR3D0BWP12T U1069 ( .A1(irdecode_inst1_N704), .B1(n1164), .B2(n1068), .ZN(
        n1151) );
  AN3D0BWP12T U1070 ( .A1(n1021), .A2(n1086), .A3(n1084), .Z(n1081) );
  AOI21D0BWP12T U1071 ( .A1(RF_MEMCTRL_address_reg[1]), .A2(n1603), .B(
        IF_RF_incremented_pc_out[1]), .ZN(n878) );
  IOA21D0BWP12T U1072 ( .A1(n1604), .A2(ALU_MISC_OUT_result[1]), .B(n878), 
        .ZN(MEMCTRL_IN_address[1]) );
  IND3D0BWP12T U1073 ( .A1(n1107), .B1(n1654), .B2(n1094), .ZN(n1101) );
  AN4D0BWP12T U1074 ( .A1(n1257), .A2(n1553), .A3(n1587), .A4(n1568), .Z(n1314) );
  IND4D0BWP12T U1075 ( .A1(n1538), .B1(n1159), .B2(n1160), .B3(n1352), .ZN(
        n1272) );
  AO222D0BWP12T U1076 ( .A1(n1512), .A2(n1002), .B1(RF_MEMCTRL_address_reg[2]), 
        .B2(n1603), .C1(ALU_MISC_OUT_result[2]), .C2(n1604), .Z(
        MEMCTRL_IN_address[2]) );
  CKND2D0BWP12T U1077 ( .A1(n1607), .A2(n1086), .ZN(n879) );
  NR2D0BWP12T U1078 ( .A1(n1063), .A2(n879), .ZN(n1729) );
  AO222D0BWP12T U1079 ( .A1(n1601), .A2(n1002), .B1(RF_MEMCTRL_address_reg[3]), 
        .B2(n1603), .C1(ALU_MISC_OUT_result[3]), .C2(n1604), .Z(
        MEMCTRL_IN_address[3]) );
  ND3D1BWP12T U1080 ( .A1(n1112), .A2(irdecode_inst1_N548), .A3(n1105), .ZN(
        n880) );
  OA31D1BWP12T U1081 ( .A1(n1669), .A2(n1107), .A3(n880), .B(n1180), .Z(n1109)
         );
  AOI21D0BWP12T U1082 ( .A1(n1152), .A2(n1155), .B(n1557), .ZN(n1312) );
  IND4D0BWP12T U1083 ( .A1(n1331), .B1(n1351), .B2(n1714), .B3(n1204), .ZN(
        n881) );
  AOI21D0BWP12T U1084 ( .A1(n1622), .A2(n881), .B(n1369), .ZN(n1349) );
  CKND2D0BWP12T U1085 ( .A1(n1655), .A2(n1608), .ZN(n882) );
  OAI21D0BWP12T U1086 ( .A1(n882), .A2(n1664), .B(n1726), .ZN(n1321) );
  AO222D0BWP12T U1087 ( .A1(n1491), .A2(n1002), .B1(RF_MEMCTRL_address_reg[4]), 
        .B2(n1603), .C1(ALU_MISC_OUT_result[4]), .C2(n1604), .Z(
        MEMCTRL_IN_address[4]) );
  IAO21D0BWP12T U1088 ( .A1(n1080), .A2(n1745), .B(n1381), .ZN(n1732) );
  MAOI22D0BWP12T U1089 ( .A1(n1086), .A2(n1084), .B1(n1086), .B2(n1084), .ZN(
        n883) );
  NR2D0BWP12T U1090 ( .A1(n1037), .A2(n883), .ZN(n1204) );
  OAI31D0BWP12T U1091 ( .A1(n1164), .A2(irdecode_inst1_N706), .A3(
        irdecode_inst1_N704), .B(n1163), .ZN(n884) );
  INR2D0BWP12T U1092 ( .A1(n1165), .B1(n884), .ZN(n885) );
  ND4D0BWP12T U1093 ( .A1(n1590), .A2(n885), .A3(n1587), .A4(n1567), .ZN(n886)
         );
  AOI211D1BWP12T U1094 ( .A1(irdecode_inst1_N548), .A2(n1168), .B(n1575), .C(
        n1167), .ZN(n887) );
  AOI21D1BWP12T U1095 ( .A1(n1182), .A2(n887), .B(n1627), .ZN(n888) );
  OAI31D0BWP12T U1096 ( .A1(n1365), .A2(n1321), .A3(n1713), .B(n1364), .ZN(
        n889) );
  AOI211D1BWP12T U1097 ( .A1(n1597), .A2(n886), .B(n888), .C(n889), .ZN(n1191)
         );
  AO222D0BWP12T U1098 ( .A1(n1602), .A2(n1002), .B1(RF_MEMCTRL_address_reg[5]), 
        .B2(n1603), .C1(ALU_MISC_OUT_result[5]), .C2(n1604), .Z(
        MEMCTRL_IN_address[5]) );
  AN2D0BWP12T U1099 ( .A1(n1002), .A2(n1223), .Z(IF_RF_incremented_pc_out[14])
         );
  IND3D0BWP12T U1100 ( .A1(n1759), .B1(n1702), .B2(n1706), .ZN(n1538) );
  AO22D0BWP12T U1101 ( .A1(n1744), .A2(n1731), .B1(n1525), .B2(n1728), .Z(
        n1612) );
  AO222D0BWP12T U1102 ( .A1(n1605), .A2(n1002), .B1(RF_MEMCTRL_address_reg[6]), 
        .B2(n1603), .C1(ALU_MISC_OUT_result[6]), .C2(n1604), .Z(
        MEMCTRL_IN_address[6]) );
  INR3D0BWP12T U1103 ( .A1(irdecode_inst1_N546), .B1(n1101), .B2(n1095), .ZN(
        n1167) );
  AOI22D0BWP12T U1104 ( .A1(RF_OUT_v), .A2(irdecode_inst1_itstate_6_), .B1(
        RF_OUT_c), .B2(n1028), .ZN(n890) );
  OAI21D0BWP12T U1105 ( .A1(n1378), .A2(irdecode_inst1_itstate_6_), .B(
        irdecode_inst1_itstate_7_), .ZN(n891) );
  IOA21D0BWP12T U1106 ( .A1(n890), .A2(n891), .B(irdecode_inst1_itstate_5_), 
        .ZN(n892) );
  OAI22D0BWP12T U1107 ( .A1(irdecode_inst1_itstate_6_), .A2(n1376), .B1(n1515), 
        .B2(n1375), .ZN(n893) );
  CKND0BWP12T U1108 ( .I(irdecode_inst1_itstate_7_), .ZN(n894) );
  OAI32D0BWP12T U1109 ( .A1(irdecode_inst1_itstate_7_), .A2(RF_OUT_n), .A3(
        n1515), .B1(n893), .B2(n894), .ZN(n895) );
  AOI211D0BWP12T U1110 ( .A1(n1028), .A2(n1027), .B(irdecode_inst1_itstate_5_), 
        .C(n895), .ZN(n896) );
  CKND0BWP12T U1111 ( .I(irdecode_inst1_itstate_4_), .ZN(n897) );
  AOI22D0BWP12T U1112 ( .A1(n1027), .A2(n1221), .B1(irdecode_inst1_itstate_7_), 
        .B2(n1376), .ZN(n898) );
  CKND0BWP12T U1113 ( .I(irdecode_inst1_itstate_6_), .ZN(n899) );
  AOI32D0BWP12T U1114 ( .A1(RF_OUT_n), .A2(irdecode_inst1_itstate_6_), .A3(
        n1221), .B1(n898), .B2(n899), .ZN(n900) );
  OR3D0BWP12T U1115 ( .A1(n1375), .A2(n899), .A3(n894), .Z(n901) );
  CKND0BWP12T U1116 ( .I(n892), .ZN(n902) );
  OAI211D0BWP12T U1117 ( .A1(irdecode_inst1_itstate_5_), .A2(n900), .B(n901), 
        .C(n892), .ZN(n903) );
  AOI21D0BWP12T U1118 ( .A1(n897), .A2(n903), .B(n1529), .ZN(n904) );
  OAI31D0BWP12T U1119 ( .A1(n902), .A2(n896), .A3(n897), .B(n904), .ZN(n1351)
         );
  AO222D0BWP12T U1120 ( .A1(n1604), .A2(ALU_MISC_OUT_result[7]), .B1(n1341), 
        .B2(n1002), .C1(n1603), .C2(RF_MEMCTRL_address_reg[7]), .Z(
        MEMCTRL_IN_address[7]) );
  NR4D0BWP12T U1121 ( .A1(n1155), .A2(irdecode_inst1_N707), .A3(
        irdecode_inst1_N710), .A4(irdecode_inst1_N708), .ZN(n905) );
  ND2D1BWP12T U1122 ( .A1(n905), .A2(n1072), .ZN(n1163) );
  CKND2D0BWP12T U1123 ( .A1(RF_pc_out[9]), .A2(RF_pc_out[10]), .ZN(n906) );
  TPNR2D1BWP12T U1124 ( .A1(n1234), .A2(n906), .ZN(n1238) );
  IOA21D0BWP12T U1125 ( .A1(n1384), .A2(n1416), .B(n1652), .ZN(n1668) );
  AN3D0BWP12T U1126 ( .A1(n1023), .A2(n1727), .A3(n1019), .Z(n1754) );
  IND2D0BWP12T U1127 ( .A1(n1178), .B1(n1315), .ZN(n907) );
  AN4D0BWP12T U1128 ( .A1(n1188), .A2(n1181), .A3(n1580), .A4(n1182), .Z(n908)
         );
  CKND0BWP12T U1129 ( .I(n1179), .ZN(n909) );
  AOI31D0BWP12T U1130 ( .A1(n1180), .A2(n908), .A3(n909), .B(n1627), .ZN(n910)
         );
  AOI211D0BWP12T U1131 ( .A1(n1597), .A2(n907), .B(n1369), .C(n910), .ZN(n1323) );
  INR2D0BWP12T U1132 ( .A1(n1220), .B1(n1700), .ZN(n1419) );
  AO222D0BWP12T U1133 ( .A1(n1604), .A2(ALU_MISC_OUT_result[8]), .B1(n1342), 
        .B2(n1002), .C1(n1603), .C2(RF_MEMCTRL_address_reg[8]), .Z(
        MEMCTRL_IN_address[8]) );
  MAOI22D0BWP12T U1134 ( .A1(n1286), .A2(n1285), .B1(n1286), .B2(n1285), .ZN(
        n911) );
  INR2D1BWP12T U1135 ( .A1(n1002), .B1(n911), .ZN(IF_RF_incremented_pc_out[15]) );
  AN2D1BWP12T U1136 ( .A1(irdecode_inst1_N707), .A2(n1071), .Z(n1156) );
  IND2D0BWP12T U1137 ( .A1(n1739), .B1(n1029), .ZN(n1712) );
  NR2D0BWP12T U1138 ( .A1(n1380), .A2(n1418), .ZN(n1544) );
  OA31D1BWP12T U1139 ( .A1(n1363), .A2(n1623), .A3(n1091), .B(n1622), .Z(n912)
         );
  AO211D1BWP12T U1140 ( .A1(n1586), .A2(n1562), .B(n912), .C(n1369), .Z(n1124)
         );
  AO222D0BWP12T U1141 ( .A1(n1604), .A2(ALU_MISC_OUT_result[9]), .B1(n1002), 
        .B2(n1340), .C1(RF_MEMCTRL_address_reg[9]), .C2(n1603), .Z(
        MEMCTRL_IN_address[9]) );
  IND2D0BWP12T U1142 ( .A1(n1147), .B1(n1149), .ZN(n1580) );
  IND2XD2BWP12T U1143 ( .A1(irdecode_inst1_N707), .B1(n1071), .ZN(n1164) );
  INR3D0BWP12T U1144 ( .A1(n1697), .B1(n1272), .B2(n1161), .ZN(n1355) );
  AN2D0BWP12T U1145 ( .A1(n1021), .A2(n1020), .Z(n1381) );
  AO222D0BWP12T U1146 ( .A1(ALU_MISC_OUT_result[10]), .A2(n1604), .B1(n1344), 
        .B2(n1002), .C1(RF_MEMCTRL_address_reg[10]), .C2(n1603), .Z(
        MEMCTRL_IN_address[10]) );
  MAOI22D0BWP12T U1147 ( .A1(n1669), .A2(n1206), .B1(n1205), .B2(n1643), .ZN(
        n913) );
  CKND0BWP12T U1148 ( .I(n1760), .ZN(n914) );
  OAI221D0BWP12T U1149 ( .A1(n1760), .A2(n913), .B1(n914), .B2(n1771), .C(
        n1349), .ZN(n773) );
  IND2D0BWP12T U1150 ( .A1(n1077), .B1(n1166), .ZN(n1324) );
  CKND2D0BWP12T U1151 ( .A1(n1283), .A2(RF_pc_out[13]), .ZN(n915) );
  NR2D0BWP12T U1152 ( .A1(n1284), .A2(n915), .ZN(n1286) );
  INR2D1BWP12T U1153 ( .A1(irdecode_inst1_N914), .B1(n1704), .ZN(n1715) );
  NR3D0BWP12T U1154 ( .A1(irdecode_inst1_itstate_3_), .A2(
        irdecode_inst1_itstate_5_), .A3(irdecode_inst1_itstate_4_), .ZN(n916)
         );
  AN3D0BWP12T U1155 ( .A1(n1028), .A2(n916), .A3(n1219), .Z(n1529) );
  CKND0BWP12T U1156 ( .I(n1023), .ZN(n917) );
  OR4D0BWP12T U1157 ( .A1(n1608), .A2(n1607), .A3(n1549), .A4(n917), .Z(n1701)
         );
  MAOI22D0BWP12T U1158 ( .A1(IF_DEC_instruction[6]), .A2(n1206), .B1(n1205), 
        .B2(n1653), .ZN(n918) );
  CKND0BWP12T U1159 ( .I(n1760), .ZN(n919) );
  OAI221D0BWP12T U1160 ( .A1(n1760), .A2(n918), .B1(n919), .B2(n1001), .C(
        n1349), .ZN(n775) );
  IND4D0BWP12T U1161 ( .A1(DEC_ALU_alu_opcode[0]), .B1(DEC_ALU_alu_opcode[2]), 
        .B2(DEC_ALU_alu_opcode[1]), .B3(n1423), .ZN(n920) );
  MAOI22D0BWP12T U1162 ( .A1(DEC_ALU_alu_opcode[4]), .A2(n920), .B1(
        DEC_ALU_alu_opcode[4]), .B2(RF_OUT_c), .ZN(ALU_IN_c) );
  CKND0BWP12T U1163 ( .I(n1164), .ZN(n921) );
  AOI31D0BWP12T U1164 ( .A1(n1078), .A2(IF_DEC_instruction[7]), .A3(n921), .B(
        n1079), .ZN(n1553) );
  INR2D0BWP12T U1165 ( .A1(n1183), .B1(n1745), .ZN(n1189) );
  OR4D0BWP12T U1166 ( .A1(n1339), .A2(n1512), .A3(n1602), .A4(n1601), .Z(n922)
         );
  OR4D0BWP12T U1167 ( .A1(n1491), .A2(n1605), .A3(n1341), .A4(n922), .Z(n923)
         );
  OR4XD1BWP12T U1168 ( .A1(n1340), .A2(n1342), .A3(n1344), .A4(n923), .Z(n924)
         );
  OR4XD1BWP12T U1169 ( .A1(n1343), .A2(n1345), .A3(RF_pc_out[13]), .A4(n924), 
        .Z(n925) );
  OR4XD1BWP12T U1170 ( .A1(RF_pc_out[15]), .A2(RF_pc_out[14]), .A3(
        RF_pc_out[16]), .A4(n925), .Z(n926) );
  OR4XD1BWP12T U1171 ( .A1(RF_pc_out[18]), .A2(RF_pc_out[17]), .A3(
        RF_pc_out[19]), .A4(n926), .Z(n927) );
  OR4D0BWP12T U1172 ( .A1(RF_pc_out[21]), .A2(RF_pc_out[20]), .A3(
        RF_pc_out[22]), .A4(n927), .Z(n928) );
  OR4D0BWP12T U1173 ( .A1(RF_pc_out[27]), .A2(RF_pc_out[24]), .A3(
        RF_pc_out[23]), .A4(n928), .Z(n929) );
  OR4D0BWP12T U1174 ( .A1(RF_pc_out[30]), .A2(RF_pc_out[26]), .A3(
        RF_pc_out[25]), .A4(n929), .Z(n930) );
  OR4D0BWP12T U1175 ( .A1(RF_pc_out[29]), .A2(RF_pc_out[28]), .A3(
        RF_pc_out[31]), .A4(n930), .Z(n1631) );
  OAI32D0BWP12T U1176 ( .A1(n1369), .A2(n1363), .A3(n1272), .B1(n1622), .B2(
        n1369), .ZN(n1583) );
  CKND0BWP12T U1177 ( .I(n1664), .ZN(n931) );
  OAI222D0BWP12T U1178 ( .A1(n931), .A2(n1549), .B1(n1712), .B2(n1747), .C1(
        n1541), .C2(n1647), .ZN(n932) );
  AOI21D0BWP12T U1179 ( .A1(n1250), .A2(IF_DEC_instruction[5]), .B(n932), .ZN(
        n933) );
  MOAI22D0BWP12T U1180 ( .A1(n1761), .A2(n933), .B1(n1760), .B2(
        DEC_RF_offset_b[6]), .ZN(n847) );
  ND2D1BWP12T U1181 ( .A1(irdecode_inst1_N914), .A2(n1759), .ZN(n934) );
  ND3D1BWP12T U1182 ( .A1(n934), .A2(n1159), .A3(n1352), .ZN(n1091) );
  IND4D1BWP12T U1183 ( .A1(n1145), .B1(irdecode_inst1_N546), .B2(n1141), .B3(
        n1307), .ZN(n1579) );
  ND3D0BWP12T U1184 ( .A1(n1587), .A2(n1568), .A3(n1588), .ZN(n935) );
  OAI31D0BWP12T U1185 ( .A1(n1176), .A2(n1312), .A3(n935), .B(n1556), .ZN(
        n1559) );
  MOAI22D0BWP12T U1186 ( .A1(RF_OUT_v), .A2(RF_OUT_n), .B1(RF_OUT_v), .B2(
        RF_OUT_n), .ZN(n1378) );
  OAI21D0BWP12T U1187 ( .A1(n1238), .A2(RF_pc_out[11]), .B(n1002), .ZN(n936)
         );
  AOI21D0BWP12T U1188 ( .A1(n1238), .A2(RF_pc_out[11]), .B(n936), .ZN(
        IF_RF_incremented_pc_out[11]) );
  NR2D0BWP12T U1189 ( .A1(n1240), .A2(n1241), .ZN(n937) );
  OAI21D0BWP12T U1190 ( .A1(RF_pc_out[6]), .A2(n937), .B(n1002), .ZN(n938) );
  AOI21D0BWP12T U1191 ( .A1(RF_pc_out[6]), .A2(n937), .B(n938), .ZN(
        IF_RF_incremented_pc_out[6]) );
  INR2D0BWP12T U1192 ( .A1(n1636), .B1(DEC_IF_stall_to_instructionfetch), .ZN(
        n939) );
  OA31D0BWP12T U1193 ( .A1(n1638), .A2(n1637), .A3(n939), .B(n1783), .Z(
        Instruction_Fetch_v2_inst1_N80) );
  INR2D0BWP12T U1194 ( .A1(n1321), .B1(n1544), .ZN(n940) );
  CKND0BWP12T U1195 ( .I(n1354), .ZN(n941) );
  AOI211D0BWP12T U1196 ( .A1(n1416), .A2(n941), .B(n1322), .C(n1745), .ZN(n942) );
  OAI211D0BWP12T U1197 ( .A1(n940), .A2(n1666), .B(n1355), .C(n942), .ZN(n943)
         );
  AOI22D0BWP12T U1198 ( .A1(DEC_RF_memory_store_data_reg[2]), .A2(n1760), .B1(
        n1622), .B2(n943), .ZN(n944) );
  CKND2D0BWP12T U1199 ( .A1(n1323), .A2(n944), .ZN(n814) );
  ND3D0BWP12T U1200 ( .A1(irdecode_inst1_N547), .A2(n1102), .A3(n1168), .ZN(
        n945) );
  IIND4D1BWP12T U1201 ( .A1(n1167), .A2(n1100), .B1(n1181), .B2(n945), .ZN(
        n1254) );
  AN2D0BWP12T U1202 ( .A1(n1002), .A2(n1265), .Z(IF_RF_incremented_pc_out[30])
         );
  CKND2D0BWP12T U1203 ( .A1(n1283), .A2(RF_pc_out[13]), .ZN(n946) );
  MAOI22D0BWP12T U1204 ( .A1(n1284), .A2(n946), .B1(n1284), .B2(n946), .ZN(
        n1223) );
  IND2D0BWP12T U1205 ( .A1(n1704), .B1(n1150), .ZN(n1661) );
  IOA21D0BWP12T U1206 ( .A1(n1702), .A2(n1248), .B(n1740), .ZN(n1642) );
  INR2D0BWP12T U1207 ( .A1(n1523), .B1(n1332), .ZN(n1520) );
  IND4D1BWP12T U1208 ( .A1(n1164), .B1(irdecode_inst1_N705), .B2(n1153), .B3(
        n1166), .ZN(n1590) );
  AO222D0BWP12T U1209 ( .A1(ALU_MISC_OUT_result[11]), .A2(n1604), .B1(n1345), 
        .B2(n1002), .C1(RF_MEMCTRL_address_reg[11]), .C2(n1603), .Z(
        MEMCTRL_IN_address[11]) );
  OAI21D0BWP12T U1210 ( .A1(RF_pc_out[3]), .A2(n1246), .B(n1002), .ZN(n947) );
  AOI21D0BWP12T U1211 ( .A1(RF_pc_out[3]), .A2(n1246), .B(n947), .ZN(
        IF_RF_incremented_pc_out[3]) );
  OAI21D0BWP12T U1212 ( .A1(n1239), .A2(RF_pc_out[9]), .B(n1002), .ZN(n948) );
  AOI21D0BWP12T U1213 ( .A1(n1239), .A2(RF_pc_out[9]), .B(n948), .ZN(
        IF_RF_incremented_pc_out[9]) );
  NR3D0BWP12T U1214 ( .A1(n1350), .A2(n1416), .A3(n1608), .ZN(n949) );
  AOI21D0BWP12T U1215 ( .A1(n1607), .A2(n1664), .B(n949), .ZN(n950) );
  ND4D0BWP12T U1216 ( .A1(n1351), .A2(n1352), .A3(n950), .A4(n1353), .ZN(n951)
         );
  AOI211D0BWP12T U1217 ( .A1(DEC_MEMCTRL_load_store_width[1]), .A2(n1760), .B(
        n1597), .C(n1369), .ZN(n952) );
  IOA21D0BWP12T U1218 ( .A1(n1622), .A2(n951), .B(n952), .ZN(n823) );
  IND2D1BWP12T U1219 ( .A1(irdecode_inst1_N909), .B1(irdecode_inst1_N915), 
        .ZN(n1150) );
  AN2D0BWP12T U1220 ( .A1(n1002), .A2(n1271), .Z(n1779) );
  IND2D0BWP12T U1221 ( .A1(DEC_CPSR_update_flag_c), .B1(RF_OUT_c), .ZN(n1294)
         );
  INR2D0BWP12T U1222 ( .A1(n1780), .B1(reset), .ZN(n1694) );
  INR2D0BWP12T U1223 ( .A1(n1561), .B1(n1562), .ZN(n1572) );
  AN3D0BWP12T U1224 ( .A1(n1587), .A2(n1588), .A3(n1589), .Z(n1594) );
  OAI21D0BWP12T U1225 ( .A1(RF_pc_out[2]), .A2(RF_pc_out[1]), .B(n1002), .ZN(
        n953) );
  AOI21D0BWP12T U1226 ( .A1(RF_pc_out[2]), .A2(RF_pc_out[1]), .B(n953), .ZN(
        IF_RF_incremented_pc_out[2]) );
  AN2D0BWP12T U1227 ( .A1(n1239), .A2(RF_pc_out[9]), .Z(n954) );
  OAI21D0BWP12T U1228 ( .A1(RF_pc_out[10]), .A2(n954), .B(n1002), .ZN(n955) );
  AOI21D0BWP12T U1229 ( .A1(RF_pc_out[10]), .A2(n954), .B(n955), .ZN(
        IF_RF_incremented_pc_out[10]) );
  OAI21D0BWP12T U1230 ( .A1(n1283), .A2(RF_pc_out[13]), .B(n1002), .ZN(n956)
         );
  AOI21D0BWP12T U1231 ( .A1(n1283), .A2(RF_pc_out[13]), .B(n956), .ZN(
        IF_RF_incremented_pc_out[13]) );
  CKND0BWP12T U1232 ( .I(n1556), .ZN(n957) );
  OAI222D0BWP12T U1233 ( .A1(n957), .A2(n1553), .B1(n1761), .B2(n1555), .C1(
        n1650), .C2(n1554), .ZN(n958) );
  AOI31D0BWP12T U1234 ( .A1(n1558), .A2(n1557), .A3(n1729), .B(n958), .ZN(n959) );
  ND3D0BWP12T U1235 ( .A1(n1617), .A2(n1559), .A3(n959), .ZN(n827) );
  MOAI22D0BWP12T U1236 ( .A1(n1643), .A2(n1712), .B1(IF_DEC_instruction[3]), 
        .B2(n1670), .ZN(n960) );
  AO22D0BWP12T U1237 ( .A1(n1608), .A2(n1664), .B1(n1416), .B2(n1675), .Z(n961) );
  AOI211D0BWP12T U1238 ( .A1(n1250), .A2(IF_DEC_instruction[4]), .B(n960), .C(
        n961), .ZN(n962) );
  MOAI22D0BWP12T U1239 ( .A1(n1761), .A2(n962), .B1(DEC_RF_offset_b[5]), .B2(
        n1760), .ZN(n848) );
  OAI211D0BWP12T U1240 ( .A1(n1607), .A2(n1749), .B(n1719), .C(n1518), .ZN(
        n963) );
  INR4D0BWP12T U1241 ( .A1(n1361), .B1(n1372), .B2(n1363), .B3(n963), .ZN(n964) );
  CKND2D0BWP12T U1242 ( .A1(DEC_ALU_alu_opcode[2]), .A2(n1760), .ZN(n965) );
  OAI211D0BWP12T U1243 ( .A1(n964), .A2(n1365), .B(n1364), .C(n965), .ZN(n832)
         );
  CKND0BWP12T U1244 ( .I(RF_pc_out[26]), .ZN(n966) );
  OAI21D0BWP12T U1245 ( .A1(n1201), .A2(n966), .B(n1002), .ZN(n967) );
  AOI21D0BWP12T U1246 ( .A1(n1201), .A2(n966), .B(n967), .ZN(
        IF_RF_incremented_pc_out[26]) );
  ND3D0BWP12T U1247 ( .A1(n1155), .A2(irdecode_inst1_N708), .A3(n1166), .ZN(
        n1568) );
  IND2D0BWP12T U1248 ( .A1(n1148), .B1(n1149), .ZN(n1578) );
  AN2D0BWP12T U1249 ( .A1(n1002), .A2(n1383), .Z(n1773) );
  OAI21D0BWP12T U1250 ( .A1(n1253), .A2(RF_pc_out[31]), .B(n1002), .ZN(n968)
         );
  AOI21D0BWP12T U1251 ( .A1(n1253), .A2(RF_pc_out[31]), .B(n968), .ZN(
        IF_RF_incremented_pc_out[31]) );
  IND3D0BWP12T U1252 ( .A1(n1224), .B1(n1283), .B2(RF_pc_out[14]), .ZN(n969)
         );
  OAI21D0BWP12T U1253 ( .A1(n1225), .A2(n969), .B(n1002), .ZN(n970) );
  AOI21D0BWP12T U1254 ( .A1(n1225), .A2(n969), .B(n970), .ZN(
        IF_RF_incremented_pc_out[16]) );
  OAI21D0BWP12T U1255 ( .A1(n1280), .A2(n1279), .B(n1002), .ZN(n971) );
  AOI21D0BWP12T U1256 ( .A1(n1280), .A2(n1279), .B(n971), .ZN(
        IF_RF_incremented_pc_out[18]) );
  CKND0BWP12T U1257 ( .I(RF_pc_out[20]), .ZN(n972) );
  OAI21D0BWP12T U1258 ( .A1(n1413), .A2(n972), .B(n1002), .ZN(n973) );
  AOI21D0BWP12T U1259 ( .A1(n1413), .A2(n972), .B(n973), .ZN(
        IF_RF_incremented_pc_out[20]) );
  AOI21D0BWP12T U1260 ( .A1(n1570), .A2(n1597), .B(n1124), .ZN(n1119) );
  OAI21D0BWP12T U1261 ( .A1(n1241), .A2(n1240), .B(n1002), .ZN(n974) );
  AOI21D0BWP12T U1262 ( .A1(n1241), .A2(n1240), .B(n974), .ZN(
        IF_RF_incremented_pc_out[5]) );
  INR3D0BWP12T U1263 ( .A1(n1387), .B1(n1520), .B2(n1715), .ZN(n975) );
  AO31D0BWP12T U1264 ( .A1(n1333), .A2(n975), .A3(n1361), .B(n1365), .Z(n976)
         );
  OAI211D0BWP12T U1265 ( .A1(n1423), .A2(n1650), .B(n1334), .C(n976), .ZN(n829) );
  NR3D0BWP12T U1266 ( .A1(n1759), .A2(n1373), .A3(n1372), .ZN(n977) );
  CKND0BWP12T U1267 ( .I(n1377), .ZN(n978) );
  MOAI22D0BWP12T U1268 ( .A1(RF_OUT_c), .A2(n978), .B1(RF_OUT_c), .B2(n1374), 
        .ZN(n979) );
  NR2D0BWP12T U1269 ( .A1(n1528), .A2(RF_OUT_z), .ZN(n980) );
  AOI211D0BWP12T U1270 ( .A1(RF_OUT_z), .A2(n1525), .B(n1380), .C(n980), .ZN(
        n981) );
  CKND0BWP12T U1271 ( .I(n1549), .ZN(n982) );
  CKND0BWP12T U1272 ( .I(n1376), .ZN(n983) );
  MAOI22D0BWP12T U1273 ( .A1(n1378), .A2(n1377), .B1(n1378), .B2(n1379), .ZN(
        n984) );
  AOI221D0BWP12T U1274 ( .A1(n1525), .A2(n1376), .B1(n1727), .B2(n983), .C(
        n984), .ZN(n985) );
  MUX2ND0BWP12T U1275 ( .I0(n1374), .I1(n1377), .S(RF_OUT_v), .ZN(n986) );
  MAOI22D0BWP12T U1276 ( .A1(RF_OUT_n), .A2(n1528), .B1(RF_OUT_n), .B2(n1525), 
        .ZN(n987) );
  CKND0BWP12T U1277 ( .I(n1745), .ZN(n988) );
  CKND0BWP12T U1278 ( .I(n1525), .ZN(n989) );
  MAOI22D0BWP12T U1279 ( .A1(n1375), .A2(n989), .B1(n1375), .B2(n1727), .ZN(
        n990) );
  OAI32D0BWP12T U1280 ( .A1(n1745), .A2(n986), .A3(n987), .B1(n988), .B2(n990), 
        .ZN(n991) );
  OAI32D0BWP12T U1281 ( .A1(n982), .A2(n1756), .A3(n985), .B1(n1549), .B2(n991), .ZN(n992) );
  AOI32D0BWP12T U1282 ( .A1(n979), .A2(n1381), .A3(n981), .B1(n992), .B2(n1381), .ZN(n993) );
  AOI31D0BWP12T U1283 ( .A1(n1702), .A2(n977), .A3(n993), .B(n1761), .ZN(
        irdecode_inst1_next_alu_write_to_reg_enable) );
  MOAI22D0BWP12T U1284 ( .A1(n1780), .A2(n1691), .B1(n1636), .B2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_3_), .ZN(
        IF_DEC_instruction[3]) );
  AO222D0BWP12T U1285 ( .A1(n1543), .A2(n1740), .B1(n1542), .B2(n1558), .C1(
        n1760), .C2(DEC_RF_operand_a[1]), .Z(n780) );
  TPND2D2BWP12T U1286 ( .A1(RF_ALU_operand_b[6]), .A2(n1496), .ZN(n1404) );
  AO22D1BWP12T U1287 ( .A1(n1040), .A2(RF_ALU_operand_b[21]), .B1(n1039), .B2(
        RF_ALU_operand_b[5]), .Z(n1681) );
  TPND2D1BWP12T U1288 ( .A1(RF_ALU_operand_b[21]), .A2(n1763), .ZN(n1499) );
  IOA21D2BWP12T U1289 ( .A1(RF_ALU_operand_b[20]), .A2(n1763), .B(n1045), .ZN(
        n1049) );
  ND2D3BWP12T U1290 ( .A1(RF_ALU_operand_b[12]), .A2(n1039), .ZN(n1045) );
  TPND2D3BWP12T U1291 ( .A1(n1395), .A2(n1394), .ZN(
        RF_ALU_operand_b_modified[26]) );
  TPNR2D2BWP12T U1292 ( .A1(n1124), .A2(n1123), .ZN(n1785) );
  TPOAI21D4BWP12T U1293 ( .A1(n1736), .A2(n1365), .B(n1120), .ZN(
        irdecode_inst1_next_step_1_) );
  CKND2D2BWP12T U1294 ( .A1(n1759), .A2(n1150), .ZN(n1736) );
  NR2D0BWP12T U1295 ( .A1(n1178), .A2(n1557), .ZN(n1122) );
  TPND2D1BWP12T U1296 ( .A1(RF_ALU_operand_b[28]), .A2(n1040), .ZN(n1046) );
  CKND2D2BWP12T U1297 ( .A1(RF_ALU_operand_b[0]), .A2(n1496), .ZN(n1486) );
  ND2D1BWP12T U1298 ( .A1(RF_ALU_operand_b[0]), .A2(n1501), .ZN(n1056) );
  CKND2D2BWP12T U1299 ( .A1(RF_ALU_operand_b[9]), .A2(n1040), .ZN(n1440) );
  TPND2D2BWP12T U1300 ( .A1(RF_ALU_operand_b[23]), .A2(n1039), .ZN(n1448) );
  AOI22D2BWP12T U1301 ( .A1(RF_ALU_operand_b[2]), .A2(n1040), .B1(
        RF_ALU_operand_b[18]), .B2(n1039), .ZN(n1507) );
  TPND2D2BWP12T U1302 ( .A1(RF_ALU_operand_b[2]), .A2(n1496), .ZN(n1441) );
  AOI22D0BWP12T U1303 ( .A1(RF_ALU_operand_b[2]), .A2(n1501), .B1(
        RF_ALU_operand_b[18]), .B2(n1763), .ZN(n1450) );
  CKND0BWP12T U1304 ( .I(RF_ALU_operand_b[28]), .ZN(n996) );
  INVD1BWP12T U1305 ( .I(n996), .ZN(n997) );
  TPND2D3BWP12T U1306 ( .A1(RF_ALU_operand_b[27]), .A2(n1039), .ZN(n1482) );
  CKND2D2BWP12T U1307 ( .A1(RF_ALU_operand_b[5]), .A2(n1496), .ZN(n1434) );
  TPND2D2BWP12T U1308 ( .A1(RF_ALU_operand_b[14]), .A2(n1040), .ZN(n1405) );
  CKND0BWP12T U1309 ( .I(n998), .ZN(n1000) );
  CKND2D2BWP12T U1310 ( .A1(RF_ALU_operand_b[31]), .A2(n1040), .ZN(n1462) );
  TPAOI22D2BWP12T U1311 ( .A1(RF_ALU_operand_b[21]), .A2(n1039), .B1(
        RF_ALU_operand_b[5]), .B2(n1040), .ZN(n1469) );
  CKND2D4BWP12T U1312 ( .A1(RF_ALU_operand_b[7]), .A2(n1042), .ZN(n1510) );
  TPND2D2BWP12T U1313 ( .A1(n1055), .A2(n1505), .ZN(
        RF_ALU_operand_b_modified[20]) );
  TPND2D2BWP12T U1314 ( .A1(RF_ALU_operand_b[13]), .A2(n1039), .ZN(n1500) );
  ND2XD0BWP12T U1315 ( .A1(RF_ALU_operand_b[2]), .A2(n1039), .ZN(n1393) );
  TPNR2D2BWP12T U1316 ( .A1(n1456), .A2(n1457), .ZN(n1458) );
  TPND2D2BWP12T U1317 ( .A1(n1453), .A2(n1452), .ZN(n1457) );
  TPNR2D2BWP12T U1318 ( .A1(n1503), .A2(n1502), .ZN(n1504) );
  ND3D4BWP12T U1319 ( .A1(n1435), .A2(n1433), .A3(n1434), .ZN(
        RF_ALU_operand_b_modified[5]) );
  ND3D2BWP12T U1320 ( .A1(n1437), .A2(n1510), .A3(n1436), .ZN(
        RF_ALU_operand_b_modified[11]) );
  TPND2D1BWP12T U1321 ( .A1(n1475), .A2(n1474), .ZN(n1476) );
  TPND2D1BWP12T U1322 ( .A1(RF_ALU_operand_b[14]), .A2(n1039), .ZN(n1474) );
  ND3XD3BWP12T U1323 ( .A1(n1511), .A2(n1510), .A3(n1509), .ZN(
        RF_ALU_operand_b_modified[12]) );
  ND3XD4BWP12T U1324 ( .A1(n1044), .A2(n1510), .A3(n1043), .ZN(
        RF_ALU_operand_b_modified[8]) );
  CKND2D2BWP12T U1325 ( .A1(RF_ALU_operand_b[7]), .A2(n1388), .ZN(n1460) );
  TPND2D3BWP12T U1326 ( .A1(RF_ALU_operand_b[25]), .A2(n1039), .ZN(n1439) );
  ND3D2BWP12T U1327 ( .A1(n1507), .A2(n1506), .A3(n1510), .ZN(
        RF_ALU_operand_b_modified[10]) );
  ND2D1BWP12T U1328 ( .A1(n1455), .A2(n1454), .ZN(n1456) );
  TPAOI22D4BWP12T U1329 ( .A1(RF_ALU_operand_b[16]), .A2(n1039), .B1(
        RF_ALU_operand_b[0]), .B2(n1040), .ZN(n1044) );
  ND3XD4BWP12T U1330 ( .A1(n1445), .A2(n1444), .A3(n1510), .ZN(
        RF_ALU_operand_b_modified[9]) );
  ND3D2BWP12T U1331 ( .A1(n1490), .A2(n1510), .A3(n1489), .ZN(
        RF_ALU_operand_b_modified[14]) );
  TPND2D2BWP12T U1332 ( .A1(n1458), .A2(n1505), .ZN(
        RF_ALU_operand_b_modified[17]) );
  CKAN2D4BWP12T U1333 ( .A1(n1459), .A2(
        DEC_MISC_OUT_operator_b_modification[0]), .Z(n1039) );
  TPNR3D8BWP12T U1334 ( .A1(n1484), .A2(
        DEC_MISC_OUT_operator_b_modification[0]), .A3(
        DEC_MISC_OUT_operator_b_modification[1]), .ZN(n1040) );
  ND2D1BWP12T U1335 ( .A1(n1654), .A2(n1093), .ZN(n1181) );
  TPNR2D2BWP12T U1336 ( .A1(n1146), .A2(n1116), .ZN(n1179) );
  TPND2D1BWP12T U1337 ( .A1(n1147), .A2(n1115), .ZN(n1116) );
  AOI211D0BWP12T U1338 ( .A1(n1670), .A2(IF_DEC_instruction[2]), .B(n1130), 
        .C(n1129), .ZN(n1131) );
  TPNR2D1BWP12T U1339 ( .A1(n1673), .A2(n1653), .ZN(n1130) );
  NR2D2BWP12T U1340 ( .A1(n1095), .A2(irdecode_inst1_N546), .ZN(n1112) );
  ND3D4BWP12T U1341 ( .A1(n1440), .A2(n1438), .A3(n1439), .ZN(
        RF_ALU_operand_b_modified[1]) );
  INVD1BWP12T U1342 ( .I(n1002), .ZN(n1632) );
  INR2D2BWP12T U1343 ( .A1(Instruction_Fetch_v2_inst1_currentState_1_), .B1(
        Instruction_Fetch_v2_inst1_currentState_0_), .ZN(n1002) );
  TPND2D2BWP12T U1344 ( .A1(RF_ALU_operand_b[15]), .A2(n1392), .ZN(n1425) );
  TIEHBWP12T U1345 ( .Z(n1769) );
  TPOAI22D2BWP12T U1346 ( .A1(n1554), .A2(MEMCTRL_write_finished), .B1(n1319), 
        .B2(MEMCTRL_read_finished), .ZN(n1031) );
  TPND2D2BWP12T U1347 ( .A1(n1031), .A2(n1783), .ZN(n1650) );
  INVD6BWP12T U1348 ( .I(n1650), .ZN(n1760) );
  AOI22D1BWP12T U1349 ( .A1(n1636), .A2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_12_), .B1(n1002), 
        .B2(MEMCTRL_RF_IF_data_in[12]), .ZN(n1003) );
  ND2D4BWP12T U1350 ( .A1(n1002), .A2(MEMCTRL_read_finished), .ZN(n1780) );
  INR2D4BWP12T U1351 ( .A1(n1780), .B1(n1636), .ZN(n1638) );
  INR2D4BWP12T U1352 ( .A1(n1003), .B1(n1638), .ZN(n1607) );
  AOI22D1BWP12T U1353 ( .A1(n1636), .A2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_9_), .B1(n1002), 
        .B2(MEMCTRL_RF_IF_data_in[9]), .ZN(n1004) );
  INVD1P75BWP12T U1354 ( .I(n1746), .ZN(n1608) );
  CKND2D0BWP12T U1355 ( .A1(n1730), .A2(n1608), .ZN(n1009) );
  AOI22D1BWP12T U1356 ( .A1(n1636), .A2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_11_), .B1(n1002), 
        .B2(MEMCTRL_RF_IF_data_in[11]), .ZN(n1005) );
  NR2D1BWP12T U1357 ( .A1(n1607), .A2(n1756), .ZN(n1609) );
  AOI22D1BWP12T U1358 ( .A1(n1636), .A2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_8_), .B1(n1002), 
        .B2(MEMCTRL_RF_IF_data_in[8]), .ZN(n1006) );
  INR2D2BWP12T U1359 ( .A1(n1006), .B1(n1638), .ZN(n1654) );
  INVD1BWP12T U1360 ( .I(n1654), .ZN(n1669) );
  AOI22D0BWP12T U1361 ( .A1(n1746), .A2(n1609), .B1(n1730), .B2(n1669), .ZN(
        n1008) );
  AOI22D1BWP12T U1362 ( .A1(n1636), .A2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_10_), .B1(n1002), 
        .B2(MEMCTRL_RF_IF_data_in[10]), .ZN(n1007) );
  MUX2XD0BWP12T U1363 ( .I0(n1009), .I1(n1008), .S(n1549), .Z(n1016) );
  AOI22D1BWP12T U1364 ( .A1(n1636), .A2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_13_), .B1(n1002), 
        .B2(MEMCTRL_RF_IF_data_in[13]), .ZN(n1010) );
  ND2D1BWP12T U1365 ( .A1(n1636), .A2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_14_), .ZN(n1012) );
  INR2D1BWP12T U1366 ( .A1(MEMCTRL_RF_IF_data_in[14]), .B1(n1780), .ZN(n1011)
         );
  NR2D1BWP12T U1367 ( .A1(n1086), .A2(n1021), .ZN(n1014) );
  AOI22D1BWP12T U1368 ( .A1(n1636), .A2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_15_), .B1(n1002), 
        .B2(MEMCTRL_RF_IF_data_in[15]), .ZN(n1013) );
  CKND2D2BWP12T U1369 ( .A1(n1014), .A2(n1088), .ZN(n1215) );
  ND2D1BWP12T U1370 ( .A1(n1088), .A2(n1021), .ZN(n1063) );
  NR2D1BWP12T U1371 ( .A1(n1063), .A2(n1086), .ZN(n1022) );
  NR2D1BWP12T U1372 ( .A1(n1730), .A2(n1756), .ZN(n1744) );
  TPND2D0BWP12T U1373 ( .A1(n1022), .A2(n1744), .ZN(n1015) );
  OAI21D1BWP12T U1374 ( .A1(n1016), .A2(n1215), .B(n1015), .ZN(n1331) );
  ND2D1BWP12T U1375 ( .A1(n1608), .A2(n1654), .ZN(n1377) );
  NR2D1BWP12T U1376 ( .A1(n1215), .A2(n1377), .ZN(n1018) );
  INVD1BWP12T U1377 ( .I(n1609), .ZN(n1738) );
  INVD1BWP12T U1378 ( .I(n1549), .ZN(n1416) );
  NR2D1BWP12T U1379 ( .A1(n1738), .A2(n1416), .ZN(n1017) );
  ND2D1BWP12T U1380 ( .A1(n1018), .A2(n1017), .ZN(n1415) );
  ND2D1BWP12T U1381 ( .A1(n1756), .A2(n1549), .ZN(n1380) );
  NR2D1BWP12T U1382 ( .A1(n1380), .A2(n1607), .ZN(n1019) );
  ND2D1BWP12T U1383 ( .A1(n1018), .A2(n1019), .ZN(n1329) );
  CKND2D1BWP12T U1384 ( .A1(n1415), .A2(n1329), .ZN(n1537) );
  NR2D1BWP12T U1385 ( .A1(n1331), .A2(n1537), .ZN(n1160) );
  INVD0BWP12T U1386 ( .I(n1160), .ZN(n1370) );
  INVD1BWP12T U1387 ( .I(n1086), .ZN(n1029) );
  NR3D1BWP12T U1388 ( .A1(n1029), .A2(n1607), .A3(n1084), .ZN(n1020) );
  TPND2D0BWP12T U1389 ( .A1(n1020), .A2(n1087), .ZN(n1354) );
  ND2D1BWP12T U1390 ( .A1(n1744), .A2(n1081), .ZN(n1697) );
  ND2D1BWP12T U1391 ( .A1(n1354), .A2(n1697), .ZN(n1187) );
  NR2D1BWP12T U1392 ( .A1(n1215), .A2(n1730), .ZN(n1542) );
  NR2D1BWP12T U1393 ( .A1(n1187), .A2(n1542), .ZN(n1735) );
  CKND2D1BWP12T U1394 ( .A1(n1654), .A2(n1746), .ZN(n1528) );
  INVD1BWP12T U1395 ( .I(n1528), .ZN(n1727) );
  INVD1BWP12T U1396 ( .I(n1754), .ZN(n1737) );
  ND2D1BWP12T U1397 ( .A1(n1735), .A2(n1737), .ZN(n1670) );
  INVD1BWP12T U1398 ( .I(n1670), .ZN(n1647) );
  CKND0BWP12T U1399 ( .I(n1381), .ZN(n1706) );
  CKND2D1BWP12T U1400 ( .A1(n1607), .A2(n1756), .ZN(n1030) );
  INVD1BWP12T U1401 ( .I(n1030), .ZN(n1036) );
  ND2D1BWP12T U1402 ( .A1(n1022), .A2(n1036), .ZN(n1702) );
  INVD1BWP12T U1403 ( .I(n1022), .ZN(n1080) );
  NR2D2BWP12T U1404 ( .A1(n1080), .A2(n1607), .ZN(n1759) );
  INVD1BWP12T U1405 ( .I(n1538), .ZN(n1719) );
  ND3XD0BWP12T U1406 ( .A1(n1647), .A2(n1719), .A3(n1701), .ZN(n1037) );
  NR2D1BWP12T U1407 ( .A1(n1370), .A2(n1037), .ZN(n1353) );
  CKND2D1BWP12T U1408 ( .A1(n1036), .A2(n1081), .ZN(n1534) );
  NR2D1BWP12T U1409 ( .A1(n1534), .A2(n1549), .ZN(n1728) );
  INVD1BWP12T U1410 ( .I(MEMCTRL_RF_IF_data_in[7]), .ZN(n1689) );
  ND2D1BWP12T U1411 ( .A1(n1636), .A2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_7_), .ZN(n1024) );
  CKND2D0BWP12T U1412 ( .A1(n1728), .A2(IF_DEC_instruction[7]), .ZN(n1366) );
  ND3D1BWP12T U1413 ( .A1(DEC_IF_stall_to_instructionfetch), .A2(
        irdecode_inst1_split_instruction), .A3(n1783), .ZN(n1025) );
  INVD3BWP12T U1414 ( .I(n1622), .ZN(n1365) );
  AOI21D0BWP12T U1415 ( .A1(n1353), .A2(n1366), .B(n1365), .ZN(n1034) );
  NR2D1BWP12T U1416 ( .A1(irdecode_inst1_itstate_7_), .A2(
        irdecode_inst1_itstate_6_), .ZN(n1028) );
  INVD1BWP12T U1417 ( .I(RF_OUT_z), .ZN(n1027) );
  INVD1BWP12T U1418 ( .I(irdecode_inst1_itstate_6_), .ZN(n1515) );
  CKND2D1BWP12T U1419 ( .A1(RF_OUT_c), .A2(n1027), .ZN(n1376) );
  ND2D1BWP12T U1420 ( .A1(n1378), .A2(n1027), .ZN(n1375) );
  CKND0BWP12T U1421 ( .I(irdecode_inst1_itstate_7_), .ZN(n1221) );
  NR3D1BWP12T U1422 ( .A1(irdecode_inst1_itstate_1_), .A2(
        irdecode_inst1_itstate_2_), .A3(irdecode_inst1_itstate_0_), .ZN(n1219)
         );
  CKND0BWP12T U1423 ( .I(n1351), .ZN(n1161) );
  INVD0BWP12T U1424 ( .I(n1728), .ZN(n1707) );
  CKND2D1BWP12T U1425 ( .A1(n1084), .A2(n1087), .ZN(n1739) );
  OAI22D0BWP12T U1426 ( .A1(n1707), .A2(n1746), .B1(n1030), .B2(n1712), .ZN(
        n1536) );
  NR2D1BWP12T U1427 ( .A1(n1161), .A2(n1536), .ZN(n1333) );
  INVD1BWP12T U1428 ( .I(n1031), .ZN(n1032) );
  OAI21D1BWP12T U1429 ( .A1(n1333), .A2(n1365), .B(n1364), .ZN(n1207) );
  AO211D0BWP12T U1430 ( .A1(n1760), .A2(n1770), .B(n1034), .C(n1207), .Z(n778)
         );
  INVD0BWP12T U1431 ( .I(MEMCTRL_RF_IF_data_in[4]), .ZN(n1690) );
  TPND2D0BWP12T U1432 ( .A1(n1636), .A2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_4_), .ZN(n1035) );
  OAI21D1BWP12T U1433 ( .A1(n1780), .A2(n1690), .B(n1035), .ZN(
        IF_DEC_instruction[4]) );
  INVD0BWP12T U1434 ( .I(IF_DEC_instruction[4]), .ZN(n1541) );
  NR2D0BWP12T U1435 ( .A1(n1537), .A2(n1036), .ZN(n1205) );
  INR2D1BWP12T U1436 ( .A1(n1086), .B1(n1739), .ZN(n1384) );
  ND2D1BWP12T U1437 ( .A1(n1738), .A2(n1384), .ZN(n1652) );
  INVD1BWP12T U1438 ( .I(n1668), .ZN(n1714) );
  OAI211D0BWP12T U1439 ( .A1(n1541), .A2(n1205), .B(n1204), .C(n1714), .ZN(
        n1038) );
  INVD1BWP12T U1440 ( .I(n1384), .ZN(n1749) );
  ND2D1BWP12T U1441 ( .A1(n1081), .A2(n1730), .ZN(n1350) );
  CKND2D1BWP12T U1442 ( .A1(n1749), .A2(n1350), .ZN(n1206) );
  AO222D0BWP12T U1443 ( .A1(n1038), .A2(n1740), .B1(n1206), .B2(n1674), .C1(
        n1000), .C2(n1760), .Z(n774) );
  INR2D4BWP12T U1444 ( .A1(DEC_MISC_OUT_operator_b_modification[1]), .B1(
        DEC_MISC_OUT_operator_b_modification[2]), .ZN(n1459) );
  INVD3BWP12T U1445 ( .I(DEC_MISC_OUT_operator_b_modification[2]), .ZN(n1484)
         );
  INVD1BWP12T U1446 ( .I(n1684), .ZN(n1041) );
  NR2D2BWP12T U1447 ( .A1(n1041), .A2(DEC_MISC_OUT_operator_b_modification[1]), 
        .ZN(n1042) );
  NR2D3BWP12T U1448 ( .A1(n1040), .A2(n1684), .ZN(n1508) );
  TPND2D2BWP12T U1449 ( .A1(RF_ALU_operand_b[8]), .A2(n1508), .ZN(n1043) );
  MUX2D2BWP12T U1450 ( .I0(DEC_MISC_OUT_operator_b_modification[2]), .I1(n1050), .S(n1052), .Z(n1763) );
  INVD1BWP12T U1451 ( .I(DEC_MISC_OUT_operator_b_modification[0]), .ZN(n1411)
         );
  NR3D1BWP12T U1452 ( .A1(n1411), .A2(n1484), .A3(
        DEC_MISC_OUT_operator_b_modification[1]), .ZN(n1501) );
  ND2D1BWP12T U1453 ( .A1(n1501), .A2(RF_ALU_operand_b[4]), .ZN(n1047) );
  CKND2D2BWP12T U1454 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  TPNR2D2BWP12T U1455 ( .A1(n1049), .A2(n1048), .ZN(n1055) );
  INVD1BWP12T U1456 ( .I(n1050), .ZN(n1051) );
  RCAOI22D2BWP12T U1457 ( .A1(RF_ALU_operand_b[15]), .A2(n1054), .B1(
        RF_ALU_operand_b[7]), .B2(n1053), .ZN(n1505) );
  IOA21D1BWP12T U1458 ( .A1(n1040), .A2(RF_ALU_operand_b[24]), .B(n1056), .ZN(
        n1060) );
  TPND2D2BWP12T U1459 ( .A1(RF_ALU_operand_b[16]), .A2(n1763), .ZN(n1058) );
  CKND2D2BWP12T U1460 ( .A1(RF_ALU_operand_b[8]), .A2(n1039), .ZN(n1057) );
  TPNR2D1BWP12T U1461 ( .A1(n1060), .A2(n1059), .ZN(n1061) );
  CKND2D2BWP12T U1462 ( .A1(n1061), .A2(n1505), .ZN(
        RF_ALU_operand_b_modified[16]) );
  INVD1BWP12T U1463 ( .I(MEMCTRL_RF_IF_data_in[2]), .ZN(n1693) );
  CKND2D1BWP12T U1464 ( .A1(n1636), .A2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_2_), .ZN(n1062) );
  ND2D1BWP12T U1465 ( .A1(n1729), .A2(n1622), .ZN(n1593) );
  INVD1BWP12T U1466 ( .I(n1593), .ZN(n1597) );
  NR3D1BWP12T U1467 ( .A1(irdecode_inst1_N709), .A2(irdecode_inst1_N710), .A3(
        irdecode_inst1_N708), .ZN(n1071) );
  INVD1BWP12T U1468 ( .I(irdecode_inst1_N706), .ZN(n1153) );
  INVD1BWP12T U1469 ( .I(irdecode_inst1_N705), .ZN(n1064) );
  ND2D1BWP12T U1470 ( .A1(n1153), .A2(n1064), .ZN(n1068) );
  INR2D0BWP12T U1471 ( .A1(n1151), .B1(IF_DEC_instruction[7]), .ZN(n1079) );
  NR2D1BWP12T U1472 ( .A1(n1079), .A2(irdecode_inst1_N710), .ZN(n1076) );
  NR2D1BWP12T U1473 ( .A1(n1068), .A2(irdecode_inst1_N704), .ZN(n1078) );
  INR2D1BWP12T U1474 ( .A1(n1078), .B1(IF_DEC_instruction[7]), .ZN(n1072) );
  NR2D1BWP12T U1475 ( .A1(irdecode_inst1_N707), .A2(irdecode_inst1_N709), .ZN(
        n1065) );
  ND2D1BWP12T U1476 ( .A1(n1072), .A2(n1065), .ZN(n1077) );
  CKND0BWP12T U1477 ( .I(irdecode_inst1_N708), .ZN(n1066) );
  ND2D0BWP12T U1478 ( .A1(n1066), .A2(irdecode_inst1_N710), .ZN(n1067) );
  INVD1BWP12T U1479 ( .I(irdecode_inst1_N709), .ZN(n1155) );
  OAI21D1BWP12T U1480 ( .A1(n1077), .A2(n1067), .B(n1163), .ZN(n1311) );
  CKND0BWP12T U1481 ( .I(n1068), .ZN(n1069) );
  AOI211XD0BWP12T U1482 ( .A1(irdecode_inst1_N706), .A2(irdecode_inst1_N705), 
        .B(n1069), .C(irdecode_inst1_N704), .ZN(n1070) );
  INR3D0BWP12T U1483 ( .A1(n1070), .B1(n1164), .B2(IF_DEC_instruction[7]), 
        .ZN(n1177) );
  NR2D1BWP12T U1484 ( .A1(n1311), .A2(n1177), .ZN(n1075) );
  CKND2D1BWP12T U1485 ( .A1(n1072), .A2(n1156), .ZN(n1165) );
  INVD1BWP12T U1486 ( .I(irdecode_inst1_N710), .ZN(n1152) );
  CKND2D1BWP12T U1487 ( .A1(n1152), .A2(irdecode_inst1_N708), .ZN(n1073) );
  NR2D1BWP12T U1488 ( .A1(n1077), .A2(n1073), .ZN(n1074) );
  INR2D1BWP12T U1489 ( .A1(n1165), .B1(n1074), .ZN(n1257) );
  ND2D1BWP12T U1490 ( .A1(n1075), .A2(n1257), .ZN(n1557) );
  INR2D2BWP12T U1491 ( .A1(n1076), .B1(n1557), .ZN(n1166) );
  ND2D1BWP12T U1492 ( .A1(n1324), .A2(n1553), .ZN(n1178) );
  ND2D1BWP12T U1493 ( .A1(n1122), .A2(n1152), .ZN(n1570) );
  CKND2D1BWP12T U1494 ( .A1(n1160), .A2(n1732), .ZN(n1623) );
  TPNR2D0BWP12T U1495 ( .A1(n1380), .A2(n1730), .ZN(n1082) );
  ND2D1BWP12T U1496 ( .A1(n1082), .A2(n1081), .ZN(n1748) );
  CKND2D0BWP12T U1497 ( .A1(n1748), .A2(n1739), .ZN(n1083) );
  NR2D1BWP12T U1498 ( .A1(n1728), .A2(n1083), .ZN(n1352) );
  TPNR2D0BWP12T U1499 ( .A1(n1754), .A2(n1542), .ZN(n1159) );
  CKND2D0BWP12T U1500 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
  NR3XD0BWP12T U1501 ( .A1(n1730), .A2(n1085), .A3(n1084), .ZN(n1675) );
  NR3XD0BWP12T U1502 ( .A1(n1088), .A2(n1087), .A3(n1086), .ZN(n1664) );
  TPNR2D0BWP12T U1503 ( .A1(n1675), .A2(n1664), .ZN(n1089) );
  ND2D1BWP12T U1504 ( .A1(n1089), .A2(n1350), .ZN(n1726) );
  NR2D1BWP12T U1505 ( .A1(n1726), .A2(n1187), .ZN(n1090) );
  TPND2D0BWP12T U1506 ( .A1(n1351), .A2(n1090), .ZN(n1363) );
  INVD1BWP12T U1507 ( .I(irdecode_inst1_N549), .ZN(n1168) );
  INVD1BWP12T U1508 ( .I(irdecode_inst1_N547), .ZN(n1141) );
  ND2D1BWP12T U1509 ( .A1(n1168), .A2(n1141), .ZN(n1095) );
  NR2D1BWP12T U1510 ( .A1(irdecode_inst1_N548), .A2(irdecode_inst1_N545), .ZN(
        n1094) );
  ND2D1BWP12T U1511 ( .A1(n1112), .A2(n1094), .ZN(n1098) );
  INVD1BWP12T U1512 ( .I(n1098), .ZN(n1103) );
  INVD0BWP12T U1513 ( .I(irdecode_inst1_N543), .ZN(n1096) );
  NR2XD0BWP12T U1514 ( .A1(n1096), .A2(irdecode_inst1_N544), .ZN(n1092) );
  ND2D1BWP12T U1515 ( .A1(n1103), .A2(n1092), .ZN(n1600) );
  NR2D1BWP12T U1516 ( .A1(n1600), .A2(irdecode_inst1_N542), .ZN(n1093) );
  NR2D1BWP12T U1517 ( .A1(irdecode_inst1_N542), .A2(irdecode_inst1_N543), .ZN(
        n1117) );
  INVD1BWP12T U1518 ( .I(irdecode_inst1_N544), .ZN(n1115) );
  ND2D1BWP12T U1519 ( .A1(n1117), .A2(n1115), .ZN(n1107) );
  ND3D0BWP12T U1520 ( .A1(n1096), .A2(n1115), .A3(irdecode_inst1_N542), .ZN(
        n1097) );
  TPNR2D0BWP12T U1521 ( .A1(n1098), .A2(n1097), .ZN(n1169) );
  NR2XD0BWP12T U1522 ( .A1(n1098), .A2(n1107), .ZN(n1099) );
  ND2D1BWP12T U1523 ( .A1(n1669), .A2(n1099), .ZN(n1188) );
  IOA21D0BWP12T U1524 ( .A1(n1654), .A2(n1169), .B(n1188), .ZN(n1100) );
  NR2D1BWP12T U1525 ( .A1(n1101), .A2(irdecode_inst1_N546), .ZN(n1102) );
  TPND3D0BWP12T U1526 ( .A1(n1102), .A2(irdecode_inst1_N549), .A3(n1141), .ZN(
        n1110) );
  ND2D1BWP12T U1527 ( .A1(n1103), .A2(irdecode_inst1_N544), .ZN(n1148) );
  INVD0BWP12T U1528 ( .I(n1117), .ZN(n1144) );
  NR2D1BWP12T U1529 ( .A1(n1148), .A2(n1144), .ZN(n1104) );
  CKND2D1BWP12T U1530 ( .A1(n1654), .A2(n1104), .ZN(n1170) );
  INVD1BWP12T U1531 ( .I(irdecode_inst1_N545), .ZN(n1105) );
  NR2D1BWP12T U1532 ( .A1(n1105), .A2(irdecode_inst1_N548), .ZN(n1106) );
  ND2D1BWP12T U1533 ( .A1(n1112), .A2(n1106), .ZN(n1147) );
  TPNR2D0BWP12T U1534 ( .A1(n1147), .A2(n1107), .ZN(n1108) );
  TPND2D0BWP12T U1535 ( .A1(n1654), .A2(n1108), .ZN(n1180) );
  ND3D1BWP12T U1536 ( .A1(n1110), .A2(n1170), .A3(n1109), .ZN(n1111) );
  TPNR2D2BWP12T U1537 ( .A1(n1254), .A2(n1111), .ZN(n1307) );
  INVD0BWP12T U1538 ( .I(n1112), .ZN(n1113) );
  NR2D1BWP12T U1539 ( .A1(n1113), .A2(irdecode_inst1_N548), .ZN(n1114) );
  ND2D1BWP12T U1540 ( .A1(n1307), .A2(n1114), .ZN(n1146) );
  ND2D1BWP12T U1541 ( .A1(n1179), .A2(n1117), .ZN(n1268) );
  ND2D1BWP12T U1542 ( .A1(n1268), .A2(n1307), .ZN(n1562) );
  TPNR2D2BWP12T U1543 ( .A1(n1701), .A2(n1365), .ZN(n1586) );
  AOI22D1BWP12T U1544 ( .A1(n1586), .A2(irdecode_inst1_N549), .B1(n1760), .B2(
        irdecode_inst1_step[1]), .ZN(n1118) );
  AN2XD2BWP12T U1545 ( .A1(n1119), .A2(n1118), .Z(n1120) );
  INVD1BWP12T U1546 ( .I(irdecode_inst1_step[0]), .ZN(n1121) );
  OAI22D1BWP12T U1547 ( .A1(n1122), .A2(n1593), .B1(n1650), .B2(n1121), .ZN(
        n1123) );
  INVD1P75BWP12T U1548 ( .I(n1785), .ZN(irdecode_inst1_next_step_0_) );
  ND2D1BWP12T U1549 ( .A1(n1759), .A2(n1745), .ZN(n1704) );
  TPNR2D1BWP12T U1550 ( .A1(irdecode_inst1_next_step_0_), .A2(n1704), .ZN(
        n1125) );
  CKND2D2BWP12T U1551 ( .A1(irdecode_inst1_next_step_1_), .A2(n1125), .ZN(
        n1248) );
  INR2D1BWP12T U1552 ( .A1(n1702), .B1(n1381), .ZN(n1126) );
  TPND2D2BWP12T U1553 ( .A1(n1248), .A2(n1126), .ZN(n1250) );
  INVD2BWP12T U1554 ( .I(n1250), .ZN(n1673) );
  INVD1BWP12T U1555 ( .I(MEMCTRL_RF_IF_data_in[3]), .ZN(n1691) );
  INVD1BWP12T U1556 ( .I(IF_DEC_instruction[3]), .ZN(n1653) );
  INVD1BWP12T U1557 ( .I(n1712), .ZN(n1731) );
  CKND2D0BWP12T U1558 ( .A1(n1731), .A2(IF_DEC_instruction[4]), .ZN(n1128) );
  AOI22D0BWP12T U1559 ( .A1(n1675), .A2(n1608), .B1(n1664), .B2(n1669), .ZN(
        n1127) );
  OAI211D0BWP12T U1560 ( .A1(n1549), .A2(n1652), .B(n1128), .C(n1127), .ZN(
        n1129) );
  MOAI22D1BWP12T U1561 ( .A1(n1131), .A2(n1761), .B1(n1760), .B2(
        DEC_RF_offset_b[4]), .ZN(n849) );
  NR2D1BWP12T U1562 ( .A1(DEC_MISC_OUT_memory_address_source_is_reg), .A2(
        Instruction_Fetch_v2_inst1_currentState_1_), .ZN(n1604) );
  INVD1BWP12T U1563 ( .I(DEC_MISC_OUT_memory_address_source_is_reg), .ZN(n1320) );
  NR2D1BWP12T U1564 ( .A1(n1320), .A2(
        Instruction_Fetch_v2_inst1_currentState_1_), .ZN(n1603) );
  NR4D0BWP12T U1565 ( .A1(RF_pc_out[4]), .A2(RF_pc_out[3]), .A3(RF_pc_out[2]), 
        .A4(RF_pc_out[1]), .ZN(n1338) );
  IND2D1BWP12T U1566 ( .A1(RF_pc_out[5]), .B1(n1338), .ZN(n1335) );
  NR2D1BWP12T U1567 ( .A1(RF_pc_out[6]), .A2(n1335), .ZN(n1247) );
  IND2D1BWP12T U1568 ( .A1(RF_pc_out[7]), .B1(n1247), .ZN(n1251) );
  NR2D1BWP12T U1569 ( .A1(RF_pc_out[8]), .A2(n1251), .ZN(n1297) );
  MAOI22D0BWP12T U1570 ( .A1(RF_pc_out[9]), .A2(n1297), .B1(RF_pc_out[9]), 
        .B2(n1297), .ZN(n1340) );
  INVD0BWP12T U1571 ( .I(MEMCTRL_RF_IF_data_in[5]), .ZN(n1692) );
  TPND2D0BWP12T U1572 ( .A1(n1636), .A2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_5_), .ZN(n1132) );
  OAI21D1BWP12T U1573 ( .A1(n1780), .A2(n1692), .B(n1132), .ZN(
        IF_DEC_instruction[5]) );
  INVD1BWP12T U1574 ( .I(IF_DEC_instruction[5]), .ZN(n1643) );
  CKND0BWP12T U1575 ( .I(DEC_RF_alu_write_to_reg[0]), .ZN(n1139) );
  TPNR2D0BWP12T U1576 ( .A1(n1363), .A2(n1331), .ZN(n1304) );
  NR2XD0BWP12T U1577 ( .A1(n1748), .A2(n1377), .ZN(n1523) );
  INVD1BWP12T U1578 ( .I(MEMCTRL_RF_IF_data_in[6]), .ZN(n1695) );
  CKND2D1BWP12T U1579 ( .A1(n1636), .A2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_6_), .ZN(n1133) );
  CKND2D0BWP12T U1580 ( .A1(n1753), .A2(IF_DEC_instruction[6]), .ZN(n1332) );
  NR2D1BWP12T U1581 ( .A1(n1608), .A2(n1654), .ZN(n1525) );
  AOI21D1BWP12T U1582 ( .A1(n1523), .A2(n1332), .B(n1612), .ZN(n1387) );
  INVD1BWP12T U1583 ( .I(n1701), .ZN(n1308) );
  NR2D0BWP12T U1584 ( .A1(n1754), .A2(n1308), .ZN(n1362) );
  NR2D1BWP12T U1585 ( .A1(n1654), .A2(n1746), .ZN(n1379) );
  ND2XD0BWP12T U1586 ( .A1(n1728), .A2(n1379), .ZN(n1718) );
  ND4D1BWP12T U1587 ( .A1(n1304), .A2(n1387), .A3(n1362), .A4(n1718), .ZN(
        n1357) );
  INVD1BWP12T U1588 ( .I(n1332), .ZN(n1526) );
  NR2D0BWP12T U1589 ( .A1(n1377), .A2(n1526), .ZN(n1135) );
  CKND0BWP12T U1590 ( .I(n1537), .ZN(n1134) );
  OAI211D1BWP12T U1591 ( .A1(n1135), .A2(n1748), .B(n1134), .C(n1749), .ZN(
        n1373) );
  RCAOI21D0BWP12T U1592 ( .A1(n1654), .A2(n1728), .B(n1373), .ZN(n1723) );
  INVD1BWP12T U1593 ( .I(MEMCTRL_RF_IF_data_in[0]), .ZN(n1688) );
  CKND2D1BWP12T U1594 ( .A1(n1636), .A2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_0_), .ZN(n1136) );
  INVD1BWP12T U1595 ( .I(IF_DEC_instruction[0]), .ZN(n1713) );
  NR2D0BWP12T U1596 ( .A1(n1712), .A2(n1744), .ZN(n1385) );
  NR3XD0BWP12T U1597 ( .A1(n1385), .A2(n1542), .A3(n1729), .ZN(n1720) );
  OAI22D0BWP12T U1598 ( .A1(n1723), .A2(n1713), .B1(n1654), .B2(n1720), .ZN(
        n1137) );
  TPOAI31D0BWP12T U1599 ( .A1(n1357), .A2(n1137), .A3(n1250), .B(n1622), .ZN(
        n1138) );
  OAI211D1BWP12T U1600 ( .A1(n1650), .A2(n1139), .B(n1138), .C(n1364), .ZN(
        n802) );
  INVD1BWP12T U1601 ( .I(irdecode_inst1_N548), .ZN(n1140) );
  ND2D1BWP12T U1602 ( .A1(n1140), .A2(n1168), .ZN(n1145) );
  TPNR2D0BWP12T U1603 ( .A1(n1145), .A2(n1141), .ZN(n1142) );
  CKND2D1BWP12T U1604 ( .A1(n1307), .A2(n1142), .ZN(n1571) );
  TPND2D0BWP12T U1605 ( .A1(n1579), .A2(n1571), .ZN(n1143) );
  TPAOI21D0BWP12T U1606 ( .A1(n1179), .A2(n1144), .B(n1143), .ZN(n1256) );
  CKND2D1BWP12T U1607 ( .A1(n1307), .A2(n1145), .ZN(n1561) );
  INVD1BWP12T U1608 ( .I(n1146), .ZN(n1149) );
  ND4D1BWP12T U1609 ( .A1(n1256), .A2(n1561), .A3(n1580), .A4(n1578), .ZN(
        n1310) );
  INVD1BWP12T U1610 ( .I(n1661), .ZN(n1613) );
  TPAOI21D0BWP12T U1611 ( .A1(n1310), .A2(n1308), .B(n1613), .ZN(n1158) );
  ND2XD0BWP12T U1612 ( .A1(n1166), .A2(n1151), .ZN(n1258) );
  CKND2D1BWP12T U1613 ( .A1(n1590), .A2(n1258), .ZN(n1176) );
  NR2D0BWP12T U1614 ( .A1(n1164), .A2(n1153), .ZN(n1154) );
  ND2D1BWP12T U1615 ( .A1(n1166), .A2(n1154), .ZN(n1588) );
  ND2D1BWP12T U1616 ( .A1(n1166), .A2(n1156), .ZN(n1587) );
  INVD1BWP12T U1617 ( .I(n1729), .ZN(n1705) );
  NR2D1BWP12T U1618 ( .A1(n1761), .A2(n1705), .ZN(n1556) );
  CKND2D0BWP12T U1619 ( .A1(n1760), .A2(irdecode_inst1_split_instruction), 
        .ZN(n1157) );
  OAI211D1BWP12T U1620 ( .A1(n1158), .A2(n1761), .B(n1559), .C(n1157), .ZN(
        n854) );
  OR2XD1BWP12T U1621 ( .A1(n1350), .A2(n1746), .Z(n1418) );
  INVD0BWP12T U1622 ( .I(n1675), .ZN(n1655) );
  ND2XD0BWP12T U1623 ( .A1(n1321), .A2(n1354), .ZN(n1174) );
  INR2D1BWP12T U1624 ( .A1(n1380), .B1(n1418), .ZN(n1322) );
  AOI21D1BWP12T U1625 ( .A1(n1174), .A2(n1745), .B(n1322), .ZN(n1317) );
  CKND2D1BWP12T U1626 ( .A1(n1355), .A2(n1317), .ZN(n1267) );
  NR2D0BWP12T U1627 ( .A1(n1354), .A2(n1654), .ZN(n1162) );
  AOI211D0BWP12T U1628 ( .A1(n1544), .A2(IF_DEC_instruction[0]), .B(n1267), 
        .C(n1162), .ZN(n1173) );
  CKND2D1BWP12T U1629 ( .A1(n1166), .A2(irdecode_inst1_N709), .ZN(n1567) );
  INVD1BWP12T U1630 ( .I(n1579), .ZN(n1575) );
  INVD0BWP12T U1631 ( .I(n1169), .ZN(n1171) );
  AN4D0BWP12T U1632 ( .A1(n1268), .A2(n1578), .A3(n1171), .A4(n1170), .Z(n1182) );
  CKND2D0BWP12T U1633 ( .A1(n1627), .A2(n1593), .ZN(n1183) );
  AOI22D0BWP12T U1634 ( .A1(n1183), .A2(n1745), .B1(n1760), .B2(
        DEC_RF_memory_store_data_reg[0]), .ZN(n1172) );
  OAI211D1BWP12T U1635 ( .A1(n1173), .A2(n1365), .B(n1191), .C(n1172), .ZN(
        n816) );
  AOI21D0BWP12T U1636 ( .A1(n1174), .A2(n1756), .B(n1544), .ZN(n1555) );
  IND3D0BWP12T U1637 ( .A1(n1272), .B1(n1555), .B2(n1351), .ZN(n1326) );
  INVD1BWP12T U1638 ( .I(n1322), .ZN(n1262) );
  INVD1BWP12T U1639 ( .I(IF_DEC_instruction[2]), .ZN(n1666) );
  AOI21D0BWP12T U1640 ( .A1(n1321), .A2(n1262), .B(n1666), .ZN(n1175) );
  AOI211D0BWP12T U1641 ( .A1(n1187), .A2(n1416), .B(n1326), .C(n1175), .ZN(
        n1185) );
  INR3XD0BWP12T U1642 ( .A1(n1588), .B1(n1177), .B2(n1176), .ZN(n1315) );
  AOI21D0BWP12T U1643 ( .A1(n1760), .A2(DEC_RF_memory_write_to_reg[2]), .B(
        n1189), .ZN(n1184) );
  OAI211D1BWP12T U1644 ( .A1(n1185), .A2(n1365), .B(n1323), .C(n1184), .ZN(
        n808) );
  NR2D0BWP12T U1645 ( .A1(n1262), .A2(n1713), .ZN(n1186) );
  AOI211D0BWP12T U1646 ( .A1(n1187), .A2(n1669), .B(n1326), .C(n1186), .ZN(
        n1192) );
  NR2D1BWP12T U1647 ( .A1(n1627), .A2(n1188), .ZN(n1565) );
  AOI211D0BWP12T U1648 ( .A1(n1760), .A2(DEC_RF_memory_write_to_reg[0]), .B(
        n1189), .C(n1565), .ZN(n1190) );
  OAI211D1BWP12T U1649 ( .A1(n1192), .A2(n1365), .B(n1191), .C(n1190), .ZN(
        n810) );
  INVD1BWP12T U1650 ( .I(RF_pc_out[14]), .ZN(n1284) );
  INVD0BWP12T U1651 ( .I(RF_pc_out[16]), .ZN(n1225) );
  ND2XD0BWP12T U1652 ( .A1(RF_pc_out[15]), .A2(RF_pc_out[13]), .ZN(n1224) );
  OR2XD1BWP12T U1653 ( .A1(n1225), .A2(n1224), .Z(n1197) );
  CKND2D1BWP12T U1654 ( .A1(RF_pc_out[5]), .A2(RF_pc_out[6]), .ZN(n1227) );
  CKND2D0BWP12T U1655 ( .A1(RF_pc_out[7]), .A2(RF_pc_out[8]), .ZN(n1193) );
  NR2D1BWP12T U1656 ( .A1(n1227), .A2(n1193), .ZN(n1195) );
  CKND2D1BWP12T U1657 ( .A1(RF_pc_out[2]), .A2(RF_pc_out[1]), .ZN(n1242) );
  TPND2D0BWP12T U1658 ( .A1(RF_pc_out[3]), .A2(RF_pc_out[4]), .ZN(n1194) );
  NR2XD1BWP12T U1659 ( .A1(n1242), .A2(n1194), .ZN(n1226) );
  INVD1BWP12T U1660 ( .I(RF_pc_out[12]), .ZN(n1231) );
  NR2D4BWP12T U1661 ( .A1(n1232), .A2(n1231), .ZN(n1283) );
  INVD1P75BWP12T U1662 ( .I(n1283), .ZN(n1196) );
  INR3XD2BWP12T U1663 ( .A1(RF_pc_out[14]), .B1(n1197), .B2(n1196), .ZN(n1281)
         );
  INVD1BWP12T U1664 ( .I(RF_pc_out[18]), .ZN(n1279) );
  NR2XD1BWP12T U1665 ( .A1(n1280), .A2(n1279), .ZN(n1277) );
  INR2D2BWP12T U1666 ( .A1(RF_pc_out[20]), .B1(n1413), .ZN(n1382) );
  INR2D2BWP12T U1667 ( .A1(RF_pc_out[26]), .B1(n1201), .ZN(n1199) );
  AN2D0BWP12T U1668 ( .A1(n1198), .A2(n1002), .Z(IF_RF_incremented_pc_out[28])
         );
  HICOND1BWP12T U1669 ( .A(RF_pc_out[27]), .CI(n1199), .CON(n1252), .S(n1200)
         );
  AN2XD1BWP12T U1670 ( .A1(n1200), .A2(n1002), .Z(n1775) );
  HICOND1BWP12T U1671 ( .A(RF_pc_out[25]), .CI(n1202), .CON(n1201), .S(n1203)
         );
  AN2D0BWP12T U1672 ( .A1(n1203), .A2(n1002), .Z(n1778) );
  IOA21D0BWP12T U1673 ( .A1(DEC_RF_operand_b[4]), .A2(n1760), .B(n1349), .ZN(
        n770) );
  INVD1BWP12T U1674 ( .I(n1207), .ZN(n1628) );
  NR2D0BWP12T U1675 ( .A1(n1726), .A2(n1384), .ZN(n1621) );
  CKND2D0BWP12T U1676 ( .A1(n1705), .A2(n1712), .ZN(n1619) );
  CKND0BWP12T U1677 ( .I(n1534), .ZN(n1618) );
  AOI22D0BWP12T U1678 ( .A1(n1619), .A2(n1416), .B1(n1618), .B2(
        IF_DEC_instruction[2]), .ZN(n1208) );
  OAI211D1BWP12T U1679 ( .A1(n1643), .A2(n1621), .B(n1353), .C(n1208), .ZN(
        n1209) );
  AOI22D1BWP12T U1680 ( .A1(n1209), .A2(n1622), .B1(n1760), .B2(
        DEC_RF_operand_a[2]), .ZN(n1210) );
  CKND2D1BWP12T U1681 ( .A1(n1628), .A2(n1210), .ZN(n779) );
  AN2D0BWP12T U1682 ( .A1(n1212), .A2(n1002), .Z(IF_RF_incremented_pc_out[24])
         );
  HICIND2BWP12T U1683 ( .A(RF_pc_out[22]), .CIN(n1213), .CO(n1273), .S(n1214)
         );
  CKAN2D0BWP12T U1684 ( .A1(n1214), .A2(n1002), .Z(
        IF_RF_incremented_pc_out[22]) );
  INVD1BWP12T U1685 ( .I(n1379), .ZN(n1374) );
  CKND2D1BWP12T U1686 ( .A1(n1609), .A2(n1416), .ZN(n1216) );
  NR3D1BWP12T U1687 ( .A1(n1374), .A2(n1216), .A3(n1215), .ZN(n1218) );
  CKND2D1BWP12T U1688 ( .A1(n1218), .A2(n1622), .ZN(n1700) );
  INVD1BWP12T U1689 ( .I(MEMCTRL_RF_IF_data_in[1]), .ZN(n1687) );
  CKND2D1BWP12T U1690 ( .A1(n1636), .A2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_1_), .ZN(n1217) );
  INVD1BWP12T U1691 ( .I(IF_DEC_instruction[1]), .ZN(n1722) );
  ND4D1BWP12T U1692 ( .A1(n1653), .A2(n1666), .A3(n1713), .A4(n1722), .ZN(
        n1220) );
  OAI22D1BWP12T U1693 ( .A1(n1700), .A2(n1220), .B1(reset), .B2(n1622), .ZN(
        n1699) );
  AOI211D1BWP12T U1694 ( .A1(n1219), .A2(irdecode_inst1_itstate_3_), .B(n1218), 
        .C(n1365), .ZN(n1420) );
  NR2D1BWP12T U1695 ( .A1(n1699), .A2(n1420), .ZN(n1516) );
  INVD1BWP12T U1696 ( .I(n1419), .ZN(n1514) );
  TPOAI22D0BWP12T U1697 ( .A1(n1516), .A2(n1221), .B1(n1753), .B2(n1514), .ZN(
        n833) );
  ND4D0BWP12T U1698 ( .A1(n1740), .A2(n1753), .A3(n1747), .A4(n1537), .ZN(
        n1222) );
  IOA21D0BWP12T U1699 ( .A1(DEC_MISC_OUT_operator_b_modification[1]), .A2(
        n1760), .B(n1222), .ZN(n799) );
  INVD1BWP12T U1700 ( .I(n1226), .ZN(n1241) );
  NR2D1BWP12T U1701 ( .A1(n1241), .A2(n1227), .ZN(n1236) );
  CKND2D1BWP12T U1702 ( .A1(n1236), .A2(RF_pc_out[7]), .ZN(n1229) );
  CKND0BWP12T U1703 ( .I(RF_pc_out[8]), .ZN(n1228) );
  XOR2XD1BWP12T U1704 ( .A1(n1229), .A2(n1228), .Z(n1230) );
  CKAN2D1BWP12T U1705 ( .A1(n1230), .A2(n1002), .Z(IF_RF_incremented_pc_out[8]) );
  XOR2XD1BWP12T U1706 ( .A1(n1232), .A2(n1231), .Z(n1233) );
  CKAN2D1BWP12T U1707 ( .A1(n1233), .A2(n1002), .Z(
        IF_RF_incremented_pc_out[12]) );
  INVD1BWP12T U1708 ( .I(n1234), .ZN(n1239) );
  CKND0BWP12T U1709 ( .I(RF_pc_out[7]), .ZN(n1235) );
  XNR2XD1BWP12T U1710 ( .A1(n1236), .A2(n1235), .ZN(n1237) );
  CKAN2D1BWP12T U1711 ( .A1(n1237), .A2(n1002), .Z(IF_RF_incremented_pc_out[7]) );
  CKND0BWP12T U1712 ( .I(RF_pc_out[5]), .ZN(n1240) );
  INVD1BWP12T U1713 ( .I(n1242), .ZN(n1246) );
  ND2XD0BWP12T U1714 ( .A1(n1246), .A2(RF_pc_out[3]), .ZN(n1244) );
  CKND0BWP12T U1715 ( .I(RF_pc_out[4]), .ZN(n1243) );
  XOR2XD1BWP12T U1716 ( .A1(n1244), .A2(n1243), .Z(n1245) );
  CKAN2D1BWP12T U1717 ( .A1(n1245), .A2(n1002), .Z(IF_RF_incremented_pc_out[4]) );
  INR2D1BWP12T U1718 ( .A1(Instruction_Fetch_v2_inst1_current_pc_modified_0_), 
        .B1(n1632), .ZN(IF_RF_incremented_pc_out[0]) );
  CKND0BWP12T U1719 ( .I(Instruction_Fetch_v2_inst1_currentState_1_), .ZN(
        n1629) );
  CKND2D1BWP12T U1720 ( .A1(n1319), .A2(n1629), .ZN(MEMCTRL_load_in) );
  MAOI22D0BWP12T U1721 ( .A1(RF_pc_out[7]), .A2(n1247), .B1(RF_pc_out[7]), 
        .B2(n1247), .ZN(n1341) );
  CKND2D1BWP12T U1722 ( .A1(n1760), .A2(DEC_RF_offset_b[11]), .ZN(n1249) );
  OAI211D1BWP12T U1723 ( .A1(n1549), .A2(n1642), .B(n1249), .C(n1640), .ZN(
        n842) );
  INVD1BWP12T U1724 ( .I(RF_pc_out[1]), .ZN(n1339) );
  NR2D0BWP12T U1725 ( .A1(RF_pc_out[1]), .A2(n1632), .ZN(
        IF_RF_incremented_pc_out[1]) );
  MOAI22D0BWP12T U1726 ( .A1(RF_pc_out[8]), .A2(n1251), .B1(RF_pc_out[8]), 
        .B2(n1251), .ZN(n1342) );
  HICIND1BWP12T U1727 ( .A(RF_pc_out[28]), .CIN(n1252), .CO(n1270), .S(n1198)
         );
  CKND0BWP12T U1728 ( .I(n1254), .ZN(n1255) );
  AOI21D0BWP12T U1729 ( .A1(n1256), .A2(n1255), .B(n1701), .ZN(n1261) );
  AOI21D0BWP12T U1730 ( .A1(n1314), .A2(n1258), .B(n1705), .ZN(n1260) );
  OAI22D0BWP12T U1731 ( .A1(n1321), .A2(n1722), .B1(n1746), .B2(n1354), .ZN(
        n1259) );
  NR3D1BWP12T U1732 ( .A1(n1261), .A2(n1260), .A3(n1259), .ZN(n1548) );
  OAI222D0BWP12T U1733 ( .A1(n1262), .A2(n1722), .B1(n1697), .B2(n1746), .C1(
        n1548), .C2(n1756), .ZN(n1263) );
  AO22XD0BWP12T U1734 ( .A1(n1263), .A2(n1740), .B1(n1760), .B2(
        DEC_RF_memory_write_to_reg[1]), .Z(n809) );
  HICIND1BWP12T U1735 ( .A(RF_pc_out[30]), .CIN(n1264), .CO(n1253), .S(n1265)
         );
  AOI21D0BWP12T U1736 ( .A1(n1756), .A2(n1324), .B(n1705), .ZN(n1266) );
  OAI21D0BWP12T U1737 ( .A1(n1267), .A2(n1266), .B(n1622), .ZN(n1269) );
  OA21D1BWP12T U1738 ( .A1(n1268), .A2(n1627), .B(n1364), .Z(n1334) );
  OAI211D1BWP12T U1739 ( .A1(n1756), .A2(n1627), .B(n1269), .C(n1334), .ZN(
        n1566) );
  AO21D1BWP12T U1740 ( .A1(n1760), .A2(DEC_RF_memory_store_data_reg[4]), .B(
        n1566), .Z(n812) );
  HICOND1BWP12T U1741 ( .A(RF_pc_out[29]), .CI(n1270), .CON(n1264), .S(n1271)
         );
  ND2D1BWP12T U1742 ( .A1(n1583), .A2(n1627), .ZN(n1552) );
  AO21D1BWP12T U1743 ( .A1(n1760), .A2(DEC_RF_memory_store_address_reg[3]), 
        .B(n1552), .Z(n818) );
  HICOND1BWP12T U1744 ( .A(RF_pc_out[23]), .CI(n1273), .CON(n1211), .S(n1274)
         );
  AN2D0BWP12T U1745 ( .A1(n1274), .A2(n1002), .Z(n1774) );
  IOA21D1BWP12T U1746 ( .A1(n1760), .A2(DEC_RF_offset_a[13]), .B(n1711), .ZN(
        n783) );
  IOA21D1BWP12T U1747 ( .A1(n1760), .A2(DEC_RF_offset_a[11]), .B(n1711), .ZN(
        n785) );
  NR2D8BWP12T U1748 ( .A1(n1039), .A2(n1040), .ZN(n1496) );
  AOI22D2BWP12T U1749 ( .A1(RF_ALU_operand_b[28]), .A2(n1039), .B1(
        RF_ALU_operand_b[4]), .B2(n1496), .ZN(n1276) );
  ND2D2BWP12T U1750 ( .A1(RF_ALU_operand_b[12]), .A2(n1040), .ZN(n1275) );
  TPND2D2BWP12T U1751 ( .A1(n1276), .A2(n1275), .ZN(
        RF_ALU_operand_b_modified[4]) );
  HICOND1BWP12T U1752 ( .A(RF_pc_out[19]), .CI(n1277), .CON(n1413), .S(n1278)
         );
  AN2D0BWP12T U1753 ( .A1(n1278), .A2(n1002), .Z(n1777) );
  HICOND2BWP12T U1754 ( .A(RF_pc_out[17]), .CI(n1281), .CON(n1280), .S(n1282)
         );
  AN2D0BWP12T U1755 ( .A1(n1282), .A2(n1002), .Z(n1776) );
  INVD0BWP12T U1756 ( .I(RF_pc_out[15]), .ZN(n1285) );
  TPND2D0BWP12T U1757 ( .A1(n1760), .A2(
        DEC_MEMCTRL_memorycontroller_sign_extend), .ZN(n1287) );
  OAI31D0BWP12T U1758 ( .A1(n1756), .A2(n1418), .A3(n1761), .B(n1287), .ZN(
        n825) );
  AO22XD0BWP12T U1759 ( .A1(n1694), .A2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_14_), .B1(n1634), 
        .B2(MEMCTRL_RF_IF_data_in[14]), .Z(Instruction_Fetch_v2_inst1_N97) );
  MUX2ND0BWP12T U1760 ( .I0(MEMCTRL_RF_IF_data_in[15]), .I1(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_15_), .S(n1780), 
        .ZN(n1288) );
  CKND2D1BWP12T U1761 ( .A1(n1288), .A2(n1783), .ZN(
        Instruction_Fetch_v2_inst1_N98) );
  MUX2ND0BWP12T U1762 ( .I0(MEMCTRL_RF_IF_data_in[12]), .I1(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_12_), .S(n1780), 
        .ZN(n1289) );
  CKND2D1BWP12T U1763 ( .A1(n1289), .A2(n1783), .ZN(
        Instruction_Fetch_v2_inst1_N95) );
  MUX2ND0BWP12T U1764 ( .I0(MEMCTRL_RF_IF_data_in[13]), .I1(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_13_), .S(n1780), 
        .ZN(n1290) );
  CKND2D1BWP12T U1765 ( .A1(n1290), .A2(n1783), .ZN(
        Instruction_Fetch_v2_inst1_N96) );
  MUX2ND0BWP12T U1766 ( .I0(MEMCTRL_RF_IF_data_in[10]), .I1(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_10_), .S(n1780), 
        .ZN(n1291) );
  CKND2D1BWP12T U1767 ( .A1(n1291), .A2(n1783), .ZN(
        Instruction_Fetch_v2_inst1_N93) );
  MUX2ND0BWP12T U1768 ( .I0(MEMCTRL_RF_IF_data_in[9]), .I1(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_9_), .S(n1780), 
        .ZN(n1292) );
  CKND2D1BWP12T U1769 ( .A1(n1292), .A2(n1783), .ZN(
        Instruction_Fetch_v2_inst1_N92) );
  MUX2ND0BWP12T U1770 ( .I0(MEMCTRL_RF_IF_data_in[8]), .I1(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_8_), .S(n1780), 
        .ZN(n1293) );
  CKND2D1BWP12T U1771 ( .A1(n1293), .A2(n1783), .ZN(
        Instruction_Fetch_v2_inst1_N91) );
  INVD1BWP12T U1772 ( .I(ALU_OUT_c), .ZN(n1296) );
  INVD1BWP12T U1773 ( .I(DEC_CPSR_update_flag_c), .ZN(n1295) );
  TPOAI21D1BWP12T U1774 ( .A1(n1296), .A2(n1295), .B(n1294), .ZN(new_c) );
  MUX2D1BWP12T U1775 ( .I0(RF_OUT_n), .I1(ALU_OUT_n), .S(
        DEC_CPSR_update_flag_z), .Z(new_n) );
  TPND2D0BWP12T U1776 ( .A1(ALU_MISC_OUT_result[12]), .A2(n1604), .ZN(n1300)
         );
  IND2D1BWP12T U1777 ( .A1(RF_pc_out[9]), .B1(n1297), .ZN(n1303) );
  NR2D1BWP12T U1778 ( .A1(RF_pc_out[10]), .A2(n1303), .ZN(n1301) );
  IND2XD1BWP12T U1779 ( .A1(RF_pc_out[11]), .B1(n1301), .ZN(n1298) );
  MOAI22D0BWP12T U1780 ( .A1(RF_pc_out[12]), .A2(n1298), .B1(RF_pc_out[12]), 
        .B2(n1298), .ZN(n1343) );
  AOI22D0BWP12T U1781 ( .A1(n1343), .A2(n1002), .B1(n1603), .B2(
        RF_MEMCTRL_address_reg[12]), .ZN(n1299) );
  CKND2D1BWP12T U1782 ( .A1(n1300), .A2(n1299), .ZN(MEMCTRL_IN_address[12]) );
  MAOI22D0BWP12T U1783 ( .A1(RF_pc_out[11]), .A2(n1301), .B1(RF_pc_out[11]), 
        .B2(n1301), .ZN(n1345) );
  CKND2D1BWP12T U1784 ( .A1(n1760), .A2(DEC_RF_offset_b[10]), .ZN(n1302) );
  OAI211D1BWP12T U1785 ( .A1(n1746), .A2(n1642), .B(n1302), .C(n1640), .ZN(
        n843) );
  MOAI22D0BWP12T U1786 ( .A1(RF_pc_out[10]), .A2(n1303), .B1(RF_pc_out[10]), 
        .B2(n1303), .ZN(n1344) );
  TPAOI31D0BWP12T U1787 ( .A1(n1304), .A2(n1387), .A3(n1661), .B(n1365), .ZN(
        n1305) );
  AO211D0BWP12T U1788 ( .A1(n1760), .A2(DEC_RF_alu_write_to_reg[4]), .B(n1369), 
        .C(n1305), .Z(n801) );
  AOI21D1BWP12T U1789 ( .A1(RF_MEMCTRL_address_reg[0]), .A2(n1603), .B(
        IF_RF_incremented_pc_out[0]), .ZN(n1306) );
  INVD0BWP12T U1790 ( .I(n1307), .ZN(n1309) );
  OAI21D1BWP12T U1791 ( .A1(n1310), .A2(n1309), .B(n1308), .ZN(n1757) );
  INVD1BWP12T U1792 ( .I(n1757), .ZN(n1741) );
  NR2D0BWP12T U1793 ( .A1(n1312), .A2(n1311), .ZN(n1313) );
  TPAOI31D0BWP12T U1794 ( .A1(n1315), .A2(n1314), .A3(n1313), .B(n1705), .ZN(
        n1316) );
  TPOAI21D0BWP12T U1795 ( .A1(n1741), .A2(n1316), .B(n1745), .ZN(n1318) );
  AO31D1BWP12T U1796 ( .A1(n1318), .A2(n1317), .A3(n1697), .B(n1761), .Z(n1725) );
  OAI21D0BWP12T U1797 ( .A1(n1650), .A2(n1319), .B(n1725), .ZN(n826) );
  NR2D1BWP12T U1798 ( .A1(n1761), .A2(n1745), .ZN(n1558) );
  ND2D1BWP12T U1799 ( .A1(n1741), .A2(n1558), .ZN(n1617) );
  INVD1BWP12T U1800 ( .I(n1556), .ZN(n1698) );
  OAI211D0BWP12T U1801 ( .A1(n1650), .A2(n1320), .B(n1617), .C(n1698), .ZN(
        n822) );
  AOI21D0BWP12T U1802 ( .A1(n1745), .A2(n1324), .B(n1705), .ZN(n1325) );
  OAI21D0BWP12T U1803 ( .A1(n1326), .A2(n1325), .B(n1622), .ZN(n1327) );
  OAI211D1BWP12T U1804 ( .A1(n1627), .A2(n1745), .B(n1327), .C(n1334), .ZN(
        n1328) );
  AO21D0BWP12T U1805 ( .A1(n1760), .A2(DEC_RF_memory_write_to_reg[4]), .B(
        n1328), .Z(n806) );
  AO211D0BWP12T U1806 ( .A1(n1760), .A2(DEC_RF_memory_write_to_reg[3]), .B(
        n1328), .C(n1565), .Z(n807) );
  CKND0BWP12T U1807 ( .I(DEC_ALU_alu_opcode[3]), .ZN(n1423) );
  CKND0BWP12T U1808 ( .I(n1329), .ZN(n1409) );
  OAI21D0BWP12T U1809 ( .A1(n1748), .A2(n1374), .B(n1415), .ZN(n1330) );
  AOI211D0BWP12T U1810 ( .A1(n1409), .A2(n1753), .B(n1331), .C(n1330), .ZN(
        n1361) );
  MOAI22D0BWP12T U1811 ( .A1(RF_pc_out[6]), .A2(n1335), .B1(RF_pc_out[6]), 
        .B2(n1335), .ZN(n1605) );
  NR2D0BWP12T U1812 ( .A1(RF_pc_out[2]), .A2(RF_pc_out[1]), .ZN(n1336) );
  MAOI22D0BWP12T U1813 ( .A1(RF_pc_out[3]), .A2(n1336), .B1(RF_pc_out[3]), 
        .B2(n1336), .ZN(n1601) );
  NR3D0BWP12T U1814 ( .A1(RF_pc_out[3]), .A2(RF_pc_out[2]), .A3(RF_pc_out[1]), 
        .ZN(n1337) );
  MAOI22D0BWP12T U1815 ( .A1(RF_pc_out[4]), .A2(n1337), .B1(RF_pc_out[4]), 
        .B2(n1337), .ZN(n1491) );
  MAOI22D0BWP12T U1816 ( .A1(RF_pc_out[2]), .A2(n1339), .B1(RF_pc_out[2]), 
        .B2(n1339), .ZN(n1512) );
  MAOI22D0BWP12T U1817 ( .A1(RF_pc_out[5]), .A2(n1338), .B1(RF_pc_out[5]), 
        .B2(n1338), .ZN(n1602) );
  CKND0BWP12T U1818 ( .I(n1631), .ZN(n1346) );
  TPAOI21D0BWP12T U1819 ( .A1(MEMCTRL_read_finished), .A2(n1346), .B(
        Instruction_Fetch_v2_inst1_first_instruction_fetched), .ZN(n1347) );
  NR2XD0BWP12T U1820 ( .A1(n1347), .A2(reset), .ZN(n874) );
  ND3D0BWP12T U1821 ( .A1(n1728), .A2(n1622), .A3(IF_DEC_instruction[6]), .ZN(
        n1348) );
  OAI211D0BWP12T U1822 ( .A1(n1650), .A2(n995), .B(n1349), .C(n1348), .ZN(n772) );
  CKND0BWP12T U1823 ( .I(n1726), .ZN(n1703) );
  AOI31D0BWP12T U1824 ( .A1(n1355), .A2(n1703), .A3(n1354), .B(n1365), .ZN(
        n1356) );
  AO211D0BWP12T U1825 ( .A1(n1760), .A2(DEC_RF_memory_store_address_reg[4]), 
        .B(n1369), .C(n1356), .Z(n817) );
  NR2XD0BWP12T U1826 ( .A1(n1357), .A2(n1538), .ZN(n1367) );
  CKND0BWP12T U1827 ( .I(n1720), .ZN(n1358) );
  MAOI22D0BWP12T U1828 ( .A1(n1416), .A2(n1358), .B1(n1723), .B2(n1666), .ZN(
        n1359) );
  AOI21D0BWP12T U1829 ( .A1(n1367), .A2(n1359), .B(n1365), .ZN(n1360) );
  AO211D0BWP12T U1830 ( .A1(n1760), .A2(DEC_RF_alu_write_to_reg[2]), .B(n1360), 
        .C(n1369), .Z(n804) );
  OAI211D0BWP12T U1831 ( .A1(n1525), .A2(n1707), .B(n1362), .C(n1720), .ZN(
        n1372) );
  INVD1BWP12T U1832 ( .I(n1748), .ZN(n1606) );
  CKND2D0BWP12T U1833 ( .A1(n1606), .A2(n1525), .ZN(n1518) );
  TPAOI21D0BWP12T U1834 ( .A1(n1367), .A2(n1366), .B(n1760), .ZN(n1368) );
  AO211D0BWP12T U1835 ( .A1(n1760), .A2(DEC_RF_alu_write_to_reg[3]), .B(n1369), 
        .C(n1368), .Z(n803) );
  OAI21D0BWP12T U1836 ( .A1(n1370), .A2(n1715), .B(n1622), .ZN(n1371) );
  OAI211D0BWP12T U1837 ( .A1(n1650), .A2(n1781), .B(n1628), .C(n1371), .ZN(
        n776) );
  HICOND1BWP12T U1838 ( .A(RF_pc_out[21]), .CI(n1382), .CON(n1213), .S(n1383)
         );
  NR3D0BWP12T U1839 ( .A1(n1385), .A2(n1606), .A3(n1384), .ZN(n1386) );
  CKND2D0BWP12T U1840 ( .A1(n1622), .A2(n1529), .ZN(n1533) );
  OAI22D0BWP12T U1841 ( .A1(n1761), .A2(n1387), .B1(n1386), .B2(n1533), .ZN(
        irdecode_inst1_next_update_flag_n) );
  NR2D1BWP12T U1842 ( .A1(n1411), .A2(DEC_MISC_OUT_operator_b_modification[1]), 
        .ZN(n1388) );
  IOA21D1BWP12T U1843 ( .A1(RF_ALU_operand_b[18]), .A2(n1040), .B(n1389), .ZN(
        n1390) );
  INR2D1BWP12T U1844 ( .A1(n1460), .B1(n1390), .ZN(n1395) );
  TPNR2D1BWP12T U1845 ( .A1(DEC_MISC_OUT_operator_b_modification[0]), .A2(
        n1391), .ZN(n1392) );
  AN2XD2BWP12T U1846 ( .A1(n1425), .A2(n1393), .Z(n1394) );
  ND2D1BWP12T U1847 ( .A1(n1558), .A2(n1759), .ZN(n1471) );
  TPND2D0BWP12T U1848 ( .A1(n1760), .A2(DEC_RF_offset_b[12]), .ZN(n1396) );
  OAI211D0BWP12T U1849 ( .A1(n1713), .A2(n1471), .B(n1396), .C(n1640), .ZN(
        n855) );
  TPND2D0BWP12T U1850 ( .A1(n1760), .A2(DEC_RF_offset_b[20]), .ZN(n1397) );
  OAI211D0BWP12T U1851 ( .A1(n1654), .A2(n1471), .B(n1397), .C(n1640), .ZN(
        n863) );
  TPND2D0BWP12T U1852 ( .A1(n1760), .A2(DEC_RF_offset_b[22]), .ZN(n1398) );
  OAI211D0BWP12T U1853 ( .A1(n1549), .A2(n1471), .B(n1398), .C(n1640), .ZN(
        n865) );
  TPND2D0BWP12T U1854 ( .A1(n1760), .A2(DEC_RF_offset_b[19]), .ZN(n1399) );
  OAI211D0BWP12T U1855 ( .A1(n1753), .A2(n1471), .B(n1399), .C(n1640), .ZN(
        n862) );
  TPND2D0BWP12T U1856 ( .A1(n1760), .A2(DEC_RF_offset_b[18]), .ZN(n1400) );
  OAI211D0BWP12T U1857 ( .A1(n1747), .A2(n1471), .B(n1400), .C(n1640), .ZN(
        n861) );
  TPND2D0BWP12T U1858 ( .A1(n1760), .A2(DEC_RF_offset_b[17]), .ZN(n1401) );
  OAI211D0BWP12T U1859 ( .A1(n1643), .A2(n1471), .B(n1401), .C(n1640), .ZN(
        n860) );
  TPND2D0BWP12T U1860 ( .A1(n1760), .A2(DEC_RF_offset_b[16]), .ZN(n1402) );
  OAI211D0BWP12T U1861 ( .A1(n1541), .A2(n1471), .B(n1402), .C(n1640), .ZN(
        n859) );
  TPND2D0BWP12T U1862 ( .A1(n1760), .A2(DEC_RF_offset_b[13]), .ZN(n1403) );
  OAI211D0BWP12T U1863 ( .A1(n1722), .A2(n1471), .B(n1403), .C(n1640), .ZN(
        n856) );
  TPND2D2BWP12T U1864 ( .A1(RF_ALU_operand_b[30]), .A2(n1039), .ZN(n1406) );
  ND3D2BWP12T U1865 ( .A1(n1406), .A2(n1405), .A3(n1404), .ZN(
        RF_ALU_operand_b_modified[6]) );
  CKND2D0BWP12T U1866 ( .A1(n1760), .A2(DEC_RF_offset_b[15]), .ZN(n1407) );
  OAI211D0BWP12T U1867 ( .A1(n1653), .A2(n1471), .B(n1407), .C(n1640), .ZN(
        n858) );
  TPND2D0BWP12T U1868 ( .A1(n1760), .A2(DEC_RF_offset_b[14]), .ZN(n1408) );
  OAI211D0BWP12T U1869 ( .A1(n1666), .A2(n1471), .B(n1408), .C(n1640), .ZN(
        n857) );
  CKND0BWP12T U1870 ( .I(n1415), .ZN(n1410) );
  AOI21D0BWP12T U1871 ( .A1(n1747), .A2(IF_DEC_instruction[7]), .B(n1526), 
        .ZN(n1517) );
  AOI22D1BWP12T U1872 ( .A1(n1410), .A2(n1517), .B1(n1409), .B2(n1526), .ZN(
        n1412) );
  OAI22D0BWP12T U1873 ( .A1(n1761), .A2(n1412), .B1(n1650), .B2(n1411), .ZN(
        n800) );
  AO21D0BWP12T U1874 ( .A1(n1760), .A2(DEC_RF_offset_a[4]), .B(n1414), .Z(n792) );
  AO21D0BWP12T U1875 ( .A1(n1760), .A2(DEC_RF_offset_a[5]), .B(n1414), .Z(n791) );
  AO21D0BWP12T U1876 ( .A1(n1760), .A2(DEC_RF_offset_a[3]), .B(n1414), .Z(n793) );
  AO21D0BWP12T U1877 ( .A1(n1760), .A2(DEC_RF_offset_a[7]), .B(n1414), .Z(n789) );
  AO21D0BWP12T U1878 ( .A1(n1760), .A2(DEC_RF_offset_a[2]), .B(n1414), .Z(n794) );
  AO21D0BWP12T U1879 ( .A1(n1760), .A2(DEC_RF_offset_a[1]), .B(n1414), .Z(n795) );
  AO21D0BWP12T U1880 ( .A1(n1760), .A2(DEC_RF_offset_a[0]), .B(n1414), .Z(n796) );
  AO21D0BWP12T U1881 ( .A1(n1760), .A2(DEC_RF_offset_a[6]), .B(n1414), .Z(n790) );
  CKND2D1BWP12T U1882 ( .A1(n1740), .A2(IF_DEC_instruction[6]), .ZN(n1648) );
  OAI22D0BWP12T U1883 ( .A1(n1648), .A2(n1415), .B1(n1650), .B2(n1484), .ZN(
        n798) );
  IOA21D0BWP12T U1884 ( .A1(n1760), .A2(DEC_RF_offset_b[31]), .B(n1640), .ZN(
        n875) );
  IOA21D0BWP12T U1885 ( .A1(n1760), .A2(DEC_RF_offset_b[30]), .B(n1640), .ZN(
        n873) );
  IOA21D0BWP12T U1886 ( .A1(n1760), .A2(DEC_RF_offset_b[29]), .B(n1640), .ZN(
        n872) );
  IOA21D0BWP12T U1887 ( .A1(n1760), .A2(DEC_RF_offset_b[28]), .B(n1640), .ZN(
        n871) );
  IOA21D0BWP12T U1888 ( .A1(n1760), .A2(DEC_RF_offset_b[27]), .B(n1640), .ZN(
        n870) );
  IOA21D0BWP12T U1889 ( .A1(n1760), .A2(DEC_RF_offset_b[26]), .B(n1640), .ZN(
        n869) );
  IOA21D0BWP12T U1890 ( .A1(n1760), .A2(DEC_RF_offset_b[25]), .B(n1640), .ZN(
        n868) );
  IOA21D0BWP12T U1891 ( .A1(n1760), .A2(DEC_RF_offset_b[24]), .B(n1640), .ZN(
        n867) );
  IOA21D0BWP12T U1892 ( .A1(n1760), .A2(DEC_RF_offset_b[23]), .B(n1640), .ZN(
        n866) );
  AOI21D0BWP12T U1893 ( .A1(n1740), .A2(n1416), .B(n1558), .ZN(n1417) );
  INVD1BWP12T U1894 ( .I(DEC_MEMCTRL_load_store_width[0]), .ZN(n1630) );
  OAI222D0BWP12T U1895 ( .A1(n1655), .A2(n1761), .B1(n1418), .B2(n1417), .C1(
        n1650), .C2(n1630), .ZN(n824) );
  AO222D0BWP12T U1896 ( .A1(n1699), .A2(irdecode_inst1_itstate_4_), .B1(
        IF_DEC_instruction[4]), .B2(n1419), .C1(irdecode_inst1_itstate_3_), 
        .C2(n1420), .Z(n836) );
  INVD1BWP12T U1897 ( .I(n1700), .ZN(n1421) );
  AO222D0BWP12T U1898 ( .A1(IF_DEC_instruction[1]), .A2(n1421), .B1(n1699), 
        .B2(irdecode_inst1_itstate_1_), .C1(n1420), .C2(
        irdecode_inst1_itstate_0_), .Z(n839) );
  AO222D0BWP12T U1899 ( .A1(n1699), .A2(irdecode_inst1_itstate_3_), .B1(
        IF_DEC_instruction[3]), .B2(n1421), .C1(irdecode_inst1_itstate_2_), 
        .C2(n1420), .Z(n837) );
  AO222D0BWP12T U1900 ( .A1(IF_DEC_instruction[2]), .A2(n1421), .B1(n1699), 
        .B2(irdecode_inst1_itstate_2_), .C1(n1420), .C2(
        irdecode_inst1_itstate_1_), .Z(n838) );
  AN2D4BWP12T U1901 ( .A1(RF_ALU_operand_a[1]), .A2(n1422), .Z(n1772) );
  INVD1BWP12T U1902 ( .I(DEC_MEMCTRL_load_store_width[1]), .ZN(n1424) );
  NR2XD0BWP12T U1903 ( .A1(n1424), .A2(
        Instruction_Fetch_v2_inst1_currentState_1_), .ZN(
        MEMCTRL_IN_load_store_width[1]) );
  AOI22D1BWP12T U1904 ( .A1(n1040), .A2(RF_ALU_operand_b[16]), .B1(
        RF_ALU_operand_b[0]), .B2(n1039), .ZN(n1429) );
  INVD1P75BWP12T U1905 ( .I(n1425), .ZN(n1427) );
  INVD2P3BWP12T U1906 ( .I(n1460), .ZN(n1426) );
  NR2XD3BWP12T U1907 ( .A1(n1427), .A2(n1426), .ZN(n1766) );
  CKND2D0BWP12T U1908 ( .A1(n1763), .A2(RF_ALU_operand_b[24]), .ZN(n1428) );
  ND3D2BWP12T U1909 ( .A1(n1429), .A2(n1766), .A3(n1428), .ZN(
        RF_ALU_operand_b_modified[24]) );
  TPND2D2BWP12T U1910 ( .A1(ALU_OUT_z), .A2(DEC_CPSR_update_flag_z), .ZN(n1432) );
  INVD0BWP12T U1911 ( .I(DEC_CPSR_update_flag_z), .ZN(n1430) );
  CKND2D1BWP12T U1912 ( .A1(n1430), .A2(RF_OUT_z), .ZN(n1431) );
  ND2D2BWP12T U1913 ( .A1(n1432), .A2(n1431), .ZN(new_z) );
  TPND2D3BWP12T U1914 ( .A1(RF_ALU_operand_b[13]), .A2(n1040), .ZN(n1435) );
  ND2D3BWP12T U1915 ( .A1(RF_ALU_operand_b[29]), .A2(n1039), .ZN(n1433) );
  AOI22D2BWP12T U1916 ( .A1(RF_ALU_operand_b[19]), .A2(n1039), .B1(
        RF_ALU_operand_b[3]), .B2(n1040), .ZN(n1437) );
  ND2D1BWP12T U1917 ( .A1(RF_ALU_operand_b[11]), .A2(n1508), .ZN(n1436) );
  TPND2D2BWP12T U1918 ( .A1(RF_ALU_operand_b[1]), .A2(n1496), .ZN(n1438) );
  CKND2D2BWP12T U1919 ( .A1(RF_ALU_operand_b[10]), .A2(n1040), .ZN(n1443) );
  ND2XD3BWP12T U1920 ( .A1(RF_ALU_operand_b[26]), .A2(n1039), .ZN(n1442) );
  ND3XD4BWP12T U1921 ( .A1(n1443), .A2(n1441), .A3(n1442), .ZN(
        RF_ALU_operand_b_modified[2]) );
  AOI22D2BWP12T U1922 ( .A1(n1040), .A2(RF_ALU_operand_b[1]), .B1(
        RF_ALU_operand_b[17]), .B2(n1039), .ZN(n1445) );
  ND2D1BWP12T U1923 ( .A1(RF_ALU_operand_b[9]), .A2(n1508), .ZN(n1444) );
  ND2D1BWP12T U1924 ( .A1(RF_ALU_operand_b[15]), .A2(n1508), .ZN(n1449) );
  NR2D1BWP12T U1925 ( .A1(n1508), .A2(n1459), .ZN(n1446) );
  ND3XD3BWP12T U1926 ( .A1(n1449), .A2(n1448), .A3(n1447), .ZN(
        RF_ALU_operand_b_modified[15]) );
  AOI22D1BWP12T U1927 ( .A1(n1040), .A2(RF_ALU_operand_b[26]), .B1(
        RF_ALU_operand_b[10]), .B2(n1039), .ZN(n1451) );
  ND3D1BWP12T U1928 ( .A1(n1451), .A2(n1505), .A3(n1450), .ZN(
        RF_ALU_operand_b_modified[18]) );
  TPND2D1BWP12T U1929 ( .A1(RF_ALU_operand_b[1]), .A2(n1501), .ZN(n1454) );
  BUFFD6BWP12T U1930 ( .I(RF_ALU_operand_a[27]), .Z(n1784) );
  ND2D1BWP12T U1931 ( .A1(RF_ALU_operand_b[15]), .A2(n1459), .ZN(n1463) );
  ND2D2BWP12T U1932 ( .A1(RF_ALU_operand_b[23]), .A2(n1763), .ZN(n1461) );
  ND4D2BWP12T U1933 ( .A1(n1463), .A2(n1462), .A3(n1461), .A4(n1460), .ZN(
        RF_ALU_operand_b_modified[23]) );
  ND2D1BWP12T U1934 ( .A1(RF_ALU_operand_b[30]), .A2(n1763), .ZN(n1464) );
  IOA21D1BWP12T U1935 ( .A1(RF_ALU_operand_b[6]), .A2(n1039), .B(n1464), .ZN(
        n1465) );
  INR2D1BWP12T U1936 ( .A1(n1466), .B1(n1465), .ZN(n1467) );
  ND2D1BWP12T U1937 ( .A1(n1467), .A2(n1766), .ZN(
        RF_ALU_operand_b_modified[30]) );
  ND2D2BWP12T U1938 ( .A1(RF_ALU_operand_b[13]), .A2(n1508), .ZN(n1468) );
  ND3XD3BWP12T U1939 ( .A1(n1469), .A2(n1510), .A3(n1468), .ZN(
        RF_ALU_operand_b_modified[13]) );
  TPND2D0BWP12T U1940 ( .A1(n1760), .A2(DEC_RF_offset_b[21]), .ZN(n1470) );
  OAI211D0BWP12T U1941 ( .A1(n1746), .A2(n1471), .B(n1470), .C(n1640), .ZN(
        n864) );
  ND2D1BWP12T U1942 ( .A1(RF_ALU_operand_b[22]), .A2(n1763), .ZN(n1473) );
  ND2D1BWP12T U1943 ( .A1(RF_ALU_operand_b[30]), .A2(n1040), .ZN(n1472) );
  TPND2D1BWP12T U1944 ( .A1(n1473), .A2(n1472), .ZN(n1477) );
  ND2D1BWP12T U1945 ( .A1(RF_ALU_operand_b[6]), .A2(n1501), .ZN(n1475) );
  TPNR2D1BWP12T U1946 ( .A1(n1477), .A2(n1476), .ZN(n1478) );
  TPND2D2BWP12T U1947 ( .A1(n1478), .A2(n1505), .ZN(
        RF_ALU_operand_b_modified[22]) );
  AOI22D1BWP12T U1948 ( .A1(RF_ALU_operand_b[27]), .A2(n1040), .B1(n1039), 
        .B2(RF_ALU_operand_b[11]), .ZN(n1480) );
  AOI22D0BWP12T U1949 ( .A1(RF_ALU_operand_b[19]), .A2(n1763), .B1(
        RF_ALU_operand_b[3]), .B2(n1501), .ZN(n1479) );
  ND3D1BWP12T U1950 ( .A1(n1480), .A2(n1505), .A3(n1479), .ZN(
        RF_ALU_operand_b_modified[19]) );
  CKND2D2BWP12T U1951 ( .A1(RF_ALU_operand_b[11]), .A2(n1040), .ZN(n1483) );
  TPND2D2BWP12T U1952 ( .A1(RF_ALU_operand_b[3]), .A2(n1496), .ZN(n1481) );
  ND3XD8BWP12T U1953 ( .A1(n1483), .A2(n1482), .A3(n1481), .ZN(
        RF_ALU_operand_b_modified[3]) );
  NR2D2BWP12T U1954 ( .A1(RF_ALU_operand_b[8]), .A2(n1484), .ZN(n1488) );
  TPOAI21D2BWP12T U1955 ( .A1(RF_ALU_operand_b[24]), .A2(
        DEC_MISC_OUT_operator_b_modification[2]), .B(n1485), .ZN(n1487) );
  TPOAI21D4BWP12T U1956 ( .A1(n1488), .A2(n1487), .B(n1486), .ZN(
        RF_ALU_operand_b_modified[0]) );
  AOI22D1BWP12T U1957 ( .A1(n1040), .A2(RF_ALU_operand_b[6]), .B1(
        RF_ALU_operand_b[14]), .B2(n1508), .ZN(n1490) );
  INVD1P75BWP12T U1958 ( .I(ALU_OUT_v), .ZN(n1495) );
  INVD1BWP12T U1959 ( .I(DEC_CPSR_update_flag_v), .ZN(n1494) );
  INR2D1BWP12T U1960 ( .A1(RF_OUT_v), .B1(DEC_CPSR_update_flag_v), .ZN(n1492)
         );
  INVD1BWP12T U1961 ( .I(n1492), .ZN(n1493) );
  TPOAI21D1BWP12T U1962 ( .A1(n1495), .A2(n1494), .B(n1493), .ZN(new_v) );
  AOI22D1BWP12T U1963 ( .A1(RF_ALU_operand_b[15]), .A2(n1040), .B1(
        RF_ALU_operand_b[7]), .B2(n1496), .ZN(n1498) );
  ND2D1BWP12T U1964 ( .A1(RF_ALU_operand_b[31]), .A2(n1039), .ZN(n1497) );
  TPND2D1BWP12T U1965 ( .A1(n1498), .A2(n1497), .ZN(
        RF_ALU_operand_b_modified[7]) );
  IOA21D2BWP12T U1966 ( .A1(RF_ALU_operand_b[29]), .A2(n1040), .B(n1499), .ZN(
        n1503) );
  IOA21D2BWP12T U1967 ( .A1(RF_ALU_operand_b[5]), .A2(n1501), .B(n1500), .ZN(
        n1502) );
  TPND2D2BWP12T U1968 ( .A1(n1505), .A2(n1504), .ZN(
        RF_ALU_operand_b_modified[21]) );
  ND2D1BWP12T U1969 ( .A1(RF_ALU_operand_b[10]), .A2(n1508), .ZN(n1506) );
  AOI22D1BWP12T U1970 ( .A1(RF_ALU_operand_b[20]), .A2(n1039), .B1(
        RF_ALU_operand_b[4]), .B2(n1040), .ZN(n1511) );
  INVD1BWP12T U1971 ( .I(irdecode_inst1_next_step_1_), .ZN(irdecode_inst1_N910) );
  CKND0BWP12T U1972 ( .I(irdecode_inst1_itstate_5_), .ZN(n1513) );
  OAI22D1BWP12T U1973 ( .A1(n1516), .A2(n1513), .B1(n1643), .B2(n1514), .ZN(
        n835) );
  OAI22D1BWP12T U1974 ( .A1(n1516), .A2(n1515), .B1(n1747), .B2(n1514), .ZN(
        n834) );
  OAI22D0BWP12T U1975 ( .A1(n1518), .A2(n1517), .B1(n1738), .B2(n1749), .ZN(
        n1519) );
  NR2D1BWP12T U1976 ( .A1(n1520), .A2(n1519), .ZN(n1524) );
  TPND2D0BWP12T U1977 ( .A1(n1740), .A2(n1612), .ZN(n1521) );
  OAI31D0BWP12T U1978 ( .A1(n1607), .A2(n1712), .A3(n1533), .B(n1521), .ZN(
        n1522) );
  RCAOI21D0BWP12T U1979 ( .A1(n1674), .A2(n1523), .B(n1522), .ZN(n1532) );
  OAI21D1BWP12T U1980 ( .A1(n1524), .A2(n1533), .B(n1532), .ZN(
        irdecode_inst1_next_update_flag_v) );
  AOI21D0BWP12T U1981 ( .A1(n1526), .A2(n1654), .B(n1525), .ZN(n1527) );
  OAI22D0BWP12T U1982 ( .A1(n1649), .A2(n1528), .B1(n1527), .B2(n1761), .ZN(
        n1530) );
  ND3XD0BWP12T U1983 ( .A1(n1530), .A2(n1606), .A3(n1529), .ZN(n1531) );
  OAI211D1BWP12T U1984 ( .A1(n1749), .A2(n1533), .B(n1532), .C(n1531), .ZN(
        irdecode_inst1_next_update_flag_c) );
  OAI21D0BWP12T U1985 ( .A1(n1534), .A2(n1722), .B(n1697), .ZN(n1535) );
  AOI211D0BWP12T U1986 ( .A1(n1608), .A2(n1619), .B(n1536), .C(n1535), .ZN(
        n1540) );
  NR2D0BWP12T U1987 ( .A1(n1538), .A2(n1537), .ZN(n1539) );
  OAI211D1BWP12T U1988 ( .A1(n1541), .A2(n1621), .B(n1540), .C(n1539), .ZN(
        n1543) );
  CKND0BWP12T U1989 ( .I(n1558), .ZN(n1547) );
  ND3XD0BWP12T U1990 ( .A1(n1740), .A2(n1544), .A3(IF_DEC_instruction[1]), 
        .ZN(n1546) );
  ND2XD0BWP12T U1991 ( .A1(n1760), .A2(DEC_RF_memory_store_data_reg[1]), .ZN(
        n1545) );
  OAI211D1BWP12T U1992 ( .A1(n1548), .A2(n1547), .B(n1546), .C(n1545), .ZN(
        n815) );
  NR2D0BWP12T U1993 ( .A1(n1593), .A2(n1549), .ZN(n1550) );
  AO211D1BWP12T U1994 ( .A1(n1760), .A2(DEC_RF_memory_store_address_reg[2]), 
        .B(n1552), .C(n1550), .Z(n819) );
  NR2D0BWP12T U1995 ( .A1(n1593), .A2(n1654), .ZN(n1551) );
  AO211D1BWP12T U1996 ( .A1(n1760), .A2(DEC_RF_memory_store_address_reg[0]), 
        .B(n1552), .C(n1551), .Z(n821) );
  CKND0BWP12T U1997 ( .I(n1567), .ZN(n1560) );
  TPNR2D0BWP12T U1998 ( .A1(n1570), .A2(n1560), .ZN(n1564) );
  MAOI22D0BWP12T U1999 ( .A1(n1760), .A2(irdecode_inst1_step[2]), .B1(n1572), 
        .B2(n1627), .ZN(n1563) );
  OAI211D1BWP12T U2000 ( .A1(n1564), .A2(n1593), .B(n1563), .C(n1583), .ZN(
        irdecode_inst1_next_step_2_) );
  AO211D1BWP12T U2001 ( .A1(n1760), .A2(DEC_RF_memory_store_data_reg[3]), .B(
        n1566), .C(n1565), .Z(n813) );
  CKND2D1BWP12T U2002 ( .A1(n1568), .A2(n1567), .ZN(n1569) );
  NR2D1BWP12T U2003 ( .A1(n1570), .A2(n1569), .ZN(n1589) );
  ND2D1BWP12T U2004 ( .A1(n1572), .A2(n1571), .ZN(n1582) );
  ND2XD0BWP12T U2005 ( .A1(n1582), .A2(n1586), .ZN(n1573) );
  OAI211D1BWP12T U2006 ( .A1(n1589), .A2(n1593), .B(n1573), .C(n1583), .ZN(
        n1574) );
  AO21D1BWP12T U2007 ( .A1(n1760), .A2(irdecode_inst1_step[3]), .B(n1574), .Z(
        irdecode_inst1_next_step_3_) );
  INVD1BWP12T U2008 ( .I(n1574), .ZN(n1577) );
  AOI22D0BWP12T U2009 ( .A1(n1575), .A2(n1586), .B1(n1760), .B2(
        irdecode_inst1_step[4]), .ZN(n1576) );
  OAI211D1BWP12T U2010 ( .A1(n1593), .A2(n1587), .B(n1577), .C(n1576), .ZN(
        irdecode_inst1_next_step_4_) );
  INVD1BWP12T U2011 ( .I(n1578), .ZN(n1585) );
  TPND2D0BWP12T U2012 ( .A1(n1580), .A2(n1579), .ZN(n1581) );
  TPOAI21D0BWP12T U2013 ( .A1(n1582), .A2(n1581), .B(n1586), .ZN(n1584) );
  CKND2D1BWP12T U2014 ( .A1(n1584), .A2(n1583), .ZN(n1596) );
  AOI21D1BWP12T U2015 ( .A1(n1586), .A2(n1585), .B(n1596), .ZN(n1599) );
  TPND2D0BWP12T U2016 ( .A1(n1594), .A2(n1590), .ZN(n1591) );
  AOI22D1BWP12T U2017 ( .A1(n1591), .A2(n1597), .B1(n1760), .B2(
        irdecode_inst1_step[6]), .ZN(n1592) );
  ND2D1BWP12T U2018 ( .A1(n1599), .A2(n1592), .ZN(irdecode_inst1_next_step_6_)
         );
  NR2D0BWP12T U2019 ( .A1(n1594), .A2(n1593), .ZN(n1595) );
  AO211D1BWP12T U2020 ( .A1(n1760), .A2(irdecode_inst1_step[5]), .B(n1596), 
        .C(n1595), .Z(irdecode_inst1_next_step_5_) );
  AOI21D0BWP12T U2021 ( .A1(n1760), .A2(irdecode_inst1_step[7]), .B(n1597), 
        .ZN(n1598) );
  OAI211D1BWP12T U2022 ( .A1(n1627), .A2(n1600), .B(n1599), .C(n1598), .ZN(
        irdecode_inst1_next_step_7_) );
  OAI21D0BWP12T U2023 ( .A1(n1606), .A2(n1754), .B(n1674), .ZN(n1616) );
  CKND2D0BWP12T U2024 ( .A1(n1760), .A2(DEC_ALU_alu_opcode[1]), .ZN(n1615) );
  AOI21D0BWP12T U2025 ( .A1(n1609), .A2(n1608), .B(n1607), .ZN(n1610) );
  OAI22D0BWP12T U2026 ( .A1(n1749), .A2(n1610), .B1(n1712), .B2(n1738), .ZN(
        n1611) );
  TPOAI31D0BWP12T U2027 ( .A1(n1613), .A2(n1612), .A3(n1611), .B(n1740), .ZN(
        n1614) );
  ND4D1BWP12T U2028 ( .A1(n1617), .A2(n1616), .A3(n1615), .A4(n1614), .ZN(n830) );
  AOI22D0BWP12T U2029 ( .A1(n1619), .A2(n1669), .B1(n1618), .B2(
        IF_DEC_instruction[0]), .ZN(n1620) );
  OAI211D0BWP12T U2030 ( .A1(n1653), .A2(n1621), .B(n1620), .C(n1736), .ZN(
        n1624) );
  OAI31D0BWP12T U2031 ( .A1(n1670), .A2(n1624), .A3(n1623), .B(n1622), .ZN(
        n1626) );
  ND2D1BWP12T U2032 ( .A1(n1760), .A2(DEC_RF_operand_a[0]), .ZN(n1625) );
  ND4D1BWP12T U2033 ( .A1(n1628), .A2(n1627), .A3(n1626), .A4(n1625), .ZN(n777) );
  ND2D1BWP12T U2034 ( .A1(n1630), .A2(n1629), .ZN(
        MEMCTRL_IN_load_store_width[0]) );
  INR3D0BWP12T U2035 ( .A1(
        Instruction_Fetch_v2_inst1_first_instruction_fetched), .B1(n1632), 
        .B2(n1631), .ZN(n1637) );
  OA21XD0BWP12T U2036 ( .A1(Instruction_Fetch_v2_inst1_currentState_1_), .A2(
        DEC_IF_stall_to_instructionfetch), .B(
        Instruction_Fetch_v2_inst1_currentState_0_), .Z(n1633) );
  TPOAI21D0BWP12T U2037 ( .A1(n1637), .A2(n1633), .B(n1783), .ZN(n1635) );
  INVD1BWP12T U2038 ( .I(n1634), .ZN(n1696) );
  ND2D1BWP12T U2039 ( .A1(n1635), .A2(n1696), .ZN(
        Instruction_Fetch_v2_inst1_N79) );
  CKND0BWP12T U2040 ( .I(n1735), .ZN(n1639) );
  AOI22D0BWP12T U2041 ( .A1(n1674), .A2(n1639), .B1(n1760), .B2(
        DEC_RF_offset_b[9]), .ZN(n1641) );
  OAI211D1BWP12T U2042 ( .A1(n1654), .A2(n1642), .B(n1641), .C(n1640), .ZN(
        n844) );
  TPNR2D0BWP12T U2043 ( .A1(n1647), .A2(n1643), .ZN(n1644) );
  AOI22D0BWP12T U2044 ( .A1(n1740), .A2(n1644), .B1(n1760), .B2(
        DEC_RF_offset_b[7]), .ZN(n1646) );
  TPND2D0BWP12T U2045 ( .A1(n1674), .A2(n1731), .ZN(n1645) );
  OAI211D1BWP12T U2046 ( .A1(n1648), .A2(n1673), .B(n1646), .C(n1645), .ZN(
        n846) );
  INVD1BWP12T U2047 ( .I(DEC_RF_offset_b[8]), .ZN(n1651) );
  OAI222D1BWP12T U2048 ( .A1(n1651), .A2(n1650), .B1(n1649), .B2(n1673), .C1(
        n1648), .C2(n1647), .ZN(n845) );
  NR2D0BWP12T U2049 ( .A1(n1652), .A2(n1746), .ZN(n1657) );
  OAI22D0BWP12T U2050 ( .A1(n1655), .A2(n1654), .B1(n1653), .B2(n1712), .ZN(
        n1656) );
  RCAOI211D0BWP12T U2051 ( .A1(n1670), .A2(IF_DEC_instruction[1]), .B(n1657), 
        .C(n1656), .ZN(n1658) );
  OAI21D1BWP12T U2052 ( .A1(n1673), .A2(n1666), .B(n1658), .ZN(n1659) );
  AO222D1BWP12T U2053 ( .A1(n1659), .A2(n1740), .B1(n1664), .B2(n1674), .C1(
        n1760), .C2(DEC_RF_offset_b[3]), .Z(n850) );
  NR2D0BWP12T U2054 ( .A1(n1712), .A2(n1722), .ZN(n1660) );
  AOI211D0BWP12T U2055 ( .A1(n1675), .A2(IF_DEC_instruction[6]), .B(n1660), 
        .C(n1729), .ZN(n1662) );
  OAI211D1BWP12T U2056 ( .A1(n1713), .A2(n1673), .B(n1662), .C(n1661), .ZN(
        n1663) );
  AO222D1BWP12T U2057 ( .A1(n1663), .A2(n1740), .B1(n1668), .B2(n1674), .C1(
        DEC_RF_offset_b[1]), .C2(n1760), .Z(n852) );
  CKND2D0BWP12T U2058 ( .A1(n1664), .A2(IF_DEC_instruction[6]), .ZN(n1665) );
  OAI211D0BWP12T U2059 ( .A1(n1666), .A2(n1712), .B(n1701), .C(n1665), .ZN(
        n1667) );
  AOI21D0BWP12T U2060 ( .A1(n1669), .A2(n1668), .B(n1667), .ZN(n1672) );
  CKND2D0BWP12T U2061 ( .A1(n1670), .A2(IF_DEC_instruction[0]), .ZN(n1671) );
  OAI211D1BWP12T U2062 ( .A1(n1722), .A2(n1673), .B(n1672), .C(n1671), .ZN(
        n1676) );
  AO222D1BWP12T U2063 ( .A1(n1676), .A2(n1740), .B1(n1675), .B2(n1674), .C1(
        n1760), .C2(DEC_RF_offset_b[2]), .Z(n851) );
  AOI22D0BWP12T U2064 ( .A1(n1040), .A2(RF_ALU_operand_b[19]), .B1(n1039), 
        .B2(RF_ALU_operand_b[3]), .ZN(n1678) );
  CKND2D0BWP12T U2065 ( .A1(RF_ALU_operand_b[27]), .A2(n1763), .ZN(n1677) );
  ND3D1BWP12T U2066 ( .A1(n1766), .A2(n1678), .A3(n1677), .ZN(
        RF_ALU_operand_b_modified[27]) );
  AOI22D1BWP12T U2067 ( .A1(RF_ALU_operand_b[20]), .A2(n1040), .B1(n1039), 
        .B2(RF_ALU_operand_b[4]), .ZN(n1680) );
  ND2D1BWP12T U2068 ( .A1(n997), .A2(n1763), .ZN(n1679) );
  ND3D1BWP12T U2069 ( .A1(n1766), .A2(n1680), .A3(n1679), .ZN(
        RF_ALU_operand_b_modified[28]) );
  ND2D1BWP12T U2070 ( .A1(RF_ALU_operand_b[29]), .A2(n1763), .ZN(n1682) );
  ND2D1BWP12T U2071 ( .A1(n1766), .A2(n1683), .ZN(
        RF_ALU_operand_b_modified[29]) );
  AOI22D1BWP12T U2072 ( .A1(n1763), .A2(RF_ALU_operand_b[31]), .B1(
        RF_ALU_operand_b[23]), .B2(n1040), .ZN(n1686) );
  CKND2D0BWP12T U2073 ( .A1(n1684), .A2(RF_ALU_operand_b[7]), .ZN(n1685) );
  MUX2ND0BWP12T U2074 ( .I0(MEMCTRL_RF_IF_data_in[11]), .I1(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_11_), .S(n1780), 
        .ZN(n1782) );
  MOAI22D0BWP12T U2075 ( .A1(n1696), .A2(n1687), .B1(n1694), .B2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_1_), .ZN(
        Instruction_Fetch_v2_inst1_N84) );
  MOAI22D0BWP12T U2076 ( .A1(n1696), .A2(n1688), .B1(n1694), .B2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_0_), .ZN(
        Instruction_Fetch_v2_inst1_N83) );
  MOAI22D0BWP12T U2077 ( .A1(n1696), .A2(n1689), .B1(n1694), .B2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_7_), .ZN(
        Instruction_Fetch_v2_inst1_N90) );
  MOAI22D0BWP12T U2078 ( .A1(n1696), .A2(n1690), .B1(n1694), .B2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_4_), .ZN(
        Instruction_Fetch_v2_inst1_N87) );
  MOAI22D0BWP12T U2079 ( .A1(n1696), .A2(n1691), .B1(n1694), .B2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_3_), .ZN(
        Instruction_Fetch_v2_inst1_N86) );
  MOAI22D0BWP12T U2080 ( .A1(n1696), .A2(n1692), .B1(n1694), .B2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_5_), .ZN(
        Instruction_Fetch_v2_inst1_N88) );
  MOAI22D0BWP12T U2081 ( .A1(n1696), .A2(n1693), .B1(n1694), .B2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_2_), .ZN(
        Instruction_Fetch_v2_inst1_N85) );
  MOAI22D0BWP12T U2082 ( .A1(n1696), .A2(n1695), .B1(n1694), .B2(
        Instruction_Fetch_v2_inst1_fetched_instruction_reg_6_), .ZN(
        Instruction_Fetch_v2_inst1_N89) );
  MOAI22D0BWP12T U2083 ( .A1(n1761), .A2(n1697), .B1(n1760), .B2(
        DEC_MISC_OUT_pc_mask_bit), .ZN(n797) );
  MOAI22D0BWP12T U2084 ( .A1(n1698), .A2(n1746), .B1(n1760), .B2(
        DEC_RF_memory_store_address_reg[1]), .ZN(n820) );
  MOAI22D0BWP12T U2085 ( .A1(n1713), .A2(n1700), .B1(n1699), .B2(
        irdecode_inst1_itstate_0_), .ZN(n840) );
  ND4D0BWP12T U2086 ( .A1(n1735), .A2(n1703), .A3(n1702), .A4(n1701), .ZN(
        n1709) );
  ND4D0BWP12T U2087 ( .A1(n1707), .A2(n1706), .A3(n1705), .A4(n1704), .ZN(
        n1708) );
  NR2XD0BWP12T U2088 ( .A1(n1709), .A2(n1708), .ZN(n1710) );
  MOAI22D0BWP12T U2089 ( .A1(n1761), .A2(n1710), .B1(n1760), .B2(
        DEC_IF_stall_to_instructionfetch), .ZN(n841) );
  IOA21D1BWP12T U2090 ( .A1(n1760), .A2(DEC_RF_offset_a[10]), .B(n1711), .ZN(
        n786) );
  IOA21D1BWP12T U2091 ( .A1(n1760), .A2(DEC_RF_offset_a[12]), .B(n1711), .ZN(
        n784) );
  IOA21D1BWP12T U2092 ( .A1(n1760), .A2(DEC_RF_offset_a[9]), .B(n1711), .ZN(
        n787) );
  IOA21D1BWP12T U2093 ( .A1(n1760), .A2(DEC_RF_offset_a[15]), .B(n1711), .ZN(
        n781) );
  IOA21D1BWP12T U2094 ( .A1(n1760), .A2(DEC_RF_offset_a[14]), .B(n1711), .ZN(
        n782) );
  IOA21D1BWP12T U2095 ( .A1(n1760), .A2(DEC_RF_offset_a[8]), .B(n1711), .ZN(
        n788) );
  OAI22D0BWP12T U2096 ( .A1(n1714), .A2(n1747), .B1(n1713), .B2(n1712), .ZN(
        n1716) );
  NR2D1BWP12T U2097 ( .A1(n1716), .A2(n1715), .ZN(n1717) );
  MOAI22D0BWP12T U2098 ( .A1(n1761), .A2(n1717), .B1(n1760), .B2(
        DEC_RF_offset_b[0]), .ZN(n853) );
  OAI211D0BWP12T U2099 ( .A1(n1746), .A2(n1720), .B(n1719), .C(n1718), .ZN(
        n1721) );
  IAO21D0BWP12T U2100 ( .A1(n1723), .A2(n1722), .B(n1721), .ZN(n1724) );
  MOAI22D0BWP12T U2101 ( .A1(n1724), .A2(n1761), .B1(n1760), .B2(
        DEC_RF_alu_write_to_reg[1]), .ZN(n805) );
  IOA21D1BWP12T U2102 ( .A1(n1760), .A2(DEC_RF_memory_write_to_reg_enable), 
        .B(n1725), .ZN(n811) );
  AOI21D0BWP12T U2103 ( .A1(n1728), .A2(n1727), .B(n1726), .ZN(n1734) );
  AOI31D0BWP12T U2104 ( .A1(n1731), .A2(n1756), .A3(n1730), .B(n1729), .ZN(
        n1733) );
  ND4D0BWP12T U2105 ( .A1(n1735), .A2(n1734), .A3(n1733), .A4(n1732), .ZN(
        n1752) );
  OAI211D0BWP12T U2106 ( .A1(n1739), .A2(n1738), .B(n1737), .C(n1736), .ZN(
        n1742) );
  TPOAI31D0BWP12T U2107 ( .A1(n1752), .A2(n1742), .A3(n1741), .B(n1740), .ZN(
        n1743) );
  IOA21D1BWP12T U2108 ( .A1(DEC_ALU_alu_opcode[4]), .A2(n1760), .B(n1743), 
        .ZN(n828) );
  AOI21D0BWP12T U2109 ( .A1(n1746), .A2(n1745), .B(n1744), .ZN(n1750) );
  OAI22D0BWP12T U2110 ( .A1(n1750), .A2(n1749), .B1(n1748), .B2(n1747), .ZN(
        n1751) );
  AOI211D0BWP12T U2111 ( .A1(n1754), .A2(n1753), .B(n1752), .C(n1751), .ZN(
        n1755) );
  TPOAI21D0BWP12T U2112 ( .A1(n1757), .A2(n1756), .B(n1755), .ZN(n1758) );
  TPAOI31D0BWP12T U2113 ( .A1(irdecode_inst1_next_step_1_), .A2(n1759), .A3(
        n1785), .B(n1758), .ZN(n1762) );
  MOAI22D0BWP12T U2114 ( .A1(n1762), .A2(n1761), .B1(n1760), .B2(
        DEC_ALU_alu_opcode[0]), .ZN(n831) );
  CKND0BWP12T U2115 ( .I(RF_ALU_operand_b[25]), .ZN(n1765) );
  INVD1BWP12T U2116 ( .I(n1763), .ZN(n1764) );
  AOI22D0BWP12T U2117 ( .A1(n1040), .A2(RF_ALU_operand_b[17]), .B1(n1039), 
        .B2(RF_ALU_operand_b[1]), .ZN(n1767) );
  IND3D1BWP12T U2118 ( .A1(n1768), .B1(n1767), .B2(n1766), .ZN(
        RF_ALU_operand_b_modified[25]) );
endmodule

