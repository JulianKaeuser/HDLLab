
module memory_interface_simple ( clock, reset, interface_cpu_sign_extend, 
        interface_cpu_word_type, interface_cpu_load_request, 
        interface_cpu_store_request, interface_cpu_address_in, 
        interface_cpu_data_in, from_mem_data_out, interface_cpu_read_finished, 
        interface_cpu_write_finished, interface_cpu_data_out, to_mem_address, 
        to_mem_data_in, to_mem_read_enable, to_mem_write_enable, to_mem_enable
 );
  input [1:0] interface_cpu_word_type;
  input [12:0] interface_cpu_address_in;
  input [31:0] interface_cpu_data_in;
  input [15:0] from_mem_data_out;
  output [31:0] interface_cpu_data_out;
  output [11:0] to_mem_address;
  output [15:0] to_mem_data_in;
  input clock, reset, interface_cpu_sign_extend, interface_cpu_load_request,
         interface_cpu_store_request;
  output interface_cpu_read_finished, interface_cpu_write_finished,
         to_mem_read_enable, to_mem_write_enable, to_mem_enable;
  wire   sign_extend, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76,
         N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90,
         N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N183, N184, N185, N186, N187, N188, N189, N190, N191,
         N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202,
         N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, n351,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796;
  wire   [5:0] state;
  wire   [15:0] tmp_value_1;
  wire   [15:0] tmp_value_2;
  wire   [31:0] cpu_data_in;
  wire   [12:1] cpu_address_in;

  DFQD1BWP12T to_mem_write_enable_reg ( .D(N212), .CP(clock), .Q(
        to_mem_write_enable) );
  DFQD1BWP12T interface_cpu_read_finished_reg ( .D(N72), .CP(clock), .Q(
        interface_cpu_read_finished) );
  DFQD1BWP12T interface_cpu_write_finished_reg ( .D(N73), .CP(clock), .Q(
        interface_cpu_write_finished) );
  DFQD1BWP12T tmp_value_1_reg_15_ ( .D(n428), .CP(clock), .Q(tmp_value_1[15])
         );
  DFQD1BWP12T tmp_value_1_reg_14_ ( .D(n427), .CP(clock), .Q(tmp_value_1[14])
         );
  DFQD1BWP12T tmp_value_1_reg_13_ ( .D(n426), .CP(clock), .Q(tmp_value_1[13])
         );
  DFQD1BWP12T tmp_value_1_reg_12_ ( .D(n425), .CP(clock), .Q(tmp_value_1[12])
         );
  DFQD1BWP12T tmp_value_1_reg_11_ ( .D(n424), .CP(clock), .Q(tmp_value_1[11])
         );
  DFQD1BWP12T tmp_value_1_reg_10_ ( .D(n423), .CP(clock), .Q(tmp_value_1[10])
         );
  DFQD1BWP12T tmp_value_1_reg_9_ ( .D(n422), .CP(clock), .Q(tmp_value_1[9]) );
  DFQD1BWP12T tmp_value_1_reg_8_ ( .D(n421), .CP(clock), .Q(tmp_value_1[8]) );
  DFQD1BWP12T tmp_value_1_reg_7_ ( .D(n420), .CP(clock), .Q(tmp_value_1[7]) );
  DFQD1BWP12T interface_cpu_data_out_reg_7_ ( .D(N81), .CP(clock), .Q(
        interface_cpu_data_out[7]) );
  DFQD1BWP12T tmp_value_1_reg_6_ ( .D(n419), .CP(clock), .Q(tmp_value_1[6]) );
  DFQD1BWP12T interface_cpu_data_out_reg_6_ ( .D(N80), .CP(clock), .Q(
        interface_cpu_data_out[6]) );
  DFQD1BWP12T tmp_value_1_reg_5_ ( .D(n418), .CP(clock), .Q(tmp_value_1[5]) );
  DFQD1BWP12T interface_cpu_data_out_reg_5_ ( .D(N79), .CP(clock), .Q(
        interface_cpu_data_out[5]) );
  DFQD1BWP12T tmp_value_1_reg_4_ ( .D(n417), .CP(clock), .Q(tmp_value_1[4]) );
  DFQD1BWP12T interface_cpu_data_out_reg_4_ ( .D(N78), .CP(clock), .Q(
        interface_cpu_data_out[4]) );
  DFQD1BWP12T tmp_value_1_reg_3_ ( .D(n416), .CP(clock), .Q(tmp_value_1[3]) );
  DFQD1BWP12T interface_cpu_data_out_reg_3_ ( .D(N77), .CP(clock), .Q(
        interface_cpu_data_out[3]) );
  DFQD1BWP12T tmp_value_1_reg_2_ ( .D(n415), .CP(clock), .Q(tmp_value_1[2]) );
  DFQD1BWP12T interface_cpu_data_out_reg_2_ ( .D(N76), .CP(clock), .Q(
        interface_cpu_data_out[2]) );
  DFQD1BWP12T tmp_value_1_reg_1_ ( .D(n414), .CP(clock), .Q(tmp_value_1[1]) );
  DFQD1BWP12T interface_cpu_data_out_reg_1_ ( .D(N75), .CP(clock), .Q(
        interface_cpu_data_out[1]) );
  DFQD1BWP12T tmp_value_1_reg_0_ ( .D(n413), .CP(clock), .Q(tmp_value_1[0]) );
  DFQD1BWP12T interface_cpu_data_out_reg_0_ ( .D(N74), .CP(clock), .Q(
        interface_cpu_data_out[0]) );
  DFQD1BWP12T tmp_value_2_reg_15_ ( .D(n412), .CP(clock), .Q(tmp_value_2[15])
         );
  DFQD1BWP12T tmp_value_2_reg_14_ ( .D(n411), .CP(clock), .Q(tmp_value_2[14])
         );
  DFQD1BWP12T tmp_value_2_reg_13_ ( .D(n410), .CP(clock), .Q(tmp_value_2[13])
         );
  DFQD1BWP12T tmp_value_2_reg_12_ ( .D(n409), .CP(clock), .Q(tmp_value_2[12])
         );
  DFQD1BWP12T tmp_value_2_reg_11_ ( .D(n408), .CP(clock), .Q(tmp_value_2[11])
         );
  DFQD1BWP12T tmp_value_2_reg_10_ ( .D(n407), .CP(clock), .Q(tmp_value_2[10])
         );
  DFQD1BWP12T tmp_value_2_reg_9_ ( .D(n406), .CP(clock), .Q(tmp_value_2[9]) );
  DFQD1BWP12T tmp_value_2_reg_8_ ( .D(n405), .CP(clock), .Q(tmp_value_2[8]) );
  DFQD1BWP12T tmp_value_2_reg_7_ ( .D(n404), .CP(clock), .Q(tmp_value_2[7]) );
  DFQD1BWP12T tmp_value_2_reg_6_ ( .D(n403), .CP(clock), .Q(tmp_value_2[6]) );
  DFQD1BWP12T tmp_value_2_reg_5_ ( .D(n402), .CP(clock), .Q(tmp_value_2[5]) );
  DFQD1BWP12T tmp_value_2_reg_4_ ( .D(n401), .CP(clock), .Q(tmp_value_2[4]) );
  DFQD1BWP12T tmp_value_2_reg_3_ ( .D(n400), .CP(clock), .Q(tmp_value_2[3]) );
  DFQD1BWP12T tmp_value_2_reg_2_ ( .D(n399), .CP(clock), .Q(tmp_value_2[2]) );
  DFQD1BWP12T tmp_value_2_reg_1_ ( .D(n398), .CP(clock), .Q(tmp_value_2[1]) );
  DFQD1BWP12T tmp_value_2_reg_0_ ( .D(n397), .CP(clock), .Q(tmp_value_2[0]) );
  DFQD1BWP12T cpu_data_in_reg_31_ ( .D(n396), .CP(clock), .Q(cpu_data_in[31])
         );
  DFQD1BWP12T cpu_data_in_reg_30_ ( .D(n395), .CP(clock), .Q(cpu_data_in[30])
         );
  DFQD1BWP12T cpu_data_in_reg_29_ ( .D(n394), .CP(clock), .Q(cpu_data_in[29])
         );
  DFQD1BWP12T cpu_data_in_reg_28_ ( .D(n393), .CP(clock), .Q(cpu_data_in[28])
         );
  DFQD1BWP12T cpu_data_in_reg_27_ ( .D(n392), .CP(clock), .Q(cpu_data_in[27])
         );
  DFQD1BWP12T cpu_data_in_reg_26_ ( .D(n391), .CP(clock), .Q(cpu_data_in[26])
         );
  DFQD1BWP12T cpu_data_in_reg_25_ ( .D(n390), .CP(clock), .Q(cpu_data_in[25])
         );
  DFQD1BWP12T cpu_data_in_reg_24_ ( .D(n389), .CP(clock), .Q(cpu_data_in[24])
         );
  DFQD1BWP12T cpu_data_in_reg_23_ ( .D(n388), .CP(clock), .Q(cpu_data_in[23])
         );
  DFQD1BWP12T cpu_data_in_reg_22_ ( .D(n387), .CP(clock), .Q(cpu_data_in[22])
         );
  DFQD1BWP12T cpu_data_in_reg_21_ ( .D(n386), .CP(clock), .Q(cpu_data_in[21])
         );
  DFQD1BWP12T cpu_data_in_reg_20_ ( .D(n385), .CP(clock), .Q(cpu_data_in[20])
         );
  DFQD1BWP12T cpu_data_in_reg_19_ ( .D(n384), .CP(clock), .Q(cpu_data_in[19])
         );
  DFQD1BWP12T cpu_data_in_reg_18_ ( .D(n383), .CP(clock), .Q(cpu_data_in[18])
         );
  DFQD1BWP12T cpu_data_in_reg_17_ ( .D(n382), .CP(clock), .Q(cpu_data_in[17])
         );
  DFQD1BWP12T cpu_data_in_reg_16_ ( .D(n381), .CP(clock), .Q(cpu_data_in[16])
         );
  DFQD1BWP12T cpu_data_in_reg_15_ ( .D(n380), .CP(clock), .Q(cpu_data_in[15])
         );
  DFQD1BWP12T cpu_data_in_reg_14_ ( .D(n379), .CP(clock), .Q(cpu_data_in[14])
         );
  DFQD1BWP12T cpu_data_in_reg_13_ ( .D(n378), .CP(clock), .Q(cpu_data_in[13])
         );
  DFQD1BWP12T cpu_data_in_reg_12_ ( .D(n377), .CP(clock), .Q(cpu_data_in[12])
         );
  DFQD1BWP12T cpu_data_in_reg_11_ ( .D(n376), .CP(clock), .Q(cpu_data_in[11])
         );
  DFQD1BWP12T cpu_data_in_reg_10_ ( .D(n375), .CP(clock), .Q(cpu_data_in[10])
         );
  DFQD1BWP12T cpu_data_in_reg_9_ ( .D(n374), .CP(clock), .Q(cpu_data_in[9]) );
  DFQD1BWP12T cpu_data_in_reg_8_ ( .D(n373), .CP(clock), .Q(cpu_data_in[8]) );
  DFQD1BWP12T cpu_data_in_reg_7_ ( .D(n372), .CP(clock), .Q(cpu_data_in[7]) );
  DFQD1BWP12T cpu_data_in_reg_6_ ( .D(n371), .CP(clock), .Q(cpu_data_in[6]) );
  DFQD1BWP12T cpu_data_in_reg_5_ ( .D(n370), .CP(clock), .Q(cpu_data_in[5]) );
  DFQD1BWP12T cpu_data_in_reg_4_ ( .D(n369), .CP(clock), .Q(cpu_data_in[4]) );
  DFQD1BWP12T cpu_data_in_reg_3_ ( .D(n368), .CP(clock), .Q(cpu_data_in[3]) );
  DFQD1BWP12T cpu_data_in_reg_2_ ( .D(n367), .CP(clock), .Q(cpu_data_in[2]) );
  DFQD1BWP12T cpu_data_in_reg_1_ ( .D(n366), .CP(clock), .Q(cpu_data_in[1]) );
  DFQD1BWP12T cpu_data_in_reg_0_ ( .D(n365), .CP(clock), .Q(cpu_data_in[0]) );
  DFQD1BWP12T cpu_address_in_reg_12_ ( .D(n364), .CP(clock), .Q(
        cpu_address_in[12]) );
  DFQD1BWP12T cpu_address_in_reg_11_ ( .D(n363), .CP(clock), .Q(
        cpu_address_in[11]) );
  DFQD1BWP12T cpu_address_in_reg_10_ ( .D(n362), .CP(clock), .Q(
        cpu_address_in[10]) );
  DFQD1BWP12T cpu_address_in_reg_9_ ( .D(n361), .CP(clock), .Q(
        cpu_address_in[9]) );
  DFQD1BWP12T cpu_address_in_reg_8_ ( .D(n360), .CP(clock), .Q(
        cpu_address_in[8]) );
  DFQD1BWP12T cpu_address_in_reg_7_ ( .D(n359), .CP(clock), .Q(
        cpu_address_in[7]) );
  DFQD1BWP12T cpu_address_in_reg_6_ ( .D(n358), .CP(clock), .Q(
        cpu_address_in[6]) );
  DFQD1BWP12T cpu_address_in_reg_5_ ( .D(n357), .CP(clock), .Q(
        cpu_address_in[5]) );
  DFQD1BWP12T cpu_address_in_reg_4_ ( .D(n356), .CP(clock), .Q(
        cpu_address_in[4]) );
  DFQD1BWP12T cpu_address_in_reg_3_ ( .D(n355), .CP(clock), .Q(
        cpu_address_in[3]) );
  DFQD1BWP12T cpu_address_in_reg_2_ ( .D(n354), .CP(clock), .Q(
        cpu_address_in[2]) );
  DFQD1BWP12T cpu_address_in_reg_1_ ( .D(n353), .CP(clock), .Q(
        cpu_address_in[1]) );
  DFQD1BWP12T sign_extend_reg ( .D(n351), .CP(clock), .Q(sign_extend) );
  DFQD1BWP12T interface_cpu_data_out_reg_8_ ( .D(N82), .CP(clock), .Q(
        interface_cpu_data_out[8]) );
  DFQD1BWP12T interface_cpu_data_out_reg_9_ ( .D(N83), .CP(clock), .Q(
        interface_cpu_data_out[9]) );
  DFQD1BWP12T interface_cpu_data_out_reg_10_ ( .D(N84), .CP(clock), .Q(
        interface_cpu_data_out[10]) );
  DFQD1BWP12T interface_cpu_data_out_reg_11_ ( .D(N85), .CP(clock), .Q(
        interface_cpu_data_out[11]) );
  DFQD1BWP12T interface_cpu_data_out_reg_12_ ( .D(N86), .CP(clock), .Q(
        interface_cpu_data_out[12]) );
  DFQD1BWP12T interface_cpu_data_out_reg_13_ ( .D(N87), .CP(clock), .Q(
        interface_cpu_data_out[13]) );
  DFQD1BWP12T interface_cpu_data_out_reg_14_ ( .D(N88), .CP(clock), .Q(
        interface_cpu_data_out[14]) );
  DFQD1BWP12T interface_cpu_data_out_reg_15_ ( .D(N89), .CP(clock), .Q(
        interface_cpu_data_out[15]) );
  DFQD1BWP12T interface_cpu_data_out_reg_16_ ( .D(N90), .CP(clock), .Q(
        interface_cpu_data_out[16]) );
  DFQD1BWP12T interface_cpu_data_out_reg_17_ ( .D(N91), .CP(clock), .Q(
        interface_cpu_data_out[17]) );
  DFQD1BWP12T interface_cpu_data_out_reg_18_ ( .D(N92), .CP(clock), .Q(
        interface_cpu_data_out[18]) );
  DFQD1BWP12T interface_cpu_data_out_reg_19_ ( .D(N93), .CP(clock), .Q(
        interface_cpu_data_out[19]) );
  DFQD1BWP12T interface_cpu_data_out_reg_20_ ( .D(N94), .CP(clock), .Q(
        interface_cpu_data_out[20]) );
  DFQD1BWP12T interface_cpu_data_out_reg_21_ ( .D(N95), .CP(clock), .Q(
        interface_cpu_data_out[21]) );
  DFQD1BWP12T interface_cpu_data_out_reg_22_ ( .D(N96), .CP(clock), .Q(
        interface_cpu_data_out[22]) );
  DFQD1BWP12T interface_cpu_data_out_reg_23_ ( .D(N97), .CP(clock), .Q(
        interface_cpu_data_out[23]) );
  DFQD1BWP12T interface_cpu_data_out_reg_24_ ( .D(N98), .CP(clock), .Q(
        interface_cpu_data_out[24]) );
  DFQD1BWP12T interface_cpu_data_out_reg_25_ ( .D(N99), .CP(clock), .Q(
        interface_cpu_data_out[25]) );
  DFQD1BWP12T interface_cpu_data_out_reg_26_ ( .D(N100), .CP(clock), .Q(
        interface_cpu_data_out[26]) );
  DFQD1BWP12T interface_cpu_data_out_reg_27_ ( .D(N101), .CP(clock), .Q(
        interface_cpu_data_out[27]) );
  DFQD1BWP12T interface_cpu_data_out_reg_28_ ( .D(N102), .CP(clock), .Q(
        interface_cpu_data_out[28]) );
  DFQD1BWP12T interface_cpu_data_out_reg_29_ ( .D(N103), .CP(clock), .Q(
        interface_cpu_data_out[29]) );
  DFQD1BWP12T interface_cpu_data_out_reg_30_ ( .D(N104), .CP(clock), .Q(
        interface_cpu_data_out[30]) );
  DFQD1BWP12T interface_cpu_data_out_reg_31_ ( .D(N105), .CP(clock), .Q(
        interface_cpu_data_out[31]) );
  DFQD1BWP12T to_mem_address_reg_10_ ( .D(N193), .CP(clock), .Q(
        to_mem_address[10]) );
  DFQD1BWP12T to_mem_address_reg_9_ ( .D(N192), .CP(clock), .Q(
        to_mem_address[9]) );
  DFQD1BWP12T to_mem_address_reg_8_ ( .D(N191), .CP(clock), .Q(
        to_mem_address[8]) );
  DFQD1BWP12T to_mem_address_reg_7_ ( .D(N190), .CP(clock), .Q(
        to_mem_address[7]) );
  DFQD1BWP12T to_mem_address_reg_6_ ( .D(N189), .CP(clock), .Q(
        to_mem_address[6]) );
  DFQD1BWP12T to_mem_address_reg_5_ ( .D(N188), .CP(clock), .Q(
        to_mem_address[5]) );
  DFQD1BWP12T to_mem_address_reg_4_ ( .D(N187), .CP(clock), .Q(
        to_mem_address[4]) );
  DFQD1BWP12T to_mem_address_reg_3_ ( .D(N186), .CP(clock), .Q(
        to_mem_address[3]) );
  DFQD1BWP12T to_mem_address_reg_2_ ( .D(N185), .CP(clock), .Q(
        to_mem_address[2]) );
  DFQD1BWP12T to_mem_address_reg_1_ ( .D(N184), .CP(clock), .Q(
        to_mem_address[1]) );
  DFQD1BWP12T to_mem_address_reg_0_ ( .D(N183), .CP(clock), .Q(
        to_mem_address[0]) );
  DFQD1BWP12T to_mem_data_in_reg_15_ ( .D(N210), .CP(clock), .Q(
        to_mem_data_in[15]) );
  DFQD1BWP12T to_mem_data_in_reg_14_ ( .D(N209), .CP(clock), .Q(
        to_mem_data_in[14]) );
  DFQD1BWP12T to_mem_data_in_reg_13_ ( .D(N208), .CP(clock), .Q(
        to_mem_data_in[13]) );
  DFQD1BWP12T to_mem_data_in_reg_12_ ( .D(N207), .CP(clock), .Q(
        to_mem_data_in[12]) );
  DFQD1BWP12T to_mem_data_in_reg_11_ ( .D(N206), .CP(clock), .Q(
        to_mem_data_in[11]) );
  DFQD1BWP12T to_mem_data_in_reg_10_ ( .D(N205), .CP(clock), .Q(
        to_mem_data_in[10]) );
  DFQD1BWP12T to_mem_data_in_reg_9_ ( .D(N204), .CP(clock), .Q(
        to_mem_data_in[9]) );
  DFQD1BWP12T to_mem_data_in_reg_8_ ( .D(N203), .CP(clock), .Q(
        to_mem_data_in[8]) );
  DFQD1BWP12T to_mem_data_in_reg_7_ ( .D(N202), .CP(clock), .Q(
        to_mem_data_in[7]) );
  DFQD1BWP12T to_mem_data_in_reg_6_ ( .D(N201), .CP(clock), .Q(
        to_mem_data_in[6]) );
  DFQD1BWP12T to_mem_data_in_reg_5_ ( .D(N200), .CP(clock), .Q(
        to_mem_data_in[5]) );
  DFQD1BWP12T to_mem_data_in_reg_4_ ( .D(N199), .CP(clock), .Q(
        to_mem_data_in[4]) );
  DFQD1BWP12T to_mem_data_in_reg_3_ ( .D(N198), .CP(clock), .Q(
        to_mem_data_in[3]) );
  DFQD1BWP12T to_mem_data_in_reg_2_ ( .D(N197), .CP(clock), .Q(
        to_mem_data_in[2]) );
  DFQD1BWP12T to_mem_data_in_reg_1_ ( .D(N196), .CP(clock), .Q(
        to_mem_data_in[1]) );
  DFQD1BWP12T to_mem_data_in_reg_0_ ( .D(N195), .CP(clock), .Q(
        to_mem_data_in[0]) );
  DFQD1BWP12T to_mem_read_enable_reg ( .D(N211), .CP(clock), .Q(
        to_mem_read_enable) );
  DFQD1BWP12T to_mem_address_reg_11_ ( .D(N194), .CP(clock), .Q(
        to_mem_address[11]) );
  DFQD2BWP12T state_reg_3_ ( .D(N69), .CP(clock), .Q(state[3]) );
  DFQD2BWP12T state_reg_5_ ( .D(N71), .CP(clock), .Q(state[5]) );
  DFQD1BWP12T state_reg_0_ ( .D(N66), .CP(clock), .Q(state[0]) );
  DFQD1BWP12T state_reg_2_ ( .D(N68), .CP(clock), .Q(state[2]) );
  DFQD1BWP12T state_reg_1_ ( .D(N67), .CP(clock), .Q(state[1]) );
  DFQD1BWP12T state_reg_4_ ( .D(N70), .CP(clock), .Q(state[4]) );
  TIELBWP12T U503 ( .ZN(n432) );
  INVD1BWP12T U504 ( .I(n432), .ZN(to_mem_enable) );
  IND2D1BWP12T U505 ( .A1(state[4]), .B1(state[5]), .ZN(n592) );
  HA1D1BWP12T U506 ( .A(n692), .B(cpu_address_in[10]), .CO(n694), .S(n693) );
  NR2D1BWP12T U507 ( .A1(n686), .A2(reset), .ZN(n687) );
  INVD1BWP12T U508 ( .I(n684), .ZN(n517) );
  AOI21D1BWP12T U509 ( .A1(n474), .A2(n497), .B(reset), .ZN(n626) );
  AN2D0BWP12T U510 ( .A1(state[2]), .A2(state[3]), .Z(n509) );
  MOAI22D0BWP12T U511 ( .A1(n758), .A2(n737), .B1(tmp_value_2[3]), .B2(n752), 
        .ZN(n433) );
  AO22D0BWP12T U512 ( .A1(n753), .A2(cpu_data_in[19]), .B1(
        from_mem_data_out[3]), .B2(n754), .Z(n434) );
  AOI211D0BWP12T U513 ( .A1(n760), .A2(cpu_data_in[3]), .B(n433), .C(n434), 
        .ZN(n435) );
  MOAI22D0BWP12T U514 ( .A1(reset), .A2(n435), .B1(cpu_data_in[27]), .B2(n761), 
        .ZN(N198) );
  IND3D0BWP12T U515 ( .A1(interface_cpu_load_request), .B1(n524), .B2(
        interface_cpu_store_request), .ZN(n673) );
  AN3D0BWP12T U516 ( .A1(n562), .A2(n563), .A3(n763), .Z(n768) );
  MOAI22D0BWP12T U517 ( .A1(n758), .A2(n738), .B1(tmp_value_2[4]), .B2(n752), 
        .ZN(n436) );
  AO22D0BWP12T U518 ( .A1(n753), .A2(cpu_data_in[20]), .B1(
        from_mem_data_out[4]), .B2(n754), .Z(n437) );
  AOI211D0BWP12T U519 ( .A1(n760), .A2(cpu_data_in[4]), .B(n436), .C(n437), 
        .ZN(n438) );
  MOAI22D0BWP12T U520 ( .A1(reset), .A2(n438), .B1(cpu_data_in[28]), .B2(n761), 
        .ZN(N199) );
  NR3D0BWP12T U521 ( .A1(state[3]), .A2(state[5]), .A3(n507), .ZN(n618) );
  MOAI22D0BWP12T U522 ( .A1(n758), .A2(n739), .B1(tmp_value_2[5]), .B2(n752), 
        .ZN(n439) );
  AO22D0BWP12T U523 ( .A1(n753), .A2(cpu_data_in[21]), .B1(
        from_mem_data_out[5]), .B2(n754), .Z(n440) );
  AOI211D0BWP12T U524 ( .A1(n760), .A2(cpu_data_in[5]), .B(n439), .C(n440), 
        .ZN(n441) );
  MOAI22D0BWP12T U525 ( .A1(reset), .A2(n441), .B1(cpu_data_in[29]), .B2(n761), 
        .ZN(N200) );
  NR3D0BWP12T U526 ( .A1(reset), .A2(n562), .A3(n666), .ZN(n625) );
  INR4D0BWP12T U527 ( .A1(n551), .B1(n678), .B2(n618), .B3(n560), .ZN(n589) );
  MOAI22D0BWP12T U528 ( .A1(n758), .A2(n745), .B1(tmp_value_2[6]), .B2(n752), 
        .ZN(n442) );
  AO22D0BWP12T U529 ( .A1(n753), .A2(cpu_data_in[22]), .B1(
        from_mem_data_out[6]), .B2(n754), .Z(n443) );
  AOI211D0BWP12T U530 ( .A1(n760), .A2(cpu_data_in[6]), .B(n442), .C(n443), 
        .ZN(n444) );
  MOAI22D0BWP12T U531 ( .A1(reset), .A2(n444), .B1(cpu_data_in[30]), .B2(n761), 
        .ZN(N201) );
  NR3D0BWP12T U532 ( .A1(state[5]), .A2(n562), .A3(n507), .ZN(n495) );
  MOAI22D0BWP12T U533 ( .A1(n758), .A2(n751), .B1(tmp_value_2[7]), .B2(n752), 
        .ZN(n445) );
  AO22D0BWP12T U534 ( .A1(n753), .A2(cpu_data_in[23]), .B1(
        from_mem_data_out[7]), .B2(n754), .Z(n446) );
  AOI211D0BWP12T U535 ( .A1(n760), .A2(cpu_data_in[7]), .B(n445), .C(n446), 
        .ZN(n447) );
  MOAI22D0BWP12T U536 ( .A1(reset), .A2(n447), .B1(cpu_data_in[31]), .B2(n761), 
        .ZN(N202) );
  AO211D0BWP12T U537 ( .A1(n763), .A2(n679), .B(n654), .C(n625), .Z(n448) );
  OAI21D0BWP12T U538 ( .A1(n682), .A2(n448), .B(sign_extend), .ZN(n449) );
  IOA21D0BWP12T U539 ( .A1(interface_cpu_sign_extend), .A2(n626), .B(n449), 
        .ZN(n351) );
  AN2D1BWP12T U540 ( .A1(n453), .A2(n512), .Z(n450) );
  ND2D1BWP12T U541 ( .A1(state[0]), .A2(state[1]), .ZN(n465) );
  INVD1BWP12T U542 ( .I(n465), .ZN(n463) );
  NR2D1BWP12T U543 ( .A1(state[2]), .A2(state[4]), .ZN(n452) );
  ND2D1BWP12T U544 ( .A1(n463), .A2(n452), .ZN(n507) );
  INR2D1BWP12T U545 ( .A1(state[5]), .B1(n507), .ZN(n563) );
  ND2D1BWP12T U546 ( .A1(n563), .A2(state[3]), .ZN(n698) );
  NR2D1BWP12T U547 ( .A1(state[2]), .A2(state[3]), .ZN(n531) );
  INR2D1BWP12T U548 ( .A1(n531), .B1(n592), .ZN(n665) );
  INR2D2BWP12T U549 ( .A1(state[1]), .B1(state[0]), .ZN(n613) );
  ND2D1BWP12T U550 ( .A1(n665), .A2(n613), .ZN(n544) );
  NR2D1BWP12T U551 ( .A1(state[1]), .A2(state[0]), .ZN(n511) );
  INR2D1BWP12T U552 ( .A1(n511), .B1(n592), .ZN(n478) );
  IND2D1BWP12T U553 ( .A1(state[2]), .B1(state[3]), .ZN(n482) );
  INVD1BWP12T U554 ( .I(n482), .ZN(n669) );
  ND2D1BWP12T U555 ( .A1(n478), .A2(n669), .ZN(n773) );
  ND3D1BWP12T U556 ( .A1(n698), .A2(n544), .A3(n773), .ZN(n595) );
  IND2D1BWP12T U557 ( .A1(state[5]), .B1(state[4]), .ZN(n483) );
  INVD1BWP12T U558 ( .I(n483), .ZN(n451) );
  ND2D1BWP12T U559 ( .A1(n613), .A2(n451), .ZN(n603) );
  INR2D2BWP12T U560 ( .A1(n669), .B1(n603), .ZN(n486) );
  INVD1BWP12T U561 ( .I(n613), .ZN(n476) );
  TPNR3D3BWP12T U562 ( .A1(n482), .A2(n476), .A3(n592), .ZN(n753) );
  NR2D2BWP12T U563 ( .A1(n486), .A2(n753), .ZN(n731) );
  ND2D1BWP12T U564 ( .A1(n451), .A2(n511), .ZN(n616) );
  INVD1BWP12T U565 ( .I(state[3]), .ZN(n562) );
  INR2D2BWP12T U566 ( .A1(state[0]), .B1(state[1]), .ZN(n619) );
  CKND2D1BWP12T U567 ( .A1(n619), .A2(n452), .ZN(n454) );
  INR2XD0BWP12T U568 ( .A1(n562), .B1(n454), .ZN(n525) );
  ND2D1BWP12T U569 ( .A1(n525), .A2(state[5]), .ZN(n545) );
  TPNR2D1BWP12T U570 ( .A1(n483), .A2(n465), .ZN(n602) );
  CKND2D1BWP12T U571 ( .A1(n602), .A2(n531), .ZN(n548) );
  OA211D1BWP12T U572 ( .A1(n616), .A2(n482), .B(n545), .C(n548), .Z(n774) );
  IND2D1BWP12T U573 ( .A1(state[3]), .B1(state[2]), .ZN(n660) );
  NR2D1BWP12T U574 ( .A1(n592), .A2(n660), .ZN(n475) );
  ND2D1BWP12T U575 ( .A1(n475), .A2(n619), .ZN(n453) );
  INVD1BWP12T U576 ( .I(n619), .ZN(n490) );
  NR2D1BWP12T U577 ( .A1(n490), .A2(n483), .ZN(n456) );
  CKND2D1BWP12T U578 ( .A1(n456), .A2(n509), .ZN(n512) );
  ND3D2BWP12T U579 ( .A1(n731), .A2(n774), .A3(n450), .ZN(n538) );
  INVD1BWP12T U580 ( .I(reset), .ZN(n763) );
  OA21XD0BWP12T U581 ( .A1(n538), .A2(n595), .B(n763), .Z(n696) );
  INVD1BWP12T U582 ( .I(n454), .ZN(n455) );
  ND2D1BWP12T U583 ( .A1(n455), .A2(state[3]), .ZN(n457) );
  INR2D1BWP12T U584 ( .A1(state[5]), .B1(n457), .ZN(n594) );
  INVD1BWP12T U585 ( .I(n456), .ZN(n504) );
  INR2D1BWP12T U586 ( .A1(n669), .B1(n504), .ZN(n606) );
  NR2D1BWP12T U587 ( .A1(n594), .A2(n606), .ZN(n729) );
  INVD1BWP12T U588 ( .I(n457), .ZN(n458) );
  INVD1BWP12T U589 ( .I(state[5]), .ZN(n530) );
  ND2D1BWP12T U590 ( .A1(n458), .A2(n530), .ZN(n730) );
  ND2D1BWP12T U591 ( .A1(n729), .A2(n730), .ZN(n760) );
  INVD1BWP12T U592 ( .I(n660), .ZN(n462) );
  INR2D1BWP12T U593 ( .A1(n462), .B1(n504), .ZN(n605) );
  INVD1BWP12T U594 ( .I(n478), .ZN(n467) );
  INR2D1BWP12T U595 ( .A1(n462), .B1(n467), .ZN(n459) );
  NR2D1BWP12T U596 ( .A1(n605), .A2(n459), .ZN(n758) );
  NR2D1BWP12T U597 ( .A1(state[4]), .A2(state[5]), .ZN(n629) );
  CKND1BWP12T U598 ( .I(n509), .ZN(n503) );
  INR2D1BWP12T U599 ( .A1(n629), .B1(n503), .ZN(n464) );
  ND2D1BWP12T U600 ( .A1(n464), .A2(n619), .ZN(n736) );
  ND2D1BWP12T U601 ( .A1(n758), .A2(n736), .ZN(n727) );
  NR2D1BWP12T U602 ( .A1(n760), .A2(n727), .ZN(n489) );
  ND2D1BWP12T U603 ( .A1(n511), .A2(n629), .ZN(n666) );
  NR2D1BWP12T U604 ( .A1(n666), .A2(n660), .ZN(n460) );
  AOI21D1BWP12T U605 ( .A1(n525), .A2(n530), .B(n460), .ZN(n621) );
  INVD1BWP12T U606 ( .I(n616), .ZN(n668) );
  ND2D0BWP12T U607 ( .A1(n668), .A2(n509), .ZN(n600) );
  ND2D1BWP12T U608 ( .A1(state[4]), .A2(state[5]), .ZN(n461) );
  ND3D1BWP12T U609 ( .A1(n463), .A2(n462), .A3(n461), .ZN(n627) );
  TPND2D0BWP12T U610 ( .A1(n600), .A2(n627), .ZN(n468) );
  CKND0BWP12T U611 ( .I(n531), .ZN(n614) );
  CKND0BWP12T U612 ( .I(n464), .ZN(n466) );
  OAI22D1BWP12T U613 ( .A1(n603), .A2(n614), .B1(n466), .B2(n465), .ZN(n547)
         );
  NR2D1BWP12T U614 ( .A1(n467), .A2(n614), .ZN(n542) );
  NR4D0BWP12T U615 ( .A1(n468), .A2(n547), .A3(n542), .A4(n495), .ZN(n469) );
  AOI31D1BWP12T U616 ( .A1(n489), .A2(n621), .A3(n469), .B(reset), .ZN(n695)
         );
  AO22XD1BWP12T U617 ( .A1(n470), .A2(n696), .B1(n695), .B2(cpu_address_in[7]), 
        .Z(N189) );
  HA1D2BWP12T U618 ( .A(n471), .B(cpu_address_in[6]), .CO(n584), .S(n472) );
  AO22XD1BWP12T U619 ( .A1(n472), .A2(n696), .B1(n695), .B2(cpu_address_in[6]), 
        .Z(N188) );
  NR2D1BWP12T U620 ( .A1(n503), .A2(n511), .ZN(n473) );
  OAI21D0BWP12T U621 ( .A1(n473), .A2(state[4]), .B(state[5]), .ZN(n474) );
  INR2D1BWP12T U622 ( .A1(n531), .B1(n666), .ZN(n524) );
  INVD1BWP12T U623 ( .I(n524), .ZN(n497) );
  AOI21D1BWP12T U624 ( .A1(n629), .A2(state[3]), .B(n475), .ZN(n477) );
  OAI22D1BWP12T U625 ( .A1(n477), .A2(n476), .B1(n660), .B2(n603), .ZN(n481)
         );
  ND2D1BWP12T U626 ( .A1(n602), .A2(n669), .ZN(n480) );
  ND2D1BWP12T U627 ( .A1(n478), .A2(n509), .ZN(n479) );
  ND2D1BWP12T U628 ( .A1(n480), .A2(n479), .ZN(n765) );
  NR2D1BWP12T U629 ( .A1(n481), .A2(n765), .ZN(n508) );
  INR2D1BWP12T U630 ( .A1(n763), .B1(n508), .ZN(N73) );
  INVD1BWP12T U631 ( .I(n511), .ZN(n661) );
  AOI211D1BWP12T U632 ( .A1(n483), .A2(n592), .B(n661), .C(n482), .ZN(n631) );
  INR3D0BWP12T U633 ( .A1(n627), .B1(n495), .B2(n631), .ZN(n549) );
  INVD1BWP12T U634 ( .I(n625), .ZN(n484) );
  OAI21D1BWP12T U635 ( .A1(n549), .A2(reset), .B(n484), .ZN(n485) );
  NR2D1BWP12T U636 ( .A1(N73), .A2(n485), .ZN(n492) );
  INVD1BWP12T U637 ( .I(n753), .ZN(n488) );
  INVD1BWP12T U638 ( .I(n486), .ZN(n487) );
  ND2D1BWP12T U639 ( .A1(n698), .A2(n487), .ZN(n752) );
  INR2D1BWP12T U640 ( .A1(n488), .B1(n752), .ZN(n767) );
  CKND2D1BWP12T U641 ( .A1(n489), .A2(n767), .ZN(n491) );
  NR4D0BWP12T U642 ( .A1(n490), .A2(reset), .A3(n660), .A4(n592), .ZN(n761) );
  AO21D1BWP12T U643 ( .A1(n491), .A2(n763), .B(n761), .Z(N212) );
  INR2D1BWP12T U644 ( .A1(n492), .B1(N212), .ZN(n684) );
  AO22XD1BWP12T U645 ( .A1(interface_cpu_data_in[2]), .A2(n626), .B1(
        cpu_data_in[2]), .B2(n517), .Z(n367) );
  AO22XD1BWP12T U646 ( .A1(interface_cpu_data_in[3]), .A2(n626), .B1(
        cpu_data_in[3]), .B2(n517), .Z(n368) );
  AO22XD1BWP12T U647 ( .A1(interface_cpu_data_in[16]), .A2(n626), .B1(
        cpu_data_in[16]), .B2(n517), .Z(n381) );
  AO22XD1BWP12T U648 ( .A1(interface_cpu_data_in[4]), .A2(n626), .B1(
        cpu_data_in[4]), .B2(n517), .Z(n369) );
  AO22XD1BWP12T U649 ( .A1(interface_cpu_data_in[31]), .A2(n626), .B1(
        cpu_data_in[31]), .B2(n517), .Z(n396) );
  INVD1BWP12T U650 ( .I(interface_cpu_word_type[1]), .ZN(n597) );
  ND2D0BWP12T U651 ( .A1(interface_cpu_address_in[0]), .A2(n597), .ZN(n632) );
  INVD1BWP12T U652 ( .I(interface_cpu_word_type[0]), .ZN(n494) );
  CKND2D1BWP12T U653 ( .A1(interface_cpu_word_type[0]), .A2(n597), .ZN(n674)
         );
  CKND0BWP12T U654 ( .I(n674), .ZN(n493) );
  AOI21D1BWP12T U655 ( .A1(n632), .A2(n494), .B(n493), .ZN(n502) );
  INVD1BWP12T U656 ( .I(n548), .ZN(n496) );
  NR2D0BWP12T U657 ( .A1(n496), .A2(n495), .ZN(n501) );
  INR2D1BWP12T U658 ( .A1(n629), .B1(n660), .ZN(n620) );
  CKND0BWP12T U659 ( .I(state[1]), .ZN(n499) );
  INR2XD0BWP12T U660 ( .A1(interface_cpu_load_request), .B1(n497), .ZN(n591)
         );
  ND2D1BWP12T U661 ( .A1(n591), .A2(n597), .ZN(n513) );
  TPNR2D0BWP12T U662 ( .A1(n513), .A2(interface_cpu_word_type[0]), .ZN(n498)
         );
  AOI22D0BWP12T U663 ( .A1(n620), .A2(n499), .B1(n498), .B2(
        interface_cpu_address_in[0]), .ZN(n500) );
  OAI211D1BWP12T U664 ( .A1(n502), .A2(n673), .B(n501), .C(n500), .ZN(n515) );
  NR2D1BWP12T U665 ( .A1(n503), .A2(state[5]), .ZN(n510) );
  CKND2D1BWP12T U666 ( .A1(n620), .A2(n613), .ZN(n565) );
  INR2D1BWP12T U667 ( .A1(n531), .B1(n504), .ZN(n636) );
  INR2D1BWP12T U668 ( .A1(n565), .B1(n636), .ZN(n623) );
  INVD1BWP12T U669 ( .I(n623), .ZN(n560) );
  NR2D1BWP12T U670 ( .A1(n616), .A2(n660), .ZN(n624) );
  CKND0BWP12T U671 ( .I(n624), .ZN(n506) );
  CKND2D0BWP12T U672 ( .A1(n563), .A2(n562), .ZN(n505) );
  ND2D1BWP12T U673 ( .A1(n506), .A2(n505), .ZN(n678) );
  ND2D1BWP12T U674 ( .A1(n602), .A2(n509), .ZN(n551) );
  CKND2D0BWP12T U675 ( .A1(n589), .A2(n508), .ZN(n598) );
  INR2D1BWP12T U676 ( .A1(n509), .B1(n603), .ZN(n771) );
  AOI211D0BWP12T U677 ( .A1(n511), .A2(n510), .B(n598), .C(n771), .ZN(n677) );
  NR2XD0BWP12T U678 ( .A1(interface_cpu_address_in[0]), .A2(n597), .ZN(n533)
         );
  INVD1BWP12T U679 ( .I(n512), .ZN(n543) );
  AOI31D1BWP12T U680 ( .A1(n591), .A2(n494), .A3(n533), .B(n543), .ZN(n609) );
  NR2D1BWP12T U681 ( .A1(interface_cpu_address_in[0]), .A2(n513), .ZN(n667) );
  CKND2D1BWP12T U682 ( .A1(n667), .A2(interface_cpu_word_type[0]), .ZN(n514)
         );
  ND4D1BWP12T U683 ( .A1(n677), .A2(n609), .A3(n698), .A4(n514), .ZN(n633) );
  TPOAI31D0BWP12T U684 ( .A1(n727), .A2(n515), .A3(n633), .B(n763), .ZN(n516)
         );
  CKND0BWP12T U685 ( .I(n761), .ZN(n536) );
  CKND2D1BWP12T U686 ( .A1(n516), .A2(n536), .ZN(N68) );
  AO22XD1BWP12T U687 ( .A1(interface_cpu_data_in[8]), .A2(n626), .B1(
        cpu_data_in[8]), .B2(n517), .Z(n373) );
  AO22XD1BWP12T U688 ( .A1(interface_cpu_data_in[1]), .A2(n626), .B1(
        cpu_data_in[1]), .B2(n517), .Z(n366) );
  AO22XD1BWP12T U689 ( .A1(interface_cpu_data_in[19]), .A2(n626), .B1(
        cpu_data_in[19]), .B2(n517), .Z(n384) );
  AO22XD1BWP12T U690 ( .A1(interface_cpu_data_in[18]), .A2(n626), .B1(
        cpu_data_in[18]), .B2(n517), .Z(n383) );
  AO22XD1BWP12T U691 ( .A1(interface_cpu_data_in[29]), .A2(n626), .B1(
        cpu_data_in[29]), .B2(n517), .Z(n394) );
  AO22XD1BWP12T U692 ( .A1(interface_cpu_data_in[24]), .A2(n626), .B1(
        cpu_data_in[24]), .B2(n517), .Z(n389) );
  AO22XD1BWP12T U693 ( .A1(interface_cpu_data_in[26]), .A2(n626), .B1(
        cpu_data_in[26]), .B2(n517), .Z(n391) );
  AO22XD1BWP12T U694 ( .A1(interface_cpu_data_in[28]), .A2(n626), .B1(
        cpu_data_in[28]), .B2(n517), .Z(n393) );
  AO22XD1BWP12T U695 ( .A1(interface_cpu_data_in[23]), .A2(n626), .B1(
        cpu_data_in[23]), .B2(n517), .Z(n388) );
  AO22XD1BWP12T U696 ( .A1(interface_cpu_data_in[27]), .A2(n626), .B1(
        cpu_data_in[27]), .B2(n517), .Z(n392) );
  AO22XD1BWP12T U697 ( .A1(interface_cpu_data_in[22]), .A2(n626), .B1(
        cpu_data_in[22]), .B2(n517), .Z(n387) );
  AO22XD1BWP12T U698 ( .A1(interface_cpu_data_in[12]), .A2(n626), .B1(
        cpu_data_in[12]), .B2(n517), .Z(n377) );
  AO22XD1BWP12T U699 ( .A1(interface_cpu_data_in[5]), .A2(n626), .B1(
        cpu_data_in[5]), .B2(n517), .Z(n370) );
  AO22XD1BWP12T U700 ( .A1(interface_cpu_data_in[15]), .A2(n626), .B1(
        cpu_data_in[15]), .B2(n517), .Z(n380) );
  AO22XD1BWP12T U701 ( .A1(interface_cpu_data_in[25]), .A2(n626), .B1(
        cpu_data_in[25]), .B2(n517), .Z(n390) );
  AO22XD1BWP12T U702 ( .A1(interface_cpu_data_in[7]), .A2(n626), .B1(
        cpu_data_in[7]), .B2(n517), .Z(n372) );
  AO22XD1BWP12T U703 ( .A1(interface_cpu_data_in[30]), .A2(n626), .B1(
        cpu_data_in[30]), .B2(n517), .Z(n395) );
  AO22XD1BWP12T U704 ( .A1(interface_cpu_data_in[0]), .A2(n626), .B1(
        cpu_data_in[0]), .B2(n517), .Z(n365) );
  AO22XD1BWP12T U705 ( .A1(interface_cpu_data_in[20]), .A2(n626), .B1(
        cpu_data_in[20]), .B2(n517), .Z(n385) );
  AO22XD1BWP12T U706 ( .A1(interface_cpu_data_in[13]), .A2(n626), .B1(
        cpu_data_in[13]), .B2(n517), .Z(n378) );
  AO22XD1BWP12T U707 ( .A1(interface_cpu_data_in[14]), .A2(n626), .B1(
        cpu_data_in[14]), .B2(n517), .Z(n379) );
  AO22XD1BWP12T U708 ( .A1(interface_cpu_data_in[9]), .A2(n626), .B1(
        cpu_data_in[9]), .B2(n517), .Z(n374) );
  AO22XD1BWP12T U709 ( .A1(interface_cpu_data_in[21]), .A2(n626), .B1(
        cpu_data_in[21]), .B2(n517), .Z(n386) );
  AO22XD1BWP12T U710 ( .A1(interface_cpu_data_in[17]), .A2(n626), .B1(
        cpu_data_in[17]), .B2(n517), .Z(n382) );
  AO22XD1BWP12T U711 ( .A1(interface_cpu_data_in[6]), .A2(n626), .B1(
        cpu_data_in[6]), .B2(n517), .Z(n371) );
  AO22XD1BWP12T U712 ( .A1(interface_cpu_data_in[11]), .A2(n626), .B1(
        cpu_data_in[11]), .B2(n517), .Z(n376) );
  AO22XD1BWP12T U713 ( .A1(interface_cpu_data_in[10]), .A2(n626), .B1(
        cpu_data_in[10]), .B2(n517), .Z(n375) );
  HA1D2BWP12T U714 ( .A(n518), .B(cpu_address_in[5]), .CO(n471), .S(n519) );
  AO22XD1BWP12T U715 ( .A1(n519), .A2(n696), .B1(n695), .B2(cpu_address_in[5]), 
        .Z(N187) );
  HA1D2BWP12T U716 ( .A(n520), .B(cpu_address_in[4]), .CO(n518), .S(n521) );
  AO22D0BWP12T U717 ( .A1(n521), .A2(n696), .B1(n695), .B2(cpu_address_in[4]), 
        .Z(N186) );
  HA1D2BWP12T U718 ( .A(n522), .B(cpu_address_in[3]), .CO(n520), .S(n523) );
  AO22D0BWP12T U719 ( .A1(n523), .A2(n696), .B1(n695), .B2(cpu_address_in[3]), 
        .Z(N185) );
  ND2D1BWP12T U720 ( .A1(n729), .A2(n544), .ZN(n764) );
  AOI31D0BWP12T U721 ( .A1(n524), .A2(interface_cpu_store_request), .A3(
        interface_cpu_address_in[0]), .B(n591), .ZN(n528) );
  NR2D0BWP12T U722 ( .A1(n543), .A2(n771), .ZN(n527) );
  AOI211D1BWP12T U723 ( .A1(n629), .A2(n619), .B(n605), .C(n525), .ZN(n526) );
  OAI211D1BWP12T U724 ( .A1(n674), .A2(n528), .B(n527), .C(n526), .ZN(n535) );
  INVD1BWP12T U725 ( .I(n731), .ZN(n529) );
  AOI31D0BWP12T U726 ( .A1(n531), .A2(n613), .A3(n530), .B(n529), .ZN(n532) );
  OA31D1BWP12T U727 ( .A1(n533), .A2(interface_cpu_word_type[0]), .A3(n673), 
        .B(n532), .Z(n676) );
  INVD1BWP12T U728 ( .I(n676), .ZN(n534) );
  OAI31D0BWP12T U729 ( .A1(n764), .A2(n535), .A3(n534), .B(n763), .ZN(n537) );
  CKND2D1BWP12T U730 ( .A1(n537), .A2(n536), .ZN(N67) );
  HA1D0BWP12T U731 ( .A(n538), .B(cpu_address_in[1]), .CO(n540), .S(n539) );
  AO22D0BWP12T U732 ( .A1(n539), .A2(n696), .B1(n695), .B2(cpu_address_in[1]), 
        .Z(N183) );
  FA1D2BWP12T U733 ( .A(n595), .B(cpu_address_in[2]), .CI(n540), .CO(n522), 
        .S(n541) );
  AO22D0BWP12T U734 ( .A1(n541), .A2(n696), .B1(n695), .B2(cpu_address_in[2]), 
        .Z(N184) );
  NR2D0BWP12T U735 ( .A1(n543), .A2(n542), .ZN(n546) );
  ND4D1BWP12T U736 ( .A1(n546), .A2(n600), .A3(n545), .A4(n544), .ZN(n680) );
  INVD1BWP12T U737 ( .I(n547), .ZN(n601) );
  CKND2D1BWP12T U738 ( .A1(n601), .A2(n548), .ZN(n679) );
  NR2D0BWP12T U739 ( .A1(n680), .A2(n679), .ZN(n550) );
  AOI31D0BWP12T U740 ( .A1(n550), .A2(n621), .A3(n549), .B(reset), .ZN(N211)
         );
  AOI222D0BWP12T U741 ( .A1(n678), .A2(tmp_value_1[3]), .B1(
        from_mem_data_out[3]), .B2(n618), .C1(n560), .C2(from_mem_data_out[11]), .ZN(n552) );
  INVD1BWP12T U742 ( .I(tmp_value_1[11]), .ZN(n728) );
  INR2D1BWP12T U743 ( .A1(n763), .B1(n551), .ZN(n681) );
  INVD1BWP12T U744 ( .I(n681), .ZN(n777) );
  OAI22D0BWP12T U745 ( .A1(n552), .A2(reset), .B1(n728), .B2(n777), .ZN(N77)
         );
  AOI222D0BWP12T U746 ( .A1(n678), .A2(tmp_value_1[0]), .B1(
        from_mem_data_out[0]), .B2(n618), .C1(n560), .C2(from_mem_data_out[8]), 
        .ZN(n553) );
  INVD1BWP12T U747 ( .I(tmp_value_1[8]), .ZN(n699) );
  OAI22D0BWP12T U748 ( .A1(n553), .A2(reset), .B1(n699), .B2(n777), .ZN(N74)
         );
  AOI222D0BWP12T U749 ( .A1(n678), .A2(tmp_value_1[1]), .B1(
        from_mem_data_out[1]), .B2(n618), .C1(n560), .C2(from_mem_data_out[9]), 
        .ZN(n554) );
  INVD1BWP12T U750 ( .I(tmp_value_1[9]), .ZN(n715) );
  OAI22D0BWP12T U751 ( .A1(n554), .A2(reset), .B1(n715), .B2(n777), .ZN(N75)
         );
  INVD1BWP12T U752 ( .I(from_mem_data_out[15]), .ZN(n795) );
  ND2D1BWP12T U753 ( .A1(n618), .A2(from_mem_data_out[7]), .ZN(n564) );
  OAI21D0BWP12T U754 ( .A1(n623), .A2(n795), .B(n564), .ZN(n555) );
  AOI21D0BWP12T U755 ( .A1(tmp_value_1[7]), .A2(n678), .B(n555), .ZN(n556) );
  INVD1BWP12T U756 ( .I(tmp_value_1[15]), .ZN(n703) );
  OAI22D0BWP12T U757 ( .A1(n556), .A2(reset), .B1(n703), .B2(n777), .ZN(N81)
         );
  AOI222D0BWP12T U758 ( .A1(n678), .A2(tmp_value_1[5]), .B1(
        from_mem_data_out[5]), .B2(n618), .C1(n560), .C2(from_mem_data_out[13]), .ZN(n557) );
  INVD1BWP12T U759 ( .I(tmp_value_1[13]), .ZN(n711) );
  OAI22D0BWP12T U760 ( .A1(n557), .A2(reset), .B1(n711), .B2(n777), .ZN(N79)
         );
  AOI222D0BWP12T U761 ( .A1(n678), .A2(tmp_value_1[6]), .B1(
        from_mem_data_out[6]), .B2(n618), .C1(n560), .C2(from_mem_data_out[14]), .ZN(n558) );
  INVD1BWP12T U762 ( .I(tmp_value_1[14]), .ZN(n707) );
  OAI22D0BWP12T U763 ( .A1(n558), .A2(reset), .B1(n707), .B2(n777), .ZN(N80)
         );
  AOI222D0BWP12T U764 ( .A1(n678), .A2(tmp_value_1[4]), .B1(
        from_mem_data_out[4]), .B2(n618), .C1(n560), .C2(from_mem_data_out[12]), .ZN(n559) );
  INVD1BWP12T U765 ( .I(tmp_value_1[12]), .ZN(n719) );
  OAI22D0BWP12T U766 ( .A1(n559), .A2(reset), .B1(n719), .B2(n777), .ZN(N78)
         );
  AOI222D0BWP12T U767 ( .A1(n678), .A2(tmp_value_1[2]), .B1(
        from_mem_data_out[2]), .B2(n618), .C1(n560), .C2(from_mem_data_out[10]), .ZN(n561) );
  INVD1BWP12T U768 ( .I(tmp_value_1[10]), .ZN(n723) );
  OAI22D0BWP12T U769 ( .A1(n561), .A2(reset), .B1(n723), .B2(n777), .ZN(N76)
         );
  AOI22D0BWP12T U770 ( .A1(n768), .A2(from_mem_data_out[8]), .B1(n681), .B2(
        from_mem_data_out[0]), .ZN(n567) );
  OA21D1BWP12T U771 ( .A1(n565), .A2(n795), .B(n564), .Z(n638) );
  TPAOI22D0BWP12T U772 ( .A1(n636), .A2(from_mem_data_out[7]), .B1(n624), .B2(
        from_mem_data_out[15]), .ZN(n566) );
  ND2D1BWP12T U773 ( .A1(sign_extend), .A2(n763), .ZN(n637) );
  AO21D1BWP12T U774 ( .A1(n638), .A2(n566), .B(n637), .Z(n582) );
  TPND2D0BWP12T U775 ( .A1(n567), .A2(n582), .ZN(N98) );
  AOI22D0BWP12T U776 ( .A1(n768), .A2(from_mem_data_out[13]), .B1(n681), .B2(
        from_mem_data_out[5]), .ZN(n568) );
  TPND2D0BWP12T U777 ( .A1(n568), .A2(n582), .ZN(N103) );
  AOI22D0BWP12T U778 ( .A1(n768), .A2(from_mem_data_out[11]), .B1(n681), .B2(
        from_mem_data_out[3]), .ZN(n569) );
  TPND2D0BWP12T U779 ( .A1(n569), .A2(n582), .ZN(N101) );
  AOI22D0BWP12T U780 ( .A1(n768), .A2(from_mem_data_out[14]), .B1(n681), .B2(
        from_mem_data_out[6]), .ZN(n570) );
  TPND2D0BWP12T U781 ( .A1(n570), .A2(n582), .ZN(N104) );
  AOI22D0BWP12T U782 ( .A1(n768), .A2(from_mem_data_out[12]), .B1(n681), .B2(
        from_mem_data_out[4]), .ZN(n571) );
  TPND2D0BWP12T U783 ( .A1(n571), .A2(n582), .ZN(N102) );
  AOI22D0BWP12T U784 ( .A1(n768), .A2(from_mem_data_out[9]), .B1(n681), .B2(
        from_mem_data_out[1]), .ZN(n572) );
  TPND2D0BWP12T U785 ( .A1(n572), .A2(n582), .ZN(N99) );
  AOI22D0BWP12T U786 ( .A1(n768), .A2(from_mem_data_out[10]), .B1(n681), .B2(
        from_mem_data_out[2]), .ZN(n573) );
  TPND2D0BWP12T U787 ( .A1(n573), .A2(n582), .ZN(N100) );
  AOI22D0BWP12T U788 ( .A1(n768), .A2(tmp_value_2[7]), .B1(n681), .B2(
        from_mem_data_out[15]), .ZN(n574) );
  TPND2D0BWP12T U789 ( .A1(n574), .A2(n582), .ZN(N97) );
  AOI22D0BWP12T U790 ( .A1(n768), .A2(tmp_value_2[6]), .B1(n681), .B2(
        from_mem_data_out[14]), .ZN(n575) );
  TPND2D0BWP12T U791 ( .A1(n575), .A2(n582), .ZN(N96) );
  AOI22D0BWP12T U792 ( .A1(n768), .A2(from_mem_data_out[15]), .B1(n681), .B2(
        from_mem_data_out[7]), .ZN(n576) );
  TPND2D0BWP12T U793 ( .A1(n576), .A2(n582), .ZN(N105) );
  AOI22D0BWP12T U794 ( .A1(n768), .A2(tmp_value_2[5]), .B1(n681), .B2(
        from_mem_data_out[13]), .ZN(n577) );
  TPND2D0BWP12T U795 ( .A1(n577), .A2(n582), .ZN(N95) );
  AOI22D0BWP12T U796 ( .A1(n768), .A2(tmp_value_2[4]), .B1(n681), .B2(
        from_mem_data_out[12]), .ZN(n578) );
  TPND2D0BWP12T U797 ( .A1(n578), .A2(n582), .ZN(N94) );
  AOI22D0BWP12T U798 ( .A1(n768), .A2(tmp_value_2[3]), .B1(n681), .B2(
        from_mem_data_out[11]), .ZN(n579) );
  TPND2D0BWP12T U799 ( .A1(n579), .A2(n582), .ZN(N93) );
  AOI22D0BWP12T U800 ( .A1(n768), .A2(tmp_value_2[2]), .B1(n681), .B2(
        from_mem_data_out[10]), .ZN(n580) );
  TPND2D0BWP12T U801 ( .A1(n580), .A2(n582), .ZN(N92) );
  AOI22D0BWP12T U802 ( .A1(n768), .A2(tmp_value_2[1]), .B1(n681), .B2(
        from_mem_data_out[9]), .ZN(n581) );
  TPND2D0BWP12T U803 ( .A1(n581), .A2(n582), .ZN(N91) );
  AOI22D0BWP12T U804 ( .A1(n768), .A2(tmp_value_2[0]), .B1(n681), .B2(
        from_mem_data_out[8]), .ZN(n583) );
  CKND2D1BWP12T U805 ( .A1(n583), .A2(n582), .ZN(N90) );
  INVD1BWP12T U806 ( .I(cpu_address_in[12]), .ZN(n588) );
  CKND0BWP12T U807 ( .I(n695), .ZN(n587) );
  HA1D2BWP12T U808 ( .A(n584), .B(cpu_address_in[7]), .CO(n688), .S(n470) );
  XOR2D2BWP12T U809 ( .A1(cpu_address_in[12]), .A2(n585), .Z(n586) );
  MOAI22D1BWP12T U810 ( .A1(n588), .A2(n587), .B1(n586), .B2(n696), .ZN(N194)
         );
  NR2D1BWP12T U811 ( .A1(reset), .A2(n589), .ZN(N72) );
  INVD1BWP12T U812 ( .I(n673), .ZN(n590) );
  AOI21D1BWP12T U813 ( .A1(n591), .A2(interface_cpu_address_in[0]), .B(n590), 
        .ZN(n611) );
  NR2D1BWP12T U814 ( .A1(n592), .A2(state[3]), .ZN(n593) );
  NR4D0BWP12T U815 ( .A1(n595), .A2(n594), .A3(n753), .A4(n593), .ZN(n596) );
  TPOAI31D0BWP12T U816 ( .A1(interface_cpu_word_type[0]), .A2(n611), .A3(n597), 
        .B(n596), .ZN(n599) );
  OA21D1BWP12T U817 ( .A1(n599), .A2(n598), .B(n763), .Z(N71) );
  OAI211D0BWP12T U818 ( .A1(state[2]), .A2(n616), .B(n601), .C(n600), .ZN(n608) );
  INVD1BWP12T U819 ( .I(n602), .ZN(n604) );
  MUX2ND0BWP12T U820 ( .I0(n604), .I1(n603), .S(state[3]), .ZN(n607) );
  NR4D0BWP12T U821 ( .A1(n608), .A2(n607), .A3(n606), .A4(n605), .ZN(n610) );
  OA211D1BWP12T U822 ( .A1(n674), .A2(n611), .B(n610), .C(n609), .Z(n612) );
  NR2D1BWP12T U823 ( .A1(n612), .A2(reset), .ZN(N70) );
  CKND2D0BWP12T U824 ( .A1(n613), .A2(n629), .ZN(n615) );
  AOI21D1BWP12T U825 ( .A1(n616), .A2(n615), .B(n614), .ZN(n617) );
  AOI211D1BWP12T U826 ( .A1(n620), .A2(n619), .B(n618), .C(n617), .ZN(n622) );
  AOI31D1BWP12T U827 ( .A1(n623), .A2(n622), .A3(n621), .B(reset), .ZN(n682)
         );
  ND2D1BWP12T U828 ( .A1(n624), .A2(n763), .ZN(n775) );
  INVD1BWP12T U829 ( .I(n775), .ZN(n654) );
  CKND0BWP12T U830 ( .I(n627), .ZN(n628) );
  AOI21D1BWP12T U831 ( .A1(n629), .A2(n669), .B(n628), .ZN(n630) );
  IND4D1BWP12T U832 ( .A1(n631), .B1(n630), .B2(n731), .B3(n736), .ZN(n635) );
  OAI31D0BWP12T U833 ( .A1(n632), .A2(n673), .A3(interface_cpu_word_type[0]), 
        .B(n729), .ZN(n634) );
  OA31D1BWP12T U834 ( .A1(n635), .A2(n634), .A3(n633), .B(n763), .Z(N69) );
  INVD1BWP12T U835 ( .I(from_mem_data_out[5]), .ZN(n785) );
  ND2D1BWP12T U836 ( .A1(n636), .A2(n763), .ZN(n659) );
  AOI22D0BWP12T U837 ( .A1(n654), .A2(from_mem_data_out[13]), .B1(n768), .B2(
        tmp_value_2[13]), .ZN(n641) );
  OR2XD1BWP12T U838 ( .A1(n638), .A2(n637), .Z(n639) );
  INVD1BWP12T U839 ( .I(n639), .ZN(n656) );
  ND2D1BWP12T U840 ( .A1(n639), .A2(n777), .ZN(n655) );
  OAI21D0BWP12T U841 ( .A1(tmp_value_1[5]), .A2(n656), .B(n655), .ZN(n640) );
  OAI211D1BWP12T U842 ( .A1(n785), .A2(n659), .B(n641), .C(n640), .ZN(N87) );
  INVD1BWP12T U843 ( .I(from_mem_data_out[7]), .ZN(n781) );
  AOI22D0BWP12T U844 ( .A1(n654), .A2(from_mem_data_out[15]), .B1(n768), .B2(
        tmp_value_2[15]), .ZN(n643) );
  OAI21D0BWP12T U845 ( .A1(tmp_value_1[7]), .A2(n656), .B(n655), .ZN(n642) );
  OAI211D1BWP12T U846 ( .A1(n781), .A2(n659), .B(n643), .C(n642), .ZN(N89) );
  INVD1BWP12T U847 ( .I(from_mem_data_out[6]), .ZN(n782) );
  AOI22D0BWP12T U848 ( .A1(n654), .A2(from_mem_data_out[14]), .B1(n768), .B2(
        tmp_value_2[14]), .ZN(n645) );
  OAI21D0BWP12T U849 ( .A1(tmp_value_1[6]), .A2(n656), .B(n655), .ZN(n644) );
  OAI211D1BWP12T U850 ( .A1(n782), .A2(n659), .B(n645), .C(n644), .ZN(N88) );
  INVD1BWP12T U851 ( .I(from_mem_data_out[0]), .ZN(n779) );
  AOI22D0BWP12T U852 ( .A1(n654), .A2(from_mem_data_out[8]), .B1(n768), .B2(
        tmp_value_2[8]), .ZN(n647) );
  OAI21D0BWP12T U853 ( .A1(tmp_value_1[0]), .A2(n656), .B(n655), .ZN(n646) );
  OAI211D1BWP12T U854 ( .A1(n779), .A2(n659), .B(n647), .C(n646), .ZN(N82) );
  INVD1BWP12T U855 ( .I(from_mem_data_out[4]), .ZN(n784) );
  AOI22D0BWP12T U856 ( .A1(n654), .A2(from_mem_data_out[12]), .B1(n768), .B2(
        tmp_value_2[12]), .ZN(n649) );
  OAI21D0BWP12T U857 ( .A1(tmp_value_1[4]), .A2(n656), .B(n655), .ZN(n648) );
  OAI211D1BWP12T U858 ( .A1(n784), .A2(n659), .B(n649), .C(n648), .ZN(N86) );
  INVD1BWP12T U859 ( .I(from_mem_data_out[1]), .ZN(n783) );
  AOI22D0BWP12T U860 ( .A1(n654), .A2(from_mem_data_out[9]), .B1(n768), .B2(
        tmp_value_2[9]), .ZN(n651) );
  OAI21D0BWP12T U861 ( .A1(tmp_value_1[1]), .A2(n656), .B(n655), .ZN(n650) );
  OAI211D1BWP12T U862 ( .A1(n783), .A2(n659), .B(n651), .C(n650), .ZN(N83) );
  INVD1BWP12T U863 ( .I(from_mem_data_out[3]), .ZN(n780) );
  AOI22D0BWP12T U864 ( .A1(n654), .A2(from_mem_data_out[11]), .B1(n768), .B2(
        tmp_value_2[11]), .ZN(n653) );
  OAI21D0BWP12T U865 ( .A1(tmp_value_1[3]), .A2(n656), .B(n655), .ZN(n652) );
  OAI211D1BWP12T U866 ( .A1(n780), .A2(n659), .B(n653), .C(n652), .ZN(N85) );
  INVD1BWP12T U867 ( .I(from_mem_data_out[2]), .ZN(n786) );
  AOI22D0BWP12T U868 ( .A1(n654), .A2(from_mem_data_out[10]), .B1(n768), .B2(
        tmp_value_2[10]), .ZN(n658) );
  OAI21D0BWP12T U869 ( .A1(tmp_value_1[2]), .A2(n656), .B(n655), .ZN(n657) );
  OAI211D1BWP12T U870 ( .A1(n786), .A2(n659), .B(n658), .C(n657), .ZN(N84) );
  INVD1BWP12T U871 ( .I(state[0]), .ZN(n664) );
  INVD1BWP12T U872 ( .I(n773), .ZN(n663) );
  NR3D1BWP12T U873 ( .A1(n661), .A2(state[4]), .A3(n660), .ZN(n662) );
  AOI211D0BWP12T U874 ( .A1(n665), .A2(n664), .B(n663), .C(n662), .ZN(n672) );
  CKND0BWP12T U875 ( .I(n666), .ZN(n670) );
  AOI211D1BWP12T U876 ( .A1(n670), .A2(n669), .B(n668), .C(n667), .ZN(n671) );
  OA211D1BWP12T U877 ( .A1(n674), .A2(n673), .B(n672), .C(n671), .Z(n675) );
  AOI31D1BWP12T U878 ( .A1(n677), .A2(n676), .A3(n675), .B(reset), .ZN(N66) );
  NR4D0BWP12T U879 ( .A1(n680), .A2(n771), .A3(n679), .A4(n678), .ZN(n685) );
  NR2D1BWP12T U880 ( .A1(n682), .A2(n681), .ZN(n683) );
  OAI211D1BWP12T U881 ( .A1(reset), .A2(n685), .B(n684), .C(n683), .ZN(n686)
         );
  AO22D1BWP12T U882 ( .A1(n687), .A2(interface_cpu_address_in[8]), .B1(
        cpu_address_in[8]), .B2(n686), .Z(n360) );
  AO22D1BWP12T U883 ( .A1(n687), .A2(interface_cpu_address_in[4]), .B1(
        cpu_address_in[4]), .B2(n686), .Z(n356) );
  AO22D1BWP12T U884 ( .A1(n687), .A2(interface_cpu_address_in[2]), .B1(
        cpu_address_in[2]), .B2(n686), .Z(n354) );
  AO22D1BWP12T U885 ( .A1(n687), .A2(interface_cpu_address_in[10]), .B1(
        cpu_address_in[10]), .B2(n686), .Z(n362) );
  AO22D1BWP12T U886 ( .A1(n687), .A2(interface_cpu_address_in[1]), .B1(
        cpu_address_in[1]), .B2(n686), .Z(n353) );
  AO22D1BWP12T U887 ( .A1(n687), .A2(interface_cpu_address_in[6]), .B1(
        cpu_address_in[6]), .B2(n686), .Z(n358) );
  AO22D1BWP12T U888 ( .A1(n687), .A2(interface_cpu_address_in[5]), .B1(
        cpu_address_in[5]), .B2(n686), .Z(n357) );
  AO22D1BWP12T U889 ( .A1(n687), .A2(interface_cpu_address_in[11]), .B1(
        cpu_address_in[11]), .B2(n686), .Z(n363) );
  AO22D1BWP12T U890 ( .A1(n687), .A2(interface_cpu_address_in[7]), .B1(
        cpu_address_in[7]), .B2(n686), .Z(n359) );
  AO22D1BWP12T U891 ( .A1(n687), .A2(interface_cpu_address_in[3]), .B1(
        cpu_address_in[3]), .B2(n686), .Z(n355) );
  AO22D1BWP12T U892 ( .A1(n687), .A2(interface_cpu_address_in[9]), .B1(
        cpu_address_in[9]), .B2(n686), .Z(n361) );
  AO22D1BWP12T U893 ( .A1(n687), .A2(interface_cpu_address_in[12]), .B1(
        cpu_address_in[12]), .B2(n686), .Z(n364) );
  HA1D2BWP12T U894 ( .A(n688), .B(cpu_address_in[8]), .CO(n690), .S(n689) );
  AO22D1BWP12T U895 ( .A1(n689), .A2(n696), .B1(n695), .B2(cpu_address_in[8]), 
        .Z(N190) );
  HA1D2BWP12T U896 ( .A(n690), .B(cpu_address_in[9]), .CO(n692), .S(n691) );
  AO22D1BWP12T U897 ( .A1(n691), .A2(n696), .B1(n695), .B2(cpu_address_in[9]), 
        .Z(N191) );
  AO22D1BWP12T U898 ( .A1(n693), .A2(n696), .B1(n695), .B2(cpu_address_in[10]), 
        .Z(N192) );
  HA1D1BWP12T U899 ( .A(n694), .B(cpu_address_in[11]), .CO(n585), .S(n697) );
  AO22D1BWP12T U900 ( .A1(n697), .A2(n696), .B1(n695), .B2(cpu_address_in[11]), 
        .Z(N193) );
  INVD1BWP12T U901 ( .I(n698), .ZN(n734) );
  MOAI22D0BWP12T U902 ( .A1(n729), .A2(n699), .B1(n727), .B2(cpu_data_in[0]), 
        .ZN(n701) );
  CKND1BWP12T U903 ( .I(cpu_data_in[8]), .ZN(n742) );
  INVD1BWP12T U904 ( .I(from_mem_data_out[8]), .ZN(n788) );
  OAI22D1BWP12T U905 ( .A1(n731), .A2(n742), .B1(n730), .B2(n788), .ZN(n700)
         );
  AOI211XD0BWP12T U906 ( .A1(n734), .A2(cpu_data_in[24]), .B(n701), .C(n700), 
        .ZN(n702) );
  MOAI22D0BWP12T U907 ( .A1(n702), .A2(reset), .B1(cpu_data_in[16]), .B2(n761), 
        .ZN(N203) );
  MOAI22D0BWP12T U908 ( .A1(n729), .A2(n703), .B1(n727), .B2(cpu_data_in[7]), 
        .ZN(n705) );
  CKND1BWP12T U909 ( .I(cpu_data_in[15]), .ZN(n751) );
  OAI22D1BWP12T U910 ( .A1(n731), .A2(n751), .B1(n730), .B2(n795), .ZN(n704)
         );
  AOI211XD0BWP12T U911 ( .A1(n734), .A2(cpu_data_in[31]), .B(n705), .C(n704), 
        .ZN(n706) );
  MOAI22D0BWP12T U912 ( .A1(n706), .A2(reset), .B1(cpu_data_in[23]), .B2(n761), 
        .ZN(N210) );
  MOAI22D0BWP12T U913 ( .A1(n729), .A2(n707), .B1(n727), .B2(cpu_data_in[6]), 
        .ZN(n709) );
  CKND1BWP12T U914 ( .I(cpu_data_in[14]), .ZN(n745) );
  INVD1BWP12T U915 ( .I(from_mem_data_out[14]), .ZN(n792) );
  OAI22D1BWP12T U916 ( .A1(n731), .A2(n745), .B1(n730), .B2(n792), .ZN(n708)
         );
  AOI211XD0BWP12T U917 ( .A1(n734), .A2(cpu_data_in[30]), .B(n709), .C(n708), 
        .ZN(n710) );
  MOAI22D0BWP12T U918 ( .A1(n710), .A2(reset), .B1(cpu_data_in[22]), .B2(n761), 
        .ZN(N209) );
  MOAI22D0BWP12T U919 ( .A1(n729), .A2(n711), .B1(n727), .B2(cpu_data_in[5]), 
        .ZN(n713) );
  CKND1BWP12T U920 ( .I(cpu_data_in[13]), .ZN(n739) );
  INVD1BWP12T U921 ( .I(from_mem_data_out[13]), .ZN(n791) );
  OAI22D1BWP12T U922 ( .A1(n731), .A2(n739), .B1(n730), .B2(n791), .ZN(n712)
         );
  AOI211XD0BWP12T U923 ( .A1(n734), .A2(cpu_data_in[29]), .B(n713), .C(n712), 
        .ZN(n714) );
  MOAI22D0BWP12T U924 ( .A1(n714), .A2(reset), .B1(cpu_data_in[21]), .B2(n761), 
        .ZN(N208) );
  MOAI22D0BWP12T U925 ( .A1(n729), .A2(n715), .B1(n727), .B2(cpu_data_in[1]), 
        .ZN(n717) );
  CKND1BWP12T U926 ( .I(cpu_data_in[9]), .ZN(n757) );
  INVD1BWP12T U927 ( .I(from_mem_data_out[9]), .ZN(n790) );
  OAI22D1BWP12T U928 ( .A1(n731), .A2(n757), .B1(n730), .B2(n790), .ZN(n716)
         );
  AOI211XD0BWP12T U929 ( .A1(n734), .A2(cpu_data_in[25]), .B(n717), .C(n716), 
        .ZN(n718) );
  MOAI22D0BWP12T U930 ( .A1(n718), .A2(reset), .B1(cpu_data_in[17]), .B2(n761), 
        .ZN(N204) );
  MOAI22D0BWP12T U931 ( .A1(n729), .A2(n719), .B1(n727), .B2(cpu_data_in[4]), 
        .ZN(n721) );
  CKND1BWP12T U932 ( .I(cpu_data_in[12]), .ZN(n738) );
  INVD1BWP12T U933 ( .I(from_mem_data_out[12]), .ZN(n789) );
  OAI22D1BWP12T U934 ( .A1(n731), .A2(n738), .B1(n730), .B2(n789), .ZN(n720)
         );
  AOI211XD0BWP12T U935 ( .A1(n734), .A2(cpu_data_in[28]), .B(n721), .C(n720), 
        .ZN(n722) );
  MOAI22D0BWP12T U936 ( .A1(n722), .A2(reset), .B1(cpu_data_in[20]), .B2(n761), 
        .ZN(N207) );
  MOAI22D0BWP12T U937 ( .A1(n729), .A2(n723), .B1(n727), .B2(cpu_data_in[2]), 
        .ZN(n725) );
  CKND1BWP12T U938 ( .I(cpu_data_in[10]), .ZN(n748) );
  INVD1BWP12T U939 ( .I(from_mem_data_out[10]), .ZN(n787) );
  OAI22D1BWP12T U940 ( .A1(n731), .A2(n748), .B1(n730), .B2(n787), .ZN(n724)
         );
  AOI211XD0BWP12T U941 ( .A1(n734), .A2(cpu_data_in[26]), .B(n725), .C(n724), 
        .ZN(n726) );
  MOAI22D0BWP12T U942 ( .A1(n726), .A2(reset), .B1(cpu_data_in[18]), .B2(n761), 
        .ZN(N205) );
  MOAI22D0BWP12T U943 ( .A1(n729), .A2(n728), .B1(n727), .B2(cpu_data_in[3]), 
        .ZN(n733) );
  CKND1BWP12T U944 ( .I(cpu_data_in[11]), .ZN(n737) );
  INVD1BWP12T U945 ( .I(from_mem_data_out[11]), .ZN(n793) );
  OAI22D1BWP12T U946 ( .A1(n731), .A2(n737), .B1(n730), .B2(n793), .ZN(n732)
         );
  AOI211XD0BWP12T U947 ( .A1(n734), .A2(cpu_data_in[27]), .B(n733), .C(n732), 
        .ZN(n735) );
  MOAI22D0BWP12T U948 ( .A1(n735), .A2(reset), .B1(cpu_data_in[19]), .B2(n761), 
        .ZN(N206) );
  INVD1BWP12T U949 ( .I(n736), .ZN(n754) );
  CKND2D0BWP12T U950 ( .A1(n752), .A2(tmp_value_2[0]), .ZN(n741) );
  AOI22D0BWP12T U951 ( .A1(n754), .A2(from_mem_data_out[0]), .B1(n753), .B2(
        cpu_data_in[16]), .ZN(n740) );
  OAI211D0BWP12T U952 ( .A1(n758), .A2(n742), .B(n741), .C(n740), .ZN(n743) );
  AOI21D0BWP12T U953 ( .A1(cpu_data_in[0]), .A2(n760), .B(n743), .ZN(n744) );
  MOAI22D0BWP12T U954 ( .A1(n744), .A2(reset), .B1(cpu_data_in[24]), .B2(n761), 
        .ZN(N195) );
  CKND2D0BWP12T U955 ( .A1(n752), .A2(tmp_value_2[2]), .ZN(n747) );
  AOI22D0BWP12T U956 ( .A1(n754), .A2(from_mem_data_out[2]), .B1(n753), .B2(
        cpu_data_in[18]), .ZN(n746) );
  OAI211D0BWP12T U957 ( .A1(n758), .A2(n748), .B(n747), .C(n746), .ZN(n749) );
  AOI21D0BWP12T U958 ( .A1(cpu_data_in[2]), .A2(n760), .B(n749), .ZN(n750) );
  MOAI22D0BWP12T U959 ( .A1(n750), .A2(reset), .B1(cpu_data_in[26]), .B2(n761), 
        .ZN(N197) );
  CKND2D0BWP12T U960 ( .A1(n752), .A2(tmp_value_2[1]), .ZN(n756) );
  AOI22D0BWP12T U961 ( .A1(n754), .A2(from_mem_data_out[1]), .B1(n753), .B2(
        cpu_data_in[17]), .ZN(n755) );
  OAI211D0BWP12T U962 ( .A1(n758), .A2(n757), .B(n756), .C(n755), .ZN(n759) );
  AOI21D0BWP12T U963 ( .A1(cpu_data_in[1]), .A2(n760), .B(n759), .ZN(n762) );
  MOAI22D0BWP12T U964 ( .A1(n762), .A2(reset), .B1(cpu_data_in[25]), .B2(n761), 
        .ZN(N196) );
  ND2D1BWP12T U965 ( .A1(n764), .A2(n763), .ZN(n776) );
  INVD0BWP12T U966 ( .I(n765), .ZN(n766) );
  AOI21D1BWP12T U967 ( .A1(n767), .A2(n766), .B(reset), .ZN(n769) );
  NR2D1BWP12T U968 ( .A1(n769), .A2(n768), .ZN(n778) );
  INVD1BWP12T U969 ( .I(n778), .ZN(n770) );
  MOAI22D0BWP12T U970 ( .A1(n783), .A2(n776), .B1(n770), .B2(tmp_value_2[1]), 
        .ZN(n398) );
  MOAI22D0BWP12T U971 ( .A1(n786), .A2(n776), .B1(n770), .B2(tmp_value_2[2]), 
        .ZN(n399) );
  MOAI22D0BWP12T U972 ( .A1(n784), .A2(n776), .B1(n770), .B2(tmp_value_2[4]), 
        .ZN(n401) );
  MOAI22D0BWP12T U973 ( .A1(n781), .A2(n776), .B1(n770), .B2(tmp_value_2[7]), 
        .ZN(n404) );
  MOAI22D0BWP12T U974 ( .A1(n780), .A2(n776), .B1(n770), .B2(tmp_value_2[3]), 
        .ZN(n400) );
  MOAI22D0BWP12T U975 ( .A1(n779), .A2(n776), .B1(n770), .B2(tmp_value_2[0]), 
        .ZN(n397) );
  MOAI22D0BWP12T U976 ( .A1(n785), .A2(n776), .B1(n770), .B2(tmp_value_2[5]), 
        .ZN(n402) );
  MOAI22D0BWP12T U977 ( .A1(n782), .A2(n776), .B1(n770), .B2(tmp_value_2[6]), 
        .ZN(n403) );
  MOAI22D0BWP12T U978 ( .A1(n788), .A2(n776), .B1(n770), .B2(tmp_value_2[8]), 
        .ZN(n405) );
  MOAI22D0BWP12T U979 ( .A1(n790), .A2(n776), .B1(n770), .B2(tmp_value_2[9]), 
        .ZN(n406) );
  MOAI22D0BWP12T U980 ( .A1(n791), .A2(n776), .B1(n770), .B2(tmp_value_2[13]), 
        .ZN(n410) );
  MOAI22D0BWP12T U981 ( .A1(n793), .A2(n776), .B1(n770), .B2(tmp_value_2[11]), 
        .ZN(n408) );
  MOAI22D0BWP12T U982 ( .A1(n789), .A2(n776), .B1(n770), .B2(tmp_value_2[12]), 
        .ZN(n409) );
  MOAI22D0BWP12T U983 ( .A1(n792), .A2(n776), .B1(n770), .B2(tmp_value_2[14]), 
        .ZN(n411) );
  MOAI22D0BWP12T U984 ( .A1(n787), .A2(n776), .B1(n770), .B2(tmp_value_2[10]), 
        .ZN(n407) );
  MOAI22D0BWP12T U985 ( .A1(n795), .A2(n776), .B1(n770), .B2(tmp_value_2[15]), 
        .ZN(n412) );
  INVD1BWP12T U986 ( .I(n771), .ZN(n772) );
  AO31D1BWP12T U987 ( .A1(n774), .A2(n773), .A3(n772), .B(reset), .Z(n796) );
  ND4D1BWP12T U988 ( .A1(n778), .A2(n777), .A3(n776), .A4(n775), .ZN(n794) );
  MOAI22D0BWP12T U989 ( .A1(n796), .A2(n779), .B1(tmp_value_1[0]), .B2(n794), 
        .ZN(n413) );
  MOAI22D0BWP12T U990 ( .A1(n796), .A2(n780), .B1(tmp_value_1[3]), .B2(n794), 
        .ZN(n416) );
  MOAI22D0BWP12T U991 ( .A1(n796), .A2(n781), .B1(tmp_value_1[7]), .B2(n794), 
        .ZN(n420) );
  MOAI22D0BWP12T U992 ( .A1(n796), .A2(n782), .B1(tmp_value_1[6]), .B2(n794), 
        .ZN(n419) );
  MOAI22D0BWP12T U993 ( .A1(n796), .A2(n783), .B1(tmp_value_1[1]), .B2(n794), 
        .ZN(n414) );
  MOAI22D0BWP12T U994 ( .A1(n796), .A2(n784), .B1(tmp_value_1[4]), .B2(n794), 
        .ZN(n417) );
  MOAI22D0BWP12T U995 ( .A1(n796), .A2(n785), .B1(tmp_value_1[5]), .B2(n794), 
        .ZN(n418) );
  MOAI22D0BWP12T U996 ( .A1(n796), .A2(n786), .B1(tmp_value_1[2]), .B2(n794), 
        .ZN(n415) );
  MOAI22D0BWP12T U997 ( .A1(n796), .A2(n787), .B1(tmp_value_1[10]), .B2(n794), 
        .ZN(n423) );
  MOAI22D0BWP12T U998 ( .A1(n796), .A2(n788), .B1(tmp_value_1[8]), .B2(n794), 
        .ZN(n421) );
  MOAI22D0BWP12T U999 ( .A1(n796), .A2(n789), .B1(tmp_value_1[12]), .B2(n794), 
        .ZN(n425) );
  MOAI22D0BWP12T U1000 ( .A1(n796), .A2(n790), .B1(tmp_value_1[9]), .B2(n794), 
        .ZN(n422) );
  MOAI22D0BWP12T U1001 ( .A1(n796), .A2(n791), .B1(tmp_value_1[13]), .B2(n794), 
        .ZN(n426) );
  MOAI22D0BWP12T U1002 ( .A1(n796), .A2(n792), .B1(tmp_value_1[14]), .B2(n794), 
        .ZN(n427) );
  MOAI22D0BWP12T U1003 ( .A1(n796), .A2(n793), .B1(tmp_value_1[11]), .B2(n794), 
        .ZN(n424) );
  MOAI22D0BWP12T U1004 ( .A1(n796), .A2(n795), .B1(tmp_value_1[15]), .B2(n794), 
        .ZN(n428) );
endmodule

