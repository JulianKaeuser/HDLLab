
module ALU_VARIABLE ( a, b, op, c_in, result, c_out, z, n, v );
  input [31:0] a;
  input [31:0] b;
  input [3:0] op;
  output [31:0] result;
  input c_in;
  output c_out, z, n, v;
  wire   n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909;
  tri   [3:0] op;

  MUX2ND0BWP12T U3 ( .I0(n5779), .I1(n5780), .S(n5864), .ZN(n4406) );
  MUX2ND0BWP12T U4 ( .I0(n5776), .I1(n5775), .S(b[15]), .ZN(n4350) );
  MUX2ND0BWP12T U5 ( .I0(n5813), .I1(n5812), .S(b[22]), .ZN(n4351) );
  MUX2ND0BWP12T U6 ( .I0(n5817), .I1(n5816), .S(b[12]), .ZN(n4355) );
  MUX2ND0BWP12T U7 ( .I0(n6240), .I1(n4755), .S(b[24]), .ZN(n4362) );
  MUX2ND0BWP12T U8 ( .I0(n5811), .I1(n5810), .S(b[22]), .ZN(n4365) );
  MUX2ND0BWP12T U9 ( .I0(n5779), .I1(n5780), .S(n5843), .ZN(n4345) );
  MUX2ND0BWP12T U10 ( .I0(n5870), .I1(n5869), .S(b[11]), .ZN(n4338) );
  XNR2D1BWP12T U11 ( .A1(a[19]), .A2(n4498), .ZN(n3490) );
  MUX2ND0BWP12T U12 ( .I0(n5876), .I1(n5875), .S(b[11]), .ZN(n3594) );
  MUX2ND0BWP12T U13 ( .I0(n5759), .I1(n5758), .S(n5612), .ZN(n3561) );
  IND2XD2BWP12T U14 ( .A1(n5360), .B1(a[0]), .ZN(n4755) );
  ND2D1BWP12T U15 ( .A1(a[17]), .A2(a[16]), .ZN(n6228) );
  OAI21D1BWP12T U16 ( .A1(n5144), .A2(n5142), .B(n5145), .ZN(n3973) );
  MUX2D1BWP12T U17 ( .I0(n6332), .I1(n6331), .S(n6576), .Z(n6339) );
  AOI22D1BWP12T U18 ( .A1(n6873), .A2(n6872), .B1(n6871), .B2(n6870), .ZN(
        n6901) );
  MUX2ND0BWP12T U19 ( .I0(n5817), .I1(n5816), .S(b[11]), .ZN(n4048) );
  MUX2ND0BWP12T U20 ( .I0(n5779), .I1(n5780), .S(n6782), .ZN(n4036) );
  MUX2ND0BWP12T U21 ( .I0(n4755), .I1(n6240), .S(n4758), .ZN(n3458) );
  MUX2ND0BWP12T U22 ( .I0(n4755), .I1(n6240), .S(n5467), .ZN(n3521) );
  MUX2ND0BWP12T U23 ( .I0(n5759), .I1(n5758), .S(n6782), .ZN(n3538) );
  MAOI22D0BWP12T U24 ( .A1(n5020), .A2(n4347), .B1(n4742), .B2(n4386), .ZN(
        n4424) );
  MUX2ND0BWP12T U25 ( .I0(n5804), .I1(n5805), .S(n6576), .ZN(n4407) );
  MAOI22D0BWP12T U26 ( .A1(n5807), .A2(n4348), .B1(n4744), .B2(n4385), .ZN(
        n4441) );
  MUX2ND0BWP12T U27 ( .I0(n5759), .I1(n5758), .S(n5379), .ZN(n4356) );
  MUX2ND0BWP12T U28 ( .I0(n5876), .I1(n5875), .S(b[18]), .ZN(n4354) );
  MUX2ND0BWP12T U29 ( .I0(n5876), .I1(n5875), .S(b[17]), .ZN(n4067) );
  XOR3D1BWP12T U30 ( .A1(n4065), .A2(n4063), .A3(n4062), .Z(n4054) );
  OAI21D1BWP12T U31 ( .A1(n6248), .A2(n5761), .B(n5759), .ZN(n3626) );
  MUX2ND0BWP12T U32 ( .I0(n5876), .I1(n5875), .S(b[9]), .ZN(n3685) );
  MAOI22D0BWP12T U33 ( .A1(n5845), .A2(n4480), .B1(n5382), .B2(n4432), .ZN(
        n4482) );
  MUX2ND0BWP12T U34 ( .I0(n5779), .I1(n5780), .S(n5379), .ZN(n4359) );
  MUX2ND0BWP12T U35 ( .I0(n5876), .I1(n5875), .S(b[20]), .ZN(n4367) );
  MUX2ND0BWP12T U36 ( .I0(n5870), .I1(n5869), .S(b[12]), .ZN(n4340) );
  MUX2ND0BWP12T U37 ( .I0(n5876), .I1(n5875), .S(b[21]), .ZN(n4496) );
  MAOI222D1BWP12T U38 ( .A(n3758), .B(n3756), .C(n3757), .ZN(n3730) );
  MUX2ND0BWP12T U39 ( .I0(n5776), .I1(n5775), .S(b[18]), .ZN(n4559) );
  MUX2ND0BWP12T U40 ( .I0(n4757), .I1(n4756), .S(n6334), .ZN(n3785) );
  ND2D1BWP12T U41 ( .A1(n3854), .A2(n3855), .ZN(n3864) );
  MUX2ND0BWP12T U42 ( .I0(n5876), .I1(n5875), .S(n6334), .ZN(n3857) );
  MUX2ND0BWP12T U43 ( .I0(n5779), .I1(n5780), .S(n5247), .ZN(n3416) );
  XOR3D1BWP12T U44 ( .A1(n3552), .A2(n3551), .A3(n3550), .Z(n3567) );
  OAI21D1BWP12T U45 ( .A1(n5500), .A2(n6061), .B(n5501), .ZN(n4010) );
  MUX2ND0BWP12T U46 ( .I0(n5876), .I1(n5875), .S(n5843), .ZN(n3755) );
  MUX2ND0BWP12T U47 ( .I0(n5779), .I1(n5780), .S(n5806), .ZN(n4590) );
  MUX2ND0BWP12T U48 ( .I0(n5759), .I1(n5758), .S(b[11]), .ZN(n4571) );
  MUX2ND0BWP12T U49 ( .I0(n5761), .I1(n5760), .S(b[12]), .ZN(n4570) );
  MUX2ND0BWP12T U50 ( .I0(n5870), .I1(n5869), .S(b[14]), .ZN(n4578) );
  FA1D0BWP12T U51 ( .A(n3819), .B(n3815), .CI(n3814), .CO(n3807), .S(n3829) );
  MUX2ND0BWP12T U52 ( .I0(n4755), .I1(n6240), .S(n4515), .ZN(n3858) );
  INVD1BWP12T U53 ( .I(n5238), .ZN(n4281) );
  FA1D0BWP12T U54 ( .A(n3653), .B(n3652), .CI(n3651), .CO(n4019), .S(n3654) );
  NR2D1BWP12T U55 ( .A1(n3999), .A2(n3998), .ZN(n4957) );
  ND3D2BWP12T U56 ( .A1(n5254), .A2(n5360), .A3(a[2]), .ZN(n5812) );
  CKBD1BWP12T U57 ( .I(n3911), .Z(n5811) );
  MUX2ND0BWP12T U58 ( .I0(n5876), .I1(n5875), .S(b[23]), .ZN(n4640) );
  INVD1BWP12T U59 ( .I(n4756), .ZN(n5836) );
  INVD1BWP12T U60 ( .I(n5861), .ZN(n5397) );
  NR2D1BWP12T U61 ( .A1(n3967), .A2(n3966), .ZN(n6014) );
  MUX2ND0BWP12T U62 ( .I0(n4755), .I1(n6240), .S(n6565), .ZN(n3881) );
  ND2D1BWP12T U63 ( .A1(n5812), .A2(n5813), .ZN(n3913) );
  INVD2BWP12T U64 ( .I(n3477), .ZN(n6520) );
  INVD1BWP12T U65 ( .I(n5719), .ZN(n5546) );
  NR2D1BWP12T U66 ( .A1(n5924), .A2(n4129), .ZN(n5505) );
  AOI21D1BWP12T U67 ( .A1(n5156), .A2(n4106), .B(n4105), .ZN(n5607) );
  AOI21D1BWP12T U68 ( .A1(n6172), .A2(n6095), .B(n4113), .ZN(n6171) );
  OAI21D1BWP12T U69 ( .A1(n5706), .A2(n5705), .B(n4111), .ZN(n6172) );
  OAI22D1BWP12T U70 ( .A1(n5069), .A2(n5238), .B1(n5239), .B2(n5016), .ZN(
        n4244) );
  MUX2D1BWP12T U71 ( .I0(a[20]), .I1(a[19]), .S(n6248), .Z(n5306) );
  AOI21D1BWP12T U72 ( .A1(n6155), .A2(n6504), .B(n6452), .ZN(n5052) );
  INVD1BWP12T U73 ( .I(n5058), .ZN(n4688) );
  OAI21D1BWP12T U74 ( .A1(n6055), .A2(n5497), .B(n5496), .ZN(n6063) );
  DEL025D1BWP12T U75 ( .I(a[12]), .Z(n6231) );
  AOI21D1BWP12T U76 ( .A1(n5525), .A2(n4212), .B(n6482), .ZN(n5001) );
  INVD2BWP12T U77 ( .I(n4371), .ZN(n5877) );
  ND2D1BWP12T U78 ( .A1(n3438), .A2(n6232), .ZN(n5872) );
  INVD1BWP12T U79 ( .I(n3405), .ZN(n5859) );
  INVD2BWP12T U80 ( .I(n5396), .ZN(n5860) );
  ND2D1BWP12T U81 ( .A1(n4381), .A2(a[16]), .ZN(n5758) );
  INVD1BWP12T U82 ( .I(n6066), .ZN(n4225) );
  INVD1BWP12T U83 ( .I(n6313), .ZN(n6297) );
  OR2XD1BWP12T U84 ( .A1(n3969), .A2(n3968), .Z(n5560) );
  ND2D1BWP12T U85 ( .A1(n3967), .A2(n3966), .ZN(n6015) );
  AOI21D1BWP12T U86 ( .A1(n5106), .A2(n4206), .B(n6499), .ZN(n5984) );
  NR2D1BWP12T U87 ( .A1(n3910), .A2(n3909), .ZN(n6028) );
  INVD1BWP12T U88 ( .I(n6862), .ZN(n6786) );
  OAI21D1BWP12T U89 ( .A1(n6055), .A2(n6054), .B(n6053), .ZN(n6060) );
  MUX2ND0BWP12T U90 ( .I0(n5870), .I1(n5869), .S(b[18]), .ZN(n5874) );
  MUX2ND0BWP12T U91 ( .I0(n5876), .I1(n5875), .S(b[26]), .ZN(n5880) );
  AO21D1BWP12T U92 ( .A1(n6085), .A2(n6834), .B(n4913), .Z(result[27]) );
  AO21D1BWP12T U93 ( .A1(n6072), .A2(n6834), .B(n5056), .Z(result[25]) );
  MAOI22D0BWP12T U94 ( .A1(n6355), .A2(n6387), .B1(n6396), .B2(n6584), .ZN(
        n6593) );
  XNR2D1BWP12T U95 ( .A1(n5105), .A2(n5104), .ZN(n6040) );
  ND2D1BWP12T U96 ( .A1(n3408), .A2(n5103), .ZN(n5104) );
  IOA21D1BWP12T U97 ( .A1(n6086), .A2(n6834), .B(n5701), .ZN(result[26]) );
  OAI21D1BWP12T U98 ( .A1(n6064), .A2(n6902), .B(n5521), .ZN(result[20]) );
  OAI21D1BWP12T U99 ( .A1(n6048), .A2(n6902), .B(n5646), .ZN(result[14]) );
  RCOAI21D1BWP12T U100 ( .A1(n6043), .A2(n6902), .B(n4273), .ZN(result[10]) );
  RCOAI21D1BWP12T U101 ( .A1(n6044), .A2(n6902), .B(n5221), .ZN(result[9]) );
  IOA21D1BWP12T U102 ( .A1(n6909), .A2(n6908), .B(n6907), .ZN(result[2]) );
  INVD1BWP12T U103 ( .I(b[22]), .ZN(n5467) );
  NR2D1BWP12T U104 ( .A1(b[16]), .A2(b[15]), .ZN(n4155) );
  MUX2ND0BWP12T U105 ( .I0(n5861), .I1(n5860), .S(b[17]), .ZN(n2975) );
  MUX2ND0BWP12T U106 ( .I0(n5859), .I1(n5858), .S(b[18]), .ZN(n2976) );
  NR2D0BWP12T U107 ( .A1(n2975), .A2(n2976), .ZN(n4043) );
  MUX2ND0BWP12T U108 ( .I0(n4755), .I1(n6240), .S(n3666), .ZN(n2977) );
  IAO21D0BWP12T U109 ( .A1(b[14]), .A2(n5361), .B(n2977), .ZN(n3716) );
  MUX2ND0BWP12T U110 ( .I0(n5761), .I1(n5760), .S(b[11]), .ZN(n2978) );
  MUX2ND0BWP12T U111 ( .I0(n5759), .I1(n5758), .S(n5806), .ZN(n2979) );
  NR2D0BWP12T U112 ( .A1(n2978), .A2(n2979), .ZN(n4485) );
  AO22D0BWP12T U113 ( .A1(n6552), .A2(n4893), .B1(n4894), .B2(n6553), .Z(n6517) );
  CKND0BWP12T U114 ( .I(n6576), .ZN(n2980) );
  AOI211D0BWP12T U115 ( .A1(n5767), .A2(n4868), .B(n5766), .C(n2980), .ZN(
        n6356) );
  MOAI22D0BWP12T U116 ( .A1(a[20]), .A2(n6648), .B1(a[20]), .B2(n6648), .ZN(
        n2981) );
  CKND0BWP12T U117 ( .I(n6398), .ZN(n2982) );
  AOI22D0BWP12T U118 ( .A1(n5507), .A2(n6394), .B1(n5546), .B2(n2982), .ZN(
        n2983) );
  OAI21D0BWP12T U119 ( .A1(b[20]), .A2(n6882), .B(n6874), .ZN(n2984) );
  AOI22D0BWP12T U120 ( .A1(a[20]), .A2(n2984), .B1(b[20]), .B2(n5509), .ZN(
        n2985) );
  CKND0BWP12T U121 ( .I(a[20]), .ZN(n2986) );
  AOI32D0BWP12T U122 ( .A1(b[20]), .A2(n2986), .A3(n6879), .B1(n6783), .B2(
        n2986), .ZN(n2987) );
  OAI211D0BWP12T U123 ( .A1(n5508), .A2(n6704), .B(n2985), .C(n2987), .ZN(
        n2988) );
  AOI211D0BWP12T U124 ( .A1(n5510), .A2(n6688), .B(n6661), .C(n2988), .ZN(
        n2989) );
  OAI211D0BWP12T U125 ( .A1(n5571), .A2(n5720), .B(n2983), .C(n2989), .ZN(
        n2990) );
  OAI22D0BWP12T U126 ( .A1(n6344), .A2(n6666), .B1(n6680), .B2(n6528), .ZN(
        n2991) );
  AOI211D0BWP12T U127 ( .A1(n6786), .A2(n2981), .B(n2990), .C(n2991), .ZN(
        n5517) );
  MAOI22D0BWP12T U128 ( .A1(n5605), .A2(n5608), .B1(n5605), .B2(n5608), .ZN(
        n5948) );
  OAI21D0BWP12T U129 ( .A1(n5607), .A2(n6089), .B(n5529), .ZN(n2992) );
  MAOI22D0BWP12T U130 ( .A1(n5530), .A2(n2992), .B1(n5530), .B2(n2992), .ZN(
        n6202) );
  MUX2ND0BWP12T U131 ( .I0(n4370), .I1(n4369), .S(b[19]), .ZN(n2993) );
  MUX2ND0BWP12T U132 ( .I0(n4372), .I1(n4371), .S(b[18]), .ZN(n2994) );
  CKND2D0BWP12T U133 ( .A1(n2993), .A2(n2994), .ZN(n4400) );
  MUX2ND0BWP12T U134 ( .I0(n4755), .I1(n6240), .S(n4576), .ZN(n2995) );
  IAO21D0BWP12T U135 ( .A1(b[12]), .A2(n5361), .B(n2995), .ZN(n3773) );
  MUX2ND0BWP12T U136 ( .I0(n5860), .I1(n5861), .S(n4745), .ZN(n2996) );
  MUX2ND0BWP12T U137 ( .I0(n5859), .I1(n5858), .S(b[12]), .ZN(n2997) );
  NR2D0BWP12T U138 ( .A1(n2996), .A2(n2997), .ZN(n3678) );
  CKND0BWP12T U139 ( .I(b[9]), .ZN(n2998) );
  MUX2ND0BWP12T U140 ( .I0(n5781), .I1(n5782), .S(n4515), .ZN(n2999) );
  OAI221D0BWP12T U141 ( .A1(b[9]), .A2(n5779), .B1(n2998), .B2(n5780), .C(
        n2999), .ZN(n4564) );
  AO222D0BWP12T U142 ( .A1(n6264), .A2(n4889), .B1(n6229), .B2(n5229), .C1(
        n5230), .C2(n6231), .Z(n6273) );
  OAI22D0BWP12T U143 ( .A1(n6533), .A2(n5435), .B1(n6530), .B2(n5436), .ZN(
        n3000) );
  OAI22D0BWP12T U144 ( .A1(n6246), .A2(a[30]), .B1(n5437), .B2(a[31]), .ZN(
        n3001) );
  AOI211D0BWP12T U145 ( .A1(n6556), .A2(n6551), .B(n3000), .C(n3001), .ZN(
        n3002) );
  IND2D0BWP12T U146 ( .A1(n5438), .B1(n6562), .ZN(n3003) );
  OAI211D0BWP12T U147 ( .A1(n6557), .A2(n3002), .B(n6355), .C(n3003), .ZN(
        n3004) );
  AOI21D0BWP12T U148 ( .A1(n6573), .A2(n6512), .B(n3004), .ZN(n6547) );
  MAOI22D0BWP12T U149 ( .A1(n5013), .A2(n5051), .B1(n5013), .B2(n5051), .ZN(
        n5963) );
  MOAI22D0BWP12T U150 ( .A1(n5071), .A2(n5097), .B1(n5071), .B2(n5097), .ZN(
        n6212) );
  MUX2ND0BWP12T U151 ( .I0(n5406), .I1(n5407), .S(n6576), .ZN(n3005) );
  MUX2ND0BWP12T U152 ( .I0(n5779), .I1(n5780), .S(n6573), .ZN(n3006) );
  NR2D0BWP12T U153 ( .A1(n3005), .A2(n3006), .ZN(n4042) );
  AO21D0BWP12T U154 ( .A1(n6403), .A2(n4381), .B(n3577), .Z(n3007) );
  OR2D0BWP12T U155 ( .A1(n3579), .A2(n3578), .Z(n3008) );
  CKND0BWP12T U156 ( .I(b[15]), .ZN(n3009) );
  CKND0BWP12T U157 ( .I(n5812), .ZN(n3010) );
  MAOI22D0BWP12T U158 ( .A1(b[14]), .A2(n3010), .B1(b[14]), .B2(n5813), .ZN(
        n3011) );
  OAI221D0BWP12T U159 ( .A1(b[15]), .A2(n3911), .B1(n3009), .B2(n5810), .C(
        n3011), .ZN(n3012) );
  MAOI222D0BWP12T U160 ( .A(n3007), .B(n3008), .C(n3012), .ZN(n3616) );
  MOAI22D0BWP12T U161 ( .A1(n3008), .A2(n3012), .B1(n3008), .B2(n3012), .ZN(
        n3013) );
  MAOI22D0BWP12T U162 ( .A1(n3007), .A2(n3013), .B1(n3007), .B2(n3013), .ZN(
        n3721) );
  MAOI222D0BWP12T U163 ( .A(a[26]), .B(a[25]), .C(n4829), .ZN(n3014) );
  AN2D0BWP12T U164 ( .A1(n3014), .A2(a[27]), .Z(n4563) );
  MUX2ND0BWP12T U165 ( .I0(n4646), .I1(n4647), .S(n4497), .ZN(n3015) );
  OAI21D0BWP12T U166 ( .A1(n5361), .A2(b[11]), .B(n3015), .ZN(n3782) );
  CKND0BWP12T U167 ( .I(b[23]), .ZN(n3016) );
  CKND0BWP12T U168 ( .I(n5875), .ZN(n3017) );
  MAOI22D0BWP12T U169 ( .A1(b[24]), .A2(n3017), .B1(b[24]), .B2(n5876), .ZN(
        n3018) );
  OAI221D0BWP12T U170 ( .A1(b[23]), .A2(n5878), .B1(n3016), .B2(n5877), .C(
        n3018), .ZN(n5398) );
  AOI22D0BWP12T U171 ( .A1(n5176), .A2(n5660), .B1(n5175), .B2(n5289), .ZN(
        n3019) );
  AOI22D0BWP12T U172 ( .A1(n5662), .A2(n5177), .B1(n5661), .B2(n5173), .ZN(
        n3020) );
  CKND2D0BWP12T U173 ( .A1(n3019), .A2(n3020), .ZN(n6395) );
  AOI21D0BWP12T U174 ( .A1(n6676), .A2(n6677), .B(n6857), .ZN(n3021) );
  MAOI22D0BWP12T U175 ( .A1(n6688), .A2(n6687), .B1(n6681), .B2(n6680), .ZN(
        n3022) );
  CKND0BWP12T U176 ( .I(a[18]), .ZN(n3023) );
  CKND0BWP12T U177 ( .I(n6679), .ZN(n3024) );
  OAI32D0BWP12T U178 ( .A1(n3023), .A2(n6862), .A3(n6678), .B1(a[18]), .B2(
        n3024), .ZN(n3025) );
  CKND0BWP12T U179 ( .I(n6682), .ZN(n3026) );
  OAI21D0BWP12T U180 ( .A1(b[18]), .A2(n6683), .B(n6874), .ZN(n3027) );
  AOI22D0BWP12T U181 ( .A1(n6747), .A2(n6685), .B1(n6684), .B2(n3027), .ZN(
        n3028) );
  OAI211D0BWP12T U182 ( .A1(n6813), .A2(n3026), .B(n6686), .C(n3028), .ZN(
        n3029) );
  AOI211D0BWP12T U183 ( .A1(n6870), .A2(n6690), .B(n3025), .C(n3029), .ZN(
        n3030) );
  OAI211D0BWP12T U184 ( .A1(n6689), .A2(n3021), .B(n3022), .C(n3030), .ZN(
        n3031) );
  AO21D0BWP12T U185 ( .A1(n6691), .A2(n6833), .B(n3031), .Z(n6692) );
  MAOI22D0BWP12T U186 ( .A1(n5650), .A2(n5652), .B1(n5650), .B2(n5652), .ZN(
        n5961) );
  MOAI22D0BWP12T U187 ( .A1(n4797), .A2(n4217), .B1(n4797), .B2(n4217), .ZN(
        n6210) );
  MUX2ND0BWP12T U188 ( .I0(n4755), .I1(n6240), .S(n4882), .ZN(n3032) );
  IAO21D0BWP12T U189 ( .A1(b[26]), .A2(n5361), .B(n3032), .ZN(n4484) );
  IND2D0BWP12T U190 ( .A1(n6332), .B1(n6576), .ZN(n5668) );
  AO22D0BWP12T U191 ( .A1(n3463), .A2(n5169), .B1(n4284), .B2(a[31]), .Z(n6323) );
  NR2D0BWP12T U192 ( .A1(n5515), .A2(n6624), .ZN(n3033) );
  CKND0BWP12T U193 ( .I(n4216), .ZN(n3034) );
  MOAI22D0BWP12T U194 ( .A1(n6624), .A2(n6618), .B1(n5463), .B2(n6614), .ZN(
        n3035) );
  AOI211D1BWP12T U195 ( .A1(n5459), .A2(n3033), .B(n3034), .C(n3035), .ZN(
        n5462) );
  CKND0BWP12T U196 ( .I(b[12]), .ZN(n3036) );
  MUX2ND0BWP12T U197 ( .I0(n5781), .I1(n5782), .S(n4745), .ZN(n3037) );
  OAI221D0BWP12T U198 ( .A1(b[12]), .A2(n5779), .B1(n3036), .B2(n5780), .C(
        n3037), .ZN(n5394) );
  CKND0BWP12T U199 ( .I(n5297), .ZN(n3038) );
  MAOI22D0BWP12T U200 ( .A1(n5662), .A2(n3038), .B1(n6409), .B2(n5250), .ZN(
        n3039) );
  OA211D0BWP12T U201 ( .A1(n6410), .A2(n5299), .B(n5730), .C(n3039), .Z(n6763)
         );
  MOAI22D0BWP12T U202 ( .A1(n4865), .A2(n4867), .B1(n4865), .B2(n4867), .ZN(
        n5964) );
  MOAI22D0BWP12T U203 ( .A1(n5651), .A2(n5652), .B1(n5651), .B2(n5652), .ZN(
        n6214) );
  CKND0BWP12T U204 ( .I(b[9]), .ZN(n3040) );
  CKND0BWP12T U205 ( .I(n5869), .ZN(n3041) );
  MAOI22D0BWP12T U206 ( .A1(n5806), .A2(n3041), .B1(n5806), .B2(n5870), .ZN(
        n3042) );
  OAI221D0BWP12T U207 ( .A1(b[9]), .A2(n5872), .B1(n3040), .B2(n5871), .C(
        n3042), .ZN(n4419) );
  MUX2ND0BWP12T U208 ( .I0(n4755), .I1(n6240), .S(n4343), .ZN(n3043) );
  IAO21D0BWP12T U209 ( .A1(n5864), .A2(n5361), .B(n3043), .ZN(n3924) );
  CKND0BWP12T U210 ( .I(b[14]), .ZN(n3044) );
  CKND0BWP12T U211 ( .I(n5758), .ZN(n3045) );
  MAOI22D0BWP12T U212 ( .A1(b[13]), .A2(n3045), .B1(b[13]), .B2(n5759), .ZN(
        n3046) );
  OAI221D0BWP12T U213 ( .A1(b[14]), .A2(n5761), .B1(n3044), .B2(n5760), .C(
        n3046), .ZN(n5399) );
  CKND0BWP12T U214 ( .I(n5614), .ZN(n3047) );
  AO222D0BWP12T U215 ( .A1(n3047), .A2(n5575), .B1(n6313), .B2(n5615), .C1(
        n6278), .C2(n5118), .Z(n6290) );
  MAOI22D0BWP12T U216 ( .A1(a[31]), .A2(n6248), .B1(a[31]), .B2(n6248), .ZN(
        n3048) );
  AOI22D0BWP12T U217 ( .A1(n5768), .A2(n5765), .B1(n5764), .B2(n3048), .ZN(
        n5826) );
  MAOI22D0BWP12T U218 ( .A1(n5528), .A2(n5530), .B1(n5528), .B2(n5530), .ZN(
        n5951) );
  MOAI22D0BWP12T U219 ( .A1(n4866), .A2(n4867), .B1(n4866), .B2(n4867), .ZN(
        n6215) );
  AOI211D0BWP12T U220 ( .A1(n6857), .A2(n6669), .B(n6668), .C(n6667), .ZN(
        n3049) );
  CKND2D0BWP12T U221 ( .A1(n6870), .A2(n6670), .ZN(n3050) );
  OAI211D0BWP12T U222 ( .A1(n6894), .A2(n6671), .B(n3049), .C(n3050), .ZN(
        n3051) );
  AOI31D0BWP12T U223 ( .A1(n6898), .A2(n6672), .A3(n6673), .B(n3051), .ZN(
        n3052) );
  IND2D0BWP12T U224 ( .A1(n6674), .B1(n6728), .ZN(n3053) );
  OAI211D0BWP12T U225 ( .A1(n6902), .A2(n6675), .B(n3052), .C(n3053), .ZN(
        result[19]) );
  CKND0BWP12T U226 ( .I(n6573), .ZN(n3054) );
  CKND0BWP12T U227 ( .I(n5869), .ZN(n3055) );
  MAOI22D0BWP12T U228 ( .A1(n6782), .A2(n3055), .B1(n6782), .B2(n5870), .ZN(
        n3056) );
  OAI221D0BWP12T U229 ( .A1(n6573), .A2(n5872), .B1(n3054), .B2(n5871), .C(
        n3056), .ZN(n3557) );
  CKND0BWP12T U230 ( .I(b[28]), .ZN(n3057) );
  CKND2D0BWP12T U231 ( .A1(n4882), .A2(n4557), .ZN(n3058) );
  OAI221D0BWP12T U232 ( .A1(b[28]), .A2(n6240), .B1(n3057), .B2(n4755), .C(
        n3058), .ZN(n4629) );
  CKND0BWP12T U233 ( .I(n5226), .ZN(n3059) );
  MUX2ND0BWP12T U234 ( .I0(n5813), .I1(n5812), .S(n5247), .ZN(n3060) );
  AOI21D0BWP12T U235 ( .A1(n3902), .A2(n3059), .B(n3060), .ZN(n3918) );
  MUX2ND0BWP12T U236 ( .I0(n5778), .I1(n5777), .S(b[18]), .ZN(n3061) );
  MUX2ND0BWP12T U237 ( .I0(n5776), .I1(n5775), .S(b[19]), .ZN(n3062) );
  NR2D0BWP12T U238 ( .A1(n3061), .A2(n3062), .ZN(n4753) );
  CKND0BWP12T U239 ( .I(b[25]), .ZN(n3063) );
  CKND0BWP12T U240 ( .I(n4746), .ZN(n3064) );
  MAOI22D0BWP12T U241 ( .A1(b[26]), .A2(n3064), .B1(b[26]), .B2(n4747), .ZN(
        n3065) );
  OAI221D0BWP12T U242 ( .A1(b[25]), .A2(n5861), .B1(n3063), .B2(n5860), .C(
        n3065), .ZN(n5393) );
  IND2D0BWP12T U243 ( .A1(n6202), .B1(n6870), .ZN(n5552) );
  OA222D0BWP12T U244 ( .A1(n5173), .A2(n6407), .B1(n6409), .B2(n5174), .C1(
        n6410), .C2(n5175), .Z(n6792) );
  MAOI22D0BWP12T U245 ( .A1(n5924), .A2(n6170), .B1(n5924), .B2(n6170), .ZN(
        n6671) );
  MAOI22D0BWP12T U246 ( .A1(n5281), .A2(n5321), .B1(n5281), .B2(n5321), .ZN(
        n6217) );
  CKND2D0BWP12T U247 ( .A1(n6317), .A2(n6316), .ZN(n3066) );
  IND3D0BWP12T U248 ( .A1(n6620), .B1(n6318), .B2(n6343), .ZN(n3067) );
  ND4D0BWP12T U249 ( .A1(n6665), .A2(n6314), .A3(n6740), .A4(n6315), .ZN(n3068) );
  NR4D0BWP12T U250 ( .A1(n6346), .A2(n3066), .A3(n3067), .A4(n3068), .ZN(n6377) );
  CKND2D0BWP12T U251 ( .A1(a[23]), .A2(a[21]), .ZN(n3069) );
  ND3D0BWP12T U252 ( .A1(a[31]), .A2(a[30]), .A3(n6783), .ZN(n3070) );
  NR4D0BWP12T U253 ( .A1(n6228), .A2(n6227), .A3(n3069), .A4(n3070), .ZN(n3071) );
  ND4D0BWP12T U254 ( .A1(n6247), .A2(a[29]), .A3(a[28]), .A4(n3071), .ZN(n6236) );
  MAOI22D0BWP12T U255 ( .A1(n6136), .A2(n6180), .B1(n6136), .B2(n6180), .ZN(
        n6899) );
  CKND0BWP12T U256 ( .I(b[13]), .ZN(n3072) );
  CKND0BWP12T U257 ( .I(n5875), .ZN(n3073) );
  MAOI22D0BWP12T U258 ( .A1(b[14]), .A2(n3073), .B1(b[14]), .B2(n5876), .ZN(
        n3074) );
  OAI221D0BWP12T U259 ( .A1(b[13]), .A2(n5878), .B1(n3072), .B2(n5877), .C(
        n3074), .ZN(n3484) );
  CKND0BWP12T U260 ( .I(b[24]), .ZN(n3075) );
  CKND0BWP12T U261 ( .I(n4746), .ZN(n3076) );
  MAOI22D0BWP12T U262 ( .A1(b[25]), .A2(n3076), .B1(b[25]), .B2(n4747), .ZN(
        n3077) );
  OAI221D0BWP12T U263 ( .A1(b[24]), .A2(n5861), .B1(n3075), .B2(n5860), .C(
        n3077), .ZN(n4740) );
  MUX2ND0BWP12T U264 ( .I0(n4755), .I1(n6240), .S(n5419), .ZN(n3078) );
  IAO21D0BWP12T U265 ( .A1(b[29]), .A2(n5361), .B(n3078), .ZN(n5385) );
  MAOI22D0BWP12T U266 ( .A1(n6576), .A2(n5073), .B1(n6576), .B2(n5079), .ZN(
        n6511) );
  IND2D0BWP12T U267 ( .A1(n6489), .B1(n4860), .ZN(n5320) );
  MAOI22D0BWP12T U268 ( .A1(n5769), .A2(n5771), .B1(n5769), .B2(n5771), .ZN(
        n3079) );
  MAOI22D0BWP12T U269 ( .A1(n5770), .A2(n3079), .B1(n5770), .B2(n3079), .ZN(
        n5787) );
  AN3D0BWP12T U270 ( .A1(n5383), .A2(a[31]), .A3(n5366), .Z(n5853) );
  INR2D0BWP12T U271 ( .A1(n6651), .B1(n5505), .ZN(n3080) );
  MAOI22D0BWP12T U272 ( .A1(n3080), .A2(n5515), .B1(n3080), .B2(n5515), .ZN(
        n5955) );
  AOI21D0BWP12T U273 ( .A1(n6167), .A2(n5428), .B(n5429), .ZN(n3081) );
  OAI21D0BWP12T U274 ( .A1(n5430), .A2(n6167), .B(n3081), .ZN(n6218) );
  AOI22D0BWP12T U275 ( .A1(n5660), .A2(n5680), .B1(n5662), .B2(n5681), .ZN(
        n3082) );
  CKND2D0BWP12T U276 ( .A1(n5661), .A2(n5682), .ZN(n3083) );
  OAI211D0BWP12T U277 ( .A1(n6409), .A2(n5663), .B(n3082), .C(n3083), .ZN(
        n3084) );
  AOI22D0BWP12T U278 ( .A1(n6411), .A2(n3084), .B1(n6391), .B2(n5664), .ZN(
        n3085) );
  AOI22D0BWP12T U279 ( .A1(n5659), .A2(n6378), .B1(n6893), .B2(n5666), .ZN(
        n3086) );
  IND3D0BWP12T U280 ( .A1(n5665), .B1(n3085), .B2(n3086), .ZN(n6434) );
  MAOI22D0BWP12T U281 ( .A1(n5227), .A2(n4952), .B1(n5227), .B2(n4952), .ZN(
        n6138) );
  IND2D0BWP12T U282 ( .A1(n5598), .B1(n5599), .ZN(n3087) );
  MAOI22D0BWP12T U283 ( .A1(n5600), .A2(n3087), .B1(n5600), .B2(n3087), .ZN(
        n6048) );
  MOAI22D0BWP12T U284 ( .A1(n6836), .A2(n6148), .B1(n6833), .B2(n5954), .ZN(
        n3088) );
  AO211D0BWP12T U285 ( .A1(n5728), .A2(n6679), .B(n5726), .C(n3088), .Z(n3089)
         );
  AOI211D0BWP12T U286 ( .A1(n5991), .A2(n6728), .B(n5727), .C(n3089), .ZN(
        n3090) );
  OAI21D0BWP12T U287 ( .A1(n6050), .A2(n6902), .B(n3090), .ZN(result[17]) );
  CKND0BWP12T U288 ( .I(b[12]), .ZN(n3091) );
  CKND2D0BWP12T U289 ( .A1(n5151), .A2(n4390), .ZN(n3092) );
  OAI221D0BWP12T U290 ( .A1(b[12]), .A2(n5819), .B1(n3091), .B2(n5818), .C(
        n3092), .ZN(n4429) );
  MOAI22D0BWP12T U291 ( .A1(n4748), .A2(n4585), .B1(n4584), .B2(n4874), .ZN(
        n3093) );
  CKND0BWP12T U292 ( .I(b[19]), .ZN(n3094) );
  CKND0BWP12T U293 ( .I(n5838), .ZN(n3095) );
  MAOI22D0BWP12T U294 ( .A1(b[18]), .A2(n3095), .B1(b[18]), .B2(n5839), .ZN(
        n3096) );
  OAI221D0BWP12T U295 ( .A1(b[19]), .A2(n5837), .B1(n3094), .B2(n5836), .C(
        n3096), .ZN(n3097) );
  CKND0BWP12T U296 ( .I(b[13]), .ZN(n3098) );
  CKND0BWP12T U297 ( .I(n5872), .ZN(n3099) );
  MAOI22D0BWP12T U298 ( .A1(n4497), .A2(n3099), .B1(n4497), .B2(n5871), .ZN(
        n3100) );
  OAI221D0BWP12T U299 ( .A1(b[13]), .A2(n5870), .B1(n3098), .B2(n5869), .C(
        n3100), .ZN(n3101) );
  MAOI222D0BWP12T U300 ( .A(n3093), .B(n3097), .C(n3101), .ZN(n4673) );
  MOAI22D0BWP12T U301 ( .A1(n3093), .A2(n3097), .B1(n3093), .B2(n3097), .ZN(
        n3102) );
  MAOI22D0BWP12T U302 ( .A1(n3101), .A2(n3102), .B1(n3101), .B2(n3102), .ZN(
        n4580) );
  OAI21D0BWP12T U303 ( .A1(n4650), .A2(n4649), .B(n5371), .ZN(n4777) );
  AN3D0BWP12T U304 ( .A1(n4135), .A2(n5762), .A3(n6887), .Z(n6789) );
  CKND0BWP12T U305 ( .I(n6572), .ZN(n3103) );
  AOI22D0BWP12T U306 ( .A1(n6573), .A2(n6574), .B1(n6578), .B2(n3103), .ZN(
        n3104) );
  OA211D0BWP12T U307 ( .A1(n6576), .A2(n6577), .B(n6575), .C(n3104), .Z(n6650)
         );
  CKND0BWP12T U308 ( .I(b[24]), .ZN(n3105) );
  CKND0BWP12T U309 ( .I(n5875), .ZN(n3106) );
  MAOI22D0BWP12T U310 ( .A1(b[25]), .A2(n3106), .B1(b[25]), .B2(n5876), .ZN(
        n3107) );
  OAI221D0BWP12T U311 ( .A1(b[24]), .A2(n5878), .B1(n3105), .B2(n5877), .C(
        n3107), .ZN(n5786) );
  MAOI22D0BWP12T U312 ( .A1(n4962), .A2(n5000), .B1(n4962), .B2(n5000), .ZN(
        n5953) );
  IND2D0BWP12T U313 ( .A1(n4804), .B1(n6845), .ZN(n4809) );
  MOAI22D0BWP12T U314 ( .A1(n5012), .A2(n5051), .B1(n5012), .B2(n5051), .ZN(
        n6213) );
  AOI22D0BWP12T U315 ( .A1(n5660), .A2(n5681), .B1(n5662), .B2(n5683), .ZN(
        n3108) );
  CKND2D0BWP12T U316 ( .A1(n5661), .A2(n5674), .ZN(n3109) );
  OAI211D0BWP12T U317 ( .A1(n6409), .A2(n5306), .B(n3108), .C(n3109), .ZN(
        n3110) );
  CKND0BWP12T U318 ( .I(n5081), .ZN(n3111) );
  AOI222D0BWP12T U319 ( .A1(n3110), .A2(n6411), .B1(n6742), .B2(n5666), .C1(
        n3111), .C2(n5664), .ZN(n3112) );
  IOA21D0BWP12T U320 ( .A1(n5659), .A2(n5080), .B(n3112), .ZN(n6432) );
  CKND2D0BWP12T U321 ( .A1(n6128), .A2(n6129), .ZN(n3113) );
  MAOI22D0BWP12T U322 ( .A1(n6707), .A2(n3113), .B1(n6707), .B2(n3113), .ZN(
        n6698) );
  CKND2D0BWP12T U323 ( .A1(n5647), .A2(n5648), .ZN(n3114) );
  MOAI22D0BWP12T U324 ( .A1(n6078), .A2(n3114), .B1(n6078), .B2(n3114), .ZN(
        n6086) );
  MOAI22D0BWP12T U325 ( .A1(n4942), .A2(n4952), .B1(n4942), .B2(n4952), .ZN(
        n5981) );
  OAI211D0BWP12T U326 ( .A1(n6894), .A2(n5951), .B(n5552), .C(n5551), .ZN(
        n3115) );
  AOI211D0BWP12T U327 ( .A1(n6728), .A2(n5554), .B(n5553), .C(n3115), .ZN(
        n3116) );
  OAI21D1BWP12T U328 ( .A1(n6049), .A2(n6902), .B(n3116), .ZN(result[15]) );
  MUX2ND0BWP12T U329 ( .I0(n5778), .I1(n5777), .S(b[11]), .ZN(n3117) );
  MUX2ND0BWP12T U330 ( .I0(n5776), .I1(n5775), .S(b[12]), .ZN(n3118) );
  NR2D0BWP12T U331 ( .A1(n3117), .A2(n3118), .ZN(n4041) );
  MAOI22D0BWP12T U332 ( .A1(n4776), .A2(n4777), .B1(n4776), .B2(n4777), .ZN(
        n3119) );
  MAOI22D0BWP12T U333 ( .A1(n4775), .A2(n3119), .B1(n4775), .B2(n3119), .ZN(
        n4774) );
  CKND0BWP12T U334 ( .I(b[14]), .ZN(n3120) );
  CKND2D0BWP12T U335 ( .A1(n5530), .A2(n4623), .ZN(n3121) );
  OAI221D0BWP12T U336 ( .A1(b[14]), .A2(n5872), .B1(n3120), .B2(n5871), .C(
        n3121), .ZN(n4739) );
  AOI222D0BWP12T U337 ( .A1(n6411), .A2(n6378), .B1(n6436), .B2(n6391), .C1(
        n6893), .C2(n6717), .ZN(n3122) );
  AOI21D0BWP12T U338 ( .A1(n3122), .A2(n6438), .B(n6677), .ZN(n6689) );
  IND2D0BWP12T U339 ( .A1(n4235), .B1(n4236), .ZN(n6198) );
  OA222D0BWP12T U340 ( .A1(n5175), .A2(n6534), .B1(n5174), .B2(n5677), .C1(
        n5173), .C2(n6533), .Z(n6778) );
  MAOI22D0BWP12T U341 ( .A1(n5704), .A2(n5705), .B1(n5704), .B2(n5705), .ZN(
        n5954) );
  NR3D0BWP12T U342 ( .A1(n6457), .A2(n6614), .A3(n6813), .ZN(n3123) );
  NR3D0BWP12T U343 ( .A1(n6450), .A2(n6452), .A3(n6451), .ZN(n3124) );
  ND4D0BWP12T U344 ( .A1(n6448), .A2(n6458), .A3(n6449), .A4(n3124), .ZN(n3125) );
  NR4D0BWP12T U345 ( .A1(n6453), .A2(n6454), .A3(n6455), .A4(n3125), .ZN(n3126) );
  ND3D0BWP12T U346 ( .A1(n6456), .A2(n3123), .A3(n3126), .ZN(n6475) );
  IND4D0BWP12T U347 ( .A1(n6473), .B1(n6472), .B2(n6471), .B3(n6470), .ZN(
        n3127) );
  INR4D0BWP12T U348 ( .A1(n6467), .B1(n6468), .B2(n6878), .B3(n6469), .ZN(
        n3128) );
  NR4D0BWP12T U349 ( .A1(n6464), .A2(n6463), .A3(n6465), .A4(n6743), .ZN(n3129) );
  INR4D0BWP12T U350 ( .A1(n6459), .B1(n6462), .B2(n6460), .B3(n6461), .ZN(
        n3130) );
  IND4D0BWP12T U351 ( .A1(n3127), .B1(n3128), .B2(n3129), .B3(n3130), .ZN(
        n6474) );
  IND2D0BWP12T U352 ( .A1(n4096), .B1(n4220), .ZN(n6154) );
  IND2D0BWP12T U353 ( .A1(n5522), .B1(n5523), .ZN(n3131) );
  MAOI22D0BWP12T U354 ( .A1(n5524), .A2(n3131), .B1(n5524), .B2(n3131), .ZN(
        n6049) );
  IND2D0BWP12T U355 ( .A1(n5968), .B1(n6164), .ZN(n3132) );
  MAOI22D0BWP12T U356 ( .A1(n6166), .A2(n3132), .B1(n6166), .B2(n3132), .ZN(
        n6831) );
  MUX2ND0BWP12T U357 ( .I0(n5161), .I1(n5160), .S(a[13]), .ZN(n3133) );
  AOI211D0BWP12T U358 ( .A1(n6870), .A2(n6199), .B(n5191), .C(n3133), .ZN(
        n3134) );
  OAI22D0BWP12T U359 ( .A1(n5950), .A2(n6894), .B1(n5988), .B2(n6890), .ZN(
        n3135) );
  AOI21D0BWP12T U360 ( .A1(n6145), .A2(n6898), .B(n3135), .ZN(n3136) );
  OAI211D0BWP12T U361 ( .A1(n6046), .A2(n6902), .B(n3134), .C(n3136), .ZN(
        result[13]) );
  CKND0BWP12T U362 ( .I(b[23]), .ZN(n3137) );
  CKND2D0BWP12T U363 ( .A1(n5467), .A2(n4557), .ZN(n3138) );
  OAI221D0BWP12T U364 ( .A1(b[23]), .A2(n6240), .B1(n3137), .B2(n4755), .C(
        n3138), .ZN(n4039) );
  MUX2ND0BWP12T U365 ( .I0(n5761), .I1(n5760), .S(n6782), .ZN(n3139) );
  MUX2ND0BWP12T U366 ( .I0(n5759), .I1(n5758), .S(n6573), .ZN(n3140) );
  NR2D0BWP12T U367 ( .A1(n3139), .A2(n3140), .ZN(n3459) );
  CKND0BWP12T U368 ( .I(n4745), .ZN(n3141) );
  MUX2ND0BWP12T U369 ( .I0(n5876), .I1(n5875), .S(b[12]), .ZN(n3142) );
  AOI221D0BWP12T U370 ( .A1(n4371), .A2(n3141), .B1(n4372), .B2(n4745), .C(
        n3142), .ZN(n3637) );
  IAO21D0BWP12T U371 ( .A1(n6623), .A2(n5069), .B(n5807), .ZN(n4347) );
  INR3D0BWP12T U372 ( .A1(n6247), .B1(n5360), .B2(a[2]), .ZN(n4935) );
  IOA21D0BWP12T U373 ( .A1(n4583), .A2(n4907), .B(n4584), .ZN(n5387) );
  MAOI22D0BWP12T U374 ( .A1(n6264), .A2(n5166), .B1(n4918), .B2(n6708), .ZN(
        n3143) );
  OA21D0BWP12T U375 ( .A1(n4919), .A2(n5626), .B(n3143), .Z(n6298) );
  MOAI22D0BWP12T U376 ( .A1(n6520), .A2(n6255), .B1(n6520), .B2(n4868), .ZN(
        n5537) );
  CKND0BWP12T U377 ( .I(b[16]), .ZN(n3144) );
  CKND0BWP12T U378 ( .I(n5869), .ZN(n3145) );
  MAOI22D0BWP12T U379 ( .A1(b[17]), .A2(n3145), .B1(b[17]), .B2(n5870), .ZN(
        n3146) );
  OAI221D0BWP12T U380 ( .A1(b[16]), .A2(n5872), .B1(n3144), .B2(n5871), .C(
        n3146), .ZN(n5771) );
  MUX2ND0BWP12T U381 ( .I0(n3405), .I1(n5395), .S(b[27]), .ZN(n3147) );
  MUX2ND0BWP12T U382 ( .I0(n5397), .I1(n5396), .S(b[26]), .ZN(n3148) );
  CKND2D0BWP12T U383 ( .A1(n3147), .A2(n3148), .ZN(n5792) );
  AOI211D0BWP12T U384 ( .A1(n6110), .A2(n6842), .B(n5910), .C(n6455), .ZN(
        n3149) );
  CKND2D0BWP12T U385 ( .A1(n5907), .A2(n5417), .ZN(n3150) );
  AOI21D0BWP12T U386 ( .A1(n3150), .A2(n6455), .B(n3149), .ZN(n5429) );
  MOAI22D0BWP12T U387 ( .A1(n5488), .A2(n5489), .B1(n5488), .B2(n5489), .ZN(
        n5959) );
  CKND2D0BWP12T U388 ( .A1(n5514), .A2(n6651), .ZN(n3151) );
  MAOI22D0BWP12T U389 ( .A1(n5515), .A2(n3151), .B1(n5515), .B2(n3151), .ZN(
        n6207) );
  OAI211D0BWP12T U390 ( .A1(n6440), .A2(n6439), .B(n6435), .C(n6438), .ZN(
        n3152) );
  AO21D0BWP12T U391 ( .A1(n6436), .A2(n6437), .B(n3152), .Z(n6619) );
  MOAI22D0BWP12T U392 ( .A1(n4963), .A2(n5000), .B1(n4963), .B2(n5000), .ZN(
        n6146) );
  IND2D0BWP12T U393 ( .A1(n6054), .B1(n6053), .ZN(n3153) );
  MAOI22D0BWP12T U394 ( .A1(n6055), .A2(n3153), .B1(n6055), .B2(n3153), .ZN(
        n6050) );
  CKND0BWP12T U395 ( .I(n5979), .ZN(n3154) );
  OA21D0BWP12T U396 ( .A1(n5977), .A2(n3154), .B(n5978), .Z(n6891) );
  CKND2D0BWP12T U397 ( .A1(n6279), .A2(n6905), .ZN(n3155) );
  AOI21D0BWP12T U398 ( .A1(n3155), .A2(n6840), .B(n6315), .ZN(n3156) );
  OAI21D0BWP12T U399 ( .A1(n5719), .A2(n6380), .B(n5214), .ZN(n3157) );
  AO211D0BWP12T U400 ( .A1(n5578), .A2(n6510), .B(n3156), .C(n3157), .Z(n3158)
         );
  CKND0BWP12T U401 ( .I(n5507), .ZN(n3159) );
  OAI22D0BWP12T U402 ( .A1(n6229), .A2(n5217), .B1(n6395), .B2(n3159), .ZN(
        n3160) );
  AOI211D0BWP12T U403 ( .A1(n5216), .A2(n5215), .B(n3158), .C(n3160), .ZN(
        n3161) );
  AOI22D0BWP12T U404 ( .A1(n6362), .A2(n6909), .B1(n6833), .B2(n5937), .ZN(
        n3162) );
  OAI211D0BWP12T U405 ( .A1(n6195), .A2(n6794), .B(n3161), .C(n3162), .ZN(
        n5218) );
  CKND2D0BWP12T U406 ( .A1(n6164), .A2(n6165), .ZN(n3163) );
  MOAI22D0BWP12T U407 ( .A1(n6166), .A2(n3163), .B1(n6166), .B2(n3163), .ZN(
        n6837) );
  MUX2ND0BWP12T U408 ( .I0(n4757), .I1(n4756), .S(b[12]), .ZN(n3164) );
  MUX2ND0BWP12T U409 ( .I0(n4759), .I1(n4760), .S(b[11]), .ZN(n3165) );
  CKND2D0BWP12T U410 ( .A1(n3164), .A2(n3165), .ZN(n3498) );
  CKND0BWP12T U411 ( .I(n3463), .ZN(n3166) );
  OAI221D0BWP12T U412 ( .A1(n3463), .A2(n6353), .B1(n3166), .B2(n4326), .C(
        n6520), .ZN(n5019) );
  CKND0BWP12T U413 ( .I(b[16]), .ZN(n3167) );
  CKND2D0BWP12T U414 ( .A1(n5530), .A2(n4738), .ZN(n3168) );
  OAI221D0BWP12T U415 ( .A1(b[16]), .A2(n5870), .B1(n3167), .B2(n5869), .C(
        n3168), .ZN(n5359) );
  MUX2ND0BWP12T U416 ( .I0(n5819), .I1(n5818), .S(b[17]), .ZN(n3169) );
  MUX2ND0BWP12T U417 ( .I0(n5817), .I1(n5816), .S(b[18]), .ZN(n3170) );
  NR2D0BWP12T U418 ( .A1(n3169), .A2(n3170), .ZN(n5400) );
  IND2D0BWP12T U419 ( .A1(n4611), .B1(n4610), .ZN(n3171) );
  MAOI22D0BWP12T U420 ( .A1(n4609), .A2(n3171), .B1(n4609), .B2(n3171), .ZN(
        n4708) );
  IOA21D0BWP12T U421 ( .A1(n6278), .A2(n6323), .B(n6335), .ZN(n6620) );
  CKND0BWP12T U422 ( .I(n5250), .ZN(n3172) );
  OAI21D0BWP12T U423 ( .A1(n6407), .A2(n5252), .B(n5251), .ZN(n3173) );
  AOI21D0BWP12T U424 ( .A1(n5660), .A2(n3172), .B(n3173), .ZN(n5571) );
  INR2D0BWP12T U425 ( .A1(n5082), .B1(n5095), .ZN(n6504) );
  MAOI222D0BWP12T U426 ( .A(n4773), .B(n4774), .C(n4772), .ZN(n3174) );
  MOAI22D0BWP12T U427 ( .A1(n5409), .A2(n3174), .B1(n5409), .B2(n3174), .ZN(
        n3175) );
  MAOI22D0BWP12T U428 ( .A1(n5408), .A2(n3175), .B1(n5408), .B2(n3175), .ZN(
        n5410) );
  MAOI222D0BWP12T U429 ( .A(n3174), .B(n3176), .C(n3177), .ZN(n5751) );
  CKND0BWP12T U430 ( .I(n5408), .ZN(n3176) );
  CKND0BWP12T U431 ( .I(n5409), .ZN(n3177) );
  CKND0BWP12T U432 ( .I(n5139), .ZN(n3178) );
  OA21D0BWP12T U433 ( .A1(n5117), .A2(n3178), .B(n5928), .Z(n5935) );
  MOAI22D0BWP12T U434 ( .A1(n4964), .A2(n5000), .B1(n4964), .B2(n5000), .ZN(
        n6203) );
  IND2D0BWP12T U435 ( .A1(n6127), .B1(n6126), .ZN(n3179) );
  MAOI22D0BWP12T U436 ( .A1(n6682), .A2(n3179), .B1(n6682), .B2(n3179), .ZN(
        n6693) );
  CKND2D0BWP12T U437 ( .A1(n6061), .A2(n6062), .ZN(n3180) );
  MOAI22D0BWP12T U438 ( .A1(n6063), .A2(n3180), .B1(n6063), .B2(n3180), .ZN(
        n6675) );
  NR2D0BWP12T U439 ( .A1(n5154), .A2(n5153), .ZN(n3181) );
  MOAI22D0BWP12T U440 ( .A1(n3181), .A2(n5157), .B1(n3181), .B2(n5157), .ZN(
        n5988) );
  CKND0BWP12T U441 ( .I(b[15]), .ZN(n3182) );
  CKND0BWP12T U442 ( .I(n5760), .ZN(n3183) );
  MAOI22D0BWP12T U443 ( .A1(b[16]), .A2(n3183), .B1(b[16]), .B2(n5761), .ZN(
        n3184) );
  OAI221D0BWP12T U444 ( .A1(b[15]), .A2(n5759), .B1(n3182), .B2(n5758), .C(
        n3184), .ZN(n3185) );
  NR2D0BWP12T U445 ( .A1(n5762), .A2(n5763), .ZN(n3186) );
  AO21D0BWP12T U446 ( .A1(a[31]), .A2(n5767), .B(n5766), .Z(n3187) );
  AOI22D0BWP12T U447 ( .A1(n5768), .A2(n3187), .B1(n5764), .B2(n5765), .ZN(
        n3188) );
  MAOI222D0BWP12T U448 ( .A(n5769), .B(n5770), .C(n5771), .ZN(n3189) );
  MAOI22D0BWP12T U449 ( .A1(n3188), .A2(n3189), .B1(n3188), .B2(n3189), .ZN(
        n3190) );
  MAOI22D0BWP12T U450 ( .A1(n3186), .A2(n3190), .B1(n3186), .B2(n3190), .ZN(
        n3191) );
  MAOI22D0BWP12T U451 ( .A1(n3185), .A2(n3191), .B1(n3185), .B2(n3191), .ZN(
        n3192) );
  CKND0BWP12T U452 ( .I(b[14]), .ZN(n3193) );
  MUX2ND0BWP12T U453 ( .I0(n5782), .I1(n5781), .S(b[13]), .ZN(n3194) );
  OAI221D0BWP12T U454 ( .A1(b[14]), .A2(n5779), .B1(n3193), .B2(n5780), .C(
        n3194), .ZN(n3195) );
  CKND0BWP12T U455 ( .I(b[22]), .ZN(n3196) );
  CKND0BWP12T U456 ( .I(n5777), .ZN(n3197) );
  MAOI22D0BWP12T U457 ( .A1(b[21]), .A2(n3197), .B1(b[21]), .B2(n5778), .ZN(
        n3198) );
  OAI221D0BWP12T U458 ( .A1(b[22]), .A2(n5776), .B1(n3196), .B2(n5775), .C(
        n3198), .ZN(n3199) );
  MAOI22D0BWP12T U459 ( .A1(n3195), .A2(n3199), .B1(n3195), .B2(n3199), .ZN(
        n3200) );
  MAOI222D0BWP12T U460 ( .A(n5774), .B(n5772), .C(n5773), .ZN(n3201) );
  MAOI22D0BWP12T U461 ( .A1(n3200), .A2(n3201), .B1(n3200), .B2(n3201), .ZN(
        n3202) );
  MAOI22D0BWP12T U462 ( .A1(n3192), .A2(n3202), .B1(n3192), .B2(n3202), .ZN(
        n5797) );
  OAI32D0BWP12T U463 ( .A1(n6824), .A2(n6808), .A3(n6807), .B1(n6840), .B2(
        n6824), .ZN(n3203) );
  CKND2D0BWP12T U464 ( .A1(n6811), .A2(n6810), .ZN(n3204) );
  OAI22D0BWP12T U465 ( .A1(n6814), .A2(n6813), .B1(n6882), .B2(n6812), .ZN(
        n3205) );
  AOI31D0BWP12T U466 ( .A1(n6815), .A2(n6816), .A3(n3204), .B(n3205), .ZN(
        n3206) );
  OAI211D0BWP12T U467 ( .A1(n6892), .A2(n6817), .B(n6888), .C(n3206), .ZN(
        n3207) );
  AOI211D0BWP12T U468 ( .A1(n6823), .A2(n6909), .B(n3203), .C(n3207), .ZN(
        n3208) );
  CKND0BWP12T U469 ( .I(n6819), .ZN(n3209) );
  CKND0BWP12T U470 ( .I(n6820), .ZN(n3210) );
  OAI32D0BWP12T U471 ( .A1(n3209), .A2(n6818), .A3(n6862), .B1(n6819), .B2(
        n3210), .ZN(n3211) );
  AOI21D0BWP12T U472 ( .A1(n6809), .A2(n6870), .B(n3211), .ZN(n3212) );
  OAI211D0BWP12T U473 ( .A1(n6822), .A2(n6821), .B(n3208), .C(n3212), .ZN(
        n6825) );
  MOAI22D0BWP12T U474 ( .A1(n5280), .A2(n5321), .B1(n5280), .B2(n5321), .ZN(
        n5967) );
  MUX2ND0BWP12T U475 ( .I0(n5813), .I1(n5812), .S(b[18]), .ZN(n3213) );
  MUX2ND0BWP12T U476 ( .I0(n5811), .I1(n5810), .S(b[19]), .ZN(n3214) );
  NR2D0BWP12T U477 ( .A1(n3213), .A2(n3214), .ZN(n3520) );
  MUX2ND0BWP12T U478 ( .I0(n5778), .I1(n5777), .S(n5612), .ZN(n3215) );
  MUX2ND0BWP12T U479 ( .I0(n5776), .I1(n5775), .S(n5247), .ZN(n3216) );
  NR2D0BWP12T U480 ( .A1(n3215), .A2(n3216), .ZN(n3800) );
  MUX2ND0BWP12T U481 ( .I0(n4755), .I1(n6240), .S(n4357), .ZN(n3217) );
  IAO21D0BWP12T U482 ( .A1(n6782), .A2(n5361), .B(n3217), .ZN(n3927) );
  MAOI22D0BWP12T U483 ( .A1(n6334), .A2(n6778), .B1(n6334), .B2(n6539), .ZN(
        n6566) );
  CKND0BWP12T U484 ( .I(n4552), .ZN(n3218) );
  MAOI22D0BWP12T U485 ( .A1(n4550), .A2(n3218), .B1(n4550), .B2(n4551), .ZN(
        n4709) );
  AO222D0BWP12T U486 ( .A1(n6264), .A2(n4985), .B1(a[14]), .B2(n5229), .C1(
        n5230), .C2(a[17]), .Z(n6252) );
  IOA21D0BWP12T U487 ( .A1(n6334), .A2(n6352), .B(n6335), .ZN(n6629) );
  IND2D0BWP12T U488 ( .A1(n4209), .B1(n6129), .ZN(n6450) );
  MAOI22D0BWP12T U489 ( .A1(n5345), .A2(n5348), .B1(n5345), .B2(n5348), .ZN(
        n3219) );
  MAOI22D0BWP12T U490 ( .A1(n5347), .A2(n3219), .B1(n5347), .B2(n3219), .ZN(
        n3220) );
  MAOI22D0BWP12T U491 ( .A1(n3220), .A2(n5411), .B1(n3220), .B2(n5411), .ZN(
        n3221) );
  MAOI22D0BWP12T U492 ( .A1(n5410), .A2(n3221), .B1(n5410), .B2(n3221), .ZN(
        n5341) );
  MAOI222D0BWP12T U493 ( .A(n5410), .B(n3220), .C(n5411), .ZN(n3222) );
  CKND0BWP12T U494 ( .I(n3222), .ZN(n5750) );
  MUX2ND0BWP12T U495 ( .I0(n5805), .I1(n5804), .S(b[11]), .ZN(n3223) );
  MUX2ND0BWP12T U496 ( .I0(n5803), .I1(n5802), .S(b[12]), .ZN(n3224) );
  NR2D0BWP12T U497 ( .A1(n3223), .A2(n3224), .ZN(n5825) );
  CKND0BWP12T U498 ( .I(b[22]), .ZN(n3225) );
  CKND0BWP12T U499 ( .I(n5836), .ZN(n3226) );
  MAOI22D0BWP12T U500 ( .A1(b[23]), .A2(n3226), .B1(b[23]), .B2(n5837), .ZN(
        n3227) );
  OAI221D0BWP12T U501 ( .A1(b[22]), .A2(n5839), .B1(n3225), .B2(n5838), .C(
        n3227), .ZN(n5769) );
  MOAI22D0BWP12T U502 ( .A1(n5801), .A2(n5799), .B1(n5801), .B2(n5799), .ZN(
        n3228) );
  MAOI22D0BWP12T U503 ( .A1(n5800), .A2(n3228), .B1(n5800), .B2(n3228), .ZN(
        n5785) );
  MAOI22D0BWP12T U504 ( .A1(n6419), .A2(n6420), .B1(n6419), .B2(n6421), .ZN(
        n6718) );
  OAI22D0BWP12T U505 ( .A1(n6408), .A2(n5175), .B1(n5240), .B2(n4923), .ZN(
        n3229) );
  NR2D0BWP12T U506 ( .A1(n4938), .A2(n5437), .ZN(n3230) );
  AOI211D0BWP12T U507 ( .A1(n4924), .A2(n3229), .B(n3230), .C(n6573), .ZN(
        n3231) );
  OA22D1BWP12T U508 ( .A1(n6297), .A2(n6299), .B1(n6259), .B2(n6306), .Z(n3232) );
  OA211D1BWP12T U509 ( .A1(n6298), .A2(n6308), .B(n3231), .C(n3232), .Z(n4950)
         );
  MAOI22D0BWP12T U510 ( .A1(n4333), .A2(n4217), .B1(n4333), .B2(n4217), .ZN(
        n5958) );
  MAOI22D0BWP12T U511 ( .A1(n5466), .A2(n5489), .B1(n5466), .B2(n5489), .ZN(
        n6209) );
  INR4D0BWP12T U512 ( .A1(n6480), .B1(n6481), .B2(n6482), .B3(n6483), .ZN(
        n6492) );
  AOI21D0BWP12T U513 ( .A1(n6063), .A2(n6062), .B(n5499), .ZN(n3233) );
  IND2D0BWP12T U514 ( .A1(n5500), .B1(n5501), .ZN(n3234) );
  MAOI22D0BWP12T U515 ( .A1(n3233), .A2(n3234), .B1(n3233), .B2(n3234), .ZN(
        n6064) );
  MAOI22D0BWP12T U516 ( .A1(n5525), .A2(n5530), .B1(n5525), .B2(n5530), .ZN(
        n5989) );
  IAO21D0BWP12T U517 ( .A1(n6463), .A2(n6135), .B(n5138), .ZN(n3235) );
  MOAI22D0BWP12T U518 ( .A1(n5139), .A2(n3235), .B1(n5139), .B2(n3235), .ZN(
        n6140) );
  CKND2D0BWP12T U519 ( .A1(n6843), .A2(n5911), .ZN(n3236) );
  MOAI22D0BWP12T U520 ( .A1(n4804), .A2(n3236), .B1(n4804), .B2(n3236), .ZN(
        n6600) );
  AN2D0BWP12T U521 ( .A1(n4823), .A2(n5866), .Z(n3237) );
  CKND0BWP12T U522 ( .I(b[26]), .ZN(n3238) );
  IND2D0BWP12T U523 ( .A1(b[25]), .B1(n4557), .ZN(n3239) );
  OAI221D0BWP12T U524 ( .A1(b[26]), .A2(n6240), .B1(n3238), .B2(n4755), .C(
        n3239), .ZN(n3240) );
  CKND0BWP12T U525 ( .I(b[24]), .ZN(n3241) );
  CKND0BWP12T U526 ( .I(n5812), .ZN(n3242) );
  MAOI22D0BWP12T U527 ( .A1(b[23]), .A2(n3242), .B1(b[23]), .B2(n5813), .ZN(
        n3243) );
  OAI221D0BWP12T U528 ( .A1(b[24]), .A2(n5811), .B1(n3241), .B2(n5810), .C(
        n3243), .ZN(n3244) );
  MAOI222D0BWP12T U529 ( .A(n3237), .B(n3240), .C(n3244), .ZN(n4560) );
  MOAI22D0BWP12T U530 ( .A1(n3240), .A2(n3244), .B1(n3240), .B2(n3244), .ZN(
        n3245) );
  MAOI22D0BWP12T U531 ( .A1(n3237), .A2(n3245), .B1(n3237), .B2(n3245), .ZN(
        n4475) );
  MUX2ND0BWP12T U532 ( .I0(n4757), .I1(n4756), .S(n5247), .ZN(n3246) );
  MUX2ND0BWP12T U533 ( .I0(n4759), .I1(n4760), .S(n5612), .ZN(n3247) );
  CKND2D0BWP12T U534 ( .A1(n3246), .A2(n3247), .ZN(n3840) );
  IOA21D0BWP12T U535 ( .A1(n4823), .A2(a[14]), .B(n4920), .ZN(n6531) );
  IOA21D0BWP12T U536 ( .A1(n4498), .A2(a[0]), .B(n4144), .ZN(n3896) );
  CKND0BWP12T U537 ( .I(b[13]), .ZN(n3248) );
  OAI21D0BWP12T U538 ( .A1(a[13]), .A2(n3248), .B(n5149), .ZN(n5601) );
  MUX2ND0BWP12T U539 ( .I0(n5804), .I1(n5805), .S(n5405), .ZN(n3249) );
  MUX2ND0BWP12T U540 ( .I0(n5803), .I1(n5802), .S(b[11]), .ZN(n3250) );
  NR2D0BWP12T U541 ( .A1(n3249), .A2(n3250), .ZN(n5831) );
  CKND0BWP12T U542 ( .I(b[15]), .ZN(n3251) );
  CKND0BWP12T U543 ( .I(n5758), .ZN(n3252) );
  MAOI22D0BWP12T U544 ( .A1(b[14]), .A2(n3252), .B1(b[14]), .B2(n5759), .ZN(
        n3253) );
  OAI221D0BWP12T U545 ( .A1(b[15]), .A2(n5761), .B1(n3251), .B2(n5760), .C(
        n3253), .ZN(n5770) );
  OAI222D0BWP12T U546 ( .A1(n6409), .A2(n5173), .B1(n6408), .B2(n5174), .C1(
        n6407), .C2(n5175), .ZN(n3254) );
  IAO21D0BWP12T U547 ( .A1(n6410), .A2(n5177), .B(n3254), .ZN(n6817) );
  CKND0BWP12T U548 ( .I(n6248), .ZN(n3255) );
  AOI221D0BWP12T U549 ( .A1(n6267), .A2(n6248), .B1(n6249), .B2(n3255), .C(
        n6533), .ZN(n3256) );
  AOI21D0BWP12T U550 ( .A1(n6245), .A2(n6875), .B(n6334), .ZN(n3257) );
  OAI21D0BWP12T U551 ( .A1(n6247), .A2(n6246), .B(n3257), .ZN(n3258) );
  AOI211D0BWP12T U552 ( .A1(n6520), .A2(n6250), .B(n3256), .C(n3258), .ZN(
        n3259) );
  OAI21D0BWP12T U553 ( .A1(n6251), .A2(n6308), .B(n6565), .ZN(n3260) );
  AOI211D0BWP12T U554 ( .A1(n6252), .A2(n6254), .B(n3259), .C(n3260), .ZN(
        n6333) );
  AOI21D0BWP12T U555 ( .A1(n6078), .A2(n5328), .B(n5337), .ZN(n3261) );
  CKND2D0BWP12T U556 ( .A1(n5279), .A2(n6074), .ZN(n3262) );
  MAOI22D0BWP12T U557 ( .A1(n3261), .A2(n3262), .B1(n3261), .B2(n3262), .ZN(
        n6084) );
  NR2D0BWP12T U558 ( .A1(n5971), .A2(n6127), .ZN(n3263) );
  MOAI22D0BWP12T U559 ( .A1(n3263), .A2(n6682), .B1(n3263), .B2(n6682), .ZN(
        n6694) );
  MAOI22D0BWP12T U560 ( .A1(n5753), .A2(n5754), .B1(n5753), .B2(n5754), .ZN(
        n3264) );
  MAOI22D0BWP12T U561 ( .A1(n5752), .A2(n3264), .B1(n5752), .B2(n3264), .ZN(
        n3265) );
  MAOI22D0BWP12T U562 ( .A1(n3265), .A2(n5751), .B1(n3265), .B2(n5751), .ZN(
        n3266) );
  MAOI22D0BWP12T U563 ( .A1(n5750), .A2(n3266), .B1(n5750), .B2(n3266), .ZN(
        n5412) );
  MAOI222D0BWP12T U564 ( .A(n5750), .B(n3265), .C(n5751), .ZN(n3267) );
  CKND0BWP12T U565 ( .I(n3267), .ZN(n5902) );
  CKND2D0BWP12T U566 ( .A1(n6197), .A2(n6198), .ZN(n3268) );
  MOAI22D0BWP12T U567 ( .A1(n6707), .A2(n3268), .B1(n6707), .B2(n3268), .ZN(
        n6727) );
  INR2D0BWP12T U568 ( .A1(n6811), .B1(n5944), .ZN(n3269) );
  MAOI22D0BWP12T U569 ( .A1(n3269), .A2(n6175), .B1(n3269), .B2(n6175), .ZN(
        n6772) );
  OA211D0BWP12T U570 ( .A1(n6892), .A2(n6792), .B(n6791), .C(n6790), .Z(n3270)
         );
  OAI32D0BWP12T U571 ( .A1(n6776), .A2(n6777), .A3(n6807), .B1(n6840), .B2(
        n6776), .ZN(n3271) );
  NR2D0BWP12T U572 ( .A1(n6795), .A2(n6794), .ZN(n3272) );
  AOI211D0BWP12T U573 ( .A1(n6793), .A2(n6909), .B(n3271), .C(n3272), .ZN(
        n3273) );
  OAI211D0BWP12T U574 ( .A1(n6822), .A2(n6778), .B(n3270), .C(n3273), .ZN(
        n6798) );
  AOI21D0BWP12T U575 ( .A1(n5227), .A2(n5226), .B(n6479), .ZN(n3274) );
  MAOI22D0BWP12T U576 ( .A1(n5274), .A2(n3274), .B1(n5274), .B2(n3274), .ZN(
        n6139) );
  AN2D0BWP12T U577 ( .A1(n5416), .A2(n6843), .Z(n6110) );
  IND2D0BWP12T U578 ( .A1(n5649), .B1(n5697), .ZN(n6160) );
  MAOI22D0BWP12T U579 ( .A1(n4539), .A2(n4537), .B1(n4539), .B2(n4537), .ZN(
        n3275) );
  MAOI22D0BWP12T U580 ( .A1(n4536), .A2(n3275), .B1(n4536), .B2(n3275), .ZN(
        n3276) );
  MAOI22D0BWP12T U581 ( .A1(n4679), .A2(n3276), .B1(n4679), .B2(n3276), .ZN(
        n3277) );
  MAOI22D0BWP12T U582 ( .A1(n4678), .A2(n3277), .B1(n4678), .B2(n3277), .ZN(
        n4686) );
  MAOI222D0BWP12T U583 ( .A(n4678), .B(n4679), .C(n3276), .ZN(n3278) );
  CKND0BWP12T U584 ( .I(n3278), .ZN(n4694) );
  CKND0BWP12T U585 ( .I(b[21]), .ZN(n3279) );
  CKND0BWP12T U586 ( .I(n5875), .ZN(n3280) );
  MAOI22D0BWP12T U587 ( .A1(b[22]), .A2(n3280), .B1(b[22]), .B2(n5876), .ZN(
        n3281) );
  OAI221D0BWP12T U588 ( .A1(b[21]), .A2(n5878), .B1(n3279), .B2(n5877), .C(
        n3281), .ZN(n4630) );
  INR2D0BWP12T U589 ( .A1(n6227), .B1(n5866), .ZN(n4584) );
  CKND0BWP12T U590 ( .I(n5612), .ZN(n3282) );
  CKND2D0BWP12T U591 ( .A1(n4888), .A2(n3903), .ZN(n3283) );
  OAI221D0BWP12T U592 ( .A1(n5612), .A2(n4747), .B1(n3282), .B2(n4746), .C(
        n3283), .ZN(n3919) );
  IND2D0BWP12T U593 ( .A1(n4524), .B1(n4525), .ZN(n3284) );
  MAOI22D0BWP12T U594 ( .A1(n4526), .A2(n3284), .B1(n4526), .B2(n3284), .ZN(
        n3407) );
  CKND0BWP12T U595 ( .I(b[11]), .ZN(n3285) );
  MUX2ND0BWP12T U596 ( .I0(n5781), .I1(n5782), .S(n5405), .ZN(n3286) );
  OAI221D0BWP12T U597 ( .A1(b[11]), .A2(n5779), .B1(n3285), .B2(n5780), .C(
        n3286), .ZN(n4780) );
  CKND0BWP12T U598 ( .I(n4611), .ZN(n3287) );
  MAOI22D0BWP12T U599 ( .A1(n4609), .A2(n3287), .B1(n4609), .B2(n4610), .ZN(
        n4711) );
  CKND0BWP12T U600 ( .I(n4922), .ZN(n3288) );
  AO32D0BWP12T U601 ( .A1(n4920), .A2(n4922), .A3(n4921), .B1(n3288), .B2(
        n6538), .Z(n6259) );
  IND2D0BWP12T U602 ( .A1(n5018), .B1(n5019), .ZN(n5209) );
  IAO21D0BWP12T U603 ( .A1(n4924), .A2(n6331), .B(n6324), .ZN(n6376) );
  IND2D0BWP12T U604 ( .A1(n4221), .B1(n4174), .ZN(n6680) );
  INR2D0BWP12T U605 ( .A1(c_in), .B1(n6457), .ZN(n4299) );
  MUX2ND0BWP12T U606 ( .I0(n5819), .I1(n5818), .S(b[18]), .ZN(n3289) );
  MUX2ND0BWP12T U607 ( .I0(n5817), .I1(n5816), .S(b[19]), .ZN(n3290) );
  NR2D0BWP12T U608 ( .A1(n3289), .A2(n3290), .ZN(n5827) );
  MAOI22D0BWP12T U609 ( .A1(n5385), .A2(n5383), .B1(n5385), .B2(n5383), .ZN(
        n3291) );
  MAOI22D0BWP12T U610 ( .A1(n5384), .A2(n3291), .B1(n5384), .B2(n3291), .ZN(
        n3292) );
  MAOI22D0BWP12T U611 ( .A1(n5371), .A2(n3292), .B1(n5371), .B2(n3292), .ZN(
        n3293) );
  MAOI22D0BWP12T U612 ( .A1(n5370), .A2(n3293), .B1(n5370), .B2(n3293), .ZN(
        n5350) );
  MAOI222D0BWP12T U613 ( .A(n5370), .B(n5371), .C(n3292), .ZN(n3294) );
  CKND0BWP12T U614 ( .I(n3294), .ZN(n5798) );
  IAO21D0BWP12T U615 ( .A1(n6357), .A2(n6317), .B(n4329), .ZN(n6283) );
  MOAI22D0BWP12T U616 ( .A1(n5067), .A2(n5097), .B1(n5067), .B2(n5097), .ZN(
        n5960) );
  INR4D0BWP12T U617 ( .A1(n6391), .B1(n6394), .B2(n6392), .B3(n6393), .ZN(
        n3295) );
  ND4D0BWP12T U618 ( .A1(n6395), .A2(n6763), .A3(n6396), .A4(n3295), .ZN(n3296) );
  ND4D0BWP12T U619 ( .A1(n6400), .A2(n6817), .A3(n6437), .A4(n6401), .ZN(n3297) );
  ND4D0BWP12T U620 ( .A1(n6792), .A2(n6398), .A3(n6399), .A4(n6397), .ZN(n3298) );
  NR4D0BWP12T U621 ( .A1(n6402), .A2(n3296), .A3(n3297), .A4(n3298), .ZN(n6428) );
  IND4D0BWP12T U622 ( .A1(n6510), .B1(n6738), .B2(n6513), .B3(n6512), .ZN(
        n3299) );
  AN4D0BWP12T U623 ( .A1(n6518), .A2(n6821), .A3(n6519), .A4(n6574), .Z(n3300)
         );
  IND4D0BWP12T U624 ( .A1(n6872), .B1(n6522), .B2(n6702), .B3(n3300), .ZN(
        n3301) );
  ND4D0BWP12T U625 ( .A1(n6778), .A2(n6524), .A3(n6514), .A4(n6515), .ZN(n3302) );
  NR4D0BWP12T U626 ( .A1(n6523), .A2(n3299), .A3(n3301), .A4(n3302), .ZN(n6585) );
  INR4D0BWP12T U627 ( .A1(n6494), .B1(n6495), .B2(n6624), .B3(n6496), .ZN(
        n6509) );
  INR4D0BWP12T U628 ( .A1(n6477), .B1(n6479), .B2(n6478), .B3(n6656), .ZN(
        n6493) );
  INR3D0BWP12T U629 ( .A1(n6487), .B1(n6488), .B2(n6489), .ZN(n6490) );
  MAOI222D0BWP12T U630 ( .A(n5392), .B(n5393), .C(n5394), .ZN(n5788) );
  INR2D0BWP12T U631 ( .A1(n5193), .B1(n5192), .ZN(n3303) );
  MAOI22D0BWP12T U632 ( .A1(n3303), .A2(n5194), .B1(n3303), .B2(n5194), .ZN(
        n6044) );
  MAOI22D0BWP12T U633 ( .A1(n6132), .A2(n6133), .B1(n6132), .B2(n6133), .ZN(
        n6827) );
  CKND0BWP12T U634 ( .I(n6191), .ZN(n3304) );
  CKND2D0BWP12T U635 ( .A1(n6833), .A2(n5935), .ZN(n3305) );
  OAI211D0BWP12T U636 ( .A1(n6794), .A2(n3304), .B(n5135), .C(n3305), .ZN(
        n5136) );
  IND2D0BWP12T U637 ( .A1(n5976), .B1(n5975), .ZN(n3306) );
  MAOI22D0BWP12T U638 ( .A1(n6134), .A2(n3306), .B1(n6134), .B2(n3306), .ZN(
        n6799) );
  CKND2D0BWP12T U639 ( .A1(n6881), .A2(n5266), .ZN(n3307) );
  MOAI22D0BWP12T U640 ( .A1(n4952), .A2(n3307), .B1(n4952), .B2(n3307), .ZN(
        n6186) );
  IND3D0BWP12T U641 ( .A1(n6597), .B1(n6353), .B2(n6786), .ZN(n5918) );
  CKND0BWP12T U642 ( .I(n5922), .ZN(n3308) );
  AOI21D0BWP12T U643 ( .A1(n6843), .A2(n3308), .B(n6842), .ZN(n3309) );
  MAOI22D0BWP12T U644 ( .A1(n3309), .A2(n4804), .B1(n3309), .B2(n4804), .ZN(
        n6004) );
  CKND0BWP12T U645 ( .I(b[31]), .ZN(n3310) );
  OA21D0BWP12T U646 ( .A1(a[31]), .A2(n3310), .B(n6476), .Z(n6612) );
  CKND0BWP12T U647 ( .I(n5612), .ZN(n3311) );
  ND2D1BWP12T U648 ( .A1(n6531), .A2(n4738), .ZN(n3312) );
  OAI221D1BWP12T U649 ( .A1(n5612), .A2(n5870), .B1(n3311), .B2(n5869), .C(
        n3312), .ZN(n3702) );
  MAOI22D0BWP12T U650 ( .A1(n3516), .A2(n3517), .B1(n3516), .B2(n3517), .ZN(
        n3313) );
  MAOI22D0BWP12T U651 ( .A1(n3520), .A2(n3313), .B1(n3520), .B2(n3313), .ZN(
        n3314) );
  MAOI22D0BWP12T U652 ( .A1(n3314), .A2(n3502), .B1(n3314), .B2(n3502), .ZN(
        n3315) );
  MAOI22D0BWP12T U653 ( .A1(n3501), .A2(n3315), .B1(n3501), .B2(n3315), .ZN(
        n3580) );
  MAOI222D0BWP12T U654 ( .A(n3501), .B(n3314), .C(n3502), .ZN(n3316) );
  CKND0BWP12T U655 ( .I(n3316), .ZN(n4077) );
  MAOI222D0BWP12T U656 ( .A(n4594), .B(n4596), .C(n4595), .ZN(n3317) );
  MOAI22D0BWP12T U657 ( .A1(n4652), .A2(n3317), .B1(n4652), .B2(n3317), .ZN(
        n3318) );
  MAOI22D0BWP12T U658 ( .A1(n4651), .A2(n3318), .B1(n4651), .B2(n3318), .ZN(
        n4615) );
  MAOI222D0BWP12T U659 ( .A(n3317), .B(n3319), .C(n3320), .ZN(n4722) );
  CKND0BWP12T U660 ( .I(n4651), .ZN(n3319) );
  CKND0BWP12T U661 ( .I(n4652), .ZN(n3320) );
  MUX2ND0BWP12T U662 ( .I0(n5839), .I1(n5838), .S(n5806), .ZN(n3321) );
  MUX2ND0BWP12T U663 ( .I0(n5837), .I1(n5836), .S(b[11]), .ZN(n3322) );
  NR2D0BWP12T U664 ( .A1(n3321), .A2(n3322), .ZN(n3589) );
  MOAI22D0BWP12T U665 ( .A1(n3774), .A2(n3773), .B1(n3774), .B2(n3773), .ZN(
        n3323) );
  MAOI22D0BWP12T U666 ( .A1(n3778), .A2(n3323), .B1(n3778), .B2(n3323), .ZN(
        n3324) );
  MAOI22D0BWP12T U667 ( .A1(n3795), .A2(n3324), .B1(n3795), .B2(n3324), .ZN(
        n3796) );
  CKND0BWP12T U668 ( .I(n3795), .ZN(n3325) );
  MAOI222D0BWP12T U669 ( .A(n3778), .B(n3325), .C(n3323), .ZN(n3791) );
  MUX2ND0BWP12T U670 ( .I0(n4755), .I1(n6240), .S(n4433), .ZN(n3326) );
  AOI21D0BWP12T U671 ( .A1(n6357), .A2(n4557), .B(n3326), .ZN(n3904) );
  IND2D0BWP12T U672 ( .A1(n4552), .B1(n4551), .ZN(n3327) );
  MAOI22D0BWP12T U673 ( .A1(n4550), .A2(n3327), .B1(n4550), .B2(n3327), .ZN(
        n3409) );
  AO31D0BWP12T U674 ( .A1(n3934), .A2(n6819), .A3(n6239), .B(n4372), .Z(n3328)
         );
  CKND0BWP12T U675 ( .I(n5612), .ZN(n3329) );
  CKND2D0BWP12T U676 ( .A1(n3935), .A2(n6263), .ZN(n3330) );
  OAI221D0BWP12T U677 ( .A1(n5612), .A2(n5876), .B1(n3329), .B2(n5875), .C(
        n3330), .ZN(n3331) );
  OR2D0BWP12T U678 ( .A1(n3933), .A2(n3932), .Z(n3332) );
  MAOI222D0BWP12T U679 ( .A(n3328), .B(n3331), .C(n3332), .ZN(n3959) );
  MOAI22D0BWP12T U680 ( .A1(n3328), .A2(n3331), .B1(n3328), .B2(n3331), .ZN(
        n3333) );
  MAOI22D0BWP12T U681 ( .A1(n3332), .A2(n3333), .B1(n3332), .B2(n3333), .ZN(
        n3949) );
  AOI32D0BWP12T U682 ( .A1(n6334), .A2(n5019), .A3(n4327), .B1(n6254), .B2(
        n5019), .ZN(n3334) );
  IND2D0BWP12T U683 ( .A1(n4328), .B1(n3334), .ZN(n6341) );
  INR2D0BWP12T U684 ( .A1(n5667), .B1(n6565), .ZN(n6364) );
  MOAI22D0BWP12T U685 ( .A1(n5767), .A2(n6256), .B1(n5767), .B2(n6259), .ZN(
        n6303) );
  AN2D0BWP12T U686 ( .A1(n6419), .A2(n5305), .Z(n5664) );
  MAOI22D0BWP12T U687 ( .A1(n5829), .A2(n5830), .B1(n5829), .B2(n5830), .ZN(
        n3335) );
  MAOI22D0BWP12T U688 ( .A1(n5831), .A2(n3335), .B1(n5831), .B2(n3335), .ZN(
        n5791) );
  CKND2D0BWP12T U689 ( .A1(n5213), .A2(n5202), .ZN(n3336) );
  MOAI22D0BWP12T U690 ( .A1(n4233), .A2(n3336), .B1(n4233), .B2(n3336), .ZN(
        n5946) );
  IND2D0BWP12T U691 ( .A1(n4179), .B1(n4174), .ZN(n6373) );
  OR4D0BWP12T U692 ( .A1(n6321), .A2(n6322), .A3(n6323), .A4(a[31]), .Z(n6386)
         );
  AOI22D0BWP12T U693 ( .A1(n5569), .A2(n6398), .B1(n5570), .B2(n5571), .ZN(
        n3337) );
  AOI21D0BWP12T U694 ( .A1(n6426), .A2(n3337), .B(n6292), .ZN(n6443) );
  CKND0BWP12T U695 ( .I(n5359), .ZN(n3338) );
  MAOI222D0BWP12T U696 ( .A(n5357), .B(n5358), .C(n3338), .ZN(n3339) );
  MAOI22D0BWP12T U697 ( .A1(n5885), .A2(n5887), .B1(n5885), .B2(n5887), .ZN(
        n3340) );
  MAOI22D0BWP12T U698 ( .A1(n5886), .A2(n3340), .B1(n5886), .B2(n3340), .ZN(
        n3341) );
  CKND0BWP12T U699 ( .I(n5798), .ZN(n3342) );
  MAOI222D0BWP12T U700 ( .A(n3339), .B(n3341), .C(n3342), .ZN(n5897) );
  MAOI22D0BWP12T U701 ( .A1(n3341), .A2(n3339), .B1(n3341), .B2(n3339), .ZN(
        n3343) );
  MAOI22D0BWP12T U702 ( .A1(n5798), .A2(n3343), .B1(n5798), .B2(n3343), .ZN(
        n5755) );
  INR4D0BWP12T U703 ( .A1(n6183), .B1(n6137), .B2(n6899), .B3(n6836), .ZN(
        n3344) );
  ND4D0BWP12T U704 ( .A1(n6138), .A2(n6139), .A3(n6796), .A4(n3344), .ZN(n3345) );
  NR4D0BWP12T U705 ( .A1(n6140), .A2(n6734), .A3(n6827), .A4(n3345), .ZN(n3346) );
  ND4D0BWP12T U706 ( .A1(n6698), .A2(n6141), .A3(n6142), .A4(n3346), .ZN(n3347) );
  NR4D0BWP12T U707 ( .A1(n6143), .A2(n6144), .A3(n6145), .A4(n3347), .ZN(n3348) );
  ND4D0BWP12T U708 ( .A1(n6148), .A2(n6146), .A3(n6147), .A4(n3348), .ZN(n3349) );
  AOI211D0BWP12T U709 ( .A1(n6673), .A2(n6672), .B(n6693), .C(n3349), .ZN(
        n3350) );
  ND4D0BWP12T U710 ( .A1(n6152), .A2(n6151), .A3(n6643), .A4(n3350), .ZN(n3351) );
  AOI211D0BWP12T U711 ( .A1(n6155), .A2(n6154), .B(n6153), .C(n3351), .ZN(
        n3352) );
  ND3D0BWP12T U712 ( .A1(n6156), .A2(n6165), .A3(n3352), .ZN(n6158) );
  CKND2D0BWP12T U713 ( .A1(n5899), .A2(n5900), .ZN(n3353) );
  MOAI22D0BWP12T U714 ( .A1(n5901), .A2(n3353), .B1(n5901), .B2(n3353), .ZN(
        n6608) );
  OA21D0BWP12T U715 ( .A1(n4040), .A2(n4039), .B(n4459), .Z(n4539) );
  MAOI222D0BWP12T U716 ( .A(n4506), .B(n4505), .C(n4507), .ZN(n3354) );
  MOAI22D0BWP12T U717 ( .A1(n4595), .A2(n4594), .B1(n4595), .B2(n4594), .ZN(
        n3355) );
  MAOI22D0BWP12T U718 ( .A1(n4596), .A2(n3355), .B1(n4596), .B2(n3355), .ZN(
        n3356) );
  MAOI22D0BWP12T U719 ( .A1(n3354), .A2(n3356), .B1(n3354), .B2(n3356), .ZN(
        n3357) );
  MAOI22D0BWP12T U720 ( .A1(n4553), .A2(n3357), .B1(n4553), .B2(n3357), .ZN(
        n4606) );
  CKND0BWP12T U721 ( .I(n4553), .ZN(n3358) );
  MAOI222D0BWP12T U722 ( .A(n3358), .B(n3354), .C(n3356), .ZN(n4614) );
  INR2D0BWP12T U723 ( .A1(n3588), .B1(n3589), .ZN(n3566) );
  MAOI22D0BWP12T U724 ( .A1(n3600), .A2(n3601), .B1(n3600), .B2(n3601), .ZN(
        n3359) );
  MAOI22D0BWP12T U725 ( .A1(n3599), .A2(n3359), .B1(n3599), .B2(n3359), .ZN(
        n3360) );
  CKND0BWP12T U726 ( .I(n3686), .ZN(n3361) );
  MAOI222D0BWP12T U727 ( .A(n3618), .B(n3360), .C(n3361), .ZN(n3651) );
  MAOI22D0BWP12T U728 ( .A1(n3686), .A2(n3360), .B1(n3686), .B2(n3360), .ZN(
        n3362) );
  MAOI22D0BWP12T U729 ( .A1(n3618), .A2(n3362), .B1(n3618), .B2(n3362), .ZN(
        n3687) );
  CKND0BWP12T U730 ( .I(n4730), .ZN(n3363) );
  MUX2ND0BWP12T U731 ( .I0(n5859), .I1(n5858), .S(n5806), .ZN(n3364) );
  AOI221D0BWP12T U732 ( .A1(n5396), .A2(n3363), .B1(n5397), .B2(n4730), .C(
        n3364), .ZN(n3977) );
  CKND0BWP12T U733 ( .I(n4524), .ZN(n3365) );
  MAOI22D0BWP12T U734 ( .A1(n4526), .A2(n3365), .B1(n4526), .B2(n4525), .ZN(
        n4707) );
  MAOI22D0BWP12T U735 ( .A1(n3466), .A2(n4025), .B1(n3466), .B2(n4025), .ZN(
        n3366) );
  MAOI22D0BWP12T U736 ( .A1(n3539), .A2(n3366), .B1(n3539), .B2(n3366), .ZN(
        n4024) );
  CKND0BWP12T U737 ( .I(n4025), .ZN(n3367) );
  MAOI222D0BWP12T U738 ( .A(n3466), .B(n3539), .C(n3367), .ZN(n4080) );
  CKND0BWP12T U739 ( .I(n3918), .ZN(n3368) );
  MAOI222D0BWP12T U740 ( .A(n3919), .B(n3920), .C(n3368), .ZN(n3921) );
  INR3D0BWP12T U741 ( .A1(n5762), .B1(n6887), .B2(n6862), .ZN(n6877) );
  IND2D0BWP12T U742 ( .A1(n6351), .B1(n6352), .ZN(n6851) );
  MAOI22D0BWP12T U743 ( .A1(n6334), .A2(n6516), .B1(n6334), .B2(n5434), .ZN(
        n6512) );
  MAOI22D0BWP12T U744 ( .A1(a[23]), .A2(n5806), .B1(a[23]), .B2(n5806), .ZN(
        n3369) );
  AOI22D0BWP12T U745 ( .A1(n5809), .A2(n5808), .B1(n5807), .B2(n3369), .ZN(
        n5824) );
  MUX2ND0BWP12T U746 ( .I0(n5407), .I1(n5406), .S(b[12]), .ZN(n3370) );
  MUX2ND0BWP12T U747 ( .I0(n5779), .I1(n5780), .S(b[13]), .ZN(n3371) );
  NR2D0BWP12T U748 ( .A1(n3370), .A2(n3371), .ZN(n5830) );
  AO222D0BWP12T U749 ( .A1(n6264), .A2(n5658), .B1(n6231), .B2(n5229), .C1(
        n5230), .C2(n6232), .Z(n6312) );
  INR2D0BWP12T U750 ( .A1(n6714), .B1(n6862), .ZN(n5590) );
  ND3D0BWP12T U751 ( .A1(n6343), .A2(n6344), .A3(n6342), .ZN(n3372) );
  NR4D0BWP12T U752 ( .A1(n6662), .A2(n6629), .A3(n6356), .A4(n3372), .ZN(n3373) );
  NR4D0BWP12T U753 ( .A1(n6341), .A2(n6687), .A3(n6340), .A4(n6385), .ZN(n3374) );
  ND3D0BWP12T U754 ( .A1(n6347), .A2(n3373), .A3(n3374), .ZN(n6349) );
  CKND0BWP12T U755 ( .I(n6411), .ZN(n3375) );
  OAI22D0BWP12T U756 ( .A1(n6409), .A2(n5680), .B1(n6410), .B2(n6223), .ZN(
        n3376) );
  OAI22D0BWP12T U757 ( .A1(n6408), .A2(n5681), .B1(n6407), .B2(n5291), .ZN(
        n3377) );
  NR2D0BWP12T U758 ( .A1(n3376), .A2(n3377), .ZN(n3378) );
  OA222D0BWP12T U759 ( .A1(n3375), .A2(n3378), .B1(n6400), .B2(n5441), .C1(
        n5623), .C2(n6417), .Z(n6431) );
  INR2D0BWP12T U760 ( .A1(n6504), .B1(n6505), .ZN(n6506) );
  INR3D0BWP12T U761 ( .A1(n6501), .B1(n6502), .B2(n6503), .ZN(n6507) );
  AOI21D0BWP12T U762 ( .A1(n6448), .A2(n5602), .B(n6500), .ZN(n3379) );
  MAOI22D0BWP12T U763 ( .A1(n3379), .A2(n5608), .B1(n3379), .B2(n5608), .ZN(
        n6144) );
  AOI22D0BWP12T U764 ( .A1(n4268), .A2(n6676), .B1(n6324), .B2(n6857), .ZN(
        n3380) );
  AOI211D0BWP12T U765 ( .A1(n6736), .A2(n4268), .B(n4265), .C(n4266), .ZN(
        n3381) );
  MAOI22D0BWP12T U766 ( .A1(n6833), .A2(n5946), .B1(n6193), .B2(n6794), .ZN(
        n3382) );
  OAI211D0BWP12T U767 ( .A1(n6289), .A2(n3380), .B(n3381), .C(n3382), .ZN(
        n3383) );
  AOI21D0BWP12T U768 ( .A1(n6909), .A2(n6367), .B(n3383), .ZN(n4271) );
  AOI21D0BWP12T U769 ( .A1(n6034), .A2(n6033), .B(n6035), .ZN(n6869) );
  ND4D0BWP12T U770 ( .A1(n5981), .A2(n6891), .A3(n5980), .A4(n6728), .ZN(n3384) );
  NR4D0BWP12T U771 ( .A1(n5982), .A2(n5983), .A3(n6799), .A4(n3384), .ZN(n3385) );
  ND4D0BWP12T U772 ( .A1(n6830), .A2(n3385), .A3(n6775), .A4(n5985), .ZN(n3386) );
  NR4D0BWP12T U773 ( .A1(n5987), .A2(n6729), .A3(n5986), .A4(n3386), .ZN(n3387) );
  IND4D0BWP12T U774 ( .A1(n5972), .B1(n5989), .B2(n5988), .B3(n3387), .ZN(
        n3388) );
  NR4D0BWP12T U775 ( .A1(n6694), .A2(n5991), .A3(n5990), .A4(n3388), .ZN(n3389) );
  ND4D0BWP12T U776 ( .A1(n5993), .A2(n5992), .A3(n6674), .A4(n3389), .ZN(n3390) );
  NR4D0BWP12T U777 ( .A1(n5996), .A2(n5995), .A3(n5994), .A4(n3390), .ZN(n3391) );
  ND4D0BWP12T U778 ( .A1(n5999), .A2(n5997), .A3(n5998), .A4(n3391), .ZN(n3392) );
  NR4D0BWP12T U779 ( .A1(n6000), .A2(n6001), .A3(n6831), .A4(n3392), .ZN(n6003) );
  MAOI222D0BWP12T U780 ( .A(n5752), .B(n5753), .C(n5754), .ZN(n3393) );
  MAOI22D0BWP12T U781 ( .A1(n5897), .A2(n5896), .B1(n5897), .B2(n5896), .ZN(
        n3394) );
  MAOI22D0BWP12T U782 ( .A1(n5895), .A2(n3394), .B1(n5895), .B2(n3394), .ZN(
        n3395) );
  MAOI222D0BWP12T U783 ( .A(n5788), .B(n5789), .C(n5790), .ZN(n3396) );
  MAOI22D0BWP12T U784 ( .A1(n5795), .A2(n3396), .B1(n5795), .B2(n3396), .ZN(
        n3397) );
  MAOI22D0BWP12T U785 ( .A1(n5796), .A2(n3397), .B1(n5796), .B2(n3397), .ZN(
        n3398) );
  MAOI22D0BWP12T U786 ( .A1(n5797), .A2(n3398), .B1(n5797), .B2(n3398), .ZN(
        n3399) );
  MAOI22D0BWP12T U787 ( .A1(n3395), .A2(n3399), .B1(n3395), .B2(n3399), .ZN(
        n3400) );
  MAOI22D0BWP12T U788 ( .A1(n5898), .A2(n3400), .B1(n5898), .B2(n3400), .ZN(
        n3401) );
  MAOI22D0BWP12T U789 ( .A1(n3393), .A2(n3401), .B1(n3393), .B2(n3401), .ZN(
        n3402) );
  MAOI22D0BWP12T U790 ( .A1(n5902), .A2(n3402), .B1(n5902), .B2(n3402), .ZN(
        n3403) );
  IOA21D0BWP12T U791 ( .A1(n5900), .A2(n5901), .B(n5899), .ZN(n3404) );
  MAOI22D0BWP12T U792 ( .A1(n3403), .A2(n3404), .B1(n3403), .B2(n3404), .ZN(
        n6609) );
  NR2D2BWP12T U793 ( .A1(n3613), .A2(n3431), .ZN(n4381) );
  NR2D2BWP12T U794 ( .A1(n3430), .A2(n4139), .ZN(n3613) );
  FA1D2BWP12T U795 ( .A(n3833), .B(n3832), .CI(n3831), .CO(n3828), .S(n3850)
         );
  FA1D0BWP12T U796 ( .A(n3818), .B(n3817), .CI(n3816), .CO(n3814), .S(n3833)
         );
  TPOAI21D1BWP12T U797 ( .A1(n5059), .A2(n5005), .B(n5004), .ZN(n5010) );
  ND4D1BWP12T U798 ( .A1(n4159), .A2(n4158), .A3(n4157), .A4(n4156), .ZN(n4164) );
  OAI211D1BWP12T U799 ( .A1(n4955), .A2(n6902), .B(n4954), .C(n4953), .ZN(
        result[3]) );
  INVD3BWP12T U800 ( .I(n4305), .ZN(n4829) );
  TPNR2D2BWP12T U801 ( .A1(n6239), .A2(n6819), .ZN(n4371) );
  INR2XD2BWP12T U802 ( .A1(n6239), .B1(n4136), .ZN(n3914) );
  TPAOI21D2BWP12T U803 ( .A1(n5560), .A2(n5556), .B(n3970), .ZN(n5142) );
  BUFFXD4BWP12T U804 ( .I(a[1]), .Z(n5360) );
  FA1D2BWP12T U805 ( .A(n3809), .B(n3808), .CI(n3807), .CO(n3975), .S(n3972)
         );
  FA1D2BWP12T U806 ( .A(n3830), .B(n3829), .CI(n3828), .CO(n3971), .S(n3969)
         );
  INR2XD2BWP12T U807 ( .A1(n5767), .B1(n4922), .ZN(n5661) );
  TPOAI21D1BWP12T U808 ( .A1(n6179), .A2(n6090), .B(n5267), .ZN(n5268) );
  NR2D2BWP12T U809 ( .A1(n5362), .A2(n4823), .ZN(n6488) );
  INVD2BWP12T U810 ( .I(n5237), .ZN(n6245) );
  ND2D8BWP12T U811 ( .A1(n4305), .A2(n3463), .ZN(n5237) );
  OAI211D1BWP12T U812 ( .A1(n5624), .A2(n6822), .B(n5132), .C(n5131), .ZN(
        n5133) );
  TPAOI21D1BWP12T U813 ( .A1(n5195), .A2(n4208), .B(n6460), .ZN(n4229) );
  OAI211D2BWP12T U814 ( .A1(n5101), .A2(n6836), .B(n5100), .C(n5099), .ZN(
        n5102) );
  TPNR2D3BWP12T U815 ( .A1(n4082), .A2(n6875), .ZN(n5979) );
  TPOAI21D1BWP12T U816 ( .A1(n4957), .A2(n5523), .B(n4958), .ZN(n4000) );
  ND2D4BWP12T U817 ( .A1(n4623), .A2(n6232), .ZN(n5870) );
  AN2XD2BWP12T U818 ( .A1(n3882), .A2(n6267), .Z(n3405) );
  OAI211D2BWP12T U819 ( .A1(n6891), .A2(n6890), .B(n6889), .C(n6888), .ZN(
        n6897) );
  INVD3BWP12T U820 ( .I(n6753), .ZN(n6888) );
  MUX2D1BWP12T U821 ( .I0(n5861), .I1(n5860), .S(n5612), .Z(n3915) );
  OAI211D0BWP12T U822 ( .A1(n6739), .A2(n6519), .B(n5746), .C(n6888), .ZN(
        n5748) );
  OAI211D0BWP12T U823 ( .A1(n6512), .A2(n6739), .B(n5548), .C(n5547), .ZN(
        n5549) );
  OAI22D0BWP12T U824 ( .A1(n6822), .A2(n6515), .B1(n5638), .B2(n5637), .ZN(
        n5639) );
  OAI22D0BWP12T U825 ( .A1(n6513), .A2(n6739), .B1(n6354), .B2(n6852), .ZN(
        n5190) );
  OA211D0BWP12T U826 ( .A1(n6514), .A2(n6822), .B(n5588), .C(n5587), .Z(n5592)
         );
  AOI21D0BWP12T U827 ( .A1(n6702), .A2(n6701), .B(n6739), .ZN(n6711) );
  OAI211D0BWP12T U828 ( .A1(b[12]), .A2(n6882), .B(n5579), .C(n6874), .ZN(
        n5582) );
  OA211D0BWP12T U829 ( .A1(n6518), .A2(n6822), .B(n4325), .C(n4324), .Z(n4332)
         );
  INVD2BWP12T U830 ( .I(n6822), .ZN(n6873) );
  DCCKND4BWP12T U831 ( .I(n6739), .ZN(n5578) );
  MUX2XD0BWP12T U832 ( .I0(n5878), .I1(n5877), .S(b[12]), .Z(n3469) );
  MUX2NXD1BWP12T U833 ( .I0(n5813), .I1(n5812), .S(b[12]), .ZN(n3682) );
  TPNR2D2BWP12T U834 ( .A1(b[12]), .A2(b[9]), .ZN(n4159) );
  DCCKND4BWP12T U835 ( .I(n4433), .ZN(n6782) );
  INVD3BWP12T U836 ( .I(b[5]), .ZN(n4433) );
  XNR2D2BWP12T U837 ( .A1(n4961), .A2(n4960), .ZN(n6052) );
  INVD2BWP12T U838 ( .I(n4357), .ZN(n5864) );
  AOI31D0BWP12T U839 ( .A1(n6296), .A2(n6295), .A3(n6294), .B(n6560), .ZN(
        n6375) );
  ND2XD4BWP12T U840 ( .A1(a[0]), .A2(n5360), .ZN(n6240) );
  FA1D2BWP12T U841 ( .A(n3989), .B(n3988), .CI(n3987), .CO(n3996), .S(n3976)
         );
  XOR3D2BWP12T U842 ( .A1(n3977), .A2(n3979), .A3(n3980), .Z(n3989) );
  AOI21D1BWP12T U843 ( .A1(n3974), .A2(n4226), .B(n3973), .ZN(n5600) );
  TPNR2D1BWP12T U844 ( .A1(n3940), .A2(n3939), .ZN(n6019) );
  XOR3D2BWP12T U845 ( .A1(n3569), .A2(n3568), .A3(n3567), .Z(n3650) );
  MUX2XD0BWP12T U846 ( .I0(n5759), .I1(n5758), .S(n5864), .Z(n4038) );
  MUX2XD0BWP12T U847 ( .I0(n5759), .I1(n5758), .S(b[12]), .Z(n4645) );
  MUX2XD0BWP12T U848 ( .I0(n5759), .I1(n5758), .S(n6334), .Z(n3433) );
  TPNR2D1BWP12T U849 ( .A1(n6185), .A2(n6794), .ZN(n5269) );
  INVD8BWP12T U850 ( .I(n4305), .ZN(n6248) );
  OA21D2BWP12T U851 ( .A1(n4013), .A2(n6055), .B(n4012), .Z(n3406) );
  CKND0BWP12T U852 ( .I(n3730), .ZN(n3713) );
  MUX2NXD1BWP12T U853 ( .I0(n4757), .I1(n4756), .S(b[16]), .ZN(n4422) );
  XOR3D2BWP12T U854 ( .A1(n3730), .A2(n3729), .A3(n3728), .Z(n3986) );
  MUX2NXD1BWP12T U855 ( .I0(n4757), .I1(n4756), .S(b[17]), .ZN(n4374) );
  BUFFD6BWP12T U856 ( .I(a[3]), .Z(n6247) );
  BUFFD3BWP12T U857 ( .I(n3507), .Z(n6576) );
  DCCKND4BWP12T U858 ( .I(b[1]), .ZN(n3463) );
  RCOAI22D2BWP12T U859 ( .A1(n4972), .A2(n5239), .B1(n5238), .B2(n6654), .ZN(
        n4246) );
  IND2XD8BWP12T U860 ( .A1(n5612), .B1(n6248), .ZN(n5238) );
  TPOAI21D2BWP12T U861 ( .A1(n4914), .A2(n3899), .B(n3898), .ZN(n5224) );
  TPND2D2BWP12T U862 ( .A1(n5222), .A2(n3892), .ZN(n4914) );
  TPAOI21D1BWP12T U863 ( .A1(n5105), .A2(n3408), .B(n3923), .ZN(n3940) );
  ND2XD4BWP12T U864 ( .A1(n3902), .A2(n6247), .ZN(n3911) );
  XOR2XD2BWP12T U865 ( .A1(a[2]), .A2(n5360), .Z(n3902) );
  OAI211D2BWP12T U866 ( .A1(n6902), .A2(n6732), .B(n6731), .C(n6730), .ZN(
        result[11]) );
  INVD4BWP12T U867 ( .I(n6264), .ZN(n4922) );
  TPNR2D3BWP12T U868 ( .A1(n4190), .A2(n4869), .ZN(n4186) );
  BUFFXD3BWP12T U869 ( .I(a[9]), .Z(n6229) );
  TPND2D4BWP12T U870 ( .A1(n3789), .A2(n6708), .ZN(n5775) );
  NR2XD3BWP12T U871 ( .A1(n4922), .A2(n6253), .ZN(n5662) );
  OAI222D0BWP12T U872 ( .A1(n5238), .A2(n4307), .B1(n3463), .B2(n4306), .C1(
        n4305), .C2(n5361), .ZN(n6036) );
  MUX2NXD1BWP12T U873 ( .I0(n5776), .I1(n5775), .S(n5612), .ZN(n3802) );
  MUX2XD0BWP12T U874 ( .I0(n3911), .I1(n5810), .S(n5612), .Z(n3885) );
  INVD1BWP12T U875 ( .I(b[4]), .ZN(n6357) );
  OR2XD1BWP12T U876 ( .A1(n3922), .A2(n3921), .Z(n3408) );
  INVD1BWP12T U877 ( .I(op[0]), .ZN(n4172) );
  NR2D1BWP12T U878 ( .A1(op[1]), .A2(n4172), .ZN(n4175) );
  CKAN2D0BWP12T U879 ( .A1(op[3]), .A2(op[2]), .Z(n4177) );
  ND2D1BWP12T U880 ( .A1(n4175), .A2(n4177), .ZN(n6902) );
  IND2XD2BWP12T U881 ( .A1(a[0]), .B1(n5360), .ZN(n5361) );
  INVD2BWP12T U882 ( .I(n5361), .ZN(n4557) );
  CKND0BWP12T U883 ( .I(b[19]), .ZN(n3411) );
  INVD1BWP12T U884 ( .I(b[20]), .ZN(n4494) );
  MUX2NXD0BWP12T U885 ( .I0(n4755), .I1(n6240), .S(n4494), .ZN(n3410) );
  AOI21D1BWP12T U886 ( .A1(n4557), .A2(n3411), .B(n3410), .ZN(n3449) );
  XOR2D1BWP12T U887 ( .A1(a[20]), .A2(a[19]), .Z(n3524) );
  INVD1BWP12T U888 ( .I(b[0]), .ZN(n3420) );
  BUFFD2BWP12T U889 ( .I(n3420), .Z(n3934) );
  INVD4BWP12T U890 ( .I(n3934), .ZN(n4823) );
  ND2D1BWP12T U891 ( .A1(n3524), .A2(n4823), .ZN(n3448) );
  INVD1BWP12T U892 ( .I(n6247), .ZN(n5254) );
  ND2D1BWP12T U893 ( .A1(n3902), .A2(n5254), .ZN(n3412) );
  BUFFD3BWP12T U894 ( .I(n3412), .Z(n5810) );
  MUX2ND0BWP12T U895 ( .I0(n5811), .I1(n5810), .S(b[18]), .ZN(n3414) );
  INVD2BWP12T U896 ( .I(n4935), .ZN(n5813) );
  MUX2ND0BWP12T U897 ( .I0(n5813), .I1(n5812), .S(b[17]), .ZN(n3413) );
  NR2D1BWP12T U898 ( .A1(n3414), .A2(n3413), .ZN(n3447) );
  ND2D1BWP12T U899 ( .A1(a[17]), .A2(a[18]), .ZN(n3421) );
  NR2D1BWP12T U900 ( .A1(n3421), .A2(a[19]), .ZN(n5781) );
  IND2D1BWP12T U901 ( .A1(a[18]), .B1(a[19]), .ZN(n3415) );
  NR2D1BWP12T U902 ( .A1(n3415), .A2(a[17]), .ZN(n5782) );
  NR2D1BWP12T U903 ( .A1(n5781), .A2(n5782), .ZN(n3489) );
  INVD3BWP12T U904 ( .I(n3463), .ZN(n4498) );
  XOR2D1BWP12T U905 ( .A1(a[17]), .A2(a[18]), .Z(n3487) );
  ND2D1BWP12T U906 ( .A1(n3487), .A2(a[19]), .ZN(n5779) );
  INVD1BWP12T U907 ( .I(a[19]), .ZN(n6654) );
  ND2D1BWP12T U908 ( .A1(n3487), .A2(n6654), .ZN(n5780) );
  INVD1BWP12T U909 ( .I(b[2]), .ZN(n3477) );
  BUFFD2BWP12T U910 ( .I(n3477), .Z(n5767) );
  INVD2BWP12T U911 ( .I(n5767), .ZN(n5247) );
  IAO21D1BWP12T U912 ( .A1(n3489), .A2(n3490), .B(n3416), .ZN(n3493) );
  BUFFD2BWP12T U913 ( .I(a[4]), .Z(n6249) );
  ND2D1BWP12T U914 ( .A1(n6249), .A2(n6247), .ZN(n3417) );
  TPNR2D1BWP12T U915 ( .A1(n6249), .A2(n6247), .ZN(n4135) );
  INR2D2BWP12T U916 ( .A1(n3417), .B1(n4135), .ZN(n3882) );
  BUFFD2BWP12T U917 ( .I(a[5]), .Z(n6267) );
  INVD1BWP12T U918 ( .I(n6267), .ZN(n6788) );
  AN2XD2BWP12T U919 ( .A1(n3882), .A2(n6788), .Z(n5395) );
  INVD1BWP12T U920 ( .I(n5395), .ZN(n5858) );
  MUX2ND0BWP12T U921 ( .I0(n5859), .I1(n5858), .S(b[15]), .ZN(n3419) );
  CKND2D2BWP12T U922 ( .A1(n4135), .A2(n6267), .ZN(n5861) );
  NR2D1BWP12T U923 ( .A1(n3417), .A2(n6267), .ZN(n5396) );
  MUX2ND0BWP12T U924 ( .I0(n5861), .I1(n5860), .S(b[14]), .ZN(n3418) );
  NR2D1BWP12T U925 ( .A1(n3419), .A2(n3418), .ZN(n3572) );
  BUFFD3BWP12T U926 ( .I(n3420), .Z(n4305) );
  IND2D1BWP12T U927 ( .A1(n6248), .B1(a[19]), .ZN(n3488) );
  INVD1BWP12T U928 ( .I(n3488), .ZN(n3422) );
  AOI21D1BWP12T U929 ( .A1(n3422), .A2(n3421), .B(n5782), .ZN(n3571) );
  CKND0BWP12T U930 ( .I(b[17]), .ZN(n3424) );
  INVD1BWP12T U931 ( .I(b[18]), .ZN(n4112) );
  MUX2ND0BWP12T U932 ( .I0(n4755), .I1(n6240), .S(n4112), .ZN(n3423) );
  AOI21D1BWP12T U933 ( .A1(n4557), .A2(n3424), .B(n3423), .ZN(n3575) );
  ND2D1BWP12T U934 ( .A1(n3487), .A2(n4823), .ZN(n3574) );
  MUX2ND0BWP12T U935 ( .I0(n5811), .I1(n5810), .S(b[16]), .ZN(n3426) );
  MUX2ND0BWP12T U936 ( .I0(n5813), .I1(n5812), .S(b[15]), .ZN(n3425) );
  NR2D1BWP12T U937 ( .A1(n3426), .A2(n3425), .ZN(n3573) );
  BUFFD2BWP12T U938 ( .I(a[11]), .Z(n6230) );
  XOR2XD2BWP12T U939 ( .A1(n6231), .A2(n6230), .Z(n4390) );
  ND2D1BWP12T U940 ( .A1(n4390), .A2(a[13]), .ZN(n5817) );
  INVD1BWP12T U941 ( .I(a[13]), .ZN(n4286) );
  CKND2D4BWP12T U942 ( .A1(n4390), .A2(n4286), .ZN(n5816) );
  MUX2NXD0BWP12T U943 ( .I0(n5817), .I1(n5816), .S(b[9]), .ZN(n3429) );
  TPNR2D0BWP12T U944 ( .A1(n6231), .A2(n6230), .ZN(n3427) );
  ND2D1BWP12T U945 ( .A1(n3427), .A2(a[13]), .ZN(n5819) );
  ND3D1BWP12T U946 ( .A1(n4286), .A2(n6231), .A3(n6230), .ZN(n5818) );
  BUFFD2BWP12T U947 ( .I(b[8]), .Z(n5843) );
  MUX2NXD0BWP12T U948 ( .I0(n5819), .I1(n5818), .S(n5843), .ZN(n3428) );
  NR2D1BWP12T U949 ( .A1(n3429), .A2(n3428), .ZN(n3505) );
  ND2D1BWP12T U950 ( .A1(a[6]), .A2(n6267), .ZN(n6239) );
  TPNR2D1BWP12T U951 ( .A1(a[6]), .A2(n6267), .ZN(n4136) );
  BUFFD6BWP12T U952 ( .I(a[7]), .Z(n6819) );
  TPND2D2BWP12T U953 ( .A1(n3914), .A2(n6819), .ZN(n5876) );
  INVD2BWP12T U954 ( .I(n6819), .ZN(n5236) );
  ND2XD4BWP12T U955 ( .A1(n3914), .A2(n5236), .ZN(n5875) );
  TPND2D1BWP12T U956 ( .A1(n4136), .A2(n6819), .ZN(n5878) );
  BUFFXD4BWP12T U957 ( .I(a[15]), .Z(n6232) );
  AN2XD2BWP12T U958 ( .A1(a[16]), .A2(n6232), .Z(n3430) );
  NR2D1BWP12T U959 ( .A1(a[16]), .A2(n6232), .ZN(n4139) );
  INVD1BWP12T U960 ( .I(n6228), .ZN(n3431) );
  ND2D1BWP12T U961 ( .A1(n4381), .A2(a[17]), .ZN(n5759) );
  INVD1BWP12T U962 ( .I(b[3]), .ZN(n3507) );
  BUFFD2BWP12T U963 ( .I(n3507), .Z(n4924) );
  INVD6BWP12T U964 ( .I(n4924), .ZN(n6334) );
  ND2D1BWP12T U965 ( .A1(n3613), .A2(a[17]), .ZN(n5761) );
  INVD1BWP12T U966 ( .I(a[17]), .ZN(n5728) );
  ND2D1BWP12T U967 ( .A1(n3613), .A2(n5728), .ZN(n5760) );
  INVD4BWP12T U968 ( .I(n6357), .ZN(n6573) );
  MUX2D1BWP12T U969 ( .I0(n5761), .I1(n5760), .S(n6573), .Z(n3432) );
  ND2D1BWP12T U970 ( .A1(n3433), .A2(n3432), .ZN(n3482) );
  MUX2D1BWP12T U971 ( .I0(n5817), .I1(n5816), .S(n5843), .Z(n3435) );
  BUFFD2BWP12T U972 ( .I(b[7]), .Z(n5379) );
  MUX2D1BWP12T U973 ( .I0(n5819), .I1(n5818), .S(n5379), .Z(n3434) );
  ND2D1BWP12T U974 ( .A1(n3435), .A2(n3434), .ZN(n3483) );
  MAOI222D1BWP12T U975 ( .A(n3484), .B(n3482), .C(n3483), .ZN(n3504) );
  MUX2ND0BWP12T U976 ( .I0(n5779), .I1(n5780), .S(n6334), .ZN(n3437) );
  INVD1BWP12T U977 ( .I(n5781), .ZN(n5406) );
  INVD1BWP12T U978 ( .I(n5782), .ZN(n5407) );
  MUX2NXD0BWP12T U979 ( .I0(n5406), .I1(n5407), .S(n5767), .ZN(n3436) );
  NR2D1BWP12T U980 ( .A1(n3437), .A2(n3436), .ZN(n3530) );
  ND2D1BWP12T U981 ( .A1(a[14]), .A2(a[13]), .ZN(n6238) );
  NR2D1BWP12T U982 ( .A1(a[14]), .A2(a[13]), .ZN(n3438) );
  INR2D2BWP12T U983 ( .A1(n6238), .B1(n3438), .ZN(n4623) );
  INVD1BWP12T U984 ( .I(n6232), .ZN(n5538) );
  CKND2D3BWP12T U985 ( .A1(n4623), .A2(n5538), .ZN(n5869) );
  MUX2NXD0BWP12T U986 ( .I0(n5870), .I1(n5869), .S(n5379), .ZN(n3440) );
  NR2D1BWP12T U987 ( .A1(n6238), .A2(n6232), .ZN(n3608) );
  INVD1BWP12T U988 ( .I(n3608), .ZN(n5871) );
  INVD1BWP12T U989 ( .I(b[6]), .ZN(n4357) );
  MUX2ND0BWP12T U990 ( .I0(n5871), .I1(n5872), .S(n4357), .ZN(n3439) );
  NR2D1BWP12T U991 ( .A1(n3440), .A2(n3439), .ZN(n3529) );
  MUX2ND0BWP12T U992 ( .I0(n5859), .I1(n5858), .S(b[17]), .ZN(n3442) );
  INVD1BWP12T U993 ( .I(b[16]), .ZN(n4092) );
  MUX2ND0BWP12T U994 ( .I0(n5860), .I1(n5861), .S(n4092), .ZN(n3441) );
  NR2D1BWP12T U995 ( .A1(n3442), .A2(n3441), .ZN(n3528) );
  XOR3D1BWP12T U996 ( .A1(n3505), .A2(n3504), .A3(n3503), .Z(n3581) );
  ND2D1BWP12T U997 ( .A1(n3524), .A2(a[21]), .ZN(n5803) );
  NR2D1BWP12T U998 ( .A1(a[20]), .A2(a[19]), .ZN(n3443) );
  ND2D1BWP12T U999 ( .A1(n3443), .A2(a[21]), .ZN(n5805) );
  OAI21D1BWP12T U1000 ( .A1(n5803), .A2(n4829), .B(n5805), .ZN(n3516) );
  INVD2BWP12T U1001 ( .I(n6230), .ZN(n6708) );
  INVD1BWP12T U1002 ( .I(b[11]), .ZN(n4745) );
  ND2D1BWP12T U1003 ( .A1(n6708), .A2(n4745), .ZN(n6703) );
  ND2D1BWP12T U1004 ( .A1(n6230), .A2(b[11]), .ZN(n6706) );
  ND2D1BWP12T U1005 ( .A1(n6703), .A2(n6706), .ZN(n6707) );
  INVD1BWP12T U1006 ( .I(n6707), .ZN(n5941) );
  BUFFD3BWP12T U1007 ( .I(a[10]), .Z(n6715) );
  XOR2XD8BWP12T U1008 ( .A1(n6715), .A2(n6229), .Z(n3789) );
  ND2D1BWP12T U1009 ( .A1(n5941), .A2(n3789), .ZN(n3446) );
  ND3D2BWP12T U1010 ( .A1(n6708), .A2(n6715), .A3(n6229), .ZN(n5777) );
  CKND1BWP12T U1011 ( .I(n5777), .ZN(n3444) );
  BUFFD2BWP12T U1012 ( .I(b[10]), .Z(n5806) );
  NR2D1BWP12T U1013 ( .A1(n6715), .A2(n5806), .ZN(n4259) );
  NR2D1BWP12T U1014 ( .A1(n6708), .A2(n6229), .ZN(n3454) );
  AOI22D1BWP12T U1015 ( .A1(n3444), .A2(n5806), .B1(n4259), .B2(n3454), .ZN(
        n3445) );
  ND2D1BWP12T U1016 ( .A1(n3446), .A2(n3445), .ZN(n3517) );
  FA1D0BWP12T U1017 ( .A(n3449), .B(n3448), .CI(n3447), .CO(n3502), .S(n3494)
         );
  MUX2ND0BWP12T U1018 ( .I0(n5859), .I1(n5858), .S(b[16]), .ZN(n3451) );
  INVD1BWP12T U1019 ( .I(b[15]), .ZN(n3666) );
  MUX2ND0BWP12T U1020 ( .I0(n5860), .I1(n5861), .S(n3666), .ZN(n3450) );
  NR2D1BWP12T U1021 ( .A1(n3451), .A2(n3450), .ZN(n3475) );
  MUX2NXD0BWP12T U1022 ( .I0(n5870), .I1(n5869), .S(n5864), .ZN(n3453) );
  MUX2ND0BWP12T U1023 ( .I0(n5871), .I1(n5872), .S(n4433), .ZN(n3452) );
  NR2D1BWP12T U1024 ( .A1(n3453), .A2(n3452), .ZN(n3474) );
  ND2XD8BWP12T U1025 ( .A1(n3789), .A2(n6230), .ZN(n5776) );
  MUX2ND0BWP12T U1026 ( .I0(n5776), .I1(n5775), .S(n5806), .ZN(n3456) );
  INVD1BWP12T U1027 ( .I(n6715), .ZN(n5232) );
  CKND2D2BWP12T U1028 ( .A1(n3454), .A2(n5232), .ZN(n5778) );
  MUX2ND0BWP12T U1029 ( .I0(n5778), .I1(n5777), .S(b[9]), .ZN(n3455) );
  NR2D1BWP12T U1030 ( .A1(n3456), .A2(n3455), .ZN(n3473) );
  CKND1BWP12T U1031 ( .I(b[21]), .ZN(n4758) );
  NR2D1BWP12T U1032 ( .A1(n5361), .A2(b[20]), .ZN(n3457) );
  NR2D1BWP12T U1033 ( .A1(n3458), .A2(n3457), .ZN(n3460) );
  NR2D1BWP12T U1034 ( .A1(n3459), .A2(n3460), .ZN(n4065) );
  AO21D1BWP12T U1035 ( .A1(n3460), .A2(n3459), .B(n4065), .Z(n3514) );
  MUX2NXD1BWP12T U1036 ( .I0(n5876), .I1(n5875), .S(b[15]), .ZN(n3462) );
  MUX2ND0BWP12T U1037 ( .I0(n5878), .I1(n5877), .S(b[14]), .ZN(n3461) );
  NR2D1BWP12T U1038 ( .A1(n3462), .A2(n3461), .ZN(n3512) );
  INVD1BWP12T U1039 ( .I(a[21]), .ZN(n6623) );
  ND3D1BWP12T U1040 ( .A1(n6623), .A2(a[20]), .A3(a[19]), .ZN(n5804) );
  CKND2D1BWP12T U1041 ( .A1(n5804), .A2(n5805), .ZN(n3526) );
  MUX2D1BWP12T U1042 ( .I0(a[21]), .I1(a[20]), .S(n6248), .Z(n6535) );
  CKBD1BWP12T U1043 ( .I(n3463), .Z(n4815) );
  INVD4BWP12T U1044 ( .I(n4815), .ZN(n5612) );
  CKXOR2D1BWP12T U1045 ( .A1(a[21]), .A2(n5612), .Z(n3527) );
  AOI22D1BWP12T U1046 ( .A1(n3526), .A2(n6535), .B1(n3524), .B2(n3527), .ZN(
        n3511) );
  INVD1P75BWP12T U1047 ( .I(a[8]), .ZN(n6760) );
  ND2D1BWP12T U1048 ( .A1(n5236), .A2(n6760), .ZN(n6756) );
  ND2D1BWP12T U1049 ( .A1(n6819), .A2(a[8]), .ZN(n6237) );
  ND2D1BWP12T U1050 ( .A1(n6756), .A2(n6237), .ZN(n3597) );
  INR2D2BWP12T U1051 ( .A1(n6229), .B1(n3597), .ZN(n4757) );
  INVD1BWP12T U1052 ( .I(n4757), .ZN(n5837) );
  INVD1BWP12T U1053 ( .I(n6229), .ZN(n5231) );
  INR2D2BWP12T U1054 ( .A1(n5231), .B1(n3597), .ZN(n4756) );
  MUX2ND0BWP12T U1055 ( .I0(n5837), .I1(n5836), .S(b[13]), .ZN(n3465) );
  TPNR2D1BWP12T U1056 ( .A1(n6756), .A2(n5231), .ZN(n4759) );
  INVD1BWP12T U1057 ( .I(n4759), .ZN(n5839) );
  NR2D1BWP12T U1058 ( .A1(n6237), .A2(n6229), .ZN(n4760) );
  INVD1BWP12T U1059 ( .I(n4760), .ZN(n5838) );
  INVD1BWP12T U1060 ( .I(b[12]), .ZN(n4497) );
  MUX2NXD1BWP12T U1061 ( .I0(n5839), .I1(n5838), .S(b[12]), .ZN(n3464) );
  NR2D1BWP12T U1062 ( .A1(n3465), .A2(n3464), .ZN(n3510) );
  INVD1BWP12T U1063 ( .I(n3498), .ZN(n3476) );
  MUX2D1BWP12T U1064 ( .I0(n5776), .I1(n5775), .S(b[9]), .Z(n3468) );
  INVD1BWP12T U1065 ( .I(n5843), .ZN(n4515) );
  MUX2D1BWP12T U1066 ( .I0(n5777), .I1(n5778), .S(n4515), .Z(n3467) );
  ND2D1BWP12T U1067 ( .A1(n3468), .A2(n3467), .ZN(n3552) );
  MUX2D1BWP12T U1068 ( .I0(n5876), .I1(n5875), .S(b[13]), .Z(n3470) );
  ND2D1BWP12T U1069 ( .A1(n3470), .A2(n3469), .ZN(n3551) );
  MUX2D1BWP12T U1070 ( .I0(n3911), .I1(n5810), .S(b[17]), .Z(n3472) );
  MUX2D1BWP12T U1071 ( .I0(n5813), .I1(n5812), .S(b[16]), .Z(n3471) );
  ND2D1BWP12T U1072 ( .A1(n3472), .A2(n3471), .ZN(n3550) );
  MAOI222D1BWP12T U1073 ( .A(n3552), .B(n3551), .C(n3550), .ZN(n3497) );
  FA1D0BWP12T U1074 ( .A(n3475), .B(n3474), .CI(n3473), .CO(n3515), .S(n3496)
         );
  MAOI222D1BWP12T U1075 ( .A(n3476), .B(n3497), .C(n3496), .ZN(n3542) );
  MUX2D1BWP12T U1076 ( .I0(n5759), .I1(n5758), .S(n6520), .Z(n3479) );
  MUX2D1BWP12T U1077 ( .I0(n5761), .I1(n5760), .S(n6334), .Z(n3478) );
  ND2D1BWP12T U1078 ( .A1(n3479), .A2(n3478), .ZN(n3555) );
  MUX2XD0BWP12T U1079 ( .I0(n6240), .I1(n4755), .S(b[19]), .Z(n3481) );
  ND2D1BWP12T U1080 ( .A1(n4557), .A2(n4112), .ZN(n3480) );
  ND2D1BWP12T U1081 ( .A1(n3481), .A2(n3480), .ZN(n3554) );
  ND2D1BWP12T U1082 ( .A1(n3555), .A2(n3554), .ZN(n3553) );
  XNR3D1BWP12T U1083 ( .A1(n3484), .A2(n3483), .A3(n3482), .ZN(n3499) );
  MUX2D1BWP12T U1084 ( .I0(n5817), .I1(n5816), .S(n5379), .Z(n3486) );
  MUX2D1BWP12T U1085 ( .I0(n5819), .I1(n5818), .S(n5864), .Z(n3485) );
  ND2D1BWP12T U1086 ( .A1(n3486), .A2(n3485), .ZN(n3558) );
  INVD1BWP12T U1087 ( .I(n3487), .ZN(n3491) );
  ND2D1BWP12T U1088 ( .A1(a[18]), .A2(n4823), .ZN(n4921) );
  ND2D1BWP12T U1089 ( .A1(n3488), .A2(n4921), .ZN(n6532) );
  INVD1BWP12T U1090 ( .I(n6532), .ZN(n5035) );
  OAI22D1BWP12T U1091 ( .A1(n3491), .A2(n3490), .B1(n3489), .B2(n5035), .ZN(
        n3559) );
  MAOI222D1BWP12T U1092 ( .A(n3558), .B(n3557), .C(n3559), .ZN(n3500) );
  MAOI222D1BWP12T U1093 ( .A(n3553), .B(n3499), .C(n3500), .ZN(n3541) );
  FA1D0BWP12T U1094 ( .A(n3494), .B(n3493), .CI(n3492), .CO(n3582), .S(n3495)
         );
  INVD1BWP12T U1095 ( .I(n3495), .ZN(n3586) );
  XOR3D1BWP12T U1096 ( .A1(n3498), .A2(n3497), .A3(n3496), .Z(n3585) );
  XNR3D1BWP12T U1097 ( .A1(n3553), .A2(n3500), .A3(n3499), .ZN(n3584) );
  MAOI222D1BWP12T U1098 ( .A(n3505), .B(n3504), .C(n3503), .ZN(n3506) );
  INVD1BWP12T U1099 ( .I(n3506), .ZN(n4076) );
  XOR3D1BWP12T U1100 ( .A1(n4041), .A2(n4042), .A3(n4043), .Z(n4058) );
  MUX2ND0BWP12T U1101 ( .I0(n5837), .I1(n5836), .S(b[14]), .ZN(n3509) );
  MUX2NXD0BWP12T U1102 ( .I0(n5839), .I1(n5838), .S(b[13]), .ZN(n3508) );
  NR2D1BWP12T U1103 ( .A1(n3509), .A2(n3508), .ZN(n4057) );
  FA1D0BWP12T U1104 ( .A(n3512), .B(n3511), .CI(n3510), .CO(n4056), .S(n3513)
         );
  FA1D0BWP12T U1105 ( .A(n3515), .B(n3514), .CI(n3513), .CO(n4050), .S(n3501)
         );
  CKND2D1BWP12T U1106 ( .A1(n3517), .A2(n3516), .ZN(n3519) );
  NR2D1BWP12T U1107 ( .A1(n3517), .A2(n3516), .ZN(n3518) );
  AOI21D1BWP12T U1108 ( .A1(n3520), .A2(n3519), .B(n3518), .ZN(n4063) );
  AOI21D1BWP12T U1109 ( .A1(n4557), .A2(n4758), .B(n3521), .ZN(n4028) );
  XOR2D1BWP12T U1110 ( .A1(a[22]), .A2(a[21]), .Z(n5807) );
  ND2D1BWP12T U1111 ( .A1(n5807), .A2(n4823), .ZN(n4027) );
  MUX2NXD0BWP12T U1112 ( .I0(n5870), .I1(n5869), .S(n5843), .ZN(n3523) );
  INVD1BWP12T U1113 ( .I(n5379), .ZN(n4343) );
  MUX2NXD0BWP12T U1114 ( .I0(n5871), .I1(n5872), .S(n4343), .ZN(n3522) );
  NR2D1BWP12T U1115 ( .A1(n3523), .A2(n3522), .ZN(n4026) );
  ND2D1BWP12T U1116 ( .A1(n3524), .A2(n6623), .ZN(n5802) );
  MUX2NXD0BWP12T U1117 ( .I0(n5803), .I1(n5802), .S(n5247), .ZN(n3525) );
  AOI21D1BWP12T U1118 ( .A1(n3527), .A2(n3526), .B(n3525), .ZN(n4053) );
  FA1D0BWP12T U1119 ( .A(n3530), .B(n3529), .CI(n3528), .CO(n4061), .S(n3503)
         );
  MUX2ND0BWP12T U1120 ( .I0(n5811), .I1(n5810), .S(b[20]), .ZN(n3532) );
  MUX2ND0BWP12T U1121 ( .I0(n5813), .I1(n5812), .S(b[19]), .ZN(n3531) );
  NR2D1BWP12T U1122 ( .A1(n3532), .A2(n3531), .ZN(n4060) );
  MUX2ND0BWP12T U1123 ( .I0(n5817), .I1(n5816), .S(n5806), .ZN(n3534) );
  MUX2NXD0BWP12T U1124 ( .I0(n5819), .I1(n5818), .S(b[9]), .ZN(n3533) );
  NR2D1BWP12T U1125 ( .A1(n3534), .A2(n3533), .ZN(n4072) );
  MUX2ND0BWP12T U1126 ( .I0(n5876), .I1(n5875), .S(b[16]), .ZN(n3536) );
  MUX2ND0BWP12T U1127 ( .I0(n5877), .I1(n5878), .S(n3666), .ZN(n3535) );
  NR2D1BWP12T U1128 ( .A1(n3536), .A2(n3535), .ZN(n4074) );
  MUX2ND0BWP12T U1129 ( .I0(n5761), .I1(n5760), .S(n5864), .ZN(n3537) );
  NR2D1BWP12T U1130 ( .A1(n3538), .A2(n3537), .ZN(n4073) );
  XOR3D1BWP12T U1131 ( .A1(n4072), .A2(n4074), .A3(n4073), .Z(n4059) );
  XOR3D1BWP12T U1132 ( .A1(n4054), .A2(n4053), .A3(n4052), .Z(n4049) );
  FA1D0BWP12T U1133 ( .A(n3542), .B(n3541), .CI(n3540), .CO(n4025), .S(n3543)
         );
  INVD1BWP12T U1134 ( .I(n3543), .ZN(n4016) );
  MUX2ND0BWP12T U1135 ( .I0(n5859), .I1(n5858), .S(b[14]), .ZN(n3545) );
  INVD1BWP12T U1136 ( .I(b[13]), .ZN(n4576) );
  MUX2D1BWP12T U1137 ( .I0(n5396), .I1(n5397), .S(n4576), .Z(n3544) );
  NR2D1BWP12T U1138 ( .A1(n3545), .A2(n3544), .ZN(n3600) );
  MUX2ND0BWP12T U1139 ( .I0(n5776), .I1(n5775), .S(n5843), .ZN(n3547) );
  MUX2ND0BWP12T U1140 ( .I0(n5778), .I1(n5777), .S(n5379), .ZN(n3546) );
  NR2D1BWP12T U1141 ( .A1(n3547), .A2(n3546), .ZN(n3601) );
  MUX2NXD0BWP12T U1142 ( .I0(n5870), .I1(n5869), .S(n6573), .ZN(n3549) );
  CKND1BWP12T U1143 ( .I(n5872), .ZN(n3609) );
  MUX2XD0BWP12T U1144 ( .I0(n3608), .I1(n3609), .S(n6576), .Z(n3548) );
  NR2D1BWP12T U1145 ( .A1(n3549), .A2(n3548), .ZN(n3599) );
  FCICOND1BWP12T U1146 ( .A(n3600), .B(n3601), .CI(n3599), .CON(n3568) );
  OAI21D1BWP12T U1147 ( .A1(n3555), .A2(n3554), .B(n3553), .ZN(n3569) );
  INVD1BWP12T U1148 ( .I(n3569), .ZN(n3556) );
  MAOI222D1BWP12T U1149 ( .A(n3568), .B(n3567), .C(n3556), .ZN(n3621) );
  XOR3D1BWP12T U1150 ( .A1(n3559), .A2(n3558), .A3(n3557), .Z(n3588) );
  MUX2ND0BWP12T U1151 ( .I0(n5761), .I1(n5760), .S(n5247), .ZN(n3560) );
  NR2D1BWP12T U1152 ( .A1(n3561), .A2(n3560), .ZN(n3591) );
  ND2D1BWP12T U1153 ( .A1(n6229), .A2(b[9]), .ZN(n6111) );
  NR2D1BWP12T U1154 ( .A1(n6229), .A2(b[9]), .ZN(n4238) );
  INR2D1BWP12T U1155 ( .A1(n6111), .B1(n4238), .ZN(n5204) );
  ND2D1BWP12T U1156 ( .A1(n5839), .A2(n5838), .ZN(n3845) );
  MUX2ND0BWP12T U1157 ( .I0(n5837), .I1(n5836), .S(n5806), .ZN(n3562) );
  AOI21D1BWP12T U1158 ( .A1(n5204), .A2(n3845), .B(n3562), .ZN(n3590) );
  MUX2ND0BWP12T U1159 ( .I0(n5817), .I1(n5816), .S(b[6]), .ZN(n3564) );
  MUX2ND0BWP12T U1160 ( .I0(n5819), .I1(n5818), .S(n6782), .ZN(n3563) );
  NR2D1BWP12T U1161 ( .A1(n3564), .A2(n3563), .ZN(n3592) );
  MAOI222D1BWP12T U1162 ( .A(n3591), .B(n3590), .C(n3592), .ZN(n3587) );
  INVD1BWP12T U1163 ( .I(n3589), .ZN(n3565) );
  OAI22D1BWP12T U1164 ( .A1(n3566), .A2(n3587), .B1(n3588), .B2(n3565), .ZN(
        n3620) );
  FA1D0BWP12T U1165 ( .A(n3572), .B(n3571), .CI(n3570), .CO(n3492), .S(n3649)
         );
  FA1D0BWP12T U1166 ( .A(n3575), .B(n3574), .CI(n3573), .CO(n3570), .S(n3617)
         );
  INVD1BWP12T U1167 ( .I(n6240), .ZN(n4647) );
  INVD1BWP12T U1168 ( .I(n4755), .ZN(n4646) );
  MUX2ND0BWP12T U1169 ( .I0(n4647), .I1(n4646), .S(b[17]), .ZN(n3576) );
  OAI21D1BWP12T U1170 ( .A1(b[16]), .A2(n5361), .B(n3576), .ZN(n3625) );
  ND2D1BWP12T U1171 ( .A1(n3625), .A2(n3626), .ZN(n3624) );
  MUX2D1BWP12T U1172 ( .I0(a[17]), .I1(a[16]), .S(n6248), .Z(n6403) );
  MUX2ND0BWP12T U1173 ( .I0(n5761), .I1(n5760), .S(n5612), .ZN(n3577) );
  MUX2ND0BWP12T U1174 ( .I0(n5776), .I1(n5775), .S(n5379), .ZN(n3579) );
  MUX2ND0BWP12T U1175 ( .I0(n5778), .I1(n5777), .S(n5864), .ZN(n3578) );
  FA1D0BWP12T U1176 ( .A(n3582), .B(n3581), .CI(n3580), .CO(n3466), .S(n4014)
         );
  INVD1BWP12T U1177 ( .I(n3583), .ZN(n4023) );
  NR2D1BWP12T U1178 ( .A1(n4024), .A2(n4023), .ZN(n5454) );
  FA1D0BWP12T U1179 ( .A(n3586), .B(n3585), .CI(n3584), .CO(n3540), .S(n4020)
         );
  XNR3XD2BWP12T U1180 ( .A1(n3589), .A2(n3588), .A3(n3587), .ZN(n3653) );
  INVD1BWP12T U1181 ( .I(n5878), .ZN(n4372) );
  XOR3D1BWP12T U1182 ( .A1(n3592), .A2(n3591), .A3(n3590), .Z(n3635) );
  INVD1BWP12T U1183 ( .I(n5806), .ZN(n5405) );
  MUX2D1BWP12T U1184 ( .I0(n4371), .I1(n4372), .S(n5405), .Z(n3593) );
  NR2D1BWP12T U1185 ( .A1(n3594), .A2(n3593), .ZN(n3628) );
  MUX2ND0BWP12T U1186 ( .I0(n5859), .I1(n5858), .S(b[13]), .ZN(n3596) );
  MUX2D1BWP12T U1187 ( .I0(n5396), .I1(n5397), .S(n4497), .Z(n3595) );
  NR2D1BWP12T U1188 ( .A1(n3596), .A2(n3595), .ZN(n3627) );
  ND2D1BWP12T U1189 ( .A1(n6760), .A2(n4515), .ZN(n4231) );
  ND2D1BWP12T U1190 ( .A1(a[8]), .A2(n5843), .ZN(n6093) );
  ND2D1BWP12T U1191 ( .A1(n4231), .A2(n6093), .ZN(n6175) );
  INVD1BWP12T U1192 ( .I(n3597), .ZN(n3859) );
  AOI22D1BWP12T U1193 ( .A1(n3845), .A2(n6175), .B1(n5204), .B2(n3859), .ZN(
        n3629) );
  MAOI222D1BWP12T U1194 ( .A(n3628), .B(n3627), .C(n3629), .ZN(n3636) );
  INVD1BWP12T U1195 ( .I(n3636), .ZN(n3598) );
  MAOI222D1BWP12T U1196 ( .A(n3637), .B(n3635), .C(n3598), .ZN(n3652) );
  INVD1BWP12T U1197 ( .I(n5817), .ZN(n3742) );
  CKND0BWP12T U1198 ( .I(n5816), .ZN(n3602) );
  MUX2ND0BWP12T U1199 ( .I0(n3742), .I1(n3602), .S(n6782), .ZN(n3605) );
  INVD1BWP12T U1200 ( .I(n5819), .ZN(n3741) );
  CKND1BWP12T U1201 ( .I(n5818), .ZN(n3603) );
  MUX2NXD0BWP12T U1202 ( .I0(n3741), .I1(n3603), .S(n6573), .ZN(n3604) );
  CKND2D1BWP12T U1203 ( .A1(n3605), .A2(n3604), .ZN(n3646) );
  CKND0BWP12T U1204 ( .I(n5870), .ZN(n3607) );
  CKND0BWP12T U1205 ( .I(n5869), .ZN(n3606) );
  MUX2ND0BWP12T U1206 ( .I0(n3607), .I1(n3606), .S(n6334), .ZN(n3611) );
  MUX2NXD0BWP12T U1207 ( .I0(n3609), .I1(n3608), .S(n5247), .ZN(n3610) );
  ND2D1BWP12T U1208 ( .A1(n3611), .A2(n3610), .ZN(n3645) );
  MUX2ND0BWP12T U1209 ( .I0(n4646), .I1(n4647), .S(n4092), .ZN(n3612) );
  OAI21D0BWP12T U1210 ( .A1(b[15]), .A2(n5361), .B(n3612), .ZN(n3675) );
  INVD1BWP12T U1211 ( .I(n3613), .ZN(n4394) );
  NR2D1BWP12T U1212 ( .A1(n4394), .A2(n3934), .ZN(n3674) );
  INVD1BWP12T U1213 ( .I(n5876), .ZN(n4370) );
  INVD1BWP12T U1214 ( .I(n5875), .ZN(n4369) );
  MUX2ND0BWP12T U1215 ( .I0(n4370), .I1(n4369), .S(n5806), .ZN(n3615) );
  MUX2ND0BWP12T U1216 ( .I0(n4372), .I1(n4371), .S(b[9]), .ZN(n3614) );
  CKND2D1BWP12T U1217 ( .A1(n3615), .A2(n3614), .ZN(n3673) );
  FA1D0BWP12T U1218 ( .A(n3617), .B(n3624), .CI(n3616), .CO(n3648), .S(n3618)
         );
  FA1D0BWP12T U1219 ( .A(n3621), .B(n3620), .CI(n3619), .CO(n4015), .S(n3622)
         );
  INVD1BWP12T U1220 ( .I(n3622), .ZN(n4018) );
  INVD1BWP12T U1221 ( .I(n3623), .ZN(n4009) );
  OAI21D1BWP12T U1222 ( .A1(n3626), .A2(n3625), .B(n3624), .ZN(n3672) );
  INVD1BWP12T U1223 ( .I(n3672), .ZN(n3634) );
  XNR3D1BWP12T U1224 ( .A1(n3629), .A2(n3628), .A3(n3627), .ZN(n3670) );
  MUX2NXD0BWP12T U1225 ( .I0(n5870), .I1(n5869), .S(n5247), .ZN(n3631) );
  MUX2ND0BWP12T U1226 ( .I0(n5871), .I1(n5872), .S(n3463), .ZN(n3630) );
  NR2D1BWP12T U1227 ( .A1(n3631), .A2(n3630), .ZN(n3677) );
  MUX2NXD0BWP12T U1228 ( .I0(n5817), .I1(n5816), .S(n6573), .ZN(n3633) );
  MUX2ND0BWP12T U1229 ( .I0(n5819), .I1(n5818), .S(n6334), .ZN(n3632) );
  NR2D1BWP12T U1230 ( .A1(n3633), .A2(n3632), .ZN(n3679) );
  MAOI222D1BWP12T U1231 ( .A(n3678), .B(n3677), .C(n3679), .ZN(n3671) );
  MAOI222D1BWP12T U1232 ( .A(n3634), .B(n3670), .C(n3671), .ZN(n3690) );
  XNR3D1BWP12T U1233 ( .A1(n3637), .A2(n3636), .A3(n3635), .ZN(n3689) );
  MUX2ND0BWP12T U1234 ( .I0(n3911), .I1(n5810), .S(b[14]), .ZN(n3639) );
  MUX2ND0BWP12T U1235 ( .I0(n5813), .I1(n5812), .S(b[13]), .ZN(n3638) );
  NR2D1BWP12T U1236 ( .A1(n3639), .A2(n3638), .ZN(n3660) );
  MUX2ND0BWP12T U1237 ( .I0(n5776), .I1(n5775), .S(n5864), .ZN(n3641) );
  MUX2ND0BWP12T U1238 ( .I0(n5778), .I1(n5777), .S(n6782), .ZN(n3640) );
  NR2D1BWP12T U1239 ( .A1(n3641), .A2(n3640), .ZN(n3659) );
  MUX2ND0BWP12T U1240 ( .I0(n5837), .I1(n5836), .S(n5843), .ZN(n3643) );
  MUX2NXD0BWP12T U1241 ( .I0(n5839), .I1(n5838), .S(n5379), .ZN(n3642) );
  NR2D1BWP12T U1242 ( .A1(n3643), .A2(n3642), .ZN(n3658) );
  FA1D0BWP12T U1243 ( .A(n3646), .B(n3645), .CI(n3644), .CO(n3686), .S(n3647)
         );
  INVD1BWP12T U1244 ( .I(n3647), .ZN(n3719) );
  FA1D0BWP12T U1245 ( .A(n3650), .B(n3649), .CI(n3648), .CO(n3619), .S(n3656)
         );
  INVD1BWP12T U1246 ( .I(n3654), .ZN(n3655) );
  NR2D2BWP12T U1247 ( .A1(n4009), .A2(n4008), .ZN(n5500) );
  FA1D0BWP12T U1248 ( .A(n3657), .B(n3656), .CI(n3655), .CO(n4008), .S(n4007)
         );
  FA1D0BWP12T U1249 ( .A(n3660), .B(n3659), .CI(n3658), .CO(n3720), .S(n3694)
         );
  MUX2D1BWP12T U1250 ( .I0(n5817), .I1(n5816), .S(n6334), .Z(n3662) );
  MUX2D1BWP12T U1251 ( .I0(n5819), .I1(n5818), .S(n6520), .Z(n3661) );
  ND2D1BWP12T U1252 ( .A1(n3662), .A2(n3661), .ZN(n3701) );
  CKND2D1BWP12T U1253 ( .A1(n5871), .A2(n5872), .ZN(n4738) );
  IND2D1BWP12T U1254 ( .A1(n4829), .B1(n6232), .ZN(n4920) );
  CKND0BWP12T U1255 ( .I(n6238), .ZN(n3663) );
  OAI21D1BWP12T U1256 ( .A1(n3663), .A2(n4920), .B(n5872), .ZN(n3703) );
  MAOI222D1BWP12T U1257 ( .A(n3701), .B(n3702), .C(n3703), .ZN(n3695) );
  NR2D1BWP12T U1258 ( .A1(n3694), .A2(n3695), .ZN(n3669) );
  MUX2ND0BWP12T U1259 ( .I0(n5776), .I1(n5775), .S(n6782), .ZN(n3665) );
  MUX2ND0BWP12T U1260 ( .I0(n5778), .I1(n5777), .S(n6573), .ZN(n3664) );
  NR2D1BWP12T U1261 ( .A1(n3665), .A2(n3664), .ZN(n3715) );
  NR2D1BWP12T U1262 ( .A1(n3715), .A2(n3716), .ZN(n3714) );
  INVD1BWP12T U1263 ( .I(n3694), .ZN(n3668) );
  INVD1BWP12T U1264 ( .I(n3695), .ZN(n3667) );
  OAI22D1BWP12T U1265 ( .A1(n3669), .A2(n3714), .B1(n3668), .B2(n3667), .ZN(
        n3724) );
  XOR3D1BWP12T U1266 ( .A1(n3672), .A2(n3671), .A3(n3670), .Z(n3723) );
  FA1D0BWP12T U1267 ( .A(n3675), .B(n3674), .CI(n3673), .CO(n3644), .S(n3676)
         );
  INVD1BWP12T U1268 ( .I(n3676), .ZN(n3747) );
  XOR3D1BWP12T U1269 ( .A1(n3679), .A2(n3678), .A3(n3677), .Z(n3746) );
  MUX2ND0BWP12T U1270 ( .I0(n5859), .I1(n5858), .S(b[11]), .ZN(n3681) );
  MUX2ND0BWP12T U1271 ( .I0(n5860), .I1(n5861), .S(n5405), .ZN(n3680) );
  NR2D1BWP12T U1272 ( .A1(n3681), .A2(n3680), .ZN(n3706) );
  MUX2ND0BWP12T U1273 ( .I0(n3911), .I1(n5810), .S(b[13]), .ZN(n3683) );
  NR2D1BWP12T U1274 ( .A1(n3683), .A2(n3682), .ZN(n3705) );
  MUX2D1BWP12T U1275 ( .I0(n4371), .I1(n4372), .S(n4515), .Z(n3684) );
  NR2D1BWP12T U1276 ( .A1(n3685), .A2(n3684), .ZN(n3704) );
  INVD1BWP12T U1277 ( .I(n3687), .ZN(n3692) );
  FA1D0BWP12T U1278 ( .A(n3690), .B(n3689), .CI(n3688), .CO(n3657), .S(n3691)
         );
  NR2D1BWP12T U1279 ( .A1(n4007), .A2(n4006), .ZN(n5498) );
  TPNR2D1BWP12T U1280 ( .A1(n5500), .A2(n5498), .ZN(n4011) );
  FA1D0BWP12T U1281 ( .A(n3693), .B(n3692), .CI(n3691), .CO(n4006), .S(n4005)
         );
  XNR3D1BWP12T U1282 ( .A1(n3714), .A2(n3695), .A3(n3694), .ZN(n3750) );
  MUX2ND0BWP12T U1283 ( .I0(n6240), .I1(n4755), .S(b[14]), .ZN(n3696) );
  AOI21D1BWP12T U1284 ( .A1(n4557), .A2(n4576), .B(n3696), .ZN(n3736) );
  ND2D1BWP12T U1285 ( .A1(n4623), .A2(n4823), .ZN(n3735) );
  MUX2NXD1BWP12T U1286 ( .I0(n3911), .I1(n5810), .S(b[12]), .ZN(n3698) );
  MUX2ND0BWP12T U1287 ( .I0(n5813), .I1(n5812), .S(b[11]), .ZN(n3697) );
  NR2D1BWP12T U1288 ( .A1(n3698), .A2(n3697), .ZN(n3734) );
  MUX2ND0BWP12T U1289 ( .I0(n5837), .I1(n5836), .S(n5379), .ZN(n3700) );
  MUX2NXD0BWP12T U1290 ( .I0(n5839), .I1(n5838), .S(b[6]), .ZN(n3699) );
  NR2D1BWP12T U1291 ( .A1(n3700), .A2(n3699), .ZN(n3732) );
  XNR3XD1BWP12T U1292 ( .A1(n3703), .A2(n3702), .A3(n3701), .ZN(n3731) );
  FA1D0BWP12T U1293 ( .A(n3706), .B(n3705), .CI(n3704), .CO(n3745), .S(n3728)
         );
  MUX2NXD0BWP12T U1294 ( .I0(n5817), .I1(n5816), .S(n5247), .ZN(n3708) );
  MUX2NXD0BWP12T U1295 ( .I0(n5819), .I1(n5818), .S(n5612), .ZN(n3707) );
  NR2D1BWP12T U1296 ( .A1(n3708), .A2(n3707), .ZN(n3758) );
  MUX2NXD0BWP12T U1297 ( .I0(n5837), .I1(n5836), .S(n5864), .ZN(n3710) );
  MUX2ND0BWP12T U1298 ( .I0(n5839), .I1(n5838), .S(n6782), .ZN(n3709) );
  NR2D1BWP12T U1299 ( .A1(n3710), .A2(n3709), .ZN(n3756) );
  MUX2ND0BWP12T U1300 ( .I0(n5776), .I1(n5775), .S(n6573), .ZN(n3712) );
  MUX2ND0BWP12T U1301 ( .I0(n5778), .I1(n5777), .S(n6334), .ZN(n3711) );
  NR2D1BWP12T U1302 ( .A1(n3712), .A2(n3711), .ZN(n3757) );
  NR2D1BWP12T U1303 ( .A1(n3728), .A2(n3713), .ZN(n3718) );
  AOI21D1BWP12T U1304 ( .A1(n3716), .A2(n3715), .B(n3714), .ZN(n3729) );
  INVD1BWP12T U1305 ( .I(n3728), .ZN(n3717) );
  OAI22D1BWP12T U1306 ( .A1(n3718), .A2(n3729), .B1(n3717), .B2(n3730), .ZN(
        n3748) );
  FA1D0BWP12T U1307 ( .A(n3721), .B(n3720), .CI(n3719), .CO(n3688), .S(n3726)
         );
  FA1D0BWP12T U1308 ( .A(n3724), .B(n3723), .CI(n3722), .CO(n3693), .S(n3725)
         );
  NR2D1BWP12T U1309 ( .A1(n4005), .A2(n4004), .ZN(n6056) );
  FA1D0BWP12T U1310 ( .A(n3727), .B(n3726), .CI(n3725), .CO(n4004), .S(n4003)
         );
  FA1D0BWP12T U1311 ( .A(n3733), .B(n3732), .CI(n3731), .CO(n3749), .S(n3985)
         );
  FA1D0BWP12T U1312 ( .A(n3736), .B(n3735), .CI(n3734), .CO(n3733), .S(n3761)
         );
  MUX2ND0BWP12T U1313 ( .I0(n5776), .I1(n5775), .S(n6334), .ZN(n3738) );
  MUX2ND0BWP12T U1314 ( .I0(n5778), .I1(n5777), .S(n5247), .ZN(n3737) );
  NR2D1BWP12T U1315 ( .A1(n3738), .A2(n3737), .ZN(n3774) );
  OR2XD1BWP12T U1316 ( .A1(n3774), .A2(n3773), .Z(n3760) );
  MUX2ND0BWP12T U1317 ( .I0(n3911), .I1(n5810), .S(b[11]), .ZN(n3740) );
  MUX2ND0BWP12T U1318 ( .I0(n5813), .I1(n5812), .S(n5806), .ZN(n3739) );
  NR2D1BWP12T U1319 ( .A1(n3740), .A2(n3739), .ZN(n3777) );
  AOI21D1BWP12T U1320 ( .A1(n3742), .A2(n4305), .B(n3741), .ZN(n3776) );
  MUX2ND0BWP12T U1321 ( .I0(n5859), .I1(n5858), .S(b[9]), .ZN(n3744) );
  MUX2ND0BWP12T U1322 ( .I0(n5860), .I1(n5861), .S(n4515), .ZN(n3743) );
  NR2D1BWP12T U1323 ( .A1(n3744), .A2(n3743), .ZN(n3775) );
  FA1D0BWP12T U1324 ( .A(n3747), .B(n3746), .CI(n3745), .CO(n3722), .S(n3991)
         );
  FA1D0BWP12T U1325 ( .A(n3750), .B(n3749), .CI(n3748), .CO(n3727), .S(n3990)
         );
  NR2D1BWP12T U1326 ( .A1(n4003), .A2(n4002), .ZN(n6054) );
  NR2D1BWP12T U1327 ( .A1(n6056), .A2(n6054), .ZN(n5494) );
  CKND2D1BWP12T U1328 ( .A1(n4011), .A2(n5494), .ZN(n4013) );
  INVD1BWP12T U1329 ( .I(b[9]), .ZN(n4730) );
  MUX2NXD0BWP12T U1330 ( .I0(a[13]), .I1(n6231), .S(n4829), .ZN(n5179) );
  INVD1BWP12T U1331 ( .I(n5179), .ZN(n5166) );
  ND2D1BWP12T U1332 ( .A1(n5818), .A2(n5819), .ZN(n4375) );
  MUX2NXD0BWP12T U1333 ( .I0(n5817), .I1(n5816), .S(n5612), .ZN(n3751) );
  AOI21D1BWP12T U1334 ( .A1(n5166), .A2(n4375), .B(n3751), .ZN(n3772) );
  ND2D1BWP12T U1335 ( .A1(n5236), .A2(n4343), .ZN(n6815) );
  ND2D1BWP12T U1336 ( .A1(n6819), .A2(n5379), .ZN(n6811) );
  ND2D1BWP12T U1337 ( .A1(n6815), .A2(n6811), .ZN(n6133) );
  INVD1BWP12T U1338 ( .I(n6133), .ZN(n6189) );
  MUX2ND0BWP12T U1339 ( .I0(n5877), .I1(n5878), .S(n4357), .ZN(n3752) );
  AOI21D1BWP12T U1340 ( .A1(n3914), .A2(n6189), .B(n3752), .ZN(n3771) );
  MUX2ND0BWP12T U1341 ( .I0(n5837), .I1(n5836), .S(n6782), .ZN(n3754) );
  MUX2NXD0BWP12T U1342 ( .I0(n5839), .I1(n5838), .S(n6573), .ZN(n3753) );
  NR2D1BWP12T U1343 ( .A1(n3754), .A2(n3753), .ZN(n3770) );
  ND2D1BWP12T U1344 ( .A1(n5877), .A2(n5878), .ZN(n3935) );
  AOI21D1BWP12T U1345 ( .A1(n6189), .A2(n3935), .B(n3755), .ZN(n3982) );
  XOR3D1BWP12T U1346 ( .A1(n3758), .A2(n3757), .A3(n3756), .Z(n3981) );
  FA1D0BWP12T U1347 ( .A(n3761), .B(n3760), .CI(n3759), .CO(n3984), .S(n3980)
         );
  CKND2D1BWP12T U1348 ( .A1(n4390), .A2(n4823), .ZN(n3783) );
  INVD1BWP12T U1349 ( .I(n3783), .ZN(n3765) );
  MUX2ND0BWP12T U1350 ( .I0(n3911), .I1(n5810), .S(n5806), .ZN(n3763) );
  MUX2ND0BWP12T U1351 ( .I0(n5813), .I1(n5812), .S(b[9]), .ZN(n3762) );
  NR2D1BWP12T U1352 ( .A1(n3763), .A2(n3762), .ZN(n3781) );
  INVD1BWP12T U1353 ( .I(n3781), .ZN(n3764) );
  MAOI222D1BWP12T U1354 ( .A(n3765), .B(n3764), .C(n3782), .ZN(n3794) );
  MUX2ND0BWP12T U1355 ( .I0(n5876), .I1(n5875), .S(n5864), .ZN(n3767) );
  MUX2ND0BWP12T U1356 ( .I0(n5877), .I1(n5878), .S(n4433), .ZN(n3766) );
  NR2D1BWP12T U1357 ( .A1(n3767), .A2(n3766), .ZN(n3799) );
  MUX2ND0BWP12T U1358 ( .I0(n4757), .I1(n4756), .S(n6573), .ZN(n3769) );
  MUX2ND0BWP12T U1359 ( .I0(n4759), .I1(n4760), .S(n6334), .ZN(n3768) );
  AN2XD1BWP12T U1360 ( .A1(n3769), .A2(n3768), .Z(n3798) );
  FA1D1BWP12T U1361 ( .A(n3772), .B(n3771), .CI(n3770), .CO(n3983), .S(n3792)
         );
  FA1D0BWP12T U1362 ( .A(n3777), .B(n3776), .CI(n3775), .CO(n3759), .S(n3778)
         );
  MUX2ND0BWP12T U1363 ( .I0(n3405), .I1(n5395), .S(n5843), .ZN(n3780) );
  MUX2ND0BWP12T U1364 ( .I0(n5397), .I1(n5396), .S(n5379), .ZN(n3779) );
  ND2D1BWP12T U1365 ( .A1(n3780), .A2(n3779), .ZN(n3812) );
  XOR3D2BWP12T U1366 ( .A1(n3783), .A2(n3782), .A3(n3781), .Z(n3811) );
  MUX2NXD0BWP12T U1367 ( .I0(n4759), .I1(n4760), .S(n5247), .ZN(n3784) );
  CKND2D1BWP12T U1368 ( .A1(n3785), .A2(n3784), .ZN(n3836) );
  MUX2ND0BWP12T U1369 ( .I0(n3405), .I1(n5395), .S(n5379), .ZN(n3787) );
  MUX2ND0BWP12T U1370 ( .I0(n5397), .I1(n5396), .S(n5864), .ZN(n3786) );
  ND2D1BWP12T U1371 ( .A1(n3787), .A2(n3786), .ZN(n3835) );
  MUX2ND0BWP12T U1372 ( .I0(n4646), .I1(n4647), .S(n5405), .ZN(n3788) );
  IOA21D1BWP12T U1373 ( .A1(n4557), .A2(n4730), .B(n3788), .ZN(n3842) );
  INVD1BWP12T U1374 ( .I(n3789), .ZN(n3790) );
  NR2D1BWP12T U1375 ( .A1(n3790), .A2(n3934), .ZN(n3841) );
  INVD1BWP12T U1376 ( .I(n3791), .ZN(n3987) );
  FA1D0BWP12T U1377 ( .A(n3794), .B(n3793), .CI(n3792), .CO(n3988), .S(n3809)
         );
  INVD1BWP12T U1378 ( .I(n3796), .ZN(n3808) );
  INVD1BWP12T U1379 ( .I(n5778), .ZN(n3822) );
  NR2XD0BWP12T U1380 ( .A1(n5776), .A2(n4823), .ZN(n3821) );
  MUX2ND0BWP12T U1381 ( .I0(n4646), .I1(n4647), .S(n4745), .ZN(n3797) );
  OAI21D1BWP12T U1382 ( .A1(n5806), .A2(n5361), .B(n3797), .ZN(n3820) );
  OAI21D1BWP12T U1383 ( .A1(n3822), .A2(n3821), .B(n3820), .ZN(n3819) );
  FA1D1BWP12T U1384 ( .A(n3800), .B(n3799), .CI(n3798), .CO(n3793), .S(n3815)
         );
  MUX2ND0BWP12T U1385 ( .I0(n5778), .I1(n5777), .S(n4823), .ZN(n3801) );
  NR2D1BWP12T U1386 ( .A1(n3802), .A2(n3801), .ZN(n3818) );
  MUX2ND0BWP12T U1387 ( .I0(n5876), .I1(n5875), .S(n6782), .ZN(n3804) );
  BUFFD3BWP12T U1388 ( .I(n6357), .Z(n6565) );
  MUX2ND0BWP12T U1389 ( .I0(n5877), .I1(n5878), .S(n6565), .ZN(n3803) );
  NR2D1BWP12T U1390 ( .A1(n3804), .A2(n3803), .ZN(n3817) );
  MUX2ND0BWP12T U1391 ( .I0(n3911), .I1(n5810), .S(b[9]), .ZN(n3806) );
  MUX2ND0BWP12T U1392 ( .I0(n5813), .I1(n5812), .S(n5843), .ZN(n3805) );
  NR2D1BWP12T U1393 ( .A1(n3806), .A2(n3805), .ZN(n3816) );
  NR2D1BWP12T U1394 ( .A1(n3976), .A2(n3975), .ZN(n5598) );
  FA1D0BWP12T U1395 ( .A(n3812), .B(n3811), .CI(n3810), .CO(n3795), .S(n3813)
         );
  INVD1BWP12T U1396 ( .I(n3813), .ZN(n3830) );
  OAI31D1BWP12T U1397 ( .A1(n3822), .A2(n3821), .A3(n3820), .B(n3819), .ZN(
        n3832) );
  NR2D1BWP12T U1398 ( .A1(n6267), .A2(n6782), .ZN(n5113) );
  INVD1BWP12T U1399 ( .I(n5113), .ZN(n6784) );
  ND2D1BWP12T U1400 ( .A1(n6267), .A2(n6782), .ZN(n6096) );
  ND2D1BWP12T U1401 ( .A1(n6784), .A2(n6096), .ZN(n6134) );
  CKND1BWP12T U1402 ( .I(n6134), .ZN(n6178) );
  ND2D1BWP12T U1403 ( .A1(n5860), .A2(n5861), .ZN(n3903) );
  MUX2ND0BWP12T U1404 ( .I0(n5859), .I1(n5858), .S(n5864), .ZN(n3823) );
  AOI21D1BWP12T U1405 ( .A1(n6178), .A2(n3903), .B(n3823), .ZN(n3853) );
  MUX2ND0BWP12T U1406 ( .I0(n5876), .I1(n5875), .S(n6573), .ZN(n3825) );
  MUX2ND0BWP12T U1407 ( .I0(n5877), .I1(n5878), .S(n6576), .ZN(n3824) );
  NR2D1BWP12T U1408 ( .A1(n3825), .A2(n3824), .ZN(n3852) );
  MUX2ND0BWP12T U1409 ( .I0(n3911), .I1(n5810), .S(n5843), .ZN(n3827) );
  MUX2ND0BWP12T U1410 ( .I0(n5813), .I1(n5812), .S(n5379), .ZN(n3826) );
  NR2D1BWP12T U1411 ( .A1(n3827), .A2(n3826), .ZN(n3851) );
  TPNR2D1BWP12T U1412 ( .A1(n3972), .A2(n3971), .ZN(n5144) );
  FA1D0BWP12T U1413 ( .A(n3836), .B(n3835), .CI(n3834), .CO(n3810), .S(n3837)
         );
  INVD1BWP12T U1414 ( .I(n3837), .ZN(n3849) );
  INVD1BWP12T U1415 ( .I(n3882), .ZN(n3838) );
  INVD1BWP12T U1416 ( .I(n6249), .ZN(n5253) );
  ND2D1BWP12T U1417 ( .A1(n5253), .A2(n6565), .ZN(n5259) );
  ND2D1BWP12T U1418 ( .A1(n6249), .A2(n6573), .ZN(n6097) );
  ND2D1BWP12T U1419 ( .A1(n5259), .A2(n6097), .ZN(n5274) );
  MOAI22D0BWP12T U1420 ( .A1(n3838), .A2(n6134), .B1(n3903), .B2(n5274), .ZN(
        n3854) );
  MUX2ND0BWP12T U1421 ( .I0(n4646), .I1(n4647), .S(n4730), .ZN(n3839) );
  OAI21D1BWP12T U1422 ( .A1(n5843), .A2(n5361), .B(n3839), .ZN(n3855) );
  FA1D0BWP12T U1423 ( .A(n3842), .B(n3841), .CI(n3840), .CO(n3834), .S(n3843)
         );
  INVD1BWP12T U1424 ( .I(n3843), .ZN(n3863) );
  MUX2XD0BWP12T U1425 ( .I0(n6229), .I1(a[8]), .S(n6248), .Z(n5165) );
  MUX2ND0BWP12T U1426 ( .I0(n5837), .I1(n5836), .S(n5612), .ZN(n3844) );
  AOI21D1BWP12T U1427 ( .A1(n5165), .A2(n3845), .B(n3844), .ZN(n3870) );
  AOI21D1BWP12T U1428 ( .A1(n4757), .A2(n3934), .B(n4759), .ZN(n3869) );
  MUX2ND0BWP12T U1429 ( .I0(n3911), .I1(n5810), .S(n5379), .ZN(n3847) );
  MUX2ND0BWP12T U1430 ( .I0(n5813), .I1(n5812), .S(b[6]), .ZN(n3846) );
  NR2D1BWP12T U1431 ( .A1(n3847), .A2(n3846), .ZN(n3868) );
  FA1D2BWP12T U1432 ( .A(n3850), .B(n3849), .CI(n3848), .CO(n3968), .S(n3967)
         );
  FA1D0BWP12T U1433 ( .A(n3853), .B(n3852), .CI(n3851), .CO(n3831), .S(n3867)
         );
  OAI21D1BWP12T U1434 ( .A1(n3855), .A2(n3854), .B(n3864), .ZN(n3879) );
  MUX2ND0BWP12T U1435 ( .I0(n5877), .I1(n5878), .S(n5767), .ZN(n3856) );
  NR2D1BWP12T U1436 ( .A1(n3857), .A2(n3856), .ZN(n3878) );
  AOI21D1BWP12T U1437 ( .A1(n4557), .A2(n4343), .B(n3858), .ZN(n3944) );
  ND2D1BWP12T U1438 ( .A1(n3859), .A2(n4823), .ZN(n3943) );
  MUX2ND0BWP12T U1439 ( .I0(n3911), .I1(n5810), .S(n5864), .ZN(n3861) );
  MUX2ND0BWP12T U1440 ( .I0(n5813), .I1(n5812), .S(n6782), .ZN(n3860) );
  NR2D1BWP12T U1441 ( .A1(n3861), .A2(n3860), .ZN(n3942) );
  FA1D0BWP12T U1442 ( .A(n3864), .B(n3863), .CI(n3862), .CO(n3848), .S(n3865)
         );
  FA1D0BWP12T U1443 ( .A(n3867), .B(n3866), .CI(n3865), .CO(n3966), .S(n3965)
         );
  FA1D0BWP12T U1444 ( .A(n3870), .B(n3869), .CI(n3868), .CO(n3862), .S(n3957)
         );
  MUX2ND0BWP12T U1445 ( .I0(n4370), .I1(n4369), .S(n5247), .ZN(n3872) );
  MUX2NXD0BWP12T U1446 ( .I0(n4372), .I1(n4371), .S(n5612), .ZN(n3871) );
  ND2D1BWP12T U1447 ( .A1(n3872), .A2(n3871), .ZN(n3947) );
  MUX2ND0BWP12T U1448 ( .I0(n5859), .I1(n5858), .S(n6334), .ZN(n3874) );
  MUX2D1BWP12T U1449 ( .I0(n5396), .I1(n5397), .S(n5767), .Z(n3873) );
  NR2D1BWP12T U1450 ( .A1(n3874), .A2(n3873), .ZN(n3925) );
  NR2D1BWP12T U1451 ( .A1(n3925), .A2(n3924), .ZN(n3946) );
  MUX2ND0BWP12T U1452 ( .I0(n3405), .I1(n5395), .S(n6573), .ZN(n3876) );
  MUX2ND0BWP12T U1453 ( .I0(n5397), .I1(n5396), .S(n6334), .ZN(n3875) );
  ND2D1BWP12T U1454 ( .A1(n3876), .A2(n3875), .ZN(n3945) );
  MAOI222D1BWP12T U1455 ( .A(n3947), .B(n3946), .C(n3945), .ZN(n3956) );
  FA1D0BWP12T U1456 ( .A(n3879), .B(n3878), .CI(n3877), .CO(n3866), .S(n3955)
         );
  MAOI222D1BWP12T U1457 ( .A(n3957), .B(n3956), .C(n3955), .ZN(n3880) );
  INVD1BWP12T U1458 ( .I(n3880), .ZN(n3964) );
  NR2D1BWP12T U1459 ( .A1(n3965), .A2(n3964), .ZN(n6012) );
  NR2D1BWP12T U1460 ( .A1(n6014), .A2(n6012), .ZN(n5555) );
  ND2D1BWP12T U1461 ( .A1(n5560), .A2(n5555), .ZN(n5143) );
  TPNR2D0BWP12T U1462 ( .A1(n5144), .A2(n5143), .ZN(n3974) );
  AOI21D1BWP12T U1463 ( .A1(n4557), .A2(n4924), .B(n3881), .ZN(n3908) );
  ND2D1BWP12T U1464 ( .A1(n3882), .A2(n4823), .ZN(n3907) );
  ND2D1BWP12T U1465 ( .A1(n5360), .A2(n4498), .ZN(n6098) );
  NR2D1BWP12T U1466 ( .A1(n5360), .A2(n4498), .ZN(n4309) );
  INR2D2BWP12T U1467 ( .A1(n6098), .B1(n4309), .ZN(n4303) );
  INVD2BWP12T U1468 ( .I(n4303), .ZN(n4304) );
  MUX2ND0BWP12T U1469 ( .I0(n3911), .I1(n5810), .S(n6520), .ZN(n3883) );
  AOI21D1BWP12T U1470 ( .A1(n4304), .A2(n3913), .B(n3883), .ZN(n3906) );
  MUX2XD0BWP12T U1471 ( .I0(n6247), .I1(a[2]), .S(n6248), .Z(n4894) );
  CKND2D1BWP12T U1472 ( .A1(n3913), .A2(n4894), .ZN(n3884) );
  ND2D1BWP12T U1473 ( .A1(n3885), .A2(n3884), .ZN(n3888) );
  MUX2XD0BWP12T U1474 ( .I0(n6240), .I1(n4755), .S(n6334), .Z(n3887) );
  CKND2D1BWP12T U1475 ( .A1(n4557), .A2(n5767), .ZN(n3886) );
  ND2D1BWP12T U1476 ( .A1(n3887), .A2(n3886), .ZN(n3889) );
  ND2D1BWP12T U1477 ( .A1(n3888), .A2(n3889), .ZN(n5222) );
  INVD1BWP12T U1478 ( .I(n3888), .ZN(n3891) );
  CKND0BWP12T U1479 ( .I(n3889), .ZN(n3890) );
  ND2D1BWP12T U1480 ( .A1(n3891), .A2(n3890), .ZN(n3892) );
  INVD1BWP12T U1481 ( .I(n5360), .ZN(n4307) );
  NR2D1BWP12T U1482 ( .A1(n4307), .A2(n4823), .ZN(n4144) );
  MUX2D1BWP12T U1483 ( .I0(n6240), .I1(n4755), .S(n6520), .Z(n3894) );
  ND2D1BWP12T U1484 ( .A1(n4557), .A2(n3463), .ZN(n3893) );
  ND2D1BWP12T U1485 ( .A1(n3894), .A2(n3893), .ZN(n3895) );
  INR2D1BWP12T U1486 ( .A1(n3896), .B1(n3895), .ZN(n6033) );
  ND2D1BWP12T U1487 ( .A1(n3902), .A2(n4823), .ZN(n6034) );
  INVD1BWP12T U1488 ( .I(n3895), .ZN(n3897) );
  OAI22D1BWP12T U1489 ( .A1(n6033), .A2(n6034), .B1(n3897), .B2(n3896), .ZN(
        n6035) );
  OAI21D1BWP12T U1490 ( .A1(n3911), .A2(n4829), .B(n5813), .ZN(n4915) );
  NR2D1BWP12T U1491 ( .A1(n6035), .A2(n4915), .ZN(n3899) );
  CKND2D1BWP12T U1492 ( .A1(n6035), .A2(n4915), .ZN(n3898) );
  INVD1BWP12T U1493 ( .I(n5224), .ZN(n3900) );
  OAI21D1BWP12T U1494 ( .A1(n5223), .A2(n5222), .B(n3900), .ZN(n3901) );
  IOA21D1BWP12T U1495 ( .A1(n5223), .A2(n5222), .B(n3901), .ZN(n3910) );
  IND2XD2BWP12T U1496 ( .A1(n6334), .B1(n6247), .ZN(n4938) );
  NR2D1BWP12T U1497 ( .A1(n6576), .A2(n6247), .ZN(n6462) );
  INR2D2BWP12T U1498 ( .A1(n4938), .B1(n6462), .ZN(n5226) );
  INVD1BWP12T U1499 ( .I(n3405), .ZN(n4747) );
  INVD1BWP12T U1500 ( .I(n5395), .ZN(n4746) );
  MUX2XD0BWP12T U1501 ( .I0(n6267), .I1(n6249), .S(n6248), .Z(n4888) );
  AOI21D1BWP12T U1502 ( .A1(n3405), .A2(n3934), .B(n5397), .ZN(n3905) );
  NR2D1BWP12T U1503 ( .A1(n3905), .A2(n3904), .ZN(n3937) );
  AOI21D1BWP12T U1504 ( .A1(n3905), .A2(n3904), .B(n3937), .ZN(n3920) );
  XOR3D1BWP12T U1505 ( .A1(n3918), .A2(n3919), .A3(n3920), .Z(n3909) );
  FICOND1BWP12T U1506 ( .A(n3908), .B(n3907), .CI(n3906), .CON(n6031), .S(
        n5223) );
  ND2D1BWP12T U1507 ( .A1(n3910), .A2(n3909), .ZN(n6029) );
  OAI21D1BWP12T U1508 ( .A1(n6028), .A2(n6031), .B(n6029), .ZN(n5105) );
  INVD1BWP12T U1509 ( .I(n5226), .ZN(n4952) );
  MUX2D1BWP12T U1510 ( .I0(n3911), .I1(n5810), .S(n6573), .Z(n3912) );
  IOA21D1BWP12T U1511 ( .A1(n4952), .A2(n3913), .B(n3912), .ZN(n3938) );
  ND2D1BWP12T U1512 ( .A1(n3914), .A2(n4823), .ZN(n3926) );
  INVD1BWP12T U1513 ( .I(n3926), .ZN(n3929) );
  INVD1BWP12T U1514 ( .I(n3927), .ZN(n3928) );
  MUX2D1BWP12T U1515 ( .I0(n4747), .I1(n4746), .S(n5247), .Z(n3916) );
  ND2D1BWP12T U1516 ( .A1(n3916), .A2(n3915), .ZN(n3931) );
  XOR3D1BWP12T U1517 ( .A1(n3929), .A2(n3928), .A3(n3931), .Z(n3936) );
  INVD1BWP12T U1518 ( .I(n3917), .ZN(n3922) );
  ND2D1BWP12T U1519 ( .A1(n3922), .A2(n3921), .ZN(n5103) );
  INVD1BWP12T U1520 ( .I(n5103), .ZN(n3923) );
  AO21D1BWP12T U1521 ( .A1(n3925), .A2(n3924), .B(n3946), .Z(n3951) );
  TPNR2D0BWP12T U1522 ( .A1(n3927), .A2(n3926), .ZN(n3930) );
  OAI22D1BWP12T U1523 ( .A1(n3931), .A2(n3930), .B1(n3929), .B2(n3928), .ZN(
        n3950) );
  MUX2ND0BWP12T U1524 ( .I0(n3911), .I1(n5810), .S(n6782), .ZN(n3933) );
  MUX2ND0BWP12T U1525 ( .I0(n5813), .I1(n5812), .S(n6573), .ZN(n3932) );
  MUX2D1BWP12T U1526 ( .I0(n6819), .I1(a[6]), .S(n6248), .Z(n6263) );
  XNR3D1BWP12T U1527 ( .A1(n3951), .A2(n3950), .A3(n3949), .ZN(n3939) );
  FA1D0BWP12T U1528 ( .A(n3938), .B(n3937), .CI(n3936), .CO(n6022), .S(n3917)
         );
  CKND0BWP12T U1529 ( .I(n6022), .ZN(n3941) );
  ND2D1BWP12T U1530 ( .A1(n3940), .A2(n3939), .ZN(n6020) );
  OAI21D1BWP12T U1531 ( .A1(n6019), .A2(n3941), .B(n6020), .ZN(n6026) );
  FA1D0BWP12T U1532 ( .A(n3944), .B(n3943), .CI(n3942), .CO(n3877), .S(n3960)
         );
  XNR3D1BWP12T U1533 ( .A1(n3947), .A2(n3946), .A3(n3945), .ZN(n3958) );
  INVD1BWP12T U1534 ( .I(n3948), .ZN(n3953) );
  MAOI222D1BWP12T U1535 ( .A(n3951), .B(n3950), .C(n3949), .ZN(n3952) );
  OR2D2BWP12T U1536 ( .A1(n3953), .A2(n3952), .Z(n6025) );
  ND2D1BWP12T U1537 ( .A1(n3953), .A2(n3952), .ZN(n6024) );
  INVD1BWP12T U1538 ( .I(n6024), .ZN(n3954) );
  TPAOI21D1BWP12T U1539 ( .A1(n6026), .A2(n6025), .B(n3954), .ZN(n3962) );
  XOR3D1BWP12T U1540 ( .A1(n3957), .A2(n3956), .A3(n3955), .Z(n3961) );
  TPNR2D1BWP12T U1541 ( .A1(n3962), .A2(n3961), .ZN(n5192) );
  FA1D0BWP12T U1542 ( .A(n3960), .B(n3959), .CI(n3958), .CO(n5194), .S(n3948)
         );
  CKND1BWP12T U1543 ( .I(n5194), .ZN(n3963) );
  CKND2D2BWP12T U1544 ( .A1(n3962), .A2(n3961), .ZN(n5193) );
  TPOAI21D1BWP12T U1545 ( .A1(n5192), .A2(n3963), .B(n5193), .ZN(n4226) );
  ND2D1BWP12T U1546 ( .A1(n3965), .A2(n3964), .ZN(n6011) );
  TPOAI21D1BWP12T U1547 ( .A1(n6014), .A2(n6011), .B(n6015), .ZN(n5556) );
  ND2D1BWP12T U1548 ( .A1(n3969), .A2(n3968), .ZN(n5559) );
  INVD1BWP12T U1549 ( .I(n5559), .ZN(n3970) );
  ND2D1BWP12T U1550 ( .A1(n3972), .A2(n3971), .ZN(n5145) );
  ND2D1BWP12T U1551 ( .A1(n3976), .A2(n3975), .ZN(n5599) );
  TPOAI21D1BWP12T U1552 ( .A1(n5598), .A2(n5600), .B(n5599), .ZN(n4956) );
  OAI21D1BWP12T U1553 ( .A1(n3980), .A2(n3979), .B(n3977), .ZN(n3978) );
  IOA21D1BWP12T U1554 ( .A1(n3980), .A2(n3979), .B(n3978), .ZN(n3995) );
  FA1D2BWP12T U1555 ( .A(n3983), .B(n3982), .CI(n3981), .CO(n3994), .S(n3979)
         );
  FA1D0BWP12T U1556 ( .A(n3986), .B(n3985), .CI(n3984), .CO(n3992), .S(n3993)
         );
  NR2D1BWP12T U1557 ( .A1(n3997), .A2(n3996), .ZN(n5522) );
  FA1D0BWP12T U1558 ( .A(n3992), .B(n3991), .CI(n3990), .CO(n4002), .S(n3999)
         );
  FA1D0BWP12T U1559 ( .A(n3995), .B(n3994), .CI(n3993), .CO(n3998), .S(n3997)
         );
  NR2D1BWP12T U1560 ( .A1(n5522), .A2(n4957), .ZN(n4001) );
  ND2D1BWP12T U1561 ( .A1(n3997), .A2(n3996), .ZN(n5523) );
  ND2D1BWP12T U1562 ( .A1(n3999), .A2(n3998), .ZN(n4958) );
  TPAOI21D1BWP12T U1563 ( .A1(n4956), .A2(n4001), .B(n4000), .ZN(n6055) );
  ND2D1BWP12T U1564 ( .A1(n4003), .A2(n4002), .ZN(n6053) );
  CKND2D1BWP12T U1565 ( .A1(n4005), .A2(n4004), .ZN(n6057) );
  OAI21D1BWP12T U1566 ( .A1(n6056), .A2(n6053), .B(n6057), .ZN(n5495) );
  ND2D1BWP12T U1567 ( .A1(n4007), .A2(n4006), .ZN(n6061) );
  ND2D1BWP12T U1568 ( .A1(n4009), .A2(n4008), .ZN(n5501) );
  TPAOI21D1BWP12T U1569 ( .A1(n4011), .A2(n5495), .B(n4010), .ZN(n4012) );
  FA1D0BWP12T U1570 ( .A(n4016), .B(n4015), .CI(n4014), .CO(n3583), .S(n4017)
         );
  INVD1BWP12T U1571 ( .I(n4017), .ZN(n4021) );
  NR2D2BWP12T U1572 ( .A1(n3406), .A2(n4021), .ZN(n6006) );
  FA1D0BWP12T U1573 ( .A(n4020), .B(n4019), .CI(n4018), .CO(n6009), .S(n3623)
         );
  INVD0BWP12T U1574 ( .I(n6009), .ZN(n4022) );
  TPND2D2BWP12T U1575 ( .A1(n3406), .A2(n4021), .ZN(n6007) );
  OA21D4BWP12T U1576 ( .A1(n6006), .A2(n4022), .B(n6007), .Z(n5457) );
  ND2D1BWP12T U1577 ( .A1(n4024), .A2(n4023), .ZN(n5455) );
  TPOAI21D4BWP12T U1578 ( .A1(n5454), .A2(n5457), .B(n5455), .ZN(n4705) );
  INVD2BWP12T U1579 ( .I(n4705), .ZN(n5059) );
  FA1D0BWP12T U1580 ( .A(n4028), .B(n4027), .CI(n4026), .CO(n4453), .S(n4062)
         );
  MUX2NXD0BWP12T U1581 ( .I0(n4747), .I1(n4746), .S(b[19]), .ZN(n4030) );
  MUX2ND0BWP12T U1582 ( .I0(n5860), .I1(n5861), .S(n4112), .ZN(n4029) );
  NR2D1BWP12T U1583 ( .A1(n4030), .A2(n4029), .ZN(n4452) );
  MUX2ND0BWP12T U1584 ( .I0(n5776), .I1(n5775), .S(b[13]), .ZN(n4032) );
  MUX2NXD1BWP12T U1585 ( .I0(n5778), .I1(n5777), .S(b[12]), .ZN(n4031) );
  NR2D1BWP12T U1586 ( .A1(n4032), .A2(n4031), .ZN(n4447) );
  MUX2ND0BWP12T U1587 ( .I0(n5803), .I1(n5802), .S(n6334), .ZN(n4034) );
  MUX2NXD0BWP12T U1588 ( .I0(n5804), .I1(n5805), .S(n5767), .ZN(n4033) );
  NR2D1BWP12T U1589 ( .A1(n4034), .A2(n4033), .ZN(n4446) );
  MUX2ND0BWP12T U1590 ( .I0(n5406), .I1(n5407), .S(n6565), .ZN(n4035) );
  NR2D1BWP12T U1591 ( .A1(n4036), .A2(n4035), .ZN(n4445) );
  MUX2D1BWP12T U1592 ( .I0(n5761), .I1(n5760), .S(n5379), .Z(n4037) );
  ND2D1BWP12T U1593 ( .A1(n4038), .A2(n4037), .ZN(n4040) );
  ND2D1BWP12T U1594 ( .A1(n4040), .A2(n4039), .ZN(n4459) );
  MAOI222D1BWP12T U1595 ( .A(n4043), .B(n4042), .C(n4041), .ZN(n4537) );
  MUX2ND0BWP12T U1596 ( .I0(n5811), .I1(n5810), .S(b[21]), .ZN(n4045) );
  MUX2ND0BWP12T U1597 ( .I0(n5813), .I1(n5812), .S(b[20]), .ZN(n4044) );
  NR2D1BWP12T U1598 ( .A1(n4045), .A2(n4044), .ZN(n4414) );
  INVD1BWP12T U1599 ( .I(a[22]), .ZN(n5487) );
  OAI21D0BWP12T U1600 ( .A1(a[22]), .A2(a[21]), .B(n4829), .ZN(n4046) );
  INVD1BWP12T U1601 ( .I(a[23]), .ZN(n5069) );
  OAI211D1BWP12T U1602 ( .A1(n5487), .A2(n6623), .B(n4046), .C(a[23]), .ZN(
        n4413) );
  MUX2NXD0BWP12T U1603 ( .I0(n5819), .I1(n5818), .S(n5806), .ZN(n4047) );
  NR2D1BWP12T U1604 ( .A1(n4048), .A2(n4047), .ZN(n4412) );
  FA1D0BWP12T U1605 ( .A(n4051), .B(n4050), .CI(n4049), .CO(n4678), .S(n4075)
         );
  MAOI222D1BWP12T U1606 ( .A(n4054), .B(n4053), .C(n4052), .ZN(n4055) );
  INVD1BWP12T U1607 ( .I(n4055), .ZN(n4545) );
  FA1D0BWP12T U1608 ( .A(n4058), .B(n4057), .CI(n4056), .CO(n4544), .S(n4051)
         );
  FA1D0BWP12T U1609 ( .A(n4061), .B(n4060), .CI(n4059), .CO(n4529), .S(n4052)
         );
  INVD1BWP12T U1610 ( .I(n4062), .ZN(n4064) );
  MAOI222D0BWP12T U1611 ( .A(n4065), .B(n4064), .C(n4063), .ZN(n4528) );
  MUX2D1BWP12T U1612 ( .I0(n4371), .I1(n4372), .S(n4092), .Z(n4066) );
  NR2D1BWP12T U1613 ( .A1(n4067), .A2(n4066), .ZN(n4454) );
  MUX2ND0BWP12T U1614 ( .I0(a[23]), .I1(a[22]), .S(n4823), .ZN(n6550) );
  INVD1BWP12T U1615 ( .I(n6550), .ZN(n5020) );
  INVD1BWP12T U1616 ( .I(n5807), .ZN(n4742) );
  XNR2D1BWP12T U1617 ( .A1(a[23]), .A2(n4498), .ZN(n4386) );
  MUX2NXD1BWP12T U1618 ( .I0(n4757), .I1(n4756), .S(b[15]), .ZN(n4069) );
  MUX2ND0BWP12T U1619 ( .I0(n4759), .I1(n4760), .S(b[14]), .ZN(n4068) );
  ND2D1BWP12T U1620 ( .A1(n4069), .A2(n4068), .ZN(n4423) );
  MUX2NXD0BWP12T U1621 ( .I0(n5870), .I1(n5869), .S(b[9]), .ZN(n4071) );
  MUX2NXD0BWP12T U1622 ( .I0(n5871), .I1(n5872), .S(n4515), .ZN(n4070) );
  NR2D1BWP12T U1623 ( .A1(n4071), .A2(n4070), .ZN(n4426) );
  XOR3D1BWP12T U1624 ( .A1(n4424), .A2(n4423), .A3(n4426), .Z(n4456) );
  MAOI222D1BWP12T U1625 ( .A(n4074), .B(n4073), .C(n4072), .ZN(n4455) );
  XOR3D1BWP12T U1626 ( .A1(n4454), .A2(n4456), .A3(n4455), .Z(n4527) );
  FA1D0BWP12T U1627 ( .A(n4077), .B(n4076), .CI(n4075), .CO(n4684), .S(n3539)
         );
  INVD1BWP12T U1628 ( .I(n4078), .ZN(n4079) );
  NR2D1BWP12T U1629 ( .A1(n4080), .A2(n4079), .ZN(n5058) );
  ND2D1BWP12T U1630 ( .A1(n4080), .A2(n4079), .ZN(n5057) );
  ND2D1BWP12T U1631 ( .A1(n4688), .A2(n5057), .ZN(n4081) );
  XOR2D1BWP12T U1632 ( .A1(n5059), .A2(n4081), .Z(n6066) );
  ND2D1BWP12T U1633 ( .A1(op[1]), .A2(n4172), .ZN(n4221) );
  INVD1BWP12T U1634 ( .I(op[3]), .ZN(n4134) );
  ND2D1BWP12T U1635 ( .A1(op[2]), .A2(n4134), .ZN(n4173) );
  NR2D1BWP12T U1636 ( .A1(n4221), .A2(n4173), .ZN(n6898) );
  IND2D1BWP12T U1637 ( .A1(a[14]), .B1(b[14]), .ZN(n6456) );
  IND2D1BWP12T U1638 ( .A1(b[14]), .B1(a[14]), .ZN(n6477) );
  ND2D1BWP12T U1639 ( .A1(n6456), .A2(n6477), .ZN(n5608) );
  IND2D1BWP12T U1640 ( .A1(n6231), .B1(b[12]), .ZN(n5149) );
  TPNR2D0BWP12T U1641 ( .A1(n5608), .A2(n5601), .ZN(n4090) );
  NR2D1BWP12T U1642 ( .A1(n4745), .A2(n6230), .ZN(n4209) );
  IND2D1BWP12T U1643 ( .A1(n6715), .B1(n5806), .ZN(n6129) );
  INVD1BWP12T U1644 ( .I(n6450), .ZN(n4088) );
  IND2D1BWP12T U1645 ( .A1(a[0]), .B1(n6248), .ZN(n4205) );
  INVD1BWP12T U1646 ( .I(n4205), .ZN(n6457) );
  INVD1BWP12T U1647 ( .I(a[0]), .ZN(n5362) );
  OAI21D1BWP12T U1648 ( .A1(n4299), .A2(n6488), .B(n4304), .ZN(n4300) );
  NR2D1BWP12T U1649 ( .A1(n4307), .A2(n4498), .ZN(n6498) );
  INVD1BWP12T U1650 ( .I(n6498), .ZN(n4310) );
  ND2D1BWP12T U1651 ( .A1(n4300), .A2(n4310), .ZN(n6136) );
  ND2D1BWP12T U1652 ( .A1(a[2]), .A2(n6520), .ZN(n6881) );
  INVD1BWP12T U1653 ( .I(n6881), .ZN(n4082) );
  TPNR2D1BWP12T U1654 ( .A1(a[2]), .A2(n6520), .ZN(n6875) );
  INVD1BWP12T U1655 ( .I(n5979), .ZN(n6180) );
  ND2D1BWP12T U1656 ( .A1(n6136), .A2(n6180), .ZN(n4946) );
  CKND1BWP12T U1657 ( .I(a[2]), .ZN(n6887) );
  NR2D1BWP12T U1658 ( .A1(n6887), .A2(n6520), .ZN(n6497) );
  INVD1BWP12T U1659 ( .I(n4938), .ZN(n6479) );
  IND2D1BWP12T U1660 ( .A1(n6573), .B1(n6249), .ZN(n5255) );
  INVD1BWP12T U1661 ( .I(n5255), .ZN(n5976) );
  AOI211D1BWP12T U1662 ( .A1(n5226), .A2(n6497), .B(n6479), .C(n5976), .ZN(
        n4083) );
  OAI21D1BWP12T U1663 ( .A1(n4946), .A2(n4952), .B(n4083), .ZN(n5137) );
  NR2D1BWP12T U1664 ( .A1(n4433), .A2(n6267), .ZN(n6463) );
  IND2D1BWP12T U1665 ( .A1(n6249), .B1(n6573), .ZN(n5256) );
  CKND0BWP12T U1666 ( .I(n5256), .ZN(n6468) );
  TPNR2D0BWP12T U1667 ( .A1(n6463), .A2(n6468), .ZN(n4084) );
  TPND2D0BWP12T U1668 ( .A1(n5137), .A2(n4084), .ZN(n4086) );
  INVD1BWP12T U1669 ( .I(a[6]), .ZN(n5240) );
  NR2D1BWP12T U1670 ( .A1(n5240), .A2(b[6]), .ZN(n6499) );
  NR2D1BWP12T U1671 ( .A1(n6788), .A2(n6782), .ZN(n5138) );
  TPNR2D0BWP12T U1672 ( .A1(n6499), .A2(n5138), .ZN(n4085) );
  IND2D1BWP12T U1673 ( .A1(a[6]), .B1(n5864), .ZN(n4206) );
  INVD1BWP12T U1674 ( .I(n4206), .ZN(n6464) );
  AOI21D1BWP12T U1675 ( .A1(n4086), .A2(n4085), .B(n6464), .ZN(n6132) );
  IND2D1BWP12T U1676 ( .A1(n5379), .B1(n6819), .ZN(n6812) );
  INVD1BWP12T U1677 ( .I(n6812), .ZN(n6484) );
  NR2D1BWP12T U1678 ( .A1(n4343), .A2(n6819), .ZN(n6465) );
  INVD1BWP12T U1679 ( .I(n6465), .ZN(n6814) );
  OAI21D1BWP12T U1680 ( .A1(n6132), .A2(n6484), .B(n6814), .ZN(n6130) );
  IND2D1BWP12T U1681 ( .A1(a[8]), .B1(n5843), .ZN(n4207) );
  INVD1BWP12T U1682 ( .I(n4207), .ZN(n6743) );
  NR2D1BWP12T U1683 ( .A1(n6760), .A2(n5843), .ZN(n6746) );
  INVD1BWP12T U1684 ( .I(n6746), .ZN(n4087) );
  OAI21D1BWP12T U1685 ( .A1(n6130), .A2(n6743), .B(n4087), .ZN(n5196) );
  IND2D1BWP12T U1686 ( .A1(b[9]), .B1(n6229), .ZN(n4208) );
  INVD1BWP12T U1687 ( .I(n4208), .ZN(n6485) );
  NR2D1BWP12T U1688 ( .A1(n4730), .A2(n6229), .ZN(n6460) );
  INVD1BWP12T U1689 ( .I(n6460), .ZN(n5210) );
  OAI21D1BWP12T U1690 ( .A1(n5196), .A2(n6485), .B(n5210), .ZN(n4230) );
  NR2D1BWP12T U1691 ( .A1(n5232), .A2(n5806), .ZN(n6486) );
  INVD1BWP12T U1692 ( .I(n6486), .ZN(n4260) );
  ND2D1BWP12T U1693 ( .A1(n4230), .A2(n4260), .ZN(n6128) );
  IND2D1BWP12T U1694 ( .A1(b[11]), .B1(n6230), .ZN(n4210) );
  INVD1BWP12T U1695 ( .I(n4210), .ZN(n6481) );
  AOI21D1BWP12T U1696 ( .A1(n4088), .A2(n6128), .B(n6481), .ZN(n5565) );
  IND2D1BWP12T U1697 ( .A1(b[12]), .B1(n6231), .ZN(n4211) );
  ND2D1BWP12T U1698 ( .A1(n5149), .A2(n4211), .ZN(n5567) );
  INVD1BWP12T U1699 ( .I(n5567), .ZN(n5566) );
  TPND2D1BWP12T U1700 ( .A1(n5565), .A2(n5566), .ZN(n5602) );
  IND2D1BWP12T U1701 ( .A1(b[13]), .B1(a[13]), .ZN(n5183) );
  TPOAI21D0BWP12T U1702 ( .A1(n5608), .A2(n5183), .B(n6477), .ZN(n4089) );
  AOI21D1BWP12T U1703 ( .A1(n4090), .A2(n5602), .B(n4089), .ZN(n5526) );
  NR2D1BWP12T U1704 ( .A1(n5538), .A2(b[15]), .ZN(n6482) );
  CKND0BWP12T U1705 ( .I(n6482), .ZN(n4091) );
  IND2D1BWP12T U1706 ( .A1(n6232), .B1(b[15]), .ZN(n4212) );
  INVD1BWP12T U1707 ( .I(n4212), .ZN(n6461) );
  AOI21D1BWP12T U1708 ( .A1(n5526), .A2(n4091), .B(n6461), .ZN(n4963) );
  INVD1BWP12T U1709 ( .I(a[16]), .ZN(n4967) );
  NR2D1BWP12T U1710 ( .A1(n4967), .A2(b[16]), .ZN(n6495) );
  NR2D1BWP12T U1711 ( .A1(n4092), .A2(a[16]), .ZN(n6473) );
  NR2D1BWP12T U1712 ( .A1(n6495), .A2(n6473), .ZN(n5000) );
  INVD1BWP12T U1713 ( .I(n5000), .ZN(n4214) );
  INVD0BWP12T U1714 ( .I(n6473), .ZN(n4093) );
  OAI21D1BWP12T U1715 ( .A1(n4963), .A2(n4214), .B(n4093), .ZN(n5703) );
  NR2D1BWP12T U1716 ( .A1(n5728), .A2(b[17]), .ZN(n6502) );
  INVD1BWP12T U1717 ( .I(n6502), .ZN(n5713) );
  ND2D1BWP12T U1718 ( .A1(n5703), .A2(n5713), .ZN(n6126) );
  IND2D1BWP12T U1719 ( .A1(a[17]), .B1(b[17]), .ZN(n5970) );
  IND2D1BWP12T U1720 ( .A1(a[18]), .B1(b[18]), .ZN(n5926) );
  ND2D1BWP12T U1721 ( .A1(n5970), .A2(n5926), .ZN(n4215) );
  INVD1BWP12T U1722 ( .I(n4215), .ZN(n6458) );
  IND2D1BWP12T U1723 ( .A1(b[18]), .B1(a[18]), .ZN(n5925) );
  INVD1BWP12T U1724 ( .I(n5925), .ZN(n6483) );
  AOI21D1BWP12T U1725 ( .A1(n6126), .A2(n6458), .B(n6483), .ZN(n6125) );
  IND2D1BWP12T U1726 ( .A1(a[19]), .B1(b[19]), .ZN(n6459) );
  IND2D1BWP12T U1727 ( .A1(b[19]), .B1(a[19]), .ZN(n4094) );
  ND2D1BWP12T U1728 ( .A1(n6459), .A2(n4094), .ZN(n6170) );
  NR2D1BWP12T U1729 ( .A1(n6125), .A2(n6170), .ZN(n6124) );
  INVD1BWP12T U1730 ( .I(n4094), .ZN(n6656) );
  IND2D1BWP12T U1731 ( .A1(a[20]), .B1(b[20]), .ZN(n5460) );
  IND2D1BWP12T U1732 ( .A1(b[20]), .B1(a[20]), .ZN(n6487) );
  ND2D1BWP12T U1733 ( .A1(n5460), .A2(n6487), .ZN(n5515) );
  INVD1BWP12T U1734 ( .I(n5515), .ZN(n5504) );
  OAI21D1BWP12T U1735 ( .A1(n6124), .A2(n6656), .B(n5504), .ZN(n5503) );
  CKND2D1BWP12T U1736 ( .A1(n5503), .A2(n6487), .ZN(n6150) );
  IND2D1BWP12T U1737 ( .A1(a[21]), .B1(b[21]), .ZN(n6472) );
  IND2D1BWP12T U1738 ( .A1(b[21]), .B1(a[21]), .ZN(n5463) );
  ND2D1BWP12T U1739 ( .A1(n6472), .A2(n5463), .ZN(n6168) );
  INVD1BWP12T U1740 ( .I(n6168), .ZN(n6618) );
  ND2D1BWP12T U1741 ( .A1(n6150), .A2(n6618), .ZN(n6149) );
  CKND2D1BWP12T U1742 ( .A1(n6149), .A2(n5463), .ZN(n5464) );
  IND2D1BWP12T U1743 ( .A1(a[22]), .B1(b[22]), .ZN(n6471) );
  IND2D1BWP12T U1744 ( .A1(b[22]), .B1(a[22]), .ZN(n4219) );
  ND2D1BWP12T U1745 ( .A1(n6471), .A2(n4219), .ZN(n5489) );
  INVD1BWP12T U1746 ( .I(n5489), .ZN(n4216) );
  ND2D1BWP12T U1747 ( .A1(n5464), .A2(n4216), .ZN(n4095) );
  ND2D1BWP12T U1748 ( .A1(n4095), .A2(n4219), .ZN(n4096) );
  NR2D1BWP12T U1749 ( .A1(n5069), .A2(b[23]), .ZN(n5095) );
  INVD1BWP12T U1750 ( .I(b[23]), .ZN(n4363) );
  NR2D1BWP12T U1751 ( .A1(n4363), .A2(a[23]), .ZN(n6453) );
  NR2D1BWP12T U1752 ( .A1(n5095), .A2(n6453), .ZN(n4217) );
  CKND2D2BWP12T U1753 ( .A1(n4096), .A2(n4217), .ZN(n6155) );
  CKND0BWP12T U1754 ( .I(n4217), .ZN(n4220) );
  INVD0BWP12T U1755 ( .I(n4173), .ZN(n4880) );
  ND2D1BWP12T U1756 ( .A1(n4175), .A2(n4880), .ZN(n6794) );
  ND2D1BWP12T U1757 ( .A1(a[20]), .A2(b[20]), .ZN(n5508) );
  ND2D1BWP12T U1758 ( .A1(a[19]), .A2(b[19]), .ZN(n6651) );
  ND2D1BWP12T U1759 ( .A1(n5508), .A2(n6651), .ZN(n6091) );
  INVD1BWP12T U1760 ( .I(n6091), .ZN(n4115) );
  INVD1BWP12T U1761 ( .I(n5204), .ZN(n5200) );
  ND2D1BWP12T U1762 ( .A1(n6715), .A2(n5806), .ZN(n6197) );
  CKND2D0BWP12T U1763 ( .A1(n6093), .A2(n6197), .ZN(n4104) );
  INVD1BWP12T U1764 ( .I(n6175), .ZN(n4101) );
  ND2D1BWP12T U1765 ( .A1(n5240), .A2(n4357), .ZN(n5126) );
  CKND0BWP12T U1766 ( .I(n5126), .ZN(n6190) );
  ND2D1BWP12T U1767 ( .A1(a[0]), .A2(n4823), .ZN(n6121) );
  INVD1BWP12T U1768 ( .I(n6121), .ZN(n5738) );
  ND2D1BWP12T U1769 ( .A1(n4303), .A2(n5738), .ZN(n4320) );
  ND2D1BWP12T U1770 ( .A1(n4320), .A2(n6098), .ZN(n5931) );
  INVD1BWP12T U1771 ( .I(n6488), .ZN(n5072) );
  ND2D1BWP12T U1772 ( .A1(n4205), .A2(n5072), .ZN(n6606) );
  ND2D1BWP12T U1773 ( .A1(n6606), .A2(c_in), .ZN(n5735) );
  NR2D1BWP12T U1774 ( .A1(n5735), .A2(n4304), .ZN(n4322) );
  NR2D1BWP12T U1775 ( .A1(n5931), .A2(n4322), .ZN(n6181) );
  ND2D1BWP12T U1776 ( .A1(n5254), .A2(n6576), .ZN(n5267) );
  ND2XD0BWP12T U1777 ( .A1(n5979), .A2(n5267), .ZN(n4098) );
  ND2D1BWP12T U1778 ( .A1(n6247), .A2(n6334), .ZN(n5273) );
  CKND2D1BWP12T U1779 ( .A1(n6881), .A2(n5273), .ZN(n6090) );
  AOI21D1BWP12T U1780 ( .A1(n6090), .A2(n5267), .B(n5274), .ZN(n4097) );
  OAI21D1BWP12T U1781 ( .A1(n6181), .A2(n4098), .B(n4097), .ZN(n4099) );
  CKND2D1BWP12T U1782 ( .A1(n4099), .A2(n5259), .ZN(n5107) );
  ND2D1BWP12T U1783 ( .A1(a[6]), .A2(b[6]), .ZN(n5929) );
  ND2D1BWP12T U1784 ( .A1(n5126), .A2(n5929), .ZN(n5139) );
  INVD1BWP12T U1785 ( .I(n5139), .ZN(n5116) );
  CKND2D1BWP12T U1786 ( .A1(n5116), .A2(n6096), .ZN(n5108) );
  TPAOI21D0BWP12T U1787 ( .A1(n5108), .A2(n5126), .B(n6133), .ZN(n4100) );
  OAI31D1BWP12T U1788 ( .A1(n6190), .A2(n6134), .A3(n5107), .B(n4100), .ZN(
        n6187) );
  CKND2D1BWP12T U1789 ( .A1(n6187), .A2(n6815), .ZN(n6174) );
  INR2XD0BWP12T U1790 ( .A1(n4101), .B1(n6174), .ZN(n6173) );
  INVD1BWP12T U1791 ( .I(n6197), .ZN(n4102) );
  NR2D1BWP12T U1792 ( .A1(n4102), .A2(n4259), .ZN(n4233) );
  INVD1BWP12T U1793 ( .I(n4238), .ZN(n5213) );
  CKND2D1BWP12T U1794 ( .A1(n4233), .A2(n5213), .ZN(n4235) );
  AOI21D0BWP12T U1795 ( .A1(n4235), .A2(n6197), .B(n6707), .ZN(n4103) );
  OAI31D1BWP12T U1796 ( .A1(n5200), .A2(n4104), .A3(n6173), .B(n4103), .ZN(
        n5156) );
  ND2D1BWP12T U1797 ( .A1(n6231), .A2(b[12]), .ZN(n6112) );
  AN2XD0BWP12T U1798 ( .A1(n6112), .A2(n6706), .Z(n4106) );
  ND2D1BWP12T U1799 ( .A1(a[13]), .A2(b[13]), .ZN(n4126) );
  NR2D1BWP12T U1800 ( .A1(a[13]), .A2(b[13]), .ZN(n5185) );
  INR2D1BWP12T U1801 ( .A1(n4126), .B1(n5185), .ZN(n5151) );
  NR2D1BWP12T U1802 ( .A1(n6231), .A2(b[12]), .ZN(n4125) );
  INVD1BWP12T U1803 ( .I(n4125), .ZN(n5581) );
  CKND2D1BWP12T U1804 ( .A1(n5151), .A2(n5581), .ZN(n4105) );
  ND2D1BWP12T U1805 ( .A1(n6232), .A2(b[15]), .ZN(n6094) );
  NR2D1BWP12T U1806 ( .A1(n6232), .A2(b[15]), .ZN(n5542) );
  INR2D1BWP12T U1807 ( .A1(n6094), .B1(n5542), .ZN(n5530) );
  NR2D1BWP12T U1808 ( .A1(a[14]), .A2(b[14]), .ZN(n5628) );
  INVD1BWP12T U1809 ( .I(n5628), .ZN(n5529) );
  TPND2D0BWP12T U1810 ( .A1(n5530), .A2(n5529), .ZN(n4108) );
  CKND1BWP12T U1811 ( .I(n4108), .ZN(n4110) );
  ND2D1BWP12T U1812 ( .A1(a[14]), .A2(b[14]), .ZN(n4127) );
  CKND2D1BWP12T U1813 ( .A1(n4127), .A2(n4126), .ZN(n6089) );
  INVD0BWP12T U1814 ( .I(n6089), .ZN(n4107) );
  RCOAI21D0BWP12T U1815 ( .A1(n4108), .A2(n4107), .B(n6094), .ZN(n4109) );
  AOI21D1BWP12T U1816 ( .A1(n5607), .A2(n4110), .B(n4109), .ZN(n4964) );
  ND2D1BWP12T U1817 ( .A1(a[16]), .A2(b[16]), .ZN(n6114) );
  NR2D1BWP12T U1818 ( .A1(a[16]), .A2(b[16]), .ZN(n4128) );
  TPAOI21D1BWP12T U1819 ( .A1(n4964), .A2(n6114), .B(n4128), .ZN(n5706) );
  NR2D1BWP12T U1820 ( .A1(a[17]), .A2(b[17]), .ZN(n5712) );
  INVD1BWP12T U1821 ( .I(n5712), .ZN(n4111) );
  ND2D1BWP12T U1822 ( .A1(a[17]), .A2(b[17]), .ZN(n6115) );
  ND2D1BWP12T U1823 ( .A1(n4111), .A2(n6115), .ZN(n5705) );
  ND2D1BWP12T U1824 ( .A1(a[18]), .A2(b[18]), .ZN(n6095) );
  INVD1BWP12T U1825 ( .I(a[18]), .ZN(n6646) );
  ND2D1BWP12T U1826 ( .A1(n6646), .A2(n4112), .ZN(n6684) );
  INVD1BWP12T U1827 ( .I(n6684), .ZN(n4113) );
  NR2D1BWP12T U1828 ( .A1(a[19]), .A2(b[19]), .ZN(n4129) );
  INVD1BWP12T U1829 ( .I(n4129), .ZN(n6652) );
  CKND2D1BWP12T U1830 ( .A1(n6171), .A2(n6652), .ZN(n5514) );
  INVD1BWP12T U1831 ( .I(a[20]), .ZN(n4972) );
  ND2D1BWP12T U1832 ( .A1(n4972), .A2(n4494), .ZN(n4130) );
  INVD1BWP12T U1833 ( .I(n4130), .ZN(n4114) );
  AOI21D1BWP12T U1834 ( .A1(n4115), .A2(n5514), .B(n4114), .ZN(n6169) );
  ND2D1BWP12T U1835 ( .A1(a[21]), .A2(b[21]), .ZN(n6627) );
  CKND0BWP12T U1836 ( .I(n6627), .ZN(n4116) );
  NR2D1BWP12T U1837 ( .A1(a[21]), .A2(b[21]), .ZN(n4131) );
  INVD1BWP12T U1838 ( .I(n4131), .ZN(n6622) );
  OAI21D1BWP12T U1839 ( .A1(n6169), .A2(n4116), .B(n6622), .ZN(n5466) );
  NR2D1BWP12T U1840 ( .A1(a[22]), .A2(b[22]), .ZN(n4132) );
  TPND2D0BWP12T U1841 ( .A1(a[22]), .A2(b[22]), .ZN(n4133) );
  OA21D1BWP12T U1842 ( .A1(n5466), .A2(n4132), .B(n4133), .Z(n4797) );
  CKND2D1BWP12T U1843 ( .A1(n5931), .A2(n5979), .ZN(n5930) );
  ND2D1BWP12T U1844 ( .A1(n5930), .A2(n6881), .ZN(n4932) );
  TPNR2D0BWP12T U1845 ( .A1(n5226), .A2(n5274), .ZN(n4117) );
  ND2D1BWP12T U1846 ( .A1(n4932), .A2(n4117), .ZN(n5115) );
  NR3D1BWP12T U1847 ( .A1(n6133), .A2(n5139), .A3(n5113), .ZN(n4120) );
  INVD1BWP12T U1848 ( .I(n4120), .ZN(n4122) );
  AN2XD0BWP12T U1849 ( .A1(n6097), .A2(n6096), .Z(n4118) );
  TPOAI21D0BWP12T U1850 ( .A1(n5274), .A2(n5273), .B(n4118), .ZN(n5112) );
  OAI211D1BWP12T U1851 ( .A1(n5929), .A2(n6133), .B(n6811), .C(n6093), .ZN(
        n4119) );
  TPAOI21D0BWP12T U1852 ( .A1(n5112), .A2(n4120), .B(n4119), .ZN(n4121) );
  OAI21D1BWP12T U1853 ( .A1(n5115), .A2(n4122), .B(n4121), .ZN(n4232) );
  OAI21D0BWP12T U1854 ( .A1(n5204), .A2(n4238), .B(n4233), .ZN(n4123) );
  TPAOI31D0BWP12T U1855 ( .A1(n4232), .A2(n4231), .A3(n5213), .B(n4123), .ZN(
        n4124) );
  NR2XD0BWP12T U1856 ( .A1(n4124), .A2(n4259), .ZN(n5942) );
  TPOAI21D1BWP12T U1857 ( .A1(n5942), .A2(n6707), .B(n6703), .ZN(n5568) );
  OAI21D1BWP12T U1858 ( .A1(n5568), .A2(n4125), .B(n6112), .ZN(n5155) );
  INVD1BWP12T U1859 ( .I(n4126), .ZN(n5606) );
  AOI21D1BWP12T U1860 ( .A1(n5155), .A2(n5151), .B(n5606), .ZN(n5605) );
  AO21D1BWP12T U1861 ( .A1(n5605), .A2(n4127), .B(n5628), .Z(n5528) );
  AO21D1BWP12T U1862 ( .A1(n5528), .A2(n6094), .B(n5542), .Z(n4962) );
  AO21D1BWP12T U1863 ( .A1(n4962), .A2(n6114), .B(n4128), .Z(n5704) );
  TPAOI21D1BWP12T U1864 ( .A1(n5704), .A2(n6115), .B(n5712), .ZN(n5927) );
  INVD1BWP12T U1865 ( .I(n6095), .ZN(n6685) );
  OAI21D1BWP12T U1866 ( .A1(n5927), .A2(n6685), .B(n6684), .ZN(n5924) );
  OAI21D1BWP12T U1867 ( .A1(n5505), .A2(n6091), .B(n4130), .ZN(n5923) );
  OA21D1BWP12T U1868 ( .A1(n5923), .A2(n4131), .B(n6627), .Z(n5488) );
  AO21D1BWP12T U1869 ( .A1(n5488), .A2(n4133), .B(n4132), .Z(n4333) );
  NR2D1BWP12T U1870 ( .A1(op[2]), .A2(n4134), .ZN(n5736) );
  CKND1BWP12T U1871 ( .I(n5736), .ZN(n4222) );
  ND2D1BWP12T U1872 ( .A1(op[0]), .A2(op[1]), .ZN(n4179) );
  NR2D1BWP12T U1873 ( .A1(n4222), .A2(n4179), .ZN(n6833) );
  CKND2D1BWP12T U1874 ( .A1(n5958), .A2(n6833), .ZN(n4203) );
  NR2D1BWP12T U1875 ( .A1(a[0]), .A2(n5360), .ZN(n5762) );
  ND2D1BWP12T U1876 ( .A1(n6789), .A2(n4136), .ZN(n6818) );
  NR2D1BWP12T U1877 ( .A1(n6818), .A2(n6756), .ZN(n5215) );
  ND2D1BWP12T U1878 ( .A1(n5215), .A2(n5231), .ZN(n4252) );
  TPND2D0BWP12T U1879 ( .A1(n6708), .A2(n5232), .ZN(n4137) );
  NR2D1BWP12T U1880 ( .A1(n4252), .A2(n4137), .ZN(n6714) );
  NR2D1BWP12T U1881 ( .A1(a[13]), .A2(n6231), .ZN(n4138) );
  CKND2D1BWP12T U1882 ( .A1(n6714), .A2(n4138), .ZN(n5635) );
  NR2D1BWP12T U1883 ( .A1(n5635), .A2(a[14]), .ZN(n5636) );
  INVD1BWP12T U1884 ( .I(n4139), .ZN(n5725) );
  NR2D1BWP12T U1885 ( .A1(n5725), .A2(a[17]), .ZN(n4140) );
  ND2D1BWP12T U1886 ( .A1(n5636), .A2(n4140), .ZN(n6678) );
  ND2D1BWP12T U1887 ( .A1(n6654), .A2(n6646), .ZN(n4141) );
  NR2D1BWP12T U1888 ( .A1(n6678), .A2(n4141), .ZN(n6648) );
  CKND2D1BWP12T U1889 ( .A1(n6648), .A2(n4972), .ZN(n6635) );
  NR2D1BWP12T U1890 ( .A1(n6635), .A2(a[21]), .ZN(n6634) );
  ND2D1BWP12T U1891 ( .A1(n6634), .A2(n5487), .ZN(n4811) );
  ND2D1BWP12T U1892 ( .A1(n5736), .A2(n4175), .ZN(n6862) );
  TPNR2D0BWP12T U1893 ( .A1(n4811), .A2(n6862), .ZN(n5070) );
  ND2D1BWP12T U1894 ( .A1(n4811), .A2(n6786), .ZN(n5482) );
  NR2D1BWP12T U1895 ( .A1(op[2]), .A2(op[3]), .ZN(n4174) );
  INVD1BWP12T U1896 ( .I(n6680), .ZN(n6855) );
  ND2D1BWP12T U1897 ( .A1(n5767), .A2(n3463), .ZN(n6534) );
  INVD1BWP12T U1898 ( .I(n6534), .ZN(n6553) );
  INVD1BWP12T U1899 ( .I(n6531), .ZN(n5023) );
  MUX2D1BWP12T U1900 ( .I0(n6230), .I1(n6715), .S(n6248), .Z(n4889) );
  INVD1BWP12T U1901 ( .I(n4889), .ZN(n5178) );
  NR2D1BWP12T U1902 ( .A1(n5767), .A2(n4498), .ZN(n6556) );
  AOI22D0BWP12T U1903 ( .A1(n6553), .A2(n5023), .B1(n5178), .B2(n6556), .ZN(
        n4143) );
  IND2D1BWP12T U1904 ( .A1(n6520), .B1(n5612), .ZN(n6533) );
  INVD1BWP12T U1905 ( .I(n6533), .ZN(n6552) );
  INVD1BWP12T U1906 ( .I(n5165), .ZN(n5176) );
  ND2D1BWP12T U1907 ( .A1(n6520), .A2(n4498), .ZN(n6530) );
  INVD1BWP12T U1908 ( .I(n6530), .ZN(n6549) );
  AOI22D0BWP12T U1909 ( .A1(n6552), .A2(n5179), .B1(n5176), .B2(n6549), .ZN(
        n4142) );
  ND2D1BWP12T U1910 ( .A1(n4143), .A2(n4142), .ZN(n5434) );
  OAI22D0BWP12T U1911 ( .A1(n6263), .A2(n6534), .B1(n4888), .B2(n6533), .ZN(
        n4147) );
  INVD1BWP12T U1912 ( .I(n6556), .ZN(n5677) );
  INVD1BWP12T U1913 ( .I(n4144), .ZN(n4145) );
  ND2D1BWP12T U1914 ( .A1(n4145), .A2(n6121), .ZN(n4893) );
  OAI22D1BWP12T U1915 ( .A1(n4894), .A2(n5677), .B1(n4893), .B2(n6530), .ZN(
        n4146) );
  NR2D1BWP12T U1916 ( .A1(n4147), .A2(n4146), .ZN(n6516) );
  OAI22D0BWP12T U1917 ( .A1(n6535), .A2(n6533), .B1(n5020), .B2(n6534), .ZN(
        n4149) );
  OAI22D0BWP12T U1918 ( .A1(n6403), .A2(n6530), .B1(n6532), .B2(n5677), .ZN(
        n4148) );
  NR2D1BWP12T U1919 ( .A1(n4149), .A2(n4148), .ZN(n5438) );
  NR2D1BWP12T U1920 ( .A1(n6573), .A2(n6334), .ZN(n6578) );
  INVD1BWP12T U1921 ( .I(n6578), .ZN(n6557) );
  OAI22D1BWP12T U1922 ( .A1(n6516), .A2(n6565), .B1(n5438), .B2(n6557), .ZN(
        n4168) );
  NR2D1BWP12T U1923 ( .A1(b[27]), .A2(b[25]), .ZN(n4151) );
  NR2D1BWP12T U1924 ( .A1(b[24]), .A2(b[23]), .ZN(n4150) );
  ND2D1BWP12T U1925 ( .A1(n4151), .A2(n4150), .ZN(n4166) );
  NR2D1BWP12T U1926 ( .A1(b[11]), .A2(n5843), .ZN(n4154) );
  NR2D1BWP12T U1927 ( .A1(n5379), .A2(n6782), .ZN(n4153) );
  NR2D1BWP12T U1928 ( .A1(n5806), .A2(b[6]), .ZN(n4152) );
  ND4D1BWP12T U1929 ( .A1(n4155), .A2(n4154), .A3(n4153), .A4(n4152), .ZN(
        n4165) );
  NR2D1BWP12T U1930 ( .A1(b[14]), .A2(b[13]), .ZN(n4158) );
  NR2D1BWP12T U1931 ( .A1(b[29]), .A2(b[28]), .ZN(n4157) );
  NR2D1BWP12T U1932 ( .A1(b[30]), .A2(b[31]), .ZN(n4156) );
  NR2D1BWP12T U1933 ( .A1(b[26]), .A2(b[21]), .ZN(n4162) );
  NR2D1BWP12T U1934 ( .A1(b[20]), .A2(b[19]), .ZN(n4161) );
  NR2D2BWP12T U1935 ( .A1(b[18]), .A2(b[17]), .ZN(n4160) );
  ND4D1BWP12T U1936 ( .A1(n4162), .A2(n4161), .A3(n4160), .A4(n5467), .ZN(
        n4163) );
  NR4D1BWP12T U1937 ( .A1(n4166), .A2(n4165), .A3(n4164), .A4(n4163), .ZN(
        n4167) );
  BUFFD6BWP12T U1938 ( .I(n4167), .Z(n6355) );
  ND2D1BWP12T U1939 ( .A1(n6573), .A2(n6334), .ZN(n5305) );
  ND2D1BWP12T U1940 ( .A1(n6355), .A2(n5305), .ZN(n6540) );
  AOI211D1BWP12T U1941 ( .A1(n6334), .A2(n5434), .B(n4168), .C(n6540), .ZN(
        n6542) );
  INVD1BWP12T U1942 ( .I(n6373), .ZN(n4169) );
  TPND2D2BWP12T U1943 ( .A1(n6355), .A2(n4169), .ZN(n4248) );
  NR2D1BWP12T U1944 ( .A1(n4179), .A2(n4173), .ZN(n6857) );
  INVD1BWP12T U1945 ( .I(n6857), .ZN(n6716) );
  ND2D3BWP12T U1946 ( .A1(n4248), .A2(n6716), .ZN(n6905) );
  ND2XD8BWP12T U1947 ( .A1(n6905), .A2(n6565), .ZN(n6840) );
  NR2D1BWP12T U1948 ( .A1(n5237), .A2(n6520), .ZN(n4190) );
  CKND0BWP12T U1949 ( .I(n4190), .ZN(n5437) );
  INVD1BWP12T U1950 ( .I(a[31]), .ZN(n6353) );
  ND2D1BWP12T U1951 ( .A1(a[31]), .A2(n6334), .ZN(n5667) );
  NR2D1BWP12T U1952 ( .A1(n5437), .A2(n5667), .ZN(n6288) );
  INVD1BWP12T U1953 ( .I(n6288), .ZN(n4170) );
  NR2D1BWP12T U1954 ( .A1(n6840), .A2(n4170), .ZN(n4185) );
  INVD1BWP12T U1955 ( .I(op[1]), .ZN(n4171) );
  ND2D1BWP12T U1956 ( .A1(n4172), .A2(n4171), .ZN(n6106) );
  CKND0BWP12T U1957 ( .I(n6106), .ZN(n4176) );
  INVD1BWP12T U1958 ( .I(op[2]), .ZN(n6810) );
  ND2D1BWP12T U1959 ( .A1(n4176), .A2(n6810), .ZN(n6880) );
  ND2D1BWP12T U1960 ( .A1(a[23]), .A2(b[23]), .ZN(n6107) );
  ND2D1BWP12T U1961 ( .A1(n6355), .A2(n6578), .ZN(n6351) );
  NR2D1BWP12T U1962 ( .A1(n6106), .A2(n4173), .ZN(n6909) );
  INVD1BWP12T U1963 ( .I(n6909), .ZN(n6852) );
  NR2D1BWP12T U1964 ( .A1(n6353), .A2(n6852), .ZN(n4819) );
  ND2D1BWP12T U1965 ( .A1(n6351), .A2(n4819), .ZN(n6850) );
  ND2D1BWP12T U1966 ( .A1(n4175), .A2(n4174), .ZN(n6813) );
  INVD1BWP12T U1967 ( .I(n4177), .ZN(n4178) );
  TPNR2D0BWP12T U1968 ( .A1(n4221), .A2(n4178), .ZN(n6655) );
  INVD1BWP12T U1969 ( .I(n6655), .ZN(n6683) );
  ND2D1BWP12T U1970 ( .A1(n6813), .A2(n6683), .ZN(n6745) );
  ND2D1BWP12T U1971 ( .A1(n4177), .A2(n4176), .ZN(n6874) );
  ND2D1BWP12T U1972 ( .A1(a[23]), .A2(n6874), .ZN(n4182) );
  NR2D1BWP12T U1973 ( .A1(b[23]), .A2(a[23]), .ZN(n4180) );
  ND2D1BWP12T U1974 ( .A1(n6874), .A2(n6813), .ZN(n6621) );
  INVD1BWP12T U1975 ( .I(n6621), .ZN(n6751) );
  NR2D1BWP12T U1976 ( .A1(n4179), .A2(n4178), .ZN(n6783) );
  INVD1BWP12T U1977 ( .I(n6783), .ZN(n6844) );
  OAI21D1BWP12T U1978 ( .A1(n4180), .A2(n6751), .B(n6844), .ZN(n4181) );
  AOI22D0BWP12T U1979 ( .A1(n5095), .A2(n6745), .B1(n4182), .B2(n4181), .ZN(
        n4183) );
  OAI211D0BWP12T U1980 ( .A1(n6880), .A2(n6107), .B(n6850), .C(n4183), .ZN(
        n4184) );
  RCAOI211D0BWP12T U1981 ( .A1(n6855), .A2(n6542), .B(n4185), .C(n4184), .ZN(
        n4200) );
  NR2D1BWP12T U1982 ( .A1(n6245), .A2(n5767), .ZN(n4869) );
  ND2D8BWP12T U1983 ( .A1(n4823), .A2(n4498), .ZN(n5235) );
  INR2XD2BWP12T U1984 ( .A1(n5235), .B1(n6245), .ZN(n6264) );
  ND2D1BWP12T U1985 ( .A1(n4186), .A2(n4922), .ZN(n6409) );
  INVD1BWP12T U1986 ( .I(n6409), .ZN(n5289) );
  TPND2D0BWP12T U1987 ( .A1(n5289), .A2(n5035), .ZN(n4189) );
  NR2D4BWP12T U1988 ( .A1(n4186), .A2(n6264), .ZN(n5660) );
  CKND2D0BWP12T U1989 ( .A1(n5660), .A2(n6550), .ZN(n4188) );
  INVD1BWP12T U1990 ( .I(n4869), .ZN(n6253) );
  INVD1BWP12T U1991 ( .I(n6535), .ZN(n5034) );
  INVD1BWP12T U1992 ( .I(n6403), .ZN(n6538) );
  AOI22D1BWP12T U1993 ( .A1(n5662), .A2(n5034), .B1(n5661), .B2(n6538), .ZN(
        n4187) );
  ND3D1BWP12T U1994 ( .A1(n4189), .A2(n4188), .A3(n4187), .ZN(n6397) );
  NR2D1BWP12T U1995 ( .A1(n4190), .A2(n4924), .ZN(n5569) );
  INVD1BWP12T U1996 ( .I(n5569), .ZN(n5570) );
  NR2D1BWP12T U1997 ( .A1(n5570), .A2(n6357), .ZN(n6411) );
  ND2D1BWP12T U1998 ( .A1(n5570), .A2(n6565), .ZN(n6438) );
  INVD1BWP12T U1999 ( .I(n6438), .ZN(n5666) );
  AOI211D0BWP12T U2000 ( .A1(n6397), .A2(n6411), .B(n5666), .C(n6716), .ZN(
        n4198) );
  ND2D1BWP12T U2001 ( .A1(n5767), .A2(n6576), .ZN(n6304) );
  NR2D1BWP12T U2002 ( .A1(n5237), .A2(n6304), .ZN(n6268) );
  NR2D1BWP12T U2003 ( .A1(n5569), .A2(n6268), .ZN(n6436) );
  NR2D1BWP12T U2004 ( .A1(n6409), .A2(n5178), .ZN(n4193) );
  INVD3BWP12T U2005 ( .I(n5661), .ZN(n6408) );
  INR2D1BWP12T U2006 ( .A1(n5247), .B1(n4922), .ZN(n5655) );
  INVD1BWP12T U2007 ( .I(n5655), .ZN(n4895) );
  OAI22D0BWP12T U2008 ( .A1(n6408), .A2(n5176), .B1(n4895), .B2(n5179), .ZN(
        n4192) );
  INVD1BWP12T U2009 ( .I(n5660), .ZN(n6410) );
  TPNR2D0BWP12T U2010 ( .A1(n6410), .A2(n5023), .ZN(n4191) );
  NR3D1BWP12T U2011 ( .A1(n4193), .A2(n4192), .A3(n4191), .ZN(n6401) );
  INVD1BWP12T U2012 ( .I(n4894), .ZN(n5173) );
  INVD1BWP12T U2013 ( .I(n4893), .ZN(n5174) );
  INVD2BWP12T U2014 ( .I(n5662), .ZN(n6407) );
  INVD1BWP12T U2015 ( .I(n4888), .ZN(n5175) );
  INVD1BWP12T U2016 ( .I(n6263), .ZN(n5177) );
  INVD1BWP12T U2017 ( .I(n6268), .ZN(n5533) );
  ND2D1BWP12T U2018 ( .A1(n5533), .A2(n6573), .ZN(n6717) );
  AOI22D1BWP12T U2019 ( .A1(n6436), .A2(n6401), .B1(n6817), .B2(n6717), .ZN(
        n4197) );
  ND2XD4BWP12T U2020 ( .A1(n6355), .A2(n6565), .ZN(n6584) );
  CKND6BWP12T U2021 ( .I(n6584), .ZN(n6350) );
  ND2D1BWP12T U2022 ( .A1(n6350), .A2(n6909), .ZN(n5470) );
  ND2D1BWP12T U2023 ( .A1(n6840), .A2(n5470), .ZN(n5479) );
  INVD1BWP12T U2024 ( .I(a[25]), .ZN(n5047) );
  IND2D4BWP12T U2025 ( .A1(n4829), .B1(n5612), .ZN(n5239) );
  INVD1BWP12T U2026 ( .I(n5239), .ZN(n4284) );
  TPAOI22D0BWP12T U2027 ( .A1(a[25]), .A2(n4284), .B1(n4281), .B2(a[24]), .ZN(
        n4195) );
  INVD1BWP12T U2028 ( .I(n5235), .ZN(n6262) );
  AOI22D1BWP12T U2029 ( .A1(n6262), .A2(a[26]), .B1(a[23]), .B2(n6245), .ZN(
        n4194) );
  ND2D1BWP12T U2030 ( .A1(n4195), .A2(n4194), .ZN(n6255) );
  MUX2D1BWP12T U2031 ( .I0(a[29]), .I1(a[30]), .S(n6248), .Z(n5169) );
  INVD1BWP12T U2032 ( .I(n5169), .ZN(n4326) );
  OAI22D1BWP12T U2033 ( .A1(n5237), .A2(a[27]), .B1(n5238), .B2(a[28]), .ZN(
        n4196) );
  AOI21D1BWP12T U2034 ( .A1(n4498), .A2(n4326), .B(n4196), .ZN(n4925) );
  INVD1BWP12T U2035 ( .I(n4925), .ZN(n4868) );
  NR2D1BWP12T U2036 ( .A1(n5537), .A2(n6334), .ZN(n6345) );
  AOI22D1BWP12T U2037 ( .A1(n4198), .A2(n4197), .B1(n5479), .B2(n6345), .ZN(
        n4199) );
  OAI211D1BWP12T U2038 ( .A1(a[23]), .A2(n5482), .B(n4200), .C(n4199), .ZN(
        n4201) );
  AOI21D1BWP12T U2039 ( .A1(a[23]), .A2(n5070), .B(n4201), .ZN(n4202) );
  OAI211D1BWP12T U2040 ( .A1(n6794), .A2(n6210), .B(n4203), .C(n4202), .ZN(
        n4204) );
  AOI31D1BWP12T U2041 ( .A1(n6898), .A2(n6155), .A3(n6154), .B(n4204), .ZN(
        n4224) );
  INVD1BWP12T U2042 ( .I(n5463), .ZN(n6624) );
  IND2D1BWP12T U2043 ( .A1(n5360), .B1(n5612), .ZN(n6467) );
  AOI21D1BWP12T U2044 ( .A1(n4205), .A2(n6467), .B(n6498), .ZN(n5977) );
  ND2D1BWP12T U2045 ( .A1(n5977), .A2(n6180), .ZN(n5978) );
  IND2D1BWP12T U2046 ( .A1(a[2]), .B1(n5247), .ZN(n6466) );
  ND2D1BWP12T U2047 ( .A1(n5978), .A2(n6466), .ZN(n4942) );
  AOI21D1BWP12T U2048 ( .A1(n4942), .A2(n5226), .B(n6462), .ZN(n5228) );
  CKND2D1BWP12T U2049 ( .A1(n5228), .A2(n5256), .ZN(n5975) );
  INR2D0BWP12T U2050 ( .A1(n5255), .B1(n5138), .ZN(n6501) );
  AOI21D1BWP12T U2051 ( .A1(n5975), .A2(n6501), .B(n6463), .ZN(n5106) );
  AOI21D1BWP12T U2052 ( .A1(n5984), .A2(n6812), .B(n6465), .ZN(n5974) );
  OAI21D1BWP12T U2053 ( .A1(n5974), .A2(n6746), .B(n4207), .ZN(n5195) );
  AOI21D1BWP12T U2054 ( .A1(n6129), .A2(n4229), .B(n6486), .ZN(n5973) );
  AOI21D1BWP12T U2055 ( .A1(n5973), .A2(n4210), .B(n4209), .ZN(n5563) );
  INVD1BWP12T U2056 ( .I(n4211), .ZN(n6478) );
  NR2D1BWP12T U2057 ( .A1(n5563), .A2(n6478), .ZN(n5154) );
  OAI21D1BWP12T U2058 ( .A1(n5154), .A2(n5601), .B(n5183), .ZN(n5603) );
  INVD1BWP12T U2059 ( .I(n5608), .ZN(n5604) );
  ND2D1BWP12T U2060 ( .A1(n5603), .A2(n5604), .ZN(n5972) );
  ND2D1BWP12T U2061 ( .A1(n5972), .A2(n6477), .ZN(n5525) );
  INVD1BWP12T U2062 ( .I(n6495), .ZN(n4213) );
  OAI21D1BWP12T U2063 ( .A1(n5001), .A2(n4214), .B(n4213), .ZN(n5702) );
  NR2D1BWP12T U2064 ( .A1(n5702), .A2(n6502), .ZN(n5971) );
  OAI21D1BWP12T U2065 ( .A1(n5971), .A2(n4215), .B(n5925), .ZN(n5969) );
  INVD1BWP12T U2066 ( .I(n6170), .ZN(n6659) );
  AOI21D1BWP12T U2067 ( .A1(n5969), .A2(n6659), .B(n6656), .ZN(n5459) );
  INVD1BWP12T U2068 ( .I(n5460), .ZN(n6614) );
  CKND0BWP12T U2069 ( .I(n5462), .ZN(n4218) );
  INVD1BWP12T U2070 ( .I(n4219), .ZN(n6496) );
  OAI21D1BWP12T U2071 ( .A1(n5462), .A2(n6496), .B(n4217), .ZN(n4791) );
  INVD1BWP12T U2072 ( .I(n4791), .ZN(n5096) );
  AOI31D1BWP12T U2073 ( .A1(n4220), .A2(n4219), .A3(n4218), .B(n5096), .ZN(
        n5994) );
  NR2D1BWP12T U2074 ( .A1(n4222), .A2(n4221), .ZN(n6728) );
  INVD1BWP12T U2075 ( .I(n6728), .ZN(n6890) );
  ND2D1BWP12T U2076 ( .A1(n5994), .A2(n6728), .ZN(n4223) );
  OAI211D2BWP12T U2077 ( .A1(n6902), .A2(n4225), .B(n4224), .C(n4223), .ZN(
        result[23]) );
  INVD1BWP12T U2078 ( .I(n4226), .ZN(n6013) );
  INVD1BWP12T U2079 ( .I(n6012), .ZN(n4227) );
  ND2D1BWP12T U2080 ( .A1(n4227), .A2(n6011), .ZN(n4228) );
  XOR2XD2BWP12T U2081 ( .A1(n6013), .A2(n4228), .Z(n6043) );
  INVD1BWP12T U2082 ( .I(n4233), .ZN(n4237) );
  XOR2XD1BWP12T U2083 ( .A1(n4229), .A2(n4237), .Z(n5986) );
  XOR2XD1BWP12T U2084 ( .A1(n4230), .A2(n4237), .Z(n6142) );
  INVD1BWP12T U2085 ( .I(n6898), .ZN(n6836) );
  CKND2D1BWP12T U2086 ( .A1(n4232), .A2(n4231), .ZN(n5203) );
  CKND2D1BWP12T U2087 ( .A1(n5203), .A2(n5204), .ZN(n5202) );
  INVD1BWP12T U2088 ( .I(n6173), .ZN(n5198) );
  INVD1BWP12T U2089 ( .I(n6093), .ZN(n6748) );
  NR2D1BWP12T U2090 ( .A1(n5200), .A2(n6748), .ZN(n4234) );
  ND2D1BWP12T U2091 ( .A1(n5198), .A2(n4234), .ZN(n4236) );
  INVD1BWP12T U2092 ( .I(n4236), .ZN(n5199) );
  TPOAI21D0BWP12T U2093 ( .A1(n5199), .A2(n4238), .B(n4237), .ZN(n4239) );
  ND2D1BWP12T U2094 ( .A1(n6198), .A2(n4239), .ZN(n6193) );
  NR2D1BWP12T U2095 ( .A1(n6264), .A2(n4823), .ZN(n5229) );
  MUX2ND0BWP12T U2096 ( .I0(a[16]), .I1(n6232), .S(n4823), .ZN(n5673) );
  INVD1BWP12T U2097 ( .I(n5673), .ZN(n4985) );
  NR2D1BWP12T U2098 ( .A1(n6264), .A2(n4305), .ZN(n5230) );
  INVD1BWP12T U2099 ( .I(n6252), .ZN(n5620) );
  NR2D1BWP12T U2100 ( .A1(n5767), .A2(n6334), .ZN(n6313) );
  OAI22D1BWP12T U2101 ( .A1(n5237), .A2(n5232), .B1(n4286), .B2(n5235), .ZN(
        n4241) );
  INVD1BWP12T U2102 ( .I(n6231), .ZN(n5589) );
  OAI22D1BWP12T U2103 ( .A1(n5589), .A2(n5239), .B1(n5238), .B2(n6708), .ZN(
        n4240) );
  NR2D1BWP12T U2104 ( .A1(n4241), .A2(n4240), .ZN(n6251) );
  INVD0BWP12T U2105 ( .I(n6251), .ZN(n4242) );
  INVD1BWP12T U2106 ( .I(n6304), .ZN(n5575) );
  TPAOI21D0BWP12T U2107 ( .A1(n4242), .A2(n5575), .B(n6573), .ZN(n4243) );
  OAI21D1BWP12T U2108 ( .A1(n5620), .A2(n6297), .B(n4243), .ZN(n6324) );
  OAI22D1BWP12T U2109 ( .A1(n5237), .A2(n5487), .B1(n5047), .B2(n5235), .ZN(
        n4245) );
  INVD1BWP12T U2110 ( .I(a[24]), .ZN(n5016) );
  NR2D1BWP12T U2111 ( .A1(n4245), .A2(n4244), .ZN(n5614) );
  OAI22D1BWP12T U2112 ( .A1(n5237), .A2(n6646), .B1(n6623), .B2(n5235), .ZN(
        n4247) );
  NR2D1BWP12T U2113 ( .A1(n4247), .A2(n4246), .ZN(n5613) );
  MUX2NXD0BWP12T U2114 ( .I0(n5614), .I1(n5613), .S(n5767), .ZN(n6325) );
  INVD1BWP12T U2115 ( .I(n6325), .ZN(n6331) );
  INVD1BWP12T U2116 ( .I(n6376), .ZN(n4268) );
  INVD0BWP12T U2117 ( .I(n4248), .ZN(n6676) );
  OAI22D1BWP12T U2118 ( .A1(n5237), .A2(a[26]), .B1(a[29]), .B2(n5235), .ZN(
        n4250) );
  OAI22D1BWP12T U2119 ( .A1(a[27]), .A2(n5238), .B1(n5239), .B2(a[28]), .ZN(
        n4249) );
  NR2D1BWP12T U2120 ( .A1(n4250), .A2(n4249), .ZN(n5615) );
  MUX2NXD0BWP12T U2121 ( .I0(a[30]), .I1(a[31]), .S(n4829), .ZN(n4251) );
  NR2D1BWP12T U2122 ( .A1(n4251), .A2(n4498), .ZN(n5118) );
  MUX2D1BWP12T U2123 ( .I0(n5615), .I1(n5118), .S(n6520), .Z(n6321) );
  ND2D1BWP12T U2124 ( .A1(n6321), .A2(n6576), .ZN(n6289) );
  INVD1BWP12T U2125 ( .I(n6840), .ZN(n6736) );
  CKND1BWP12T U2126 ( .I(n4252), .ZN(n4253) );
  NR2D1BWP12T U2127 ( .A1(n4253), .A2(n6862), .ZN(n5216) );
  NR2XD0BWP12T U2128 ( .A1(n5216), .A2(n6783), .ZN(n5217) );
  ND2D1BWP12T U2129 ( .A1(n4253), .A2(n6786), .ZN(n6713) );
  MUX2ND0BWP12T U2130 ( .I0(n5217), .I1(n6713), .S(n6715), .ZN(n4266) );
  ND2D1BWP12T U2131 ( .A1(n6411), .A2(n6857), .ZN(n6892) );
  MUX2ND0BWP12T U2132 ( .I0(a[6]), .I1(n6267), .S(n4823), .ZN(n5297) );
  ND2XD0BWP12T U2133 ( .A1(n5289), .A2(n5297), .ZN(n4256) );
  MUX2ND0BWP12T U2134 ( .I0(n6715), .I1(n6229), .S(n4829), .ZN(n5298) );
  CKND2D0BWP12T U2135 ( .A1(n5660), .A2(n5298), .ZN(n4255) );
  MUX2ND0BWP12T U2136 ( .I0(a[8]), .I1(n6819), .S(n4829), .ZN(n5299) );
  MUX2ND0BWP12T U2137 ( .I0(n6249), .I1(n6247), .S(n4829), .ZN(n5250) );
  AOI22D1BWP12T U2138 ( .A1(n5662), .A2(n5299), .B1(n5661), .B2(n5250), .ZN(
        n4254) );
  ND3D1BWP12T U2139 ( .A1(n4256), .A2(n4255), .A3(n4254), .ZN(n6391) );
  ND2XD3BWP12T U2140 ( .A1(n6350), .A2(n6855), .ZN(n6739) );
  AOI22D1BWP12T U2141 ( .A1(n6553), .A2(n5298), .B1(n5250), .B2(n6549), .ZN(
        n4258) );
  AOI22D0BWP12T U2142 ( .A1(n6556), .A2(n5297), .B1(n5299), .B2(n6552), .ZN(
        n4257) );
  ND2D1BWP12T U2143 ( .A1(n4258), .A2(n4257), .ZN(n6524) );
  MUX2XD0BWP12T U2144 ( .I0(a[2]), .I1(n5360), .S(n6248), .Z(n5249) );
  INVD1BWP12T U2145 ( .I(n5249), .ZN(n5252) );
  MUX2D1BWP12T U2146 ( .I0(n5072), .I1(n5252), .S(n3463), .Z(n6521) );
  NR2D1BWP12T U2147 ( .A1(n4924), .A2(n6520), .ZN(n6278) );
  INVD1BWP12T U2148 ( .I(n6278), .ZN(n6308) );
  OAI22D1BWP12T U2149 ( .A1(n6524), .A2(n6334), .B1(n6521), .B2(n6308), .ZN(
        n5688) );
  ND2D1BWP12T U2150 ( .A1(n5578), .A2(n5688), .ZN(n4264) );
  INVD1BWP12T U2151 ( .I(n6436), .ZN(n6419) );
  INR2D1BWP12T U2152 ( .A1(n6573), .B1(n6419), .ZN(n5659) );
  ND2D1BWP12T U2153 ( .A1(n5659), .A2(n6857), .ZN(n5719) );
  AOI22D1BWP12T U2154 ( .A1(n5660), .A2(n5249), .B1(n6488), .B2(n6549), .ZN(
        n6893) );
  INVD0BWP12T U2155 ( .I(n6893), .ZN(n6383) );
  INVD1BWP12T U2156 ( .I(n6745), .ZN(n6882) );
  OAI22D0BWP12T U2157 ( .A1(n4260), .A2(n6882), .B1(n4259), .B2(n6874), .ZN(
        n4262) );
  OAI22D0BWP12T U2158 ( .A1(n6129), .A2(n6813), .B1(n6197), .B2(n6880), .ZN(
        n4261) );
  AOI211D1BWP12T U2159 ( .A1(n5546), .A2(n6383), .B(n4262), .C(n4261), .ZN(
        n4263) );
  OAI211D1BWP12T U2160 ( .A1(n6892), .A2(n6391), .B(n4264), .C(n4263), .ZN(
        n4265) );
  NR2D1BWP12T U2161 ( .A1(n5767), .A2(a[31]), .ZN(n5766) );
  NR2D1BWP12T U2162 ( .A1(n6556), .A2(n5766), .ZN(n4267) );
  OAI22D1BWP12T U2163 ( .A1(n5118), .A2(n4267), .B1(n5615), .B2(n6520), .ZN(
        n6332) );
  INVD1BWP12T U2164 ( .I(n5668), .ZN(n4269) );
  INVD1BWP12T U2165 ( .I(n6364), .ZN(n5172) );
  OAI211D1BWP12T U2166 ( .A1(n4269), .A2(n5172), .B(n4268), .C(n6355), .ZN(
        n4270) );
  INVD1BWP12T U2167 ( .I(n6355), .ZN(n6560) );
  CKND2D2BWP12T U2168 ( .A1(n6560), .A2(a[31]), .ZN(n6336) );
  ND2D1BWP12T U2169 ( .A1(n4270), .A2(n6336), .ZN(n6367) );
  OAI21D1BWP12T U2170 ( .A1(n6142), .A2(n6836), .B(n4271), .ZN(n4272) );
  AOI21D1BWP12T U2171 ( .A1(n6728), .A2(n5986), .B(n4272), .ZN(n4273) );
  CKND1BWP12T U2172 ( .I(a[28]), .ZN(n5310) );
  OAI22D1BWP12T U2173 ( .A1(n5237), .A2(n5047), .B1(n5310), .B2(n5235), .ZN(
        n4275) );
  INVD1BWP12T U2174 ( .I(a[27]), .ZN(n4907) );
  CKND1BWP12T U2175 ( .I(a[26]), .ZN(n4583) );
  TPOAI22D0BWP12T U2176 ( .A1(n4907), .A2(n5239), .B1(n5238), .B2(n4583), .ZN(
        n4274) );
  NR2D1BWP12T U2177 ( .A1(n4275), .A2(n4274), .ZN(n6274) );
  INVD1BWP12T U2178 ( .I(n6274), .ZN(n4327) );
  INR2D1BWP12T U2179 ( .A1(n5767), .B1(n4327), .ZN(n5018) );
  NR2XD0BWP12T U2180 ( .A1(n5018), .A2(n4924), .ZN(n4285) );
  OAI22D1BWP12T U2181 ( .A1(n5237), .A2(n6623), .B1(n5238), .B2(n5487), .ZN(
        n4277) );
  OAI22D1BWP12T U2182 ( .A1(n5239), .A2(n5069), .B1(n5016), .B2(n5235), .ZN(
        n4276) );
  NR2D1BWP12T U2183 ( .A1(n4277), .A2(n4276), .ZN(n6275) );
  NR2D1BWP12T U2184 ( .A1(n5239), .A2(a[19]), .ZN(n4279) );
  NR2D1BWP12T U2185 ( .A1(n5235), .A2(a[20]), .ZN(n4278) );
  NR2D1BWP12T U2186 ( .A1(n4279), .A2(n4278), .ZN(n4283) );
  NR2D1BWP12T U2187 ( .A1(a[17]), .A2(n4498), .ZN(n4280) );
  OAI21D1BWP12T U2188 ( .A1(n4281), .A2(n4280), .B(n4921), .ZN(n4282) );
  ND2D1BWP12T U2189 ( .A1(n4283), .A2(n4282), .ZN(n6270) );
  OAI22D1BWP12T U2190 ( .A1(n6275), .A2(n6297), .B1(n6270), .B2(n6304), .ZN(
        n4328) );
  ND2D1BWP12T U2191 ( .A1(n6520), .A2(n6334), .ZN(n6306) );
  OAI22D1BWP12T U2192 ( .A1(n4285), .A2(n4328), .B1(n6306), .B2(n6323), .ZN(
        n6317) );
  INVD1BWP12T U2193 ( .I(n6306), .ZN(n6254) );
  CKND0BWP12T U2194 ( .I(a[14]), .ZN(n5626) );
  OAI22D1BWP12T U2195 ( .A1(n5237), .A2(n4286), .B1(n5238), .B2(n5626), .ZN(
        n4288) );
  OAI22D1BWP12T U2196 ( .A1(n4920), .A2(n3463), .B1(n4967), .B2(n5235), .ZN(
        n4287) );
  NR2D1BWP12T U2197 ( .A1(n4288), .A2(n4287), .ZN(n6266) );
  INVD1BWP12T U2198 ( .I(n6266), .ZN(n4289) );
  TPAOI22D0BWP12T U2199 ( .A1(n6273), .A2(n6278), .B1(n6254), .B2(n4289), .ZN(
        n4298) );
  NR2D1BWP12T U2200 ( .A1(n4895), .A2(n5177), .ZN(n4296) );
  NR2D1BWP12T U2201 ( .A1(n6530), .A2(n6760), .ZN(n4291) );
  NR2XD0BWP12T U2202 ( .A1(n6534), .A2(n4307), .ZN(n4290) );
  MUX2D1BWP12T U2203 ( .I0(n4291), .I1(n4290), .S(n4305), .Z(n4295) );
  ND3D0BWP12T U2204 ( .A1(n6245), .A2(n5247), .A3(n6267), .ZN(n4293) );
  INR2D1BWP12T U2205 ( .A1(n6248), .B1(n6533), .ZN(n5731) );
  ND2D1BWP12T U2206 ( .A1(n5731), .A2(n6249), .ZN(n4292) );
  OAI211D1BWP12T U2207 ( .A1(n5173), .A2(n6408), .B(n4293), .C(n4292), .ZN(
        n4294) );
  TPOAI31D0BWP12T U2208 ( .A1(n4296), .A2(n4295), .A3(n4294), .B(n6578), .ZN(
        n4297) );
  OAI21D1BWP12T U2209 ( .A1(n4298), .A2(n6573), .B(n4297), .ZN(n4329) );
  INVD1BWP12T U2210 ( .I(n6905), .ZN(n6807) );
  ND2D1BWP12T U2211 ( .A1(n4893), .A2(n6553), .ZN(n6518) );
  TPND2D2BWP12T U2212 ( .A1(n5578), .A2(n6576), .ZN(n6822) );
  ND2D1BWP12T U2213 ( .A1(n5660), .A2(n4893), .ZN(n6380) );
  INVD0BWP12T U2214 ( .I(n6380), .ZN(n4318) );
  INVD1BWP12T U2215 ( .I(n6892), .ZN(n5507) );
  CKXOR2D1BWP12T U2216 ( .A1(n4304), .A2(n6457), .Z(n5980) );
  CKND0BWP12T U2217 ( .I(n4299), .ZN(n4302) );
  INVD0BWP12T U2218 ( .I(n4300), .ZN(n4301) );
  TPAOI31D0BWP12T U2219 ( .A1(n4303), .A2(n5072), .A3(n4302), .B(n4301), .ZN(
        n6137) );
  MOAI22D0BWP12T U2220 ( .A1(n5980), .A2(n6890), .B1(n6137), .B2(n6898), .ZN(
        n4317) );
  INVD1BWP12T U2221 ( .I(n6833), .ZN(n6894) );
  CKND2D1BWP12T U2222 ( .A1(n4304), .A2(n6121), .ZN(n4319) );
  TPND2D0BWP12T U2223 ( .A1(n4320), .A2(n4319), .ZN(n5932) );
  NR2D0BWP12T U2224 ( .A1(n6488), .A2(n4646), .ZN(n4306) );
  INVD1BWP12T U2225 ( .I(n6902), .ZN(n6834) );
  CKND2D0BWP12T U2226 ( .A1(n6036), .A2(n6834), .ZN(n4315) );
  TPOAI21D0BWP12T U2227 ( .A1(n5762), .A2(n6862), .B(n6844), .ZN(n6886) );
  NR2D1BWP12T U2228 ( .A1(a[0]), .A2(n6862), .ZN(n4934) );
  INVD0BWP12T U2229 ( .I(n4934), .ZN(n4308) );
  ND2D1BWP12T U2230 ( .A1(n4308), .A2(n5360), .ZN(n4313) );
  OAI22D0BWP12T U2231 ( .A1(n4310), .A2(n6882), .B1(n4309), .B2(n6874), .ZN(
        n4312) );
  OAI22D0BWP12T U2232 ( .A1(n6467), .A2(n6813), .B1(n6098), .B2(n6880), .ZN(
        n4311) );
  AOI211D1BWP12T U2233 ( .A1(n6886), .A2(n4313), .B(n4312), .C(n4311), .ZN(
        n4314) );
  OAI211D1BWP12T U2234 ( .A1(n6894), .A2(n5932), .B(n4315), .C(n4314), .ZN(
        n4316) );
  AOI211D1BWP12T U2235 ( .A1(n4318), .A2(n5507), .B(n4317), .C(n4316), .ZN(
        n4325) );
  INVD1BWP12T U2236 ( .I(n6794), .ZN(n6870) );
  INVD1BWP12T U2237 ( .I(n4319), .ZN(n4323) );
  CKND0BWP12T U2238 ( .I(n4320), .ZN(n4321) );
  AOI211XD0BWP12T U2239 ( .A1(n4323), .A2(n5735), .B(n4322), .C(n4321), .ZN(
        n6182) );
  INR2D2BWP12T U2240 ( .A1(n6909), .B1(n6336), .ZN(n6753) );
  AOI21D1BWP12T U2241 ( .A1(n6870), .A2(n6182), .B(n6753), .ZN(n4324) );
  AOI21D1BWP12T U2242 ( .A1(n6573), .A2(n6341), .B(n4329), .ZN(n4330) );
  NR2D1BWP12T U2243 ( .A1(n4330), .A2(n6560), .ZN(n6348) );
  CKND2D1BWP12T U2244 ( .A1(n6348), .A2(n6909), .ZN(n4331) );
  OAI211D1BWP12T U2245 ( .A1(n6283), .A2(n6807), .B(n4332), .C(n4331), .ZN(
        result[1]) );
  NR2D1BWP12T U2246 ( .A1(a[23]), .A2(b[23]), .ZN(n4796) );
  OA21D1BWP12T U2247 ( .A1(n4333), .A2(n4796), .B(n6107), .Z(n5067) );
  CKND2D1BWP12T U2248 ( .A1(a[24]), .A2(b[24]), .ZN(n6101) );
  NR2D1BWP12T U2249 ( .A1(a[24]), .A2(b[24]), .ZN(n4798) );
  AO21D1BWP12T U2250 ( .A1(n5067), .A2(n6101), .B(n4798), .Z(n5013) );
  NR2D1BWP12T U2251 ( .A1(a[25]), .A2(b[25]), .ZN(n4799) );
  CKND2D1BWP12T U2252 ( .A1(a[25]), .A2(b[25]), .ZN(n6104) );
  OA21D1BWP12T U2253 ( .A1(n5013), .A2(n4799), .B(n6104), .Z(n5650) );
  CKND2D1BWP12T U2254 ( .A1(a[26]), .A2(b[26]), .ZN(n6116) );
  NR2D1BWP12T U2255 ( .A1(a[26]), .A2(b[26]), .ZN(n4800) );
  AO21D1BWP12T U2256 ( .A1(n5650), .A2(n6116), .B(n4800), .Z(n4865) );
  NR2D1BWP12T U2257 ( .A1(a[27]), .A2(b[27]), .ZN(n4801) );
  CKND2D1BWP12T U2258 ( .A1(a[27]), .A2(b[27]), .ZN(n4802) );
  OA21D1BWP12T U2259 ( .A1(n4865), .A2(n4801), .B(n4802), .Z(n5280) );
  CKND2D1BWP12T U2260 ( .A1(a[28]), .A2(b[28]), .ZN(n6113) );
  NR2D1BWP12T U2261 ( .A1(a[28]), .A2(b[28]), .ZN(n5311) );
  AOI21D1BWP12T U2262 ( .A1(n5280), .A2(n6113), .B(n5311), .ZN(n5922) );
  CKND2D1BWP12T U2263 ( .A1(a[29]), .A2(b[29]), .ZN(n6843) );
  NR2D1BWP12T U2264 ( .A1(a[29]), .A2(b[29]), .ZN(n6842) );
  NR2D1BWP12T U2265 ( .A1(a[30]), .A2(b[30]), .ZN(n5910) );
  INVD1BWP12T U2266 ( .I(n5910), .ZN(n5417) );
  ND2D1BWP12T U2267 ( .A1(a[30]), .A2(b[30]), .ZN(n5416) );
  ND2D1BWP12T U2268 ( .A1(n5417), .A2(n5416), .ZN(n4804) );
  MUX2ND0BWP12T U2269 ( .I0(n4747), .I1(n4746), .S(b[21]), .ZN(n4335) );
  MUX2ND0BWP12T U2270 ( .I0(n5860), .I1(n5861), .S(n4494), .ZN(n4334) );
  NR2D1BWP12T U2271 ( .A1(n4335), .A2(n4334), .ZN(n4389) );
  TPND2D0BWP12T U2272 ( .A1(n5069), .A2(n5016), .ZN(n4810) );
  CKND2D0BWP12T U2273 ( .A1(n4810), .A2(n4823), .ZN(n4336) );
  OAI211D1BWP12T U2274 ( .A1(n5016), .A2(n5069), .B(n4336), .C(a[25]), .ZN(
        n4388) );
  MUX2ND0BWP12T U2275 ( .I0(n5871), .I1(n5872), .S(n5405), .ZN(n4337) );
  NR2D1BWP12T U2276 ( .A1(n4338), .A2(n4337), .ZN(n4387) );
  MUX2ND0BWP12T U2277 ( .I0(n5871), .I1(n5872), .S(n4745), .ZN(n4339) );
  NR2D1BWP12T U2278 ( .A1(n4340), .A2(n4339), .ZN(n4517) );
  MUX2ND0BWP12T U2279 ( .I0(n4747), .I1(n4746), .S(b[22]), .ZN(n4342) );
  MUX2ND0BWP12T U2280 ( .I0(n5860), .I1(n5861), .S(n4758), .ZN(n4341) );
  NR2D1BWP12T U2281 ( .A1(n4342), .A2(n4341), .ZN(n4493) );
  MUX2ND0BWP12T U2282 ( .I0(n5406), .I1(n5407), .S(n4343), .ZN(n4344) );
  NR2D1BWP12T U2283 ( .A1(n4345), .A2(n4344), .ZN(n4492) );
  CKND2D0BWP12T U2284 ( .A1(n5069), .A2(n5487), .ZN(n4346) );
  ND2D1BWP12T U2285 ( .A1(n4347), .A2(n4346), .ZN(n4744) );
  INVD1BWP12T U2286 ( .I(n4744), .ZN(n5809) );
  XOR2D1BWP12T U2287 ( .A1(a[23]), .A2(n6334), .Z(n4348) );
  XOR2D1BWP12T U2288 ( .A1(a[23]), .A2(n6573), .Z(n4486) );
  AOI22D1BWP12T U2289 ( .A1(n5809), .A2(n4348), .B1(n5807), .B2(n4486), .ZN(
        n4491) );
  XNR2D1BWP12T U2290 ( .A1(a[23]), .A2(n6520), .ZN(n4385) );
  MUX2ND0BWP12T U2291 ( .I0(n5778), .I1(n5777), .S(b[14]), .ZN(n4349) );
  NR2D1BWP12T U2292 ( .A1(n4350), .A2(n4349), .ZN(n4440) );
  MUX2ND0BWP12T U2293 ( .I0(n5811), .I1(n5810), .S(b[23]), .ZN(n4352) );
  NR2D1BWP12T U2294 ( .A1(n4352), .A2(n4351), .ZN(n4439) );
  MUX2ND0BWP12T U2295 ( .I0(n5878), .I1(n5877), .S(b[17]), .ZN(n4353) );
  NR2D1BWP12T U2296 ( .A1(n4354), .A2(n4353), .ZN(n4450) );
  AOI21D1BWP12T U2297 ( .A1(n6707), .A2(n4375), .B(n4355), .ZN(n4449) );
  XNR2D1BWP12T U2298 ( .A1(a[17]), .A2(n5843), .ZN(n4395) );
  IAO21D1BWP12T U2299 ( .A1(n4395), .A2(n4394), .B(n4356), .ZN(n4448) );
  MUX2ND0BWP12T U2300 ( .I0(n5406), .I1(n5407), .S(n4357), .ZN(n4358) );
  NR2D1BWP12T U2301 ( .A1(n4359), .A2(n4358), .ZN(n4438) );
  MUX2ND0BWP12T U2302 ( .I0(n5803), .I1(n5802), .S(n6782), .ZN(n4361) );
  MUX2ND0BWP12T U2303 ( .I0(n5804), .I1(n5805), .S(n6565), .ZN(n4360) );
  NR2D1BWP12T U2304 ( .A1(n4361), .A2(n4360), .ZN(n4437) );
  TPAOI21D0BWP12T U2305 ( .A1(n4557), .A2(n4363), .B(n4362), .ZN(n4411) );
  XOR2D1BWP12T U2306 ( .A1(a[23]), .A2(a[24]), .Z(n5845) );
  ND2D1BWP12T U2307 ( .A1(n5845), .A2(n4823), .ZN(n4410) );
  MUX2ND0BWP12T U2308 ( .I0(n5813), .I1(n5812), .S(b[21]), .ZN(n4364) );
  NR2D1BWP12T U2309 ( .A1(n4365), .A2(n4364), .ZN(n4409) );
  MUX2ND0BWP12T U2310 ( .I0(n5878), .I1(n5877), .S(b[19]), .ZN(n4366) );
  NR2D1BWP12T U2311 ( .A1(n4367), .A2(n4366), .ZN(n4507) );
  XNR2D1BWP12T U2312 ( .A1(a[25]), .A2(a[24]), .ZN(n4368) );
  NR2D1BWP12T U2313 ( .A1(n4368), .A2(n5845), .ZN(n5847) );
  INVD1BWP12T U2314 ( .I(n5847), .ZN(n5382) );
  MUX2ND0BWP12T U2315 ( .I0(a[25]), .I1(a[24]), .S(n4829), .ZN(n6555) );
  INVD1BWP12T U2316 ( .I(n5845), .ZN(n5380) );
  XNR2D1BWP12T U2317 ( .A1(a[25]), .A2(n4498), .ZN(n4432) );
  OAI22D1BWP12T U2318 ( .A1(n5382), .A2(n6555), .B1(n5380), .B2(n4432), .ZN(
        n4402) );
  MUX2ND0BWP12T U2319 ( .I0(n4759), .I1(n4760), .S(b[16]), .ZN(n4373) );
  ND2D1BWP12T U2320 ( .A1(n4374), .A2(n4373), .ZN(n4401) );
  MAOI222D1BWP12T U2321 ( .A(n4402), .B(n4400), .C(n4401), .ZN(n4505) );
  MUX2D1BWP12T U2322 ( .I0(n5817), .I1(n5816), .S(b[14]), .Z(n4377) );
  ND2XD0BWP12T U2323 ( .A1(n4375), .A2(n5151), .ZN(n4376) );
  ND2D1BWP12T U2324 ( .A1(n4377), .A2(n4376), .ZN(n4512) );
  MUX2NXD1BWP12T U2325 ( .I0(n4757), .I1(n4756), .S(b[18]), .ZN(n4379) );
  MUX2NXD0BWP12T U2326 ( .I0(n4759), .I1(n4760), .S(b[17]), .ZN(n4378) );
  ND2D1BWP12T U2327 ( .A1(n4379), .A2(n4378), .ZN(n4511) );
  CKND2D0BWP12T U2328 ( .A1(n5728), .A2(n4967), .ZN(n4380) );
  ND2D1BWP12T U2329 ( .A1(n4381), .A2(n4380), .ZN(n4396) );
  XNR2D1BWP12T U2330 ( .A1(a[17]), .A2(b[9]), .ZN(n4393) );
  MUX2D1BWP12T U2331 ( .I0(n5761), .I1(n5760), .S(n5806), .Z(n4382) );
  OAI21D1BWP12T U2332 ( .A1(n4396), .A2(n4393), .B(n4382), .ZN(n4510) );
  XNR3D1BWP12T U2333 ( .A1(n4512), .A2(n4511), .A3(n4510), .ZN(n4506) );
  XOR3D1BWP12T U2334 ( .A1(n4507), .A2(n4505), .A3(n4506), .Z(n4501) );
  MUX2D1BWP12T U2335 ( .I0(n4747), .I1(n4746), .S(b[20]), .Z(n4384) );
  MUX2D1BWP12T U2336 ( .I0(n5861), .I1(n5860), .S(b[19]), .Z(n4383) );
  ND2D1BWP12T U2337 ( .A1(n4384), .A2(n4383), .ZN(n4418) );
  OAI22D1BWP12T U2338 ( .A1(n4744), .A2(n4386), .B1(n4742), .B2(n4385), .ZN(
        n4420) );
  MAOI222D1BWP12T U2339 ( .A(n4419), .B(n4418), .C(n4420), .ZN(n4428) );
  INVD1BWP12T U2340 ( .I(n4428), .ZN(n4392) );
  FA1D0BWP12T U2341 ( .A(n4389), .B(n4388), .CI(n4387), .CO(n4518), .S(n4427)
         );
  INVD1BWP12T U2342 ( .I(n4427), .ZN(n4391) );
  MAOI222D1BWP12T U2343 ( .A(n4392), .B(n4391), .C(n4429), .ZN(n4500) );
  OAI22D1BWP12T U2344 ( .A1(n4396), .A2(n4395), .B1(n4394), .B2(n4393), .ZN(
        n4399) );
  MUX2ND0BWP12T U2345 ( .I0(n4647), .I1(n4646), .S(b[25]), .ZN(n4397) );
  OAI21D0BWP12T U2346 ( .A1(b[24]), .A2(n5361), .B(n4397), .ZN(n4398) );
  ND2D1BWP12T U2347 ( .A1(n4398), .A2(n4399), .ZN(n4476) );
  OAI21D1BWP12T U2348 ( .A1(n4399), .A2(n4398), .B(n4476), .ZN(n4444) );
  XNR3D1BWP12T U2349 ( .A1(n4402), .A2(n4401), .A3(n4400), .ZN(n4443) );
  MUX2ND0BWP12T U2350 ( .I0(n5776), .I1(n5775), .S(b[14]), .ZN(n4404) );
  MUX2ND0BWP12T U2351 ( .I0(n5778), .I1(n5777), .S(b[13]), .ZN(n4403) );
  NR2D1BWP12T U2352 ( .A1(n4404), .A2(n4403), .ZN(n4417) );
  MUX2ND0BWP12T U2353 ( .I0(n5406), .I1(n5407), .S(n4433), .ZN(n4405) );
  NR2D1BWP12T U2354 ( .A1(n4406), .A2(n4405), .ZN(n4416) );
  MUX2NXD0BWP12T U2355 ( .I0(n5803), .I1(n5802), .S(n6573), .ZN(n4408) );
  NR2D1BWP12T U2356 ( .A1(n4408), .A2(n4407), .ZN(n4415) );
  FA1D0BWP12T U2357 ( .A(n4411), .B(n4410), .CI(n4409), .CO(n4436), .S(n4532)
         );
  FA1D0BWP12T U2358 ( .A(n4414), .B(n4413), .CI(n4412), .CO(n4531), .S(n4536)
         );
  FA1D0BWP12T U2359 ( .A(n4417), .B(n4416), .CI(n4415), .CO(n4442), .S(n4530)
         );
  XOR3D1BWP12T U2360 ( .A1(n4420), .A2(n4419), .A3(n4418), .Z(n4541) );
  MUX2ND0BWP12T U2361 ( .I0(n4759), .I1(n4760), .S(b[15]), .ZN(n4421) );
  ND2D1BWP12T U2362 ( .A1(n4422), .A2(n4421), .ZN(n4542) );
  INVD1BWP12T U2363 ( .I(n4423), .ZN(n4425) );
  MAOI222D1BWP12T U2364 ( .A(n4426), .B(n4425), .C(n4424), .ZN(n4540) );
  MAOI222D1BWP12T U2365 ( .A(n4541), .B(n4542), .C(n4540), .ZN(n4465) );
  XNR3D1BWP12T U2366 ( .A1(n4429), .A2(n4428), .A3(n4427), .ZN(n4464) );
  MUX2ND0BWP12T U2367 ( .I0(n5776), .I1(n5775), .S(b[16]), .ZN(n4431) );
  MUX2ND0BWP12T U2368 ( .I0(n5778), .I1(n5777), .S(b[15]), .ZN(n4430) );
  NR2D1BWP12T U2369 ( .A1(n4431), .A2(n4430), .ZN(n4483) );
  XOR2D1BWP12T U2370 ( .A1(a[25]), .A2(n6520), .Z(n4480) );
  MUX2NXD0BWP12T U2371 ( .I0(n5803), .I1(n5802), .S(n5864), .ZN(n4435) );
  MUX2ND0BWP12T U2372 ( .I0(n5804), .I1(n5805), .S(n4433), .ZN(n4434) );
  NR2D1BWP12T U2373 ( .A1(n4435), .A2(n4434), .ZN(n4481) );
  FA1D0BWP12T U2374 ( .A(n4438), .B(n4437), .CI(n4436), .CO(n4503), .S(n4461)
         );
  FA1D0BWP12T U2375 ( .A(n4441), .B(n4440), .CI(n4439), .CO(n4477), .S(n4463)
         );
  CKXOR2D1BWP12T U2376 ( .A1(a[26]), .A2(a[25]), .Z(n5866) );
  FA1D0BWP12T U2377 ( .A(n4444), .B(n4443), .CI(n4442), .CO(n4499), .S(n4548)
         );
  FA1D0BWP12T U2378 ( .A(n4447), .B(n4446), .CI(n4445), .CO(n4460), .S(n4451)
         );
  FA1D0BWP12T U2379 ( .A(n4450), .B(n4449), .CI(n4448), .CO(n4462), .S(n4458)
         );
  FA1D0BWP12T U2380 ( .A(n4453), .B(n4452), .CI(n4451), .CO(n4535), .S(n4679)
         );
  INVD1BWP12T U2381 ( .I(n4454), .ZN(n4457) );
  MAOI222D1BWP12T U2382 ( .A(n4457), .B(n4456), .C(n4455), .ZN(n4534) );
  FA1D0BWP12T U2383 ( .A(n4460), .B(n4459), .CI(n4458), .CO(n4547), .S(n4533)
         );
  FA1D0BWP12T U2384 ( .A(n4463), .B(n4462), .CI(n4461), .CO(n4473), .S(n4470)
         );
  FA1D0BWP12T U2385 ( .A(n4466), .B(n4465), .CI(n4464), .CO(n4522), .S(n4469)
         );
  NR2D1BWP12T U2386 ( .A1(n4468), .A2(n4467), .ZN(n4524) );
  ND2D1BWP12T U2387 ( .A1(n4468), .A2(n4467), .ZN(n4525) );
  FA1D0BWP12T U2388 ( .A(n4471), .B(n4470), .CI(n4469), .CO(n4526), .S(n4546)
         );
  FA1D0BWP12T U2389 ( .A(n4474), .B(n4473), .CI(n4472), .CO(n4520), .S(n4468)
         );
  FA1D0BWP12T U2390 ( .A(n4477), .B(n4476), .CI(n4475), .CO(n4556), .S(n4502)
         );
  MUX2ND0BWP12T U2391 ( .I0(n5776), .I1(n5775), .S(b[17]), .ZN(n4479) );
  MUX2ND0BWP12T U2392 ( .I0(n5778), .I1(n5777), .S(b[16]), .ZN(n4478) );
  NR2D1BWP12T U2393 ( .A1(n4479), .A2(n4478), .ZN(n4562) );
  XOR2D1BWP12T U2394 ( .A1(a[25]), .A2(n6334), .Z(n4586) );
  AOI22D1BWP12T U2395 ( .A1(n5847), .A2(n4480), .B1(n5845), .B2(n4586), .ZN(
        n4561) );
  FA1D0BWP12T U2396 ( .A(n4483), .B(n4482), .CI(n4481), .CO(n4599), .S(n4504)
         );
  INVD1BWP12T U2397 ( .I(b[27]), .ZN(n4882) );
  NR2D1BWP12T U2398 ( .A1(n4485), .A2(n4484), .ZN(n4662) );
  AO21D1BWP12T U2399 ( .A1(n4485), .A2(n4484), .B(n4662), .Z(n4598) );
  XOR2D1BWP12T U2400 ( .A1(a[23]), .A2(n6782), .Z(n4579) );
  AOI22D1BWP12T U2401 ( .A1(n5809), .A2(n4486), .B1(n5807), .B2(n4579), .ZN(
        n4593) );
  MUX2ND0BWP12T U2402 ( .I0(n5817), .I1(n5816), .S(b[15]), .ZN(n4488) );
  MUX2ND0BWP12T U2403 ( .I0(n5819), .I1(n5818), .S(b[14]), .ZN(n4487) );
  NR2D1BWP12T U2404 ( .A1(n4488), .A2(n4487), .ZN(n4592) );
  MUX2ND0BWP12T U2405 ( .I0(n5811), .I1(n5810), .S(b[25]), .ZN(n4490) );
  MUX2ND0BWP12T U2406 ( .I0(n5813), .I1(n5812), .S(b[24]), .ZN(n4489) );
  NR2D1BWP12T U2407 ( .A1(n4490), .A2(n4489), .ZN(n4591) );
  FA1D0BWP12T U2408 ( .A(n4493), .B(n4492), .CI(n4491), .CO(n4582), .S(n4516)
         );
  MUX2ND0BWP12T U2409 ( .I0(n5877), .I1(n5878), .S(n4494), .ZN(n4495) );
  NR2D1BWP12T U2410 ( .A1(n4496), .A2(n4495), .ZN(n4581) );
  MUX2ND0BWP12T U2411 ( .I0(a[27]), .I1(a[26]), .S(n4829), .ZN(n6551) );
  INVD1BWP12T U2412 ( .I(n6551), .ZN(n4874) );
  CKND2D1BWP12T U2413 ( .A1(a[27]), .A2(a[26]), .ZN(n6227) );
  INVD1BWP12T U2414 ( .I(n5866), .ZN(n4748) );
  XNR2D1BWP12T U2415 ( .A1(a[27]), .A2(n4498), .ZN(n4585) );
  FA1D0BWP12T U2416 ( .A(n4501), .B(n4500), .CI(n4499), .CO(n4608), .S(n4523)
         );
  FA1D0BWP12T U2417 ( .A(n4504), .B(n4503), .CI(n4502), .CO(n4607), .S(n4521)
         );
  MUX2ND0BWP12T U2418 ( .I0(n4747), .I1(n4746), .S(b[23]), .ZN(n4509) );
  MUX2ND0BWP12T U2419 ( .I0(n5860), .I1(n5861), .S(n5467), .ZN(n4508) );
  NR2D1BWP12T U2420 ( .A1(n4509), .A2(n4508), .ZN(n4595) );
  MAOI222D1BWP12T U2421 ( .A(n4512), .B(n4511), .C(n4510), .ZN(n4594) );
  MUX2D1BWP12T U2422 ( .I0(n5803), .I1(n5802), .S(n5379), .Z(n4514) );
  MUX2D1BWP12T U2423 ( .I0(n5805), .I1(n5804), .S(n5864), .Z(n4513) );
  ND2D1BWP12T U2424 ( .A1(n4514), .A2(n4513), .ZN(n4565) );
  XNR3XD1BWP12T U2425 ( .A1(n4563), .A2(n4565), .A3(n4564), .ZN(n4596) );
  FA1D0BWP12T U2426 ( .A(n4518), .B(n4517), .CI(n4516), .CO(n4553), .S(n4474)
         );
  XOR3D1BWP12T U2427 ( .A1(n4602), .A2(n4601), .A3(n4600), .Z(n4519) );
  NR2D1BWP12T U2428 ( .A1(n4520), .A2(n4519), .ZN(n4552) );
  ND2D1BWP12T U2429 ( .A1(n4520), .A2(n4519), .ZN(n4551) );
  FA1D0BWP12T U2430 ( .A(n4523), .B(n4522), .CI(n4521), .CO(n4550), .S(n4472)
         );
  NR2D1BWP12T U2431 ( .A1(n4707), .A2(n3409), .ZN(n4854) );
  FA1D0BWP12T U2432 ( .A(n4529), .B(n4528), .CI(n4527), .CO(n4682), .S(n4543)
         );
  FA1D0BWP12T U2433 ( .A(n4532), .B(n4531), .CI(n4530), .CO(n4466), .S(n4681)
         );
  FA1D0BWP12T U2434 ( .A(n4535), .B(n4534), .CI(n4533), .CO(n4471), .S(n4680)
         );
  INVD1BWP12T U2435 ( .I(n4536), .ZN(n4538) );
  MAOI222D1BWP12T U2436 ( .A(n4539), .B(n4538), .C(n4537), .ZN(n4677) );
  XNR3D1BWP12T U2437 ( .A1(n4542), .A2(n4541), .A3(n4540), .ZN(n4676) );
  FA1D0BWP12T U2438 ( .A(n4545), .B(n4544), .CI(n4543), .CO(n4675), .S(n4685)
         );
  FA1D0BWP12T U2439 ( .A(n4548), .B(n4547), .CI(n4546), .CO(n4467), .S(n4689)
         );
  INVD1BWP12T U2440 ( .I(n4549), .ZN(n4706) );
  NR2D1BWP12T U2441 ( .A1(n3407), .A2(n4706), .ZN(n4852) );
  NR2D1BWP12T U2442 ( .A1(n4854), .A2(n4852), .ZN(n5328) );
  INVD1BWP12T U2443 ( .I(n5328), .ZN(n6073) );
  FA1D0BWP12T U2444 ( .A(n4556), .B(n4555), .CI(n4554), .CO(n4613), .S(n4602)
         );
  XOR2XD1BWP12T U2445 ( .A1(a[27]), .A2(a[28]), .Z(n5849) );
  CKND2D1BWP12T U2446 ( .A1(n5849), .A2(n4823), .ZN(n4628) );
  XOR3D1BWP12T U2447 ( .A1(n4628), .A2(n4629), .A3(n4630), .Z(n4659) );
  MUX2ND0BWP12T U2448 ( .I0(n5778), .I1(n5777), .S(b[17]), .ZN(n4558) );
  NR2D1BWP12T U2449 ( .A1(n4559), .A2(n4558), .ZN(n4658) );
  FA1D0BWP12T U2450 ( .A(n4562), .B(n4561), .CI(n4560), .CO(n4657), .S(n4555)
         );
  MAOI222D1BWP12T U2451 ( .A(n4565), .B(n4564), .C(n4563), .ZN(n4660) );
  MUX2D1BWP12T U2452 ( .I0(n5817), .I1(n5816), .S(b[16]), .Z(n4567) );
  MUX2XD0BWP12T U2453 ( .I0(n5819), .I1(n5818), .S(b[15]), .Z(n4566) );
  ND2D1BWP12T U2454 ( .A1(n4567), .A2(n4566), .ZN(n4667) );
  MUX2ND0BWP12T U2455 ( .I0(n3911), .I1(n5810), .S(b[26]), .ZN(n4569) );
  MUX2ND0BWP12T U2456 ( .I0(n5813), .I1(n5812), .S(b[25]), .ZN(n4568) );
  NR2D1BWP12T U2457 ( .A1(n4569), .A2(n4568), .ZN(n4670) );
  NR2D1BWP12T U2458 ( .A1(n4571), .A2(n4570), .ZN(n4669) );
  XNR3D1BWP12T U2459 ( .A1(n4667), .A2(n4670), .A3(n4669), .ZN(n4661) );
  XNR3D1BWP12T U2460 ( .A1(n4662), .A2(n4660), .A3(n4661), .ZN(n4653) );
  MUX2ND0BWP12T U2461 ( .I0(n5837), .I1(n5836), .S(b[20]), .ZN(n4573) );
  MUX2NXD0BWP12T U2462 ( .I0(n5839), .I1(n5838), .S(b[19]), .ZN(n4572) );
  NR2D1BWP12T U2463 ( .A1(n4573), .A2(n4572), .ZN(n4672) );
  MUX2ND0BWP12T U2464 ( .I0(n4747), .I1(n4746), .S(b[24]), .ZN(n4575) );
  MUX2ND0BWP12T U2465 ( .I0(n5861), .I1(n5860), .S(b[23]), .ZN(n4574) );
  NR2D1BWP12T U2466 ( .A1(n4575), .A2(n4574), .ZN(n4620) );
  MUX2NXD0BWP12T U2467 ( .I0(n5871), .I1(n5872), .S(n4576), .ZN(n4577) );
  NR2D1BWP12T U2468 ( .A1(n4578), .A2(n4577), .ZN(n4619) );
  XOR2D1BWP12T U2469 ( .A1(a[23]), .A2(n5864), .Z(n4634) );
  AOI22D1BWP12T U2470 ( .A1(n5809), .A2(n4579), .B1(n5807), .B2(n4634), .ZN(
        n4618) );
  XOR3D1BWP12T U2471 ( .A1(n4655), .A2(n4653), .A3(n4654), .Z(n4617) );
  FA1D0BWP12T U2472 ( .A(n4582), .B(n4581), .CI(n4580), .CO(n4616), .S(n4601)
         );
  XNR2D1BWP12T U2473 ( .A1(a[27]), .A2(n6520), .ZN(n4624) );
  OAI22D1BWP12T U2474 ( .A1(n5387), .A2(n4585), .B1(n4748), .B2(n4624), .ZN(
        n4643) );
  CKXOR2D1BWP12T U2475 ( .A1(a[25]), .A2(n6573), .Z(n4664) );
  AO22D1BWP12T U2476 ( .A1(n5847), .A2(n4586), .B1(n5845), .B2(n4664), .Z(
        n4641) );
  MUX2D1BWP12T U2477 ( .I0(n5803), .I1(n5802), .S(n5843), .Z(n4588) );
  MUX2D1BWP12T U2478 ( .I0(n5805), .I1(n5804), .S(n5379), .Z(n4587) );
  ND2D1BWP12T U2479 ( .A1(n4588), .A2(n4587), .ZN(n4642) );
  XNR3D1BWP12T U2480 ( .A1(n4643), .A2(n4641), .A3(n4642), .ZN(n4627) );
  MUX2ND0BWP12T U2481 ( .I0(n5406), .I1(n5407), .S(n4730), .ZN(n4589) );
  NR2D1BWP12T U2482 ( .A1(n4590), .A2(n4589), .ZN(n4626) );
  FA1D0BWP12T U2483 ( .A(n4593), .B(n4592), .CI(n4591), .CO(n4625), .S(n4597)
         );
  FA1D0BWP12T U2484 ( .A(n4599), .B(n4598), .CI(n4597), .CO(n4651), .S(n4554)
         );
  MAOI222D1BWP12T U2485 ( .A(n4602), .B(n4601), .C(n4600), .ZN(n4603) );
  INVD1BWP12T U2486 ( .I(n4603), .ZN(n4604) );
  NR2D1BWP12T U2487 ( .A1(n4605), .A2(n4604), .ZN(n4611) );
  ND2D1BWP12T U2488 ( .A1(n4605), .A2(n4604), .ZN(n4610) );
  FA1D0BWP12T U2489 ( .A(n4608), .B(n4607), .CI(n4606), .CO(n4609), .S(n4600)
         );
  NR2D1BWP12T U2490 ( .A1(n4709), .A2(n4708), .ZN(n6075) );
  INVD1BWP12T U2491 ( .I(n6075), .ZN(n5279) );
  FA1D0BWP12T U2492 ( .A(n4614), .B(n4613), .CI(n4612), .CO(n4719), .S(n4605)
         );
  FA1D0BWP12T U2493 ( .A(n4617), .B(n4616), .CI(n4615), .CO(n4718), .S(n4612)
         );
  FA1D0BWP12T U2494 ( .A(n4620), .B(n4619), .CI(n4618), .CO(n4785), .S(n4671)
         );
  MUX2NXD0BWP12T U2495 ( .I0(n5817), .I1(n5816), .S(b[17]), .ZN(n4622) );
  MUX2ND0BWP12T U2496 ( .I0(n5819), .I1(n5818), .S(b[16]), .ZN(n4621) );
  NR2D1BWP12T U2497 ( .A1(n4622), .A2(n4621), .ZN(n4784) );
  XNR2D1BWP12T U2498 ( .A1(a[27]), .A2(n6334), .ZN(n4749) );
  OAI22D1BWP12T U2499 ( .A1(n5387), .A2(n4624), .B1(n4749), .B2(n4748), .ZN(
        n4741) );
  XNR3D1BWP12T U2500 ( .A1(n4739), .A2(n4741), .A3(n4740), .ZN(n4783) );
  FA1D0BWP12T U2501 ( .A(n4627), .B(n4626), .CI(n4625), .CO(n4767), .S(n4652)
         );
  INVD1BWP12T U2502 ( .I(n4628), .ZN(n4631) );
  MAOI222D1BWP12T U2503 ( .A(n4631), .B(n4630), .C(n4629), .ZN(n4772) );
  MUX2ND0BWP12T U2504 ( .I0(n5811), .I1(n5810), .S(b[27]), .ZN(n4633) );
  MUX2ND0BWP12T U2505 ( .I0(n5813), .I1(n5812), .S(b[26]), .ZN(n4632) );
  NR2D1BWP12T U2506 ( .A1(n4633), .A2(n4632), .ZN(n4765) );
  XNR2D1BWP12T U2507 ( .A1(a[23]), .A2(n5379), .ZN(n4743) );
  MAOI22D0BWP12T U2508 ( .A1(n5809), .A2(n4634), .B1(n4742), .B2(n4743), .ZN(
        n4764) );
  XNR2D0BWP12T U2509 ( .A1(a[29]), .A2(a[28]), .ZN(n4635) );
  NR2D1BWP12T U2510 ( .A1(n5849), .A2(n4635), .ZN(n5851) );
  MUX2NXD0BWP12T U2511 ( .I0(a[29]), .I1(a[28]), .S(n4823), .ZN(n6554) );
  INVD1BWP12T U2512 ( .I(n6554), .ZN(n5435) );
  CKXOR2D1BWP12T U2513 ( .A1(a[29]), .A2(n5612), .Z(n4733) );
  AOI22D1BWP12T U2514 ( .A1(n5851), .A2(n5435), .B1(n5849), .B2(n4733), .ZN(
        n4763) );
  MUX2ND0BWP12T U2515 ( .I0(n5837), .I1(n5836), .S(b[21]), .ZN(n4637) );
  MUX2ND0BWP12T U2516 ( .I0(n5839), .I1(n5838), .S(b[20]), .ZN(n4636) );
  NR2D1BWP12T U2517 ( .A1(n4637), .A2(n4636), .ZN(n4729) );
  OAI21D0BWP12T U2518 ( .A1(a[27]), .A2(a[28]), .B(n4829), .ZN(n4638) );
  OAI211D1BWP12T U2519 ( .A1(n5310), .A2(n4907), .B(n4638), .C(a[29]), .ZN(
        n4728) );
  MUX2ND0BWP12T U2520 ( .I0(n5877), .I1(n5878), .S(n5467), .ZN(n4639) );
  NR2D1BWP12T U2521 ( .A1(n4640), .A2(n4639), .ZN(n4727) );
  MAOI222D1BWP12T U2522 ( .A(n4643), .B(n4642), .C(n4641), .ZN(n4776) );
  MUX2D1BWP12T U2523 ( .I0(n5761), .I1(n5760), .S(b[13]), .Z(n4644) );
  ND2D1BWP12T U2524 ( .A1(n4645), .A2(n4644), .ZN(n4650) );
  MUX2ND0BWP12T U2525 ( .I0(n4647), .I1(n4646), .S(b[29]), .ZN(n4648) );
  OAI21D0BWP12T U2526 ( .A1(b[28]), .A2(n5361), .B(n4648), .ZN(n4649) );
  ND2D1BWP12T U2527 ( .A1(n4650), .A2(n4649), .ZN(n5371) );
  XOR3D1BWP12T U2528 ( .A1(n4772), .A2(n4773), .A3(n4774), .Z(n4766) );
  MAOI222D0BWP12T U2529 ( .A(n4655), .B(n4654), .C(n4653), .ZN(n4656) );
  INVD1BWP12T U2530 ( .I(n4656), .ZN(n4726) );
  FA1D0BWP12T U2531 ( .A(n4659), .B(n4658), .CI(n4657), .CO(n4725), .S(n4655)
         );
  TPNR2D0BWP12T U2532 ( .A1(n4661), .A2(n4660), .ZN(n4663) );
  MOAI22D0BWP12T U2533 ( .A1(n4663), .A2(n4662), .B1(n4661), .B2(n4660), .ZN(
        n4771) );
  XOR2D1BWP12T U2534 ( .A1(a[25]), .A2(n6782), .Z(n4735) );
  AOI22D1BWP12T U2535 ( .A1(n5847), .A2(n4664), .B1(n5845), .B2(n4735), .ZN(
        n4752) );
  MUX2NXD0BWP12T U2536 ( .I0(n5803), .I1(n5802), .S(b[9]), .ZN(n4666) );
  MUX2NXD0BWP12T U2537 ( .I0(n5805), .I1(n5804), .S(n5843), .ZN(n4665) );
  NR2D1BWP12T U2538 ( .A1(n4666), .A2(n4665), .ZN(n4754) );
  XOR3D1BWP12T U2539 ( .A1(n4752), .A2(n4754), .A3(n4753), .Z(n4779) );
  INVD1BWP12T U2540 ( .I(n4667), .ZN(n4668) );
  MAOI222D1BWP12T U2541 ( .A(n4670), .B(n4669), .C(n4668), .ZN(n4782) );
  XOR3D1BWP12T U2542 ( .A1(n4780), .A2(n4779), .A3(n4782), .Z(n4770) );
  FA1D0BWP12T U2543 ( .A(n4673), .B(n4672), .CI(n4671), .CO(n4769), .S(n4654)
         );
  INVD1BWP12T U2544 ( .I(n4674), .ZN(n4710) );
  OR2XD1BWP12T U2545 ( .A1(n4711), .A2(n4710), .Z(n6081) );
  CKND2D1BWP12T U2546 ( .A1(n5279), .A2(n6081), .ZN(n4714) );
  NR2D1BWP12T U2547 ( .A1(n6073), .A2(n4714), .ZN(n4716) );
  FA1D0BWP12T U2548 ( .A(n4677), .B(n4676), .CI(n4675), .CO(n4690), .S(n4695)
         );
  FA1D0BWP12T U2549 ( .A(n4682), .B(n4681), .CI(n4680), .CO(n4691), .S(n4693)
         );
  INVD1BWP12T U2550 ( .I(n4683), .ZN(n4698) );
  FA1D0BWP12T U2551 ( .A(n4686), .B(n4685), .CI(n4684), .CO(n4687), .S(n4078)
         );
  INVD1BWP12T U2552 ( .I(n4687), .ZN(n4697) );
  OR2D2BWP12T U2553 ( .A1(n4698), .A2(n4697), .Z(n5061) );
  ND2D1BWP12T U2554 ( .A1(n4688), .A2(n5061), .ZN(n5005) );
  FA1D0BWP12T U2555 ( .A(n4691), .B(n4690), .CI(n4689), .CO(n4549), .S(n4692)
         );
  INVD1BWP12T U2556 ( .I(n4692), .ZN(n4702) );
  FA1D0BWP12T U2557 ( .A(n4695), .B(n4694), .CI(n4693), .CO(n4696), .S(n4683)
         );
  INVD1BWP12T U2558 ( .I(n4696), .ZN(n4701) );
  NR2D1BWP12T U2559 ( .A1(n4702), .A2(n4701), .ZN(n5006) );
  NR2D1BWP12T U2560 ( .A1(n5005), .A2(n5006), .ZN(n4704) );
  INVD1BWP12T U2561 ( .I(n5057), .ZN(n4700) );
  ND2D1BWP12T U2562 ( .A1(n4698), .A2(n4697), .ZN(n5060) );
  INVD1BWP12T U2563 ( .I(n5060), .ZN(n4699) );
  TPAOI21D2BWP12T U2564 ( .A1(n4700), .A2(n5061), .B(n4699), .ZN(n5004) );
  ND2D1BWP12T U2565 ( .A1(n4702), .A2(n4701), .ZN(n5007) );
  TPOAI21D1BWP12T U2566 ( .A1(n5004), .A2(n5006), .B(n5007), .ZN(n4703) );
  TPAOI21D2BWP12T U2567 ( .A1(n4705), .A2(n4704), .B(n4703), .ZN(n5339) );
  INVD2BWP12T U2568 ( .I(n5339), .ZN(n6078) );
  ND2D1BWP12T U2569 ( .A1(n3407), .A2(n4706), .ZN(n5647) );
  ND2D1BWP12T U2570 ( .A1(n4707), .A2(n3409), .ZN(n4855) );
  OAI21D1BWP12T U2571 ( .A1(n4854), .A2(n5647), .B(n4855), .ZN(n5337) );
  INVD1BWP12T U2572 ( .I(n5337), .ZN(n6076) );
  ND2D1BWP12T U2573 ( .A1(n4709), .A2(n4708), .ZN(n6074) );
  INVD0BWP12T U2574 ( .I(n6074), .ZN(n4712) );
  ND2D1BWP12T U2575 ( .A1(n4711), .A2(n4710), .ZN(n6080) );
  INVD1BWP12T U2576 ( .I(n6080), .ZN(n5331) );
  AOI21D1BWP12T U2577 ( .A1(n4712), .A2(n6081), .B(n5331), .ZN(n4713) );
  OAI21D1BWP12T U2578 ( .A1(n6076), .A2(n4714), .B(n4713), .ZN(n4715) );
  AOI21D1BWP12T U2579 ( .A1(n4716), .A2(n6078), .B(n4715), .ZN(n4790) );
  FA1D0BWP12T U2580 ( .A(n4719), .B(n4718), .CI(n4717), .CO(n4720), .S(n4674)
         );
  INVD1BWP12T U2581 ( .I(n4720), .ZN(n4788) );
  FA1D0BWP12T U2582 ( .A(n4723), .B(n4722), .CI(n4721), .CO(n5343), .S(n4717)
         );
  FA1D0BWP12T U2583 ( .A(n4726), .B(n4725), .CI(n4724), .CO(n5342), .S(n4721)
         );
  FA1D0BWP12T U2584 ( .A(n4729), .B(n4728), .CI(n4727), .CO(n5356), .S(n4775)
         );
  MUX2ND0BWP12T U2585 ( .I0(n5803), .I1(n5802), .S(n5806), .ZN(n4732) );
  MUX2NXD0BWP12T U2586 ( .I0(n5804), .I1(n5805), .S(n4730), .ZN(n4731) );
  NR2D1BWP12T U2587 ( .A1(n4732), .A2(n4731), .ZN(n5355) );
  XOR2D1BWP12T U2588 ( .A1(a[29]), .A2(n6520), .Z(n5386) );
  AOI22D1BWP12T U2589 ( .A1(n5851), .A2(n4733), .B1(n5849), .B2(n5386), .ZN(
        n5365) );
  XNR2D1BWP12T U2590 ( .A1(a[25]), .A2(b[6]), .ZN(n5381) );
  INVD1BWP12T U2591 ( .I(n5381), .ZN(n4734) );
  AOI22D1BWP12T U2592 ( .A1(n5847), .A2(n4735), .B1(n5845), .B2(n4734), .ZN(
        n5363) );
  MUX2ND0BWP12T U2593 ( .I0(n5776), .I1(n5775), .S(b[20]), .ZN(n4737) );
  MUX2ND0BWP12T U2594 ( .I0(n5778), .I1(n5777), .S(b[19]), .ZN(n4736) );
  NR2D1BWP12T U2595 ( .A1(n4737), .A2(n4736), .ZN(n5364) );
  XOR3D1BWP12T U2596 ( .A1(n5365), .A2(n5363), .A3(n5364), .Z(n5354) );
  MAOI222D1BWP12T U2597 ( .A(n4741), .B(n4740), .C(n4739), .ZN(n5357) );
  XNR2D1BWP12T U2598 ( .A1(a[23]), .A2(n5843), .ZN(n5403) );
  OAI22D1BWP12T U2599 ( .A1(n4744), .A2(n4743), .B1(n4742), .B2(n5403), .ZN(
        n5392) );
  XNR3D1BWP12T U2600 ( .A1(n5392), .A2(n5394), .A3(n5393), .ZN(n5358) );
  XOR3D1BWP12T U2601 ( .A1(n5359), .A2(n5357), .A3(n5358), .Z(n5348) );
  XNR2XD1BWP12T U2602 ( .A1(a[27]), .A2(n6573), .ZN(n5388) );
  OAI22D1BWP12T U2603 ( .A1(n5387), .A2(n4749), .B1(n4748), .B2(n5388), .ZN(
        n5351) );
  MUX2ND0BWP12T U2604 ( .I0(n5811), .I1(n5810), .S(b[28]), .ZN(n4751) );
  MUX2ND0BWP12T U2605 ( .I0(n5813), .I1(n5812), .S(b[27]), .ZN(n4750) );
  NR2D1BWP12T U2606 ( .A1(n4751), .A2(n4750), .ZN(n5375) );
  MAOI222D1BWP12T U2607 ( .A(n4754), .B(n4753), .C(n4752), .ZN(n5378) );
  XNR3D1BWP12T U2608 ( .A1(n5398), .A2(n5400), .A3(n5399), .ZN(n5377) );
  XOR3D1BWP12T U2609 ( .A1(n5375), .A2(n5378), .A3(n5377), .Z(n5349) );
  INVD1BWP12T U2610 ( .I(b[30]), .ZN(n5419) );
  XOR2XD1BWP12T U2611 ( .A1(a[30]), .A2(a[29]), .Z(n5768) );
  ND2D1BWP12T U2612 ( .A1(n5768), .A2(n4823), .ZN(n5383) );
  MUX2XD0BWP12T U2613 ( .I0(n4757), .I1(n4756), .S(b[22]), .Z(n4762) );
  CKMUX2D1BWP12T U2614 ( .I0(n4760), .I1(n4759), .S(n4758), .Z(n4761) );
  NR2D1BWP12T U2615 ( .A1(n4762), .A2(n4761), .ZN(n5384) );
  FA1D0BWP12T U2616 ( .A(n4765), .B(n4764), .CI(n4763), .CO(n5370), .S(n4773)
         );
  XOR3D1BWP12T U2617 ( .A1(n5351), .A2(n5349), .A3(n5350), .Z(n5347) );
  FA1D0BWP12T U2618 ( .A(n4768), .B(n4767), .CI(n4766), .CO(n5411), .S(n4723)
         );
  FA1D0BWP12T U2619 ( .A(n4771), .B(n4770), .CI(n4769), .CO(n5409), .S(n4724)
         );
  MAOI222D1BWP12T U2620 ( .A(n4777), .B(n4776), .C(n4775), .ZN(n4778) );
  INVD1BWP12T U2621 ( .I(n4778), .ZN(n5374) );
  INVD1BWP12T U2622 ( .I(n4779), .ZN(n4781) );
  MAOI222D1BWP12T U2623 ( .A(n4782), .B(n4781), .C(n4780), .ZN(n5373) );
  FA1D0BWP12T U2624 ( .A(n4785), .B(n4784), .CI(n4783), .CO(n5372), .S(n4768)
         );
  INVD1BWP12T U2625 ( .I(n4786), .ZN(n4787) );
  OR2XD1BWP12T U2626 ( .A1(n4788), .A2(n4787), .Z(n5332) );
  ND2D1BWP12T U2627 ( .A1(n4788), .A2(n4787), .ZN(n5329) );
  ND2D1BWP12T U2628 ( .A1(n5332), .A2(n5329), .ZN(n4789) );
  XOR2XD1BWP12T U2629 ( .A1(n4790), .A2(n4789), .Z(n6069) );
  IND2D1BWP12T U2630 ( .A1(b[26]), .B1(a[26]), .ZN(n4863) );
  INVD1BWP12T U2631 ( .I(n4863), .ZN(n6503) );
  IND2D1BWP12T U2632 ( .A1(a[25]), .B1(b[25]), .ZN(n5693) );
  IND2D1BWP12T U2633 ( .A1(b[25]), .B1(a[25]), .ZN(n6494) );
  ND2D1BWP12T U2634 ( .A1(n5693), .A2(n6494), .ZN(n5051) );
  IND2XD1BWP12T U2635 ( .A1(b[24]), .B1(a[24]), .ZN(n5082) );
  IND2D1BWP12T U2636 ( .A1(a[24]), .B1(b[24]), .ZN(n5065) );
  INVD1BWP12T U2637 ( .I(n5065), .ZN(n6452) );
  AOI21D1BWP12T U2638 ( .A1(n4791), .A2(n6504), .B(n6452), .ZN(n5011) );
  IND2D1BWP12T U2639 ( .A1(a[26]), .B1(b[26]), .ZN(n6470) );
  ND2D1BWP12T U2640 ( .A1(n6470), .A2(n4863), .ZN(n5652) );
  INVD1BWP12T U2641 ( .I(n5652), .ZN(n5697) );
  CKND2D1BWP12T U2642 ( .A1(n5697), .A2(n5693), .ZN(n4859) );
  NR2D1BWP12T U2643 ( .A1(n4907), .A2(b[27]), .ZN(n6489) );
  NR2D1BWP12T U2644 ( .A1(n4882), .A2(a[27]), .ZN(n6454) );
  NR2D1BWP12T U2645 ( .A1(n6489), .A2(n6454), .ZN(n4867) );
  INVD1BWP12T U2646 ( .I(n4867), .ZN(n4862) );
  AOI21D1BWP12T U2647 ( .A1(n4859), .A2(n4863), .B(n4862), .ZN(n4792) );
  OAI31D1BWP12T U2648 ( .A1(n6503), .A2(n5051), .A3(n5011), .B(n4792), .ZN(
        n4860) );
  IND2D1BWP12T U2649 ( .A1(a[28]), .B1(b[28]), .ZN(n6164) );
  IND2D1BWP12T U2650 ( .A1(b[28]), .B1(a[28]), .ZN(n6480) );
  ND2D1BWP12T U2651 ( .A1(n6164), .A2(n6480), .ZN(n5321) );
  NR2D1BWP12T U2652 ( .A1(n5320), .A2(n5321), .ZN(n5968) );
  IND2D1BWP12T U2653 ( .A1(b[29]), .B1(a[29]), .ZN(n6845) );
  CKND0BWP12T U2654 ( .I(n4809), .ZN(n4795) );
  IND2XD1BWP12T U2655 ( .A1(a[29]), .B1(b[29]), .ZN(n6841) );
  ND2D1BWP12T U2656 ( .A1(n6841), .A2(n6164), .ZN(n5422) );
  NR2D1BWP12T U2657 ( .A1(n5968), .A2(n5422), .ZN(n4793) );
  INVD1BWP12T U2658 ( .I(n6845), .ZN(n4805) );
  OAI21D1BWP12T U2659 ( .A1(n4793), .A2(n4805), .B(n4804), .ZN(n5327) );
  INVD1BWP12T U2660 ( .I(n5327), .ZN(n4794) );
  INVD1BWP12T U2661 ( .I(n5422), .ZN(n6449) );
  NR2D1BWP12T U2662 ( .A1(n4809), .A2(n6449), .ZN(n4806) );
  AOI211D1BWP12T U2663 ( .A1(n5968), .A2(n4795), .B(n4794), .C(n4806), .ZN(
        n6001) );
  AOI22D1BWP12T U2664 ( .A1(n6069), .A2(n6834), .B1(n6001), .B2(n6728), .ZN(
        n4851) );
  AO21D1BWP12T U2665 ( .A1(n4797), .A2(n6107), .B(n4796), .Z(n5071) );
  OA21D1BWP12T U2666 ( .A1(n5071), .A2(n4798), .B(n6101), .Z(n5012) );
  AO21D1BWP12T U2667 ( .A1(n5012), .A2(n6104), .B(n4799), .Z(n5651) );
  OA21D1BWP12T U2668 ( .A1(n5651), .A2(n4800), .B(n6116), .Z(n4866) );
  AO21D1BWP12T U2669 ( .A1(n4866), .A2(n4802), .B(n4801), .Z(n5281) );
  AOI21D1BWP12T U2670 ( .A1(n5281), .A2(n6113), .B(n5311), .ZN(n6167) );
  INVD1BWP12T U2671 ( .I(n6842), .ZN(n5908) );
  CKND2D1BWP12T U2672 ( .A1(n6167), .A2(n5908), .ZN(n5911) );
  TPOAI21D1BWP12T U2673 ( .A1(n5052), .A2(n5051), .B(n5693), .ZN(n5649) );
  AOI211D1BWP12T U2674 ( .A1(n4867), .A2(n6503), .B(n6489), .C(n5321), .ZN(
        n4803) );
  OAI31D1BWP12T U2675 ( .A1(n4862), .A2(n5652), .A3(n5649), .B(n4803), .ZN(
        n6165) );
  INVD1BWP12T U2676 ( .I(n6165), .ZN(n5423) );
  NR2D1BWP12T U2677 ( .A1(n5423), .A2(n5422), .ZN(n5904) );
  OAI21D1BWP12T U2678 ( .A1(n5904), .A2(n4805), .B(n4804), .ZN(n4808) );
  INVD1BWP12T U2679 ( .I(n4806), .ZN(n4807) );
  OAI211D1BWP12T U2680 ( .A1(n4809), .A2(n6165), .B(n4808), .C(n4807), .ZN(
        n6162) );
  NR2D1BWP12T U2681 ( .A1(n6162), .A2(n6836), .ZN(n4849) );
  NR2D1BWP12T U2682 ( .A1(n4811), .A2(n4810), .ZN(n5015) );
  CKND2D1BWP12T U2683 ( .A1(n5015), .A2(n5047), .ZN(n5654) );
  NR2D1BWP12T U2684 ( .A1(n5654), .A2(a[26]), .ZN(n5653) );
  CKND2D1BWP12T U2685 ( .A1(n5653), .A2(n4907), .ZN(n6220) );
  NR2D1BWP12T U2686 ( .A1(n6220), .A2(a[28]), .ZN(n6224) );
  INVD1BWP12T U2687 ( .I(a[29]), .ZN(n6223) );
  ND2D1BWP12T U2688 ( .A1(n6224), .A2(n6223), .ZN(n6222) );
  NR2D1BWP12T U2689 ( .A1(n6222), .A2(a[30]), .ZN(n6597) );
  AO21D0BWP12T U2690 ( .A1(a[30]), .A2(n6222), .B(n6597), .Z(n6226) );
  ND2D1BWP12T U2691 ( .A1(n5118), .A2(n5575), .ZN(n6319) );
  INVD1BWP12T U2692 ( .I(n6319), .ZN(n4846) );
  MUX2ND0BWP12T U2693 ( .I0(a[18]), .I1(a[17]), .S(n4829), .ZN(n5674) );
  MUX2NXD0BWP12T U2694 ( .I0(a[22]), .I1(a[21]), .S(n4829), .ZN(n5683) );
  INVD1BWP12T U2695 ( .I(n5683), .ZN(n5663) );
  TPND2D0BWP12T U2696 ( .A1(n5660), .A2(n5663), .ZN(n4813) );
  AOI22D1BWP12T U2697 ( .A1(n5306), .A2(n5662), .B1(n5661), .B2(n4985), .ZN(
        n4812) );
  OAI211D1BWP12T U2698 ( .A1(n5674), .A2(n6409), .B(n4813), .C(n4812), .ZN(
        n6393) );
  INVD1BWP12T U2699 ( .I(n6393), .ZN(n5471) );
  TPND2D0BWP12T U2700 ( .A1(n5419), .A2(n6745), .ZN(n4814) );
  OAI211D0BWP12T U2701 ( .A1(a[30]), .A2(n6813), .B(n4814), .C(n6874), .ZN(
        n4818) );
  NR3D0BWP12T U2702 ( .A1(n5470), .A2(n4815), .A3(n6353), .ZN(n4817) );
  OAI22D0BWP12T U2703 ( .A1(n5416), .A2(n6880), .B1(a[30]), .B2(n6844), .ZN(
        n4816) );
  AOI211D0BWP12T U2704 ( .A1(n5417), .A2(n4818), .B(n4817), .C(n4816), .ZN(
        n4820) );
  INVD1BWP12T U2705 ( .I(n5470), .ZN(n6688) );
  ND2D1BWP12T U2706 ( .A1(n6304), .A2(a[31]), .ZN(n5585) );
  INVD1BWP12T U2707 ( .I(n5585), .ZN(n6358) );
  ND2D1BWP12T U2708 ( .A1(n6584), .A2(n4819), .ZN(n6686) );
  INVD1BWP12T U2709 ( .I(n6686), .ZN(n6661) );
  AOI21D1BWP12T U2710 ( .A1(n6688), .A2(n6358), .B(n6661), .ZN(n4886) );
  OAI211D0BWP12T U2711 ( .A1(n5471), .A2(n5719), .B(n4820), .C(n4886), .ZN(
        n4845) );
  CKND0BWP12T U2712 ( .I(n6521), .ZN(n4822) );
  AOI22D1BWP12T U2713 ( .A1(n6553), .A2(n5297), .B1(n5250), .B2(n6552), .ZN(
        n4821) );
  OAI21D1BWP12T U2714 ( .A1(n4822), .A2(n5767), .B(n4821), .ZN(n5624) );
  INVD1BWP12T U2715 ( .I(n5624), .ZN(n6523) );
  ND2D1BWP12T U2716 ( .A1(n6553), .A2(n4823), .ZN(n6246) );
  MUX2NXD0BWP12T U2717 ( .I0(a[28]), .I1(a[27]), .S(n4829), .ZN(n5291) );
  MUX2D1BWP12T U2718 ( .I0(a[24]), .I1(a[23]), .S(n6248), .Z(n5288) );
  INVD1BWP12T U2719 ( .I(n5288), .ZN(n5681) );
  AOI22D0BWP12T U2720 ( .A1(n6552), .A2(n5291), .B1(n5681), .B2(n6549), .ZN(
        n4825) );
  MUX2NXD0BWP12T U2721 ( .I0(a[26]), .I1(a[25]), .S(n4829), .ZN(n5680) );
  CKND2D0BWP12T U2722 ( .A1(n5680), .A2(n6556), .ZN(n4824) );
  OAI211D0BWP12T U2723 ( .A1(a[29]), .A2(n6246), .B(n4825), .C(n4824), .ZN(
        n4828) );
  NR2D1BWP12T U2724 ( .A1(n6576), .A2(n6573), .ZN(n6562) );
  AOI22D0BWP12T U2725 ( .A1(n6553), .A2(n5683), .B1(n5673), .B2(n6549), .ZN(
        n4827) );
  INVD1BWP12T U2726 ( .I(n5306), .ZN(n5682) );
  AOI22D0BWP12T U2727 ( .A1(n6556), .A2(n5674), .B1(n5682), .B2(n6552), .ZN(
        n4826) );
  ND2D1BWP12T U2728 ( .A1(n4827), .A2(n4826), .ZN(n5475) );
  AOI22D0BWP12T U2729 ( .A1(n4828), .A2(n6578), .B1(n6562), .B2(n5475), .ZN(
        n4834) );
  NR2D1BWP12T U2730 ( .A1(n6565), .A2(n6334), .ZN(n5302) );
  MUX2D1BWP12T U2731 ( .I0(a[14]), .I1(a[13]), .S(n6248), .Z(n5658) );
  INVD1BWP12T U2732 ( .I(n5298), .ZN(n4835) );
  RCOAI22D0BWP12T U2733 ( .A1(n5658), .A2(n6534), .B1(n4835), .B2(n5677), .ZN(
        n4831) );
  INVD1BWP12T U2734 ( .I(n5299), .ZN(n4836) );
  MUX2NXD0BWP12T U2735 ( .I0(n6231), .I1(n6230), .S(n4829), .ZN(n5675) );
  INVD1BWP12T U2736 ( .I(n5675), .ZN(n4837) );
  OAI22D0BWP12T U2737 ( .A1(n4836), .A2(n6530), .B1(n4837), .B2(n6533), .ZN(
        n4830) );
  NR2D1BWP12T U2738 ( .A1(n4831), .A2(n4830), .ZN(n5477) );
  INVD1BWP12T U2739 ( .I(n5477), .ZN(n6515) );
  ND2D1BWP12T U2740 ( .A1(n6268), .A2(n6565), .ZN(n6219) );
  NR2D0BWP12T U2741 ( .A1(n6219), .A2(a[30]), .ZN(n4832) );
  AOI211D0BWP12T U2742 ( .A1(n5302), .A2(n6515), .B(n4832), .C(n6560), .ZN(
        n4833) );
  OAI211D1BWP12T U2743 ( .A1(n6523), .A2(n5305), .B(n4834), .C(n4833), .ZN(
        n6571) );
  CKND2D1BWP12T U2744 ( .A1(n5289), .A2(n4835), .ZN(n4840) );
  TPND2D0BWP12T U2745 ( .A1(n5660), .A2(n5658), .ZN(n4839) );
  AOI22D1BWP12T U2746 ( .A1(n5662), .A2(n4837), .B1(n5661), .B2(n4836), .ZN(
        n4838) );
  ND3D1BWP12T U2747 ( .A1(n4840), .A2(n4839), .A3(n4838), .ZN(n6392) );
  INVD1BWP12T U2748 ( .I(n6392), .ZN(n5623) );
  ND2D1BWP12T U2749 ( .A1(n5664), .A2(n6219), .ZN(n6417) );
  NR2D1BWP12T U2750 ( .A1(n6409), .A2(n5252), .ZN(n4843) );
  NR2D1BWP12T U2751 ( .A1(n6410), .A2(n5297), .ZN(n4842) );
  OAI22D1BWP12T U2752 ( .A1(n6407), .A2(n5250), .B1(n5072), .B2(n6533), .ZN(
        n4841) );
  NR3D1BWP12T U2753 ( .A1(n4843), .A2(n4842), .A3(n4841), .ZN(n6400) );
  ND2D1BWP12T U2754 ( .A1(n6436), .A2(n6565), .ZN(n5441) );
  OAI22D1BWP12T U2755 ( .A1(n6571), .A2(n6680), .B1(n6431), .B2(n6716), .ZN(
        n4844) );
  AOI211D1BWP12T U2756 ( .A1(n4846), .A2(n5479), .B(n4845), .C(n4844), .ZN(
        n4847) );
  OAI21D1BWP12T U2757 ( .A1(n6226), .A2(n6862), .B(n4847), .ZN(n4848) );
  AOI211D1BWP12T U2758 ( .A1(n6600), .A2(n6870), .B(n4849), .C(n4848), .ZN(
        n4850) );
  OAI211D1BWP12T U2759 ( .A1(n6004), .A2(n6894), .B(n4851), .C(n4850), .ZN(
        result[30]) );
  INVD1BWP12T U2760 ( .I(n4852), .ZN(n5648) );
  INVD1BWP12T U2761 ( .I(n5647), .ZN(n4853) );
  AOI21D1BWP12T U2762 ( .A1(n6078), .A2(n5648), .B(n4853), .ZN(n4858) );
  INVD1BWP12T U2763 ( .I(n4854), .ZN(n4856) );
  ND2D1BWP12T U2764 ( .A1(n4856), .A2(n4855), .ZN(n4857) );
  XOR2XD2BWP12T U2765 ( .A1(n4858), .A2(n4857), .Z(n6085) );
  NR2D1BWP12T U2766 ( .A1(n5011), .A2(n5051), .ZN(n5694) );
  NR2D1BWP12T U2767 ( .A1(n5694), .A2(n4859), .ZN(n5999) );
  CKND2D0BWP12T U2768 ( .A1(n4862), .A2(n4863), .ZN(n4861) );
  TPOAI21D0BWP12T U2769 ( .A1(n5999), .A2(n4861), .B(n4860), .ZN(n5998) );
  INVD1BWP12T U2770 ( .I(n4861), .ZN(n4864) );
  AOI21D1BWP12T U2771 ( .A1(n4863), .A2(n6160), .B(n4862), .ZN(n5278) );
  AOI21D1BWP12T U2772 ( .A1(n4864), .A2(n6160), .B(n5278), .ZN(n6157) );
  CKND2D1BWP12T U2773 ( .A1(n6157), .A2(n6898), .ZN(n4912) );
  OAI21D1BWP12T U2774 ( .A1(n6840), .A2(n4869), .B(n5470), .ZN(n4906) );
  OAI22D0BWP12T U2775 ( .A1(n6263), .A2(n5677), .B1(n4888), .B2(n6530), .ZN(
        n4871) );
  OAI22D0BWP12T U2776 ( .A1(n4889), .A2(n6534), .B1(n5165), .B2(n6533), .ZN(
        n4870) );
  NR2D1BWP12T U2777 ( .A1(n4871), .A2(n4870), .ZN(n6577) );
  ND2D1BWP12T U2778 ( .A1(n6577), .A2(n6576), .ZN(n6702) );
  ND2D1BWP12T U2779 ( .A1(n6517), .A2(n6334), .ZN(n6701) );
  CKND0BWP12T U2780 ( .I(n6562), .ZN(n4878) );
  OAI22D0BWP12T U2781 ( .A1(n5677), .A2(n6531), .B1(n6532), .B2(n6534), .ZN(
        n4873) );
  NR2D0BWP12T U2782 ( .A1(n5166), .A2(n6530), .ZN(n4872) );
  AOI211D1BWP12T U2783 ( .A1(n6552), .A2(n6538), .B(n4873), .C(n4872), .ZN(
        n6572) );
  OAI22D0BWP12T U2784 ( .A1(n5020), .A2(n5677), .B1(n4874), .B2(n6534), .ZN(
        n4876) );
  CKND0BWP12T U2785 ( .I(n6555), .ZN(n5436) );
  OAI22D0BWP12T U2786 ( .A1(n5436), .A2(n6533), .B1(n6535), .B2(n6530), .ZN(
        n4875) );
  OAI21D0BWP12T U2787 ( .A1(n4876), .A2(n4875), .B(n6578), .ZN(n4877) );
  OAI211D1BWP12T U2788 ( .A1(n4878), .A2(n6572), .B(n6355), .C(n4877), .ZN(
        n4879) );
  TPAOI31D0BWP12T U2789 ( .A1(n6573), .A2(n6702), .A3(n6701), .B(n4879), .ZN(
        n6581) );
  INVD1BWP12T U2790 ( .I(n6581), .ZN(n4887) );
  INVD1BWP12T U2791 ( .I(n6813), .ZN(n6879) );
  NR2D1BWP12T U2792 ( .A1(n4880), .A2(n6106), .ZN(n6816) );
  MUX2ND0BWP12T U2793 ( .I0(n6745), .I1(n6816), .S(b[27]), .ZN(n4881) );
  AOI21D0BWP12T U2794 ( .A1(n6874), .A2(n4881), .B(n4907), .ZN(n4884) );
  ND2D1BWP12T U2795 ( .A1(op[2]), .A2(n6816), .ZN(n5629) );
  OAI22D0BWP12T U2796 ( .A1(n4882), .A2(n5629), .B1(a[27]), .B2(n6844), .ZN(
        n4883) );
  AOI211D0BWP12T U2797 ( .A1(n6879), .A2(n6454), .B(n4884), .C(n4883), .ZN(
        n4885) );
  OAI211D1BWP12T U2798 ( .A1(n6680), .A2(n4887), .B(n4886), .C(n4885), .ZN(
        n4905) );
  NR2D1BWP12T U2799 ( .A1(n6409), .A2(n6263), .ZN(n4892) );
  OAI22D1BWP12T U2800 ( .A1(n5165), .A2(n6407), .B1(n6408), .B2(n4888), .ZN(
        n4891) );
  NR2D0BWP12T U2801 ( .A1(n6410), .A2(n4889), .ZN(n4890) );
  NR3D1BWP12T U2802 ( .A1(n4892), .A2(n4891), .A3(n4890), .ZN(n6420) );
  AOI22D1BWP12T U2803 ( .A1(n5660), .A2(n4894), .B1(n5662), .B2(n4893), .ZN(
        n6421) );
  NR2D1BWP12T U2804 ( .A1(n6409), .A2(n6531), .ZN(n4898) );
  OAI22D0BWP12T U2805 ( .A1(n6403), .A2(n4895), .B1(n6408), .B2(n5166), .ZN(
        n4897) );
  NR2D0BWP12T U2806 ( .A1(n6410), .A2(n6532), .ZN(n4896) );
  NR3D1BWP12T U2807 ( .A1(n4898), .A2(n4897), .A3(n4896), .ZN(n6418) );
  INVD1BWP12T U2808 ( .I(n6418), .ZN(n4902) );
  CKND2D0BWP12T U2809 ( .A1(n5660), .A2(n6551), .ZN(n4900) );
  AOI22D1BWP12T U2810 ( .A1(n5662), .A2(n6555), .B1(n5661), .B2(n5034), .ZN(
        n4899) );
  OAI211D0BWP12T U2811 ( .A1(n5020), .A2(n6409), .B(n4900), .C(n4899), .ZN(
        n4901) );
  AOI22D1BWP12T U2812 ( .A1(n5659), .A2(n4902), .B1(n4901), .B2(n6411), .ZN(
        n6425) );
  TPND3D0BWP12T U2813 ( .A1(n6425), .A2(n6857), .A3(n6219), .ZN(n4903) );
  AOI21D1BWP12T U2814 ( .A1(n6718), .A2(n6717), .B(n4903), .ZN(n4904) );
  AOI211D1BWP12T U2815 ( .A1(n6356), .A2(n4906), .B(n4905), .C(n4904), .ZN(
        n4909) );
  OAI211D1BWP12T U2816 ( .A1(n5653), .A2(n4907), .B(n6220), .C(n6786), .ZN(
        n4908) );
  OAI211D1BWP12T U2817 ( .A1(n6794), .A2(n6215), .B(n4909), .C(n4908), .ZN(
        n4910) );
  RCIAO21D0BWP12T U2818 ( .A1(n5964), .A2(n6894), .B(n4910), .ZN(n4911) );
  OAI211D1BWP12T U2819 ( .A1(n6890), .A2(n5998), .B(n4912), .C(n4911), .ZN(
        n4913) );
  XNR3D1BWP12T U2820 ( .A1(n6035), .A2(n4915), .A3(n4914), .ZN(n6037) );
  INVD1BWP12T U2821 ( .I(n6037), .ZN(n4955) );
  INVD1BWP12T U2822 ( .I(n5229), .ZN(n4918) );
  OAI22D1BWP12T U2823 ( .A1(n4918), .A2(n5236), .B1(n4922), .B2(n5176), .ZN(
        n4917) );
  INVD1BWP12T U2824 ( .I(n5230), .ZN(n4919) );
  NR2XD0BWP12T U2825 ( .A1(n4919), .A2(n5232), .ZN(n4916) );
  NR2D1BWP12T U2826 ( .A1(n4917), .A2(n4916), .ZN(n6299) );
  CKND1BWP12T U2827 ( .I(n5731), .ZN(n4923) );
  NR2D0BWP12T U2828 ( .A1(n4925), .A2(n6308), .ZN(n4930) );
  OAI22D1BWP12T U2829 ( .A1(n5237), .A2(a[19]), .B1(a[22]), .B2(n5235), .ZN(
        n4927) );
  OAI22D1BWP12T U2830 ( .A1(a[20]), .A2(n5238), .B1(n5239), .B2(a[21]), .ZN(
        n4926) );
  NR2D1BWP12T U2831 ( .A1(n4927), .A2(n4926), .ZN(n6256) );
  OAI22D1BWP12T U2832 ( .A1(n6256), .A2(n6304), .B1(a[31]), .B2(n6306), .ZN(
        n4929) );
  NR2D1BWP12T U2833 ( .A1(n6255), .A2(n6297), .ZN(n4928) );
  NR3D1BWP12T U2834 ( .A1(n4930), .A2(n4929), .A3(n4928), .ZN(n6662) );
  AOI21D1BWP12T U2835 ( .A1(n6355), .A2(n6662), .B(n6350), .ZN(n4931) );
  OAI21D1BWP12T U2836 ( .A1(n4950), .A2(n4931), .B(n6336), .ZN(n6328) );
  ND2D1BWP12T U2837 ( .A1(n4932), .A2(n4952), .ZN(n5272) );
  TPOAI21D0BWP12T U2838 ( .A1(n4952), .A2(n4932), .B(n5272), .ZN(n5933) );
  TPNR2D0BWP12T U2839 ( .A1(n6877), .A2(n6886), .ZN(n4933) );
  MUX2ND0BWP12T U2840 ( .I0(n4933), .I1(n6874), .S(n6247), .ZN(n4940) );
  CKND2D0BWP12T U2841 ( .A1(n4935), .A2(n4934), .ZN(n4937) );
  OAI211D1BWP12T U2842 ( .A1(n6247), .A2(op[2]), .B(n6334), .C(n6816), .ZN(
        n4936) );
  OAI211D0BWP12T U2843 ( .A1(n6683), .A2(n4938), .B(n4937), .C(n4936), .ZN(
        n4939) );
  AOI211D1BWP12T U2844 ( .A1(n6879), .A2(n4952), .B(n4940), .C(n4939), .ZN(
        n4941) );
  TPOAI21D0BWP12T U2845 ( .A1(n6421), .A2(n6892), .B(n4941), .ZN(n4944) );
  NR2XD0BWP12T U2846 ( .A1(n5981), .A2(n6890), .ZN(n4943) );
  AOI211D1BWP12T U2847 ( .A1(n6873), .A2(n6517), .B(n4944), .C(n4943), .ZN(
        n4945) );
  OAI21D1BWP12T U2848 ( .A1(n5933), .A2(n6894), .B(n4945), .ZN(n4948) );
  INVD1BWP12T U2849 ( .I(n6497), .ZN(n6883) );
  ND2D1BWP12T U2850 ( .A1(n4946), .A2(n6883), .ZN(n5227) );
  NR2D1BWP12T U2851 ( .A1(n6138), .A2(n6836), .ZN(n4947) );
  AOI211D1BWP12T U2852 ( .A1(n6909), .A2(n6328), .B(n4948), .C(n4947), .ZN(
        n4954) );
  ND2D1BWP12T U2853 ( .A1(n6254), .A2(n5237), .ZN(n4949) );
  ND2D1BWP12T U2854 ( .A1(n6662), .A2(n4949), .ZN(n6665) );
  AOI21D1BWP12T U2855 ( .A1(n6573), .A2(n6665), .B(n4950), .ZN(n6287) );
  INVD1BWP12T U2856 ( .I(n6181), .ZN(n4951) );
  CKND2D1BWP12T U2857 ( .A1(n4951), .A2(n5979), .ZN(n5266) );
  MAOI22D0BWP12T U2858 ( .A1(n6287), .A2(n6905), .B1(n6186), .B2(n6794), .ZN(
        n4953) );
  INVD1BWP12T U2859 ( .I(n4956), .ZN(n5524) );
  TPOAI21D1BWP12T U2860 ( .A1(n5524), .A2(n5522), .B(n5523), .ZN(n4961) );
  INVD1BWP12T U2861 ( .I(n4957), .ZN(n4959) );
  CKND2D1BWP12T U2862 ( .A1(n4959), .A2(n4958), .ZN(n4960) );
  NR2D1BWP12T U2863 ( .A1(n6146), .A2(n6836), .ZN(n4999) );
  CKND2D1BWP12T U2864 ( .A1(n5661), .A2(n5249), .ZN(n5730) );
  INVD1BWP12T U2865 ( .I(n6763), .ZN(n5081) );
  OAI22D1BWP12T U2866 ( .A1(n5237), .A2(a[24]), .B1(a[27]), .B2(n5235), .ZN(
        n4966) );
  OAI22D1BWP12T U2867 ( .A1(a[25]), .A2(n5238), .B1(n5239), .B2(a[26]), .ZN(
        n4965) );
  NR2D1BWP12T U2868 ( .A1(n4966), .A2(n4965), .ZN(n5245) );
  INVD1BWP12T U2869 ( .I(n5245), .ZN(n5572) );
  OAI22D1BWP12T U2870 ( .A1(n5237), .A2(n4967), .B1(n6654), .B2(n5235), .ZN(
        n4969) );
  OAI22D1BWP12T U2871 ( .A1(n6646), .A2(n5239), .B1(n5238), .B2(n5728), .ZN(
        n4968) );
  NR2D1BWP12T U2872 ( .A1(n4969), .A2(n4968), .ZN(n6309) );
  OAI22D1BWP12T U2873 ( .A1(n5572), .A2(n6308), .B1(n6309), .B2(n6304), .ZN(
        n4976) );
  OAI22D1BWP12T U2874 ( .A1(n5237), .A2(a[28]), .B1(a[31]), .B2(n5235), .ZN(
        n4971) );
  OAI22D1BWP12T U2875 ( .A1(a[29]), .A2(n5238), .B1(n5239), .B2(a[30]), .ZN(
        n4970) );
  NR2D1BWP12T U2876 ( .A1(n4971), .A2(n4970), .ZN(n6322) );
  INVD1BWP12T U2877 ( .I(n6322), .ZN(n5282) );
  OAI22D1BWP12T U2878 ( .A1(n5237), .A2(n4972), .B1(n5069), .B2(n5235), .ZN(
        n4974) );
  OAI22D1BWP12T U2879 ( .A1(n5487), .A2(n5239), .B1(n5238), .B2(n6623), .ZN(
        n4973) );
  NR2D1BWP12T U2880 ( .A1(n4974), .A2(n4973), .ZN(n6307) );
  OAI22D1BWP12T U2881 ( .A1(n5282), .A2(n6306), .B1(n6307), .B2(n6297), .ZN(
        n4975) );
  NR2D1BWP12T U2882 ( .A1(n4976), .A2(n4975), .ZN(n6343) );
  INVD1BWP12T U2883 ( .I(n5479), .ZN(n6666) );
  INVD1BWP12T U2884 ( .I(n5658), .ZN(n5676) );
  AOI22D0BWP12T U2885 ( .A1(n6556), .A2(n5675), .B1(n5676), .B2(n6552), .ZN(
        n4978) );
  AOI22D0BWP12T U2886 ( .A1(n6553), .A2(n5673), .B1(n5298), .B2(n6549), .ZN(
        n4977) );
  ND2D1BWP12T U2887 ( .A1(n4978), .A2(n4977), .ZN(n5077) );
  ND2D1BWP12T U2888 ( .A1(n6268), .A2(a[0]), .ZN(n6519) );
  CKND0BWP12T U2889 ( .I(n6519), .ZN(n4987) );
  AOI22D1BWP12T U2890 ( .A1(n6556), .A2(n5250), .B1(n5252), .B2(n6549), .ZN(
        n4980) );
  AOI22D1BWP12T U2891 ( .A1(n6553), .A2(n5299), .B1(n5297), .B2(n6552), .ZN(
        n4979) );
  ND2D1BWP12T U2892 ( .A1(n4980), .A2(n4979), .ZN(n5073) );
  ND2D1BWP12T U2893 ( .A1(n5073), .A2(n6334), .ZN(n4981) );
  OAI211D1BWP12T U2894 ( .A1(n4987), .A2(n6565), .B(n4981), .C(n6355), .ZN(
        n4982) );
  RCAOI21D0BWP12T U2895 ( .A1(n6578), .A2(n5077), .B(n4982), .ZN(n6545) );
  MOAI22D0BWP12T U2896 ( .A1(n6343), .A2(n6666), .B1(n6545), .B2(n6855), .ZN(
        n4990) );
  NR2D1BWP12T U2897 ( .A1(n6409), .A2(n5675), .ZN(n4984) );
  OAI22D1BWP12T U2898 ( .A1(n6408), .A2(n5298), .B1(n6407), .B2(n5676), .ZN(
        n4983) );
  AOI211D1BWP12T U2899 ( .A1(n5660), .A2(n4985), .B(n4984), .C(n4983), .ZN(
        n5080) );
  NR2D1BWP12T U2900 ( .A1(n6565), .A2(n6716), .ZN(n6755) );
  INVD1BWP12T U2901 ( .I(n6874), .ZN(n6744) );
  TPOAI21D0BWP12T U2902 ( .A1(n6114), .A2(n6744), .B(n6621), .ZN(n4992) );
  CKND0BWP12T U2903 ( .I(n4992), .ZN(n4986) );
  AOI22D1BWP12T U2904 ( .A1(n4987), .A2(n6755), .B1(b[16]), .B2(n4986), .ZN(
        n4988) );
  OAI211D0BWP12T U2905 ( .A1(n5080), .A2(n6892), .B(n6686), .C(n4988), .ZN(
        n4989) );
  AOI211D1BWP12T U2906 ( .A1(n5546), .A2(n5081), .B(n4990), .C(n4989), .ZN(
        n4997) );
  INVD0BWP12T U2907 ( .I(n5636), .ZN(n4991) );
  AOI21D1BWP12T U2908 ( .A1(n4991), .A2(n6786), .B(n6783), .ZN(n5611) );
  OAI21D0BWP12T U2909 ( .A1(n5538), .A2(n6862), .B(n5611), .ZN(n4995) );
  ND2D1BWP12T U2910 ( .A1(n5636), .A2(n6786), .ZN(n5724) );
  INVD1BWP12T U2911 ( .I(n6880), .ZN(n6747) );
  MUX2ND0BWP12T U2912 ( .I0(n6655), .I1(n6747), .S(b[16]), .ZN(n4993) );
  OAI211D0BWP12T U2913 ( .A1(n6232), .A2(n5724), .B(n4993), .C(n4992), .ZN(
        n4994) );
  MUX2ND0BWP12T U2914 ( .I0(n4995), .I1(n4994), .S(a[16]), .ZN(n4996) );
  OAI211D1BWP12T U2915 ( .A1(n6794), .A2(n6203), .B(n4997), .C(n4996), .ZN(
        n4998) );
  AOI211D1BWP12T U2916 ( .A1(n6833), .A2(n5953), .B(n4999), .C(n4998), .ZN(
        n5003) );
  XNR2XD1BWP12T U2917 ( .A1(n5001), .A2(n5000), .ZN(n5990) );
  ND2D1BWP12T U2918 ( .A1(n5990), .A2(n6728), .ZN(n5002) );
  OAI211D4BWP12T U2919 ( .A1(n6902), .A2(n6052), .B(n5003), .C(n5002), .ZN(
        result[16]) );
  INVD1BWP12T U2920 ( .I(n5006), .ZN(n5008) );
  CKND2D1BWP12T U2921 ( .A1(n5008), .A2(n5007), .ZN(n5009) );
  XNR2D1BWP12T U2922 ( .A1(n5010), .A2(n5009), .ZN(n6072) );
  AOI21D1BWP12T U2923 ( .A1(n5011), .A2(n5051), .B(n5694), .ZN(n5997) );
  NR2D1BWP12T U2924 ( .A1(n5963), .A2(n6894), .ZN(n5050) );
  INVD1BWP12T U2925 ( .I(n5629), .ZN(n5509) );
  INVD1BWP12T U2926 ( .I(n6816), .ZN(n6704) );
  MUX2ND0BWP12T U2927 ( .I0(n6683), .I1(n6704), .S(b[25]), .ZN(n5014) );
  AOI211D1BWP12T U2928 ( .A1(n5015), .A2(n6786), .B(n5509), .C(n5014), .ZN(
        n5048) );
  AO21D0BWP12T U2929 ( .A1(n5016), .A2(n6862), .B(n5015), .Z(n5092) );
  OAI21D1BWP12T U2930 ( .A1(n5092), .A2(n6862), .B(n6844), .ZN(n5017) );
  CKND2D0BWP12T U2931 ( .A1(n5017), .A2(n5047), .ZN(n5046) );
  MUX2NXD0BWP12T U2932 ( .I0(n5209), .I1(n6353), .S(n6351), .ZN(n6327) );
  NR2D1BWP12T U2933 ( .A1(n6409), .A2(n6535), .ZN(n5022) );
  OAI22D1BWP12T U2934 ( .A1(n5020), .A2(n6407), .B1(n6408), .B2(n6532), .ZN(
        n5021) );
  AOI211D0BWP12T U2935 ( .A1(n5660), .A2(n6555), .B(n5022), .C(n5021), .ZN(
        n5029) );
  INVD1BWP12T U2936 ( .I(n6411), .ZN(n6439) );
  NR2D1BWP12T U2937 ( .A1(n6409), .A2(n5179), .ZN(n5026) );
  OAI22D1BWP12T U2938 ( .A1(n5023), .A2(n6407), .B1(n6408), .B2(n5178), .ZN(
        n5025) );
  NR2D0BWP12T U2939 ( .A1(n6410), .A2(n6538), .ZN(n5024) );
  NR3D1BWP12T U2940 ( .A1(n5026), .A2(n5025), .A3(n5024), .ZN(n6399) );
  AOI22D1BWP12T U2941 ( .A1(n5664), .A2(n6395), .B1(n6399), .B2(n5659), .ZN(
        n5028) );
  CKND0BWP12T U2942 ( .I(n6219), .ZN(n5665) );
  AOI21D0BWP12T U2943 ( .A1(n6380), .A2(n5666), .B(n5665), .ZN(n5027) );
  OAI211D1BWP12T U2944 ( .A1(n5029), .A2(n6439), .B(n5028), .C(n5027), .ZN(
        n6433) );
  AOI22D0BWP12T U2945 ( .A1(n6556), .A2(n5175), .B1(n5173), .B2(n6549), .ZN(
        n5031) );
  AOI22D0BWP12T U2946 ( .A1(n6553), .A2(n5176), .B1(n5177), .B2(n6552), .ZN(
        n5030) );
  ND2D1BWP12T U2947 ( .A1(n5031), .A2(n5030), .ZN(n5707) );
  MUX2ND0BWP12T U2948 ( .I0(n5707), .I1(n6518), .S(n6334), .ZN(n6510) );
  AOI22D0BWP12T U2949 ( .A1(n6553), .A2(n6538), .B1(n5178), .B2(n6549), .ZN(
        n5033) );
  CKND2D0BWP12T U2950 ( .A1(n5179), .A2(n6556), .ZN(n5032) );
  OAI211D0BWP12T U2951 ( .A1(n6531), .A2(n6533), .B(n5033), .C(n5032), .ZN(
        n5711) );
  AOI22D0BWP12T U2952 ( .A1(n6552), .A2(n6550), .B1(n6555), .B2(n6553), .ZN(
        n5037) );
  AOI22D0BWP12T U2953 ( .A1(n6549), .A2(n5035), .B1(n5034), .B2(n6556), .ZN(
        n5036) );
  AOI21D0BWP12T U2954 ( .A1(n5037), .A2(n5036), .B(n6557), .ZN(n5038) );
  AOI211D0BWP12T U2955 ( .A1(n5711), .A2(n6562), .B(n5038), .C(n6560), .ZN(
        n5039) );
  OAI21D1BWP12T U2956 ( .A1(n6510), .A2(n6565), .B(n5039), .ZN(n6529) );
  OAI22D1BWP12T U2957 ( .A1(n6433), .A2(n6716), .B1(n6529), .B2(n6680), .ZN(
        n5044) );
  CKND0BWP12T U2958 ( .I(n6323), .ZN(n5040) );
  OAI22D1BWP12T U2959 ( .A1(n6274), .A2(n6304), .B1(n5040), .B2(n6297), .ZN(
        n6279) );
  INVD1BWP12T U2960 ( .I(n6279), .ZN(n5042) );
  AOI22D0BWP12T U2961 ( .A1(n5051), .A2(n6879), .B1(b[25]), .B2(n6744), .ZN(
        n5041) );
  OAI21D1BWP12T U2962 ( .A1(n6840), .A2(n5042), .B(n5041), .ZN(n5043) );
  AOI211D1BWP12T U2963 ( .A1(n6909), .A2(n6327), .B(n5044), .C(n5043), .ZN(
        n5045) );
  OAI211D1BWP12T U2964 ( .A1(n5048), .A2(n5047), .B(n5046), .C(n5045), .ZN(
        n5049) );
  AOI211D1BWP12T U2965 ( .A1(n6870), .A2(n6213), .B(n5050), .C(n5049), .ZN(
        n5055) );
  XOR2XD1BWP12T U2966 ( .A1(n5052), .A2(n5051), .Z(n6156) );
  INVD1BWP12T U2967 ( .I(n6156), .ZN(n5053) );
  ND2D1BWP12T U2968 ( .A1(n5053), .A2(n6898), .ZN(n5054) );
  OAI211D1BWP12T U2969 ( .A1(n5997), .A2(n6890), .B(n5055), .C(n5054), .ZN(
        n5056) );
  TPOAI21D1BWP12T U2970 ( .A1(n5059), .A2(n5058), .B(n5057), .ZN(n5063) );
  ND2D1BWP12T U2971 ( .A1(n5061), .A2(n5060), .ZN(n5062) );
  XNR2D2BWP12T U2972 ( .A1(n5063), .A2(n5062), .ZN(n6071) );
  INVD1BWP12T U2973 ( .I(n6155), .ZN(n5064) );
  NR2D1BWP12T U2974 ( .A1(n5064), .A2(n5095), .ZN(n5066) );
  ND2D1BWP12T U2975 ( .A1(n5065), .A2(n5082), .ZN(n5097) );
  XOR2XD1BWP12T U2976 ( .A1(n5066), .A2(n5097), .Z(n6153) );
  INVD1BWP12T U2977 ( .I(n6153), .ZN(n5101) );
  CKND0BWP12T U2978 ( .I(b[24]), .ZN(n5083) );
  OAI211D0BWP12T U2979 ( .A1(n6704), .A2(n5083), .B(a[24]), .C(n5629), .ZN(
        n5068) );
  AOI21D0BWP12T U2980 ( .A1(n5070), .A2(n5069), .B(n5068), .ZN(n5093) );
  ND2D1BWP12T U2981 ( .A1(n6212), .A2(n6870), .ZN(n5091) );
  TPNR2D0BWP12T U2982 ( .A1(n6534), .A2(n5072), .ZN(n5079) );
  AOI22D0BWP12T U2983 ( .A1(n6553), .A2(n5681), .B1(n5683), .B2(n6552), .ZN(
        n5075) );
  AOI22D0BWP12T U2984 ( .A1(n6549), .A2(n5674), .B1(n5682), .B2(n6556), .ZN(
        n5074) );
  AOI21D0BWP12T U2985 ( .A1(n5075), .A2(n5074), .B(n6557), .ZN(n5076) );
  AOI211D0BWP12T U2986 ( .A1(n6562), .A2(n5077), .B(n5076), .C(n6560), .ZN(
        n5078) );
  OAI21D1BWP12T U2987 ( .A1(n6511), .A2(n6565), .B(n5078), .ZN(n6567) );
  INVD1BWP12T U2988 ( .I(n6567), .ZN(n5089) );
  ND2D1BWP12T U2989 ( .A1(n5079), .A2(n6334), .ZN(n6742) );
  NR2D1BWP12T U2990 ( .A1(n6432), .A2(n6716), .ZN(n5088) );
  AOI22D1BWP12T U2991 ( .A1(n5575), .A2(n5245), .B1(n6322), .B2(n6313), .ZN(
        n6735) );
  TPNR2D0BWP12T U2992 ( .A1(n5082), .A2(n6683), .ZN(n5085) );
  OAI22D0BWP12T U2993 ( .A1(n5083), .A2(n6874), .B1(a[24]), .B2(n6844), .ZN(
        n5084) );
  AOI211D0BWP12T U2994 ( .A1(n5097), .A2(n6879), .B(n5085), .C(n5084), .ZN(
        n5086) );
  OAI211D1BWP12T U2995 ( .A1(n6735), .A2(n6666), .B(n5086), .C(n6850), .ZN(
        n5087) );
  AOI211D1BWP12T U2996 ( .A1(n6855), .A2(n5089), .B(n5088), .C(n5087), .ZN(
        n5090) );
  OAI211D1BWP12T U2997 ( .A1(n5093), .A2(n5092), .B(n5091), .C(n5090), .ZN(
        n5094) );
  AOI21D1BWP12T U2998 ( .A1(n5960), .A2(n6833), .B(n5094), .ZN(n5100) );
  NR2D1BWP12T U2999 ( .A1(n5096), .A2(n5095), .ZN(n5098) );
  XOR2D1BWP12T U3000 ( .A1(n5098), .A2(n5097), .Z(n5996) );
  ND2D1BWP12T U3001 ( .A1(n5996), .A2(n6728), .ZN(n5099) );
  AO21D4BWP12T U3002 ( .A1(n6071), .A2(n6834), .B(n5102), .Z(result[24]) );
  XOR2XD1BWP12T U3003 ( .A1(n5106), .A2(n5139), .Z(n5983) );
  INVD1BWP12T U3004 ( .I(n5107), .ZN(n6177) );
  ND2D1BWP12T U3005 ( .A1(n6177), .A2(n6178), .ZN(n6176) );
  INVD1BWP12T U3006 ( .I(n6176), .ZN(n5109) );
  NR2D1BWP12T U3007 ( .A1(n5109), .A2(n5108), .ZN(n6188) );
  INVD1BWP12T U3008 ( .I(n6188), .ZN(n5111) );
  CKND0BWP12T U3009 ( .I(n6096), .ZN(n6779) );
  TPOAI21D0BWP12T U3010 ( .A1(n5109), .A2(n6779), .B(n5139), .ZN(n5110) );
  ND2D1BWP12T U3011 ( .A1(n5111), .A2(n5110), .ZN(n6191) );
  INVD1BWP12T U3012 ( .I(n5112), .ZN(n5114) );
  AOI21D1BWP12T U3013 ( .A1(n5115), .A2(n5114), .B(n5113), .ZN(n5117) );
  ND2D1BWP12T U3014 ( .A1(n5117), .A2(n5116), .ZN(n5928) );
  INVD1BWP12T U3015 ( .I(n6290), .ZN(n5124) );
  OAI21D1BWP12T U3016 ( .A1(n6534), .A2(n6565), .B(n5172), .ZN(n5123) );
  TPOAI22D0BWP12T U3017 ( .A1(n5613), .A2(n6306), .B1(n6251), .B2(n6297), .ZN(
        n5122) );
  OAI22D1BWP12T U3018 ( .A1(n5237), .A2(n5240), .B1(n5231), .B2(n5235), .ZN(
        n5120) );
  OAI22D1BWP12T U3019 ( .A1(n5236), .A2(n5238), .B1(n5239), .B2(n6760), .ZN(
        n5119) );
  NR2D1BWP12T U3020 ( .A1(n5120), .A2(n5119), .ZN(n6250) );
  OAI21D1BWP12T U3021 ( .A1(n6250), .A2(n6304), .B(n6565), .ZN(n5121) );
  AOI211D1BWP12T U3022 ( .A1(n6278), .A2(n6252), .B(n5122), .C(n5121), .ZN(
        n6318) );
  AOI211D1BWP12T U3023 ( .A1(n5124), .A2(n5123), .B(n6318), .C(n6560), .ZN(
        n6363) );
  AOI21D1BWP12T U3024 ( .A1(n6290), .A2(n6905), .B(n6736), .ZN(n5125) );
  NR2D1BWP12T U3025 ( .A1(n5125), .A2(n6318), .ZN(n5134) );
  ND2D1BWP12T U3026 ( .A1(n6818), .A2(n6786), .ZN(n5129) );
  ND2D1BWP12T U3027 ( .A1(n5129), .A2(n6844), .ZN(n6820) );
  CKND2D0BWP12T U3028 ( .A1(n6789), .A2(n6788), .ZN(n6787) );
  AOI22D0BWP12T U3029 ( .A1(n6464), .A2(n6879), .B1(n6499), .B2(n6745), .ZN(
        n5128) );
  TPND2D0BWP12T U3030 ( .A1(n5929), .A2(n6810), .ZN(n6092) );
  ND3D0BWP12T U3031 ( .A1(n6092), .A2(n6816), .A3(n5126), .ZN(n5127) );
  OAI211D1BWP12T U3032 ( .A1(n6787), .A2(n5129), .B(n5128), .C(n5127), .ZN(
        n5130) );
  AOI211D1BWP12T U3033 ( .A1(n5240), .A2(n6820), .B(n6753), .C(n5130), .ZN(
        n5132) );
  INVD1BWP12T U3034 ( .I(n6400), .ZN(n5474) );
  CKND2D1BWP12T U3035 ( .A1(n5474), .A2(n5507), .ZN(n5131) );
  AOI211D1BWP12T U3036 ( .A1(n6909), .A2(n6363), .B(n5134), .C(n5133), .ZN(
        n5135) );
  AOI21D1BWP12T U3037 ( .A1(n6728), .A2(n5983), .B(n5136), .ZN(n5141) );
  ND2D1BWP12T U3038 ( .A1(n5137), .A2(n5256), .ZN(n6135) );
  ND2D1BWP12T U3039 ( .A1(n6140), .A2(n6898), .ZN(n5140) );
  OAI211D4BWP12T U3040 ( .A1(n6902), .A2(n6040), .B(n5141), .C(n5140), .ZN(
        result[6]) );
  OAI21D1BWP12T U3041 ( .A1(n6013), .A2(n5143), .B(n5142), .ZN(n5148) );
  INVD1BWP12T U3042 ( .I(n5144), .ZN(n5146) );
  ND2D1BWP12T U3043 ( .A1(n5146), .A2(n5145), .ZN(n5147) );
  XNR2D1BWP12T U3044 ( .A1(n5148), .A2(n5147), .ZN(n6046) );
  CKND0BWP12T U3045 ( .I(n5602), .ZN(n5150) );
  INVD1BWP12T U3046 ( .I(n5149), .ZN(n5153) );
  NR2D1BWP12T U3047 ( .A1(n5150), .A2(n5153), .ZN(n5152) );
  INVD1BWP12T U3048 ( .I(n5151), .ZN(n5157) );
  XOR2XD1BWP12T U3049 ( .A1(n5152), .A2(n5157), .Z(n6145) );
  XOR2XD0BWP12T U3050 ( .A1(n5155), .A2(n5157), .Z(n5950) );
  ND2XD0BWP12T U3051 ( .A1(n5156), .A2(n6706), .ZN(n5564) );
  CKND0BWP12T U3052 ( .I(n6112), .ZN(n5580) );
  OAI21D0BWP12T U3053 ( .A1(n5564), .A2(n5580), .B(n5581), .ZN(n5158) );
  AOI21D0BWP12T U3054 ( .A1(n5158), .A2(n5157), .B(n5607), .ZN(n6199) );
  OAI21D1BWP12T U3055 ( .A1(n6714), .A2(n6862), .B(n6844), .ZN(n6699) );
  TPNR2D0BWP12T U3056 ( .A1(n5589), .A2(n6862), .ZN(n5159) );
  AOI211XD0BWP12T U3057 ( .A1(n6879), .A2(b[13]), .B(n6699), .C(n5159), .ZN(
        n5161) );
  CKND2D1BWP12T U3058 ( .A1(n5590), .A2(n5589), .ZN(n5160) );
  CKND2D1BWP12T U3059 ( .A1(n6323), .A2(n5575), .ZN(n6839) );
  OAI22D0BWP12T U3060 ( .A1(n6275), .A2(n6308), .B1(n6270), .B2(n6297), .ZN(
        n5164) );
  OAI21D1BWP12T U3061 ( .A1(n6274), .A2(n6306), .B(n6565), .ZN(n5163) );
  NR2D1BWP12T U3062 ( .A1(n6266), .A2(n6304), .ZN(n5162) );
  NR3D1BWP12T U3063 ( .A1(n5164), .A2(n5163), .A3(n5162), .ZN(n5170) );
  RCAOI21D0BWP12T U3064 ( .A1(n6573), .A2(n6839), .B(n5170), .ZN(n6384) );
  OAI22D0BWP12T U3065 ( .A1(n6263), .A2(n6530), .B1(n5165), .B2(n5677), .ZN(
        n5168) );
  NR2D0BWP12T U3066 ( .A1(n5166), .A2(n6534), .ZN(n5167) );
  AOI211D1BWP12T U3067 ( .A1(n6552), .A2(n5178), .B(n5168), .C(n5167), .ZN(
        n6539) );
  INVD1BWP12T U3068 ( .I(n6566), .ZN(n6513) );
  MUX2D1BWP12T U3069 ( .I0(a[31]), .I1(n5169), .S(n6553), .Z(n6352) );
  INVD0BWP12T U3070 ( .I(n5170), .ZN(n5171) );
  ND2D0BWP12T U3071 ( .A1(n6540), .A2(n6353), .ZN(n5207) );
  OAI211D1BWP12T U3072 ( .A1(n5172), .A2(n6352), .B(n5171), .C(n5207), .ZN(
        n6354) );
  NR2D1BWP12T U3073 ( .A1(n6409), .A2(n5176), .ZN(n5182) );
  OAI22D1BWP12T U3074 ( .A1(n5178), .A2(n6407), .B1(n6408), .B2(n5177), .ZN(
        n5181) );
  NR2D0BWP12T U3075 ( .A1(n6410), .A2(n5179), .ZN(n5180) );
  NR3D1BWP12T U3076 ( .A1(n5182), .A2(n5181), .A3(n5180), .ZN(n6437) );
  CKND0BWP12T U3077 ( .I(n6437), .ZN(n5187) );
  CKND1BWP12T U3078 ( .I(n5183), .ZN(n6500) );
  AOI22D0BWP12T U3079 ( .A1(n6500), .A2(n6745), .B1(n5606), .B2(n6747), .ZN(
        n5184) );
  OAI21D0BWP12T U3080 ( .A1(n5185), .A2(n6874), .B(n5184), .ZN(n5186) );
  AOI211XD0BWP12T U3081 ( .A1(n5187), .A2(n5507), .B(n6753), .C(n5186), .ZN(
        n5188) );
  OAI21D0BWP12T U3082 ( .A1(n6792), .A2(n5719), .B(n5188), .ZN(n5189) );
  AO211D1BWP12T U3083 ( .A1(n6384), .A2(n6905), .B(n5190), .C(n5189), .Z(n5191) );
  CKXOR2D1BWP12T U3084 ( .A1(n5195), .A2(n5200), .Z(n5985) );
  INVD1BWP12T U3085 ( .I(n5985), .ZN(n5220) );
  INVD1BWP12T U3086 ( .I(n5196), .ZN(n5197) );
  XOR2D1BWP12T U3087 ( .A1(n5197), .A2(n5200), .Z(n6141) );
  NR2D1BWP12T U3088 ( .A1(n6141), .A2(n6836), .ZN(n5219) );
  CKND2D0BWP12T U3089 ( .A1(n5198), .A2(n6093), .ZN(n5201) );
  AOI21D1BWP12T U3090 ( .A1(n5201), .A2(n5200), .B(n5199), .ZN(n6195) );
  OAI21D1BWP12T U3091 ( .A1(n5204), .A2(n5203), .B(n5202), .ZN(n5937) );
  OAI22D0BWP12T U3092 ( .A1(n6266), .A2(n6297), .B1(n6270), .B2(n6308), .ZN(
        n5206) );
  OAI21D1BWP12T U3093 ( .A1(n6275), .A2(n6306), .B(n6565), .ZN(n5205) );
  AOI211D1BWP12T U3094 ( .A1(n5575), .A2(n6273), .B(n5206), .C(n5205), .ZN(
        n6315) );
  INVD1BWP12T U3095 ( .I(n5207), .ZN(n5208) );
  AOI211D1BWP12T U3096 ( .A1(n6364), .A2(n5209), .B(n6315), .C(n5208), .ZN(
        n6362) );
  OAI21D0BWP12T U3097 ( .A1(b[9]), .A2(n6882), .B(n6874), .ZN(n5212) );
  OAI22D0BWP12T U3098 ( .A1(n5210), .A2(n6813), .B1(n6111), .B2(n6880), .ZN(
        n5211) );
  AOI211XD0BWP12T U3099 ( .A1(n5213), .A2(n5212), .B(n6753), .C(n5211), .ZN(
        n5214) );
  AOI211D1BWP12T U3100 ( .A1(n6728), .A2(n5220), .B(n5219), .C(n5218), .ZN(
        n5221) );
  INVD1BWP12T U3101 ( .I(n5222), .ZN(n5225) );
  XOR3D1BWP12T U3102 ( .A1(n5225), .A2(n5224), .A3(n5223), .Z(n6038) );
  XOR2XD0BWP12T U3103 ( .A1(n5228), .A2(n5274), .Z(n5982) );
  OAI22D1BWP12T U3104 ( .A1(n5237), .A2(n6760), .B1(n6708), .B2(n5235), .ZN(
        n5234) );
  OAI22D1BWP12T U3105 ( .A1(n5232), .A2(n5239), .B1(n5238), .B2(n5231), .ZN(
        n5233) );
  NR2D1BWP12T U3106 ( .A1(n5234), .A2(n5233), .ZN(n6305) );
  OAI22D1BWP12T U3107 ( .A1(n5237), .A2(n5253), .B1(n5236), .B2(n5235), .ZN(
        n5242) );
  TPOAI22D0BWP12T U3108 ( .A1(n5240), .A2(n5239), .B1(n5238), .B2(n6788), .ZN(
        n5241) );
  NR2D1BWP12T U3109 ( .A1(n5242), .A2(n5241), .ZN(n5729) );
  OAI22D1BWP12T U3110 ( .A1(n6305), .A2(n6297), .B1(n5729), .B2(n6304), .ZN(
        n5244) );
  OAI21D1BWP12T U3111 ( .A1(n6309), .A2(n6306), .B(n6565), .ZN(n5243) );
  AOI211D1BWP12T U3112 ( .A1(n6278), .A2(n6312), .B(n5244), .C(n5243), .ZN(
        n6314) );
  INVD1BWP12T U3113 ( .I(n6307), .ZN(n5246) );
  AO222D1BWP12T U3114 ( .A1(n5246), .A2(n5575), .B1(n6278), .B2(n6322), .C1(
        n6313), .C2(n5245), .Z(n6280) );
  AOI21D1BWP12T U3115 ( .A1(n6280), .A2(n6905), .B(n6736), .ZN(n5265) );
  CKND2D1BWP12T U3116 ( .A1(n6488), .A2(n6556), .ZN(n5251) );
  OAI21D1BWP12T U3117 ( .A1(n5250), .A2(n5247), .B(n5251), .ZN(n5248) );
  MUX2D1BWP12T U3118 ( .I0(n5249), .I1(n5248), .S(n6533), .Z(n5577) );
  ND2D1BWP12T U3119 ( .A1(n6873), .A2(n5577), .ZN(n5264) );
  INVD1BWP12T U3120 ( .I(n5571), .ZN(n6382) );
  AOI31D1BWP12T U3121 ( .A1(n5762), .A2(n6887), .A3(n5254), .B(n5253), .ZN(
        n5261) );
  OAI22D0BWP12T U3122 ( .A1(n5255), .A2(n6882), .B1(n6097), .B2(n6704), .ZN(
        n5258) );
  OAI22D1BWP12T U3123 ( .A1(n5256), .A2(n6813), .B1(n6249), .B2(n6844), .ZN(
        n5257) );
  AOI211D0BWP12T U3124 ( .A1(n5509), .A2(n5259), .B(n5258), .C(n5257), .ZN(
        n5260) );
  OAI31D0BWP12T U3125 ( .A1(n6789), .A2(n5261), .A3(n6862), .B(n5260), .ZN(
        n5262) );
  AOI211D1BWP12T U3126 ( .A1(n6382), .A2(n5507), .B(n6753), .C(n5262), .ZN(
        n5263) );
  OAI211D1BWP12T U3127 ( .A1(n6314), .A2(n5265), .B(n5264), .C(n5263), .ZN(
        n5270) );
  INVD1BWP12T U3128 ( .I(n5266), .ZN(n6179) );
  XNR2D1BWP12T U3129 ( .A1(n5268), .A2(n5274), .ZN(n6185) );
  AOI211D1BWP12T U3130 ( .A1(n6728), .A2(n5982), .B(n5270), .C(n5269), .ZN(
        n5276) );
  TPNR2D0BWP12T U3131 ( .A1(n6353), .A2(n6306), .ZN(n5510) );
  OAI21D1BWP12T U3132 ( .A1(n6280), .A2(n5510), .B(n6355), .ZN(n5271) );
  AOI21D1BWP12T U3133 ( .A1(n5271), .A2(n6584), .B(n6314), .ZN(n6330) );
  AOI21D1BWP12T U3134 ( .A1(n5272), .A2(n5273), .B(n5274), .ZN(n5938) );
  AOI31D1BWP12T U3135 ( .A1(n5274), .A2(n5273), .A3(n5272), .B(n5938), .ZN(
        n5936) );
  AOI22D1BWP12T U3136 ( .A1(n6330), .A2(n6909), .B1(n5936), .B2(n6833), .ZN(
        n5275) );
  OA211D1BWP12T U3137 ( .A1(n6139), .A2(n6836), .B(n5276), .C(n5275), .Z(n5277) );
  OAI21D1BWP12T U3138 ( .A1(n6038), .A2(n6902), .B(n5277), .ZN(result[4]) );
  OAI21D1BWP12T U3139 ( .A1(n5278), .A2(n6489), .B(n5321), .ZN(n6161) );
  ND2D1BWP12T U3140 ( .A1(n6084), .A2(n6834), .ZN(n5326) );
  AOI21D0BWP12T U3141 ( .A1(a[28]), .A2(n6220), .B(n6224), .ZN(n6221) );
  NR2D1BWP12T U3142 ( .A1(n6217), .A2(n6794), .ZN(n5319) );
  NR2D1BWP12T U3143 ( .A1(n5282), .A2(n6304), .ZN(n5576) );
  INVD1BWP12T U3144 ( .I(n5576), .ZN(n6342) );
  NR2D1BWP12T U3145 ( .A1(n6409), .A2(n5299), .ZN(n5285) );
  OAI22D1BWP12T U3146 ( .A1(n6408), .A2(n5297), .B1(n6407), .B2(n5298), .ZN(
        n5284) );
  NR2D0BWP12T U3147 ( .A1(n6410), .A2(n5675), .ZN(n5283) );
  NR3D1BWP12T U3148 ( .A1(n5285), .A2(n5284), .A3(n5283), .ZN(n6398) );
  NR2D0BWP12T U3149 ( .A1(n6410), .A2(n5291), .ZN(n5287) );
  OAI22D1BWP12T U3150 ( .A1(n6408), .A2(n5683), .B1(n6407), .B2(n5680), .ZN(
        n5286) );
  RCAOI211D0BWP12T U3151 ( .A1(n5289), .A2(n5288), .B(n5287), .C(n5286), .ZN(
        n5290) );
  OAI222D1BWP12T U3152 ( .A1(n5441), .A2(n5571), .B1(n6417), .B2(n6398), .C1(
        n6439), .C2(n5290), .ZN(n6388) );
  AOI22D0BWP12T U3153 ( .A1(n6556), .A2(n5681), .B1(n5291), .B2(n6553), .ZN(
        n5293) );
  AOI22D0BWP12T U3154 ( .A1(n6552), .A2(n5680), .B1(n5683), .B2(n6549), .ZN(
        n5292) );
  CKND2D1BWP12T U3155 ( .A1(n5293), .A2(n5292), .ZN(n5296) );
  AOI22D0BWP12T U3156 ( .A1(n6552), .A2(n5674), .B1(n5673), .B2(n6556), .ZN(
        n5295) );
  AOI22D0BWP12T U3157 ( .A1(n6553), .A2(n5682), .B1(n5676), .B2(n6549), .ZN(
        n5294) );
  ND2D1BWP12T U3158 ( .A1(n5295), .A2(n5294), .ZN(n5511) );
  AOI22D0BWP12T U3159 ( .A1(n6578), .A2(n5296), .B1(n5511), .B2(n6562), .ZN(
        n5304) );
  AOI22D0BWP12T U3160 ( .A1(n6552), .A2(n5298), .B1(n5297), .B2(n6549), .ZN(
        n5301) );
  AOI22D0BWP12T U3161 ( .A1(n6556), .A2(n5299), .B1(n5675), .B2(n6553), .ZN(
        n5300) );
  ND2D1BWP12T U3162 ( .A1(n5301), .A2(n5300), .ZN(n6514) );
  AOI21D0BWP12T U3163 ( .A1(n6514), .A2(n5302), .B(n6560), .ZN(n5303) );
  OAI211D1BWP12T U3164 ( .A1(n5305), .A2(n5577), .B(n5304), .C(n5303), .ZN(
        n6570) );
  MAOI22D0BWP12T U3165 ( .A1(n6857), .A2(n6388), .B1(n6570), .B2(n6680), .ZN(
        n5317) );
  TPND2D0BWP12T U3166 ( .A1(n5660), .A2(n5306), .ZN(n5309) );
  CKND0BWP12T U3167 ( .I(n5674), .ZN(n5307) );
  AOI22D1BWP12T U3168 ( .A1(n5307), .A2(n5662), .B1(n5661), .B2(n5658), .ZN(
        n5308) );
  OAI211D1BWP12T U3169 ( .A1(n6409), .A2(n5673), .B(n5309), .C(n5308), .ZN(
        n6394) );
  TPOAI21D0BWP12T U3170 ( .A1(n5310), .A2(n6744), .B(n6621), .ZN(n5312) );
  OAI22D0BWP12T U3171 ( .A1(n5312), .A2(n5311), .B1(n6480), .B2(n6882), .ZN(
        n5314) );
  OAI22D0BWP12T U3172 ( .A1(n6113), .A2(n6880), .B1(a[28]), .B2(n6844), .ZN(
        n5313) );
  AO211D1BWP12T U3173 ( .A1(n6358), .A2(n6909), .B(n5314), .C(n5313), .Z(n5315) );
  AOI211D1BWP12T U3174 ( .A1(n6394), .A2(n5546), .B(n6661), .C(n5315), .ZN(
        n5316) );
  OAI211D1BWP12T U3175 ( .A1(n6666), .A2(n6342), .B(n5317), .C(n5316), .ZN(
        n5318) );
  AOI211D1BWP12T U3176 ( .A1(n6786), .A2(n6221), .B(n5319), .C(n5318), .ZN(
        n5323) );
  AO21D1BWP12T U3177 ( .A1(n5321), .A2(n5320), .B(n5968), .Z(n6000) );
  ND2D1BWP12T U3178 ( .A1(n6000), .A2(n6728), .ZN(n5322) );
  OAI211D1BWP12T U3179 ( .A1(n6836), .A2(n6165), .B(n5323), .C(n5322), .ZN(
        n5324) );
  AOI21D1BWP12T U3180 ( .A1(n5967), .A2(n6833), .B(n5324), .ZN(n5325) );
  OAI211D2BWP12T U3181 ( .A1(n6161), .A2(n6836), .B(n5326), .C(n5325), .ZN(
        result[28]) );
  CKND2D1BWP12T U3182 ( .A1(n5419), .A2(a[30]), .ZN(n5420) );
  ND2D1BWP12T U3183 ( .A1(n5327), .A2(n5420), .ZN(n5906) );
  IND2XD1BWP12T U3184 ( .A1(b[31]), .B1(a[31]), .ZN(n6476) );
  XNR2D1BWP12T U3185 ( .A1(n5906), .A2(n6612), .ZN(n6002) );
  CKND2D1BWP12T U3186 ( .A1(n6081), .A2(n5332), .ZN(n5334) );
  NR2D1BWP12T U3187 ( .A1(n5334), .A2(n6075), .ZN(n5336) );
  CKND2D1BWP12T U3188 ( .A1(n5328), .A2(n5336), .ZN(n5340) );
  INVD1BWP12T U3189 ( .I(n5329), .ZN(n5330) );
  TPAOI21D0BWP12T U3190 ( .A1(n5332), .A2(n5331), .B(n5330), .ZN(n5333) );
  TPOAI21D0BWP12T U3191 ( .A1(n5334), .A2(n6074), .B(n5333), .ZN(n5335) );
  TPAOI21D0BWP12T U3192 ( .A1(n5337), .A2(n5336), .B(n5335), .ZN(n5338) );
  OAI21D1BWP12T U3193 ( .A1(n5340), .A2(n5339), .B(n5338), .ZN(n5901) );
  FA1D0BWP12T U3194 ( .A(n5343), .B(n5342), .CI(n5341), .CO(n5344), .S(n4786)
         );
  INVD1BWP12T U3195 ( .I(n5344), .ZN(n5414) );
  INVD0BWP12T U3196 ( .I(n5345), .ZN(n5346) );
  MAOI222D1BWP12T U3197 ( .A(n5348), .B(n5347), .C(n5346), .ZN(n5753) );
  INVD1BWP12T U3198 ( .I(n5349), .ZN(n5353) );
  INVD0BWP12T U3199 ( .I(n5350), .ZN(n5352) );
  MAOI222D1BWP12T U3200 ( .A(n5353), .B(n5352), .C(n5351), .ZN(n5757) );
  FA1D0BWP12T U3201 ( .A(n5356), .B(n5355), .CI(n5354), .CO(n5756), .S(n5345)
         );
  ND2D0BWP12T U3202 ( .A1(a[30]), .A2(a[29]), .ZN(n5366) );
  XNR2D1BWP12T U3203 ( .A1(n5360), .A2(b[31]), .ZN(n5763) );
  TPOAI22D0BWP12T U3204 ( .A1(n5763), .A2(n5362), .B1(b[30]), .B2(n5361), .ZN(
        n5852) );
  XOR2XD1BWP12T U3205 ( .A1(n5853), .A2(n5852), .Z(n5885) );
  MAOI222D1BWP12T U3206 ( .A(n5365), .B(n5364), .C(n5363), .ZN(n5887) );
  ND2D0BWP12T U3207 ( .A1(n6223), .A2(a[31]), .ZN(n5367) );
  OAI22D1BWP12T U3208 ( .A1(n5367), .A2(a[30]), .B1(n5366), .B2(a[31]), .ZN(
        n5764) );
  CKXOR2D1BWP12T U3209 ( .A1(a[31]), .A2(n5612), .Z(n5765) );
  MUX2ND0BWP12T U3210 ( .I0(n5811), .I1(n5810), .S(b[29]), .ZN(n5369) );
  MUX2ND0BWP12T U3211 ( .I0(n5813), .I1(n5812), .S(b[28]), .ZN(n5368) );
  NR2D1BWP12T U3212 ( .A1(n5369), .A2(n5368), .ZN(n5828) );
  XNR3D1BWP12T U3213 ( .A1(n5826), .A2(n5828), .A3(n5827), .ZN(n5886) );
  FA1D0BWP12T U3214 ( .A(n5374), .B(n5373), .CI(n5372), .CO(n5894), .S(n5408)
         );
  INVD0BWP12T U3215 ( .I(n5375), .ZN(n5376) );
  MAOI222D1BWP12T U3216 ( .A(n5378), .B(n5377), .C(n5376), .ZN(n5893) );
  XNR2XD1BWP12T U3217 ( .A1(a[25]), .A2(n5379), .ZN(n5842) );
  TPOAI22D0BWP12T U3218 ( .A1(n5382), .A2(n5381), .B1(n5380), .B2(n5842), .ZN(
        n5799) );
  MAOI222D1BWP12T U3219 ( .A(n5385), .B(n5384), .C(n5383), .ZN(n5801) );
  XOR2D1BWP12T U3220 ( .A1(a[29]), .A2(n6334), .Z(n5850) );
  AOI22D1BWP12T U3221 ( .A1(n5851), .A2(n5386), .B1(n5849), .B2(n5850), .ZN(
        n5772) );
  CKND0BWP12T U3222 ( .I(n5387), .ZN(n5868) );
  CKND0BWP12T U3223 ( .I(n5388), .ZN(n5389) );
  XOR2D1BWP12T U3224 ( .A1(a[27]), .A2(n6782), .Z(n5867) );
  AOI22D1BWP12T U3225 ( .A1(n5868), .A2(n5389), .B1(n5866), .B2(n5867), .ZN(
        n5774) );
  MUX2ND0BWP12T U3226 ( .I0(n5776), .I1(n5775), .S(b[21]), .ZN(n5391) );
  MUX2ND0BWP12T U3227 ( .I0(n5778), .I1(n5777), .S(b[20]), .ZN(n5390) );
  NR2D1BWP12T U3228 ( .A1(n5391), .A2(n5390), .ZN(n5773) );
  XNR3D1BWP12T U3229 ( .A1(n5772), .A2(n5774), .A3(n5773), .ZN(n5800) );
  XOR3D1BWP12T U3230 ( .A1(n5786), .A2(n5788), .A3(n5787), .Z(n5783) );
  INVD0BWP12T U3231 ( .I(n5398), .ZN(n5402) );
  INVD0BWP12T U3232 ( .I(n5399), .ZN(n5401) );
  MAOI222D1BWP12T U3233 ( .A(n5402), .B(n5401), .C(n5400), .ZN(n5794) );
  CKND0BWP12T U3234 ( .I(n5403), .ZN(n5404) );
  XOR2D1BWP12T U3235 ( .A1(a[23]), .A2(b[9]), .Z(n5808) );
  AOI22D1BWP12T U3236 ( .A1(n5809), .A2(n5404), .B1(n5807), .B2(n5808), .ZN(
        n5829) );
  XOR3D1BWP12T U3237 ( .A1(n5792), .A2(n5794), .A3(n5791), .Z(n5784) );
  XOR3D1BWP12T U3238 ( .A1(n5785), .A2(n5783), .A3(n5784), .Z(n5892) );
  INVD1BWP12T U3239 ( .I(n5412), .ZN(n5413) );
  OR2XD1BWP12T U3240 ( .A1(n5414), .A2(n5413), .Z(n5900) );
  ND2D1BWP12T U3241 ( .A1(n5414), .A2(n5413), .ZN(n5899) );
  ND2D1BWP12T U3242 ( .A1(n6608), .A2(n6834), .ZN(n5453) );
  CKND2D0BWP12T U3243 ( .A1(n5417), .A2(n5908), .ZN(n5415) );
  TPNR2D0BWP12T U3244 ( .A1(n6612), .A2(n5415), .ZN(n5428) );
  TPND2D0BWP12T U3245 ( .A1(n6612), .A2(n6110), .ZN(n5430) );
  TPNR2D0BWP12T U3246 ( .A1(n5922), .A2(n5430), .ZN(n5418) );
  INVD1BWP12T U3247 ( .I(n6612), .ZN(n6455) );
  INVD1BWP12T U3248 ( .I(n6110), .ZN(n5907) );
  AOI211D1BWP12T U3249 ( .A1(n5922), .A2(n5428), .B(n5418), .C(n5429), .ZN(
        n5966) );
  NR2D1BWP12T U3250 ( .A1(n5419), .A2(a[30]), .ZN(n6451) );
  CKND2D1BWP12T U3251 ( .A1(n5420), .A2(n6845), .ZN(n6505) );
  CKND0BWP12T U3252 ( .I(n6505), .ZN(n5421) );
  OAI21D0BWP12T U3253 ( .A1(n6451), .A2(n5421), .B(n6455), .ZN(n5427) );
  INVD1BWP12T U3254 ( .I(n6451), .ZN(n5903) );
  OAI211D0BWP12T U3255 ( .A1(n6449), .A2(n6505), .B(n6612), .C(n5903), .ZN(
        n5426) );
  NR3D1BWP12T U3256 ( .A1(n6165), .A2(n6455), .A3(n6505), .ZN(n5425) );
  NR4D0BWP12T U3257 ( .A1(n5423), .A2(n6612), .A3(n6451), .A4(n5422), .ZN(
        n5424) );
  AOI211D1BWP12T U3258 ( .A1(n5427), .A2(n5426), .B(n5425), .C(n5424), .ZN(
        n6163) );
  NR2D1BWP12T U3259 ( .A1(n6163), .A2(n6836), .ZN(n5451) );
  NR2XD0BWP12T U3260 ( .A1(n6840), .A2(n5533), .ZN(n5433) );
  TPNR2D0BWP12T U3261 ( .A1(b[31]), .A2(op[2]), .ZN(n5431) );
  TPOAI22D0BWP12T U3262 ( .A1(n5431), .A2(n6106), .B1(b[31]), .B2(n6683), .ZN(
        n5432) );
  AOI211D1BWP12T U3263 ( .A1(n6597), .A2(n6786), .B(n5433), .C(n5432), .ZN(
        n5448) );
  NR2D1BWP12T U3264 ( .A1(n6409), .A2(n6551), .ZN(n5440) );
  OAI22D1BWP12T U3265 ( .A1(n6408), .A2(n6555), .B1(n6407), .B2(n6554), .ZN(
        n5439) );
  AOI211D0BWP12T U3266 ( .A1(n5660), .A2(a[30]), .B(n5440), .C(n5439), .ZN(
        n5442) );
  OA222D1BWP12T U3267 ( .A1(n6439), .A2(n5442), .B1(n5441), .B2(n6817), .C1(
        n6417), .C2(n6401), .Z(n6441) );
  NR2D1BWP12T U3268 ( .A1(n6441), .A2(n6716), .ZN(n5446) );
  AOI22D0BWP12T U3269 ( .A1(n6353), .A2(n6783), .B1(n6744), .B2(b[31]), .ZN(
        n5444) );
  TPND2D0BWP12T U3270 ( .A1(n6455), .A2(n6879), .ZN(n5443) );
  OAI211D0BWP12T U3271 ( .A1(n5719), .A2(n6397), .B(n5444), .C(n5443), .ZN(
        n5445) );
  AOI211D1BWP12T U3272 ( .A1(n6855), .A2(n6547), .B(n5446), .C(n5445), .ZN(
        n5447) );
  OA211D1BWP12T U3273 ( .A1(n5448), .A2(n6353), .B(n5918), .C(n5447), .Z(n5449) );
  OAI21D1BWP12T U3274 ( .A1(n6218), .A2(n6794), .B(n5449), .ZN(n5450) );
  AOI211D1BWP12T U3275 ( .A1(n5966), .A2(n6833), .B(n5451), .C(n5450), .ZN(
        n5452) );
  OAI211D1BWP12T U3276 ( .A1(n6002), .A2(n6890), .B(n5453), .C(n5452), .ZN(
        result[31]) );
  BUFFXD0BWP12T U3277 ( .I(result[31]), .Z(n) );
  INVD1BWP12T U3278 ( .I(n5454), .ZN(n5456) );
  ND2D1BWP12T U3279 ( .A1(n5456), .A2(n5455), .ZN(n5458) );
  XOR2XD1BWP12T U3280 ( .A1(n5458), .A2(n5457), .Z(n6068) );
  INVD1BWP12T U3281 ( .I(n5459), .ZN(n5502) );
  NR2D1BWP12T U3282 ( .A1(n5502), .A2(n5515), .ZN(n6615) );
  CKND2D0BWP12T U3283 ( .A1(n6618), .A2(n5460), .ZN(n5461) );
  NR2D1BWP12T U3284 ( .A1(n6615), .A2(n5461), .ZN(n5992) );
  INVD1BWP12T U3285 ( .I(n5992), .ZN(n6616) );
  TPAOI31D0BWP12T U3286 ( .A1(n6616), .A2(n5489), .A3(n5463), .B(n5462), .ZN(
        n5995) );
  INVD0BWP12T U3287 ( .I(n5464), .ZN(n5465) );
  XNR2XD1BWP12T U3288 ( .A1(n5465), .A2(n5489), .ZN(n6152) );
  OAI211D1BWP12T U3289 ( .A1(n6751), .A2(n5467), .B(n5482), .C(n6844), .ZN(
        n5486) );
  NR2D1BWP12T U3290 ( .A1(n6209), .A2(n6794), .ZN(n5485) );
  CKND0BWP12T U3291 ( .I(n6634), .ZN(n5483) );
  NR2D1BWP12T U3292 ( .A1(n6417), .A2(n6716), .ZN(n5506) );
  AOI211D0BWP12T U3293 ( .A1(n5467), .A2(n6810), .B(n5487), .C(n6704), .ZN(
        n5468) );
  AOI211D0BWP12T U3294 ( .A1(n6496), .A2(n6745), .B(n6661), .C(n5468), .ZN(
        n5469) );
  TPOAI31D0BWP12T U3295 ( .A1(n6553), .A2(n5667), .A3(n5470), .B(n5469), .ZN(
        n5473) );
  OAI22D1BWP12T U3296 ( .A1(n5623), .A2(n5719), .B1(n5471), .B2(n6892), .ZN(
        n5472) );
  AOI211D1BWP12T U3297 ( .A1(n5506), .A2(n5474), .B(n5473), .C(n5472), .ZN(
        n5481) );
  CKND2D0BWP12T U3298 ( .A1(n5475), .A2(n6578), .ZN(n5476) );
  INVD1BWP12T U3299 ( .I(n6540), .ZN(n6575) );
  OAI211D0BWP12T U3300 ( .A1(n5477), .A2(n6576), .B(n5476), .C(n6575), .ZN(
        n5478) );
  AOI21D0BWP12T U3301 ( .A1(n6573), .A2(n5624), .B(n5478), .ZN(n6546) );
  AOI22D1BWP12T U3302 ( .A1(n6546), .A2(n6855), .B1(n6290), .B2(n5479), .ZN(
        n5480) );
  OAI211D1BWP12T U3303 ( .A1(n5483), .A2(n5482), .B(n5481), .C(n5480), .ZN(
        n5484) );
  AOI211D1BWP12T U3304 ( .A1(n5487), .A2(n5486), .B(n5485), .C(n5484), .ZN(
        n5491) );
  CKND2D1BWP12T U3305 ( .A1(n5959), .A2(n6833), .ZN(n5490) );
  OAI211D1BWP12T U3306 ( .A1(n6836), .A2(n6152), .B(n5491), .C(n5490), .ZN(
        n5492) );
  AOI21D1BWP12T U3307 ( .A1(n5995), .A2(n6728), .B(n5492), .ZN(n5493) );
  IOA21D2BWP12T U3308 ( .A1(n6068), .A2(n6834), .B(n5493), .ZN(result[22]) );
  INVD1BWP12T U3309 ( .I(n5494), .ZN(n5497) );
  INVD1BWP12T U3310 ( .I(n5495), .ZN(n5496) );
  INVD1BWP12T U3311 ( .I(n5498), .ZN(n6062) );
  INVD1BWP12T U3312 ( .I(n6061), .ZN(n5499) );
  AOI21D1BWP12T U3313 ( .A1(n5515), .A2(n5502), .B(n6615), .ZN(n5993) );
  INVD1BWP12T U3314 ( .I(n5993), .ZN(n5520) );
  OAI31D0BWP12T U3315 ( .A1(n5504), .A2(n6656), .A3(n6124), .B(n5503), .ZN(
        n6151) );
  NR2D1BWP12T U3316 ( .A1(n6151), .A2(n6836), .ZN(n5519) );
  INVD1BWP12T U3317 ( .I(n5506), .ZN(n5720) );
  INVD1BWP12T U3318 ( .I(n6280), .ZN(n6344) );
  AOI21D1BWP12T U3319 ( .A1(n6514), .A2(n6334), .B(n6540), .ZN(n5513) );
  CKND2D0BWP12T U3320 ( .A1(n5511), .A2(n6578), .ZN(n5512) );
  OAI211D1BWP12T U3321 ( .A1(n5577), .A2(n6565), .B(n5513), .C(n5512), .ZN(
        n6528) );
  ND2D1BWP12T U3322 ( .A1(n6207), .A2(n6870), .ZN(n5516) );
  OAI211D1BWP12T U3323 ( .A1(n6894), .A2(n5955), .B(n5517), .C(n5516), .ZN(
        n5518) );
  AOI211D1BWP12T U3324 ( .A1(n5520), .A2(n6728), .B(n5519), .C(n5518), .ZN(
        n5521) );
  INVD1BWP12T U3325 ( .I(n5989), .ZN(n5554) );
  CKND1BWP12T U3326 ( .I(n5526), .ZN(n5527) );
  XOR2D1BWP12T U3327 ( .A1(n5527), .A2(n5530), .Z(n6147) );
  NR2D1BWP12T U3328 ( .A1(n6147), .A2(n6836), .ZN(n5553) );
  INVD0BWP12T U3329 ( .I(n6303), .ZN(n5535) );
  INVD0BWP12T U3330 ( .I(n5537), .ZN(n5531) );
  TPND2D0BWP12T U3331 ( .A1(n5531), .A2(n6562), .ZN(n5532) );
  OAI31D0BWP12T U3332 ( .A1(n6353), .A2(n6357), .A3(n5533), .B(n5532), .ZN(
        n5534) );
  RCAOI21D0BWP12T U3333 ( .A1(n6578), .A2(n5535), .B(n5534), .ZN(n6442) );
  INVD1BWP12T U3334 ( .I(n6442), .ZN(n6293) );
  MUX2ND0BWP12T U3335 ( .I0(n5611), .I1(n5724), .S(n6232), .ZN(n5550) );
  ND2D1BWP12T U3336 ( .A1(n6355), .A2(n6562), .ZN(n5536) );
  OAI22D1BWP12T U3337 ( .A1(n6303), .A2(n6351), .B1(n5537), .B2(n5536), .ZN(
        n6365) );
  CKND2D1BWP12T U3338 ( .A1(n6365), .A2(n6909), .ZN(n5548) );
  INVD0BWP12T U3339 ( .I(n6817), .ZN(n5545) );
  NR2D0BWP12T U3340 ( .A1(n6401), .A2(n6892), .ZN(n5544) );
  AOI21D0BWP12T U3341 ( .A1(n5538), .A2(n6879), .B(n6744), .ZN(n5541) );
  CKND0BWP12T U3342 ( .I(n6094), .ZN(n5539) );
  AOI22D0BWP12T U3343 ( .A1(n5539), .A2(n6747), .B1(n6482), .B2(n6745), .ZN(
        n5540) );
  OAI211D0BWP12T U3344 ( .A1(n5542), .A2(n5541), .B(n6686), .C(n5540), .ZN(
        n5543) );
  AOI211D1BWP12T U3345 ( .A1(n5546), .A2(n5545), .B(n5544), .C(n5543), .ZN(
        n5547) );
  RCAOI211D0BWP12T U3346 ( .A1(n6293), .A2(n6905), .B(n5550), .C(n5549), .ZN(
        n5551) );
  INVD1BWP12T U3347 ( .I(n5555), .ZN(n5558) );
  INVD1BWP12T U3348 ( .I(n5556), .ZN(n5557) );
  OAI21D1BWP12T U3349 ( .A1(n6013), .A2(n5558), .B(n5557), .ZN(n5562) );
  ND2D1BWP12T U3350 ( .A1(n5560), .A2(n5559), .ZN(n5561) );
  XNR2D1BWP12T U3351 ( .A1(n5562), .A2(n5561), .ZN(n6045) );
  XNR2XD1BWP12T U3352 ( .A1(n5563), .A2(n5567), .ZN(n5987) );
  XNR2XD1BWP12T U3353 ( .A1(n5564), .A2(n5567), .ZN(n6196) );
  OAI21D1BWP12T U3354 ( .A1(n5566), .A2(n5565), .B(n5602), .ZN(n6143) );
  ND2D1BWP12T U3355 ( .A1(n6143), .A2(n6898), .ZN(n5595) );
  XNR2D0BWP12T U3356 ( .A1(n5568), .A2(n5567), .ZN(n5945) );
  INVD0BWP12T U3357 ( .I(n6717), .ZN(n6426) );
  OAI22D0BWP12T U3358 ( .A1(n6307), .A2(n6308), .B1(n6309), .B2(n6297), .ZN(
        n5574) );
  OAI21D1BWP12T U3359 ( .A1(n5572), .A2(n6306), .B(n6565), .ZN(n5573) );
  AOI211D1BWP12T U3360 ( .A1(n5575), .A2(n6312), .B(n5574), .C(n5573), .ZN(
        n5584) );
  NR2D1BWP12T U3361 ( .A1(n5576), .A2(n6565), .ZN(n5586) );
  NR2D1BWP12T U3362 ( .A1(n5584), .A2(n5586), .ZN(n6292) );
  CKND1BWP12T U3363 ( .I(n5577), .ZN(n6522) );
  ND2D1BWP12T U3364 ( .A1(n5578), .A2(n6334), .ZN(n5625) );
  CKND2D0BWP12T U3365 ( .A1(n5589), .A2(n6879), .ZN(n5579) );
  RCAOI22D0BWP12T U3366 ( .A1(n5582), .A2(n5581), .B1(n5580), .B2(n6747), .ZN(
        n5583) );
  OA211D1BWP12T U3367 ( .A1(n6522), .A2(n5625), .B(n5583), .C(n6888), .Z(n5588) );
  AOI211D1BWP12T U3368 ( .A1(n5586), .A2(n5585), .B(n5584), .C(n6560), .ZN(
        n6366) );
  AOI22D1BWP12T U3369 ( .A1(n6366), .A2(n6909), .B1(n6292), .B2(n6676), .ZN(
        n5587) );
  MUX2ND0BWP12T U3370 ( .I0(n5590), .I1(n6699), .S(n5589), .ZN(n5591) );
  OAI211D1BWP12T U3371 ( .A1(n6443), .A2(n6716), .B(n5592), .C(n5591), .ZN(
        n5593) );
  AOI21D1BWP12T U3372 ( .A1(n6833), .A2(n5945), .B(n5593), .ZN(n5594) );
  OAI211D1BWP12T U3373 ( .A1(n6794), .A2(n6196), .B(n5595), .C(n5594), .ZN(
        n5596) );
  AOI21D1BWP12T U3374 ( .A1(n5987), .A2(n6728), .B(n5596), .ZN(n5597) );
  RCOAI21D1BWP12T U3375 ( .A1(n6045), .A2(n6902), .B(n5597), .ZN(result[12])
         );
  CKND0BWP12T U3376 ( .I(n5601), .ZN(n6448) );
  OA211D1BWP12T U3377 ( .A1(n5604), .A2(n5603), .B(n5972), .C(n6728), .Z(n5645) );
  NR2D1BWP12T U3378 ( .A1(n5607), .A2(n5606), .ZN(n5609) );
  XNR2D0BWP12T U3379 ( .A1(n5609), .A2(n5608), .ZN(n6201) );
  ND2D1BWP12T U3380 ( .A1(b[14]), .A2(n6879), .ZN(n5610) );
  AOI21D1BWP12T U3381 ( .A1(n5611), .A2(n5610), .B(a[14]), .ZN(n5642) );
  CKND2D1BWP12T U3382 ( .A1(n6319), .A2(n6573), .ZN(n6281) );
  CKND0BWP12T U3383 ( .I(n6281), .ZN(n5622) );
  OAI21D1BWP12T U3384 ( .A1(n6304), .A2(n5612), .B(a[31]), .ZN(n5621) );
  OAI22D0BWP12T U3385 ( .A1(n5614), .A2(n6308), .B1(n5613), .B2(n6297), .ZN(
        n5618) );
  CKND0BWP12T U3386 ( .I(n5615), .ZN(n5616) );
  OAI21D1BWP12T U3387 ( .A1(n5616), .A2(n6306), .B(n6565), .ZN(n5617) );
  NR2D1BWP12T U3388 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  OAI21D1BWP12T U3389 ( .A1(n5620), .A2(n6304), .B(n5619), .ZN(n6282) );
  INVD1BWP12T U3390 ( .I(n6282), .ZN(n5638) );
  AOI211D1BWP12T U3391 ( .A1(n5622), .A2(n5621), .B(n5638), .C(n6560), .ZN(
        n6329) );
  OAI22D1BWP12T U3392 ( .A1(n5625), .A2(n5624), .B1(n5623), .B2(n6892), .ZN(
        n5633) );
  NR2D0BWP12T U3393 ( .A1(n6400), .A2(n5719), .ZN(n5632) );
  TPNR2D0BWP12T U3394 ( .A1(n5626), .A2(n6704), .ZN(n5627) );
  MUX2ND0BWP12T U3395 ( .I0(n6745), .I1(n5627), .S(b[14]), .ZN(n5630) );
  AOI21D0BWP12T U3396 ( .A1(n5630), .A2(n5629), .B(n5628), .ZN(n5631) );
  NR4D0BWP12T U3397 ( .A1(n5633), .A2(n5632), .A3(n6753), .A4(n5631), .ZN(
        n5634) );
  OAI31D0BWP12T U3398 ( .A1(n5636), .A2(n5635), .A3(n6862), .B(n5634), .ZN(
        n5640) );
  TPND2D0BWP12T U3399 ( .A1(n6905), .A2(n6281), .ZN(n5637) );
  AO211D1BWP12T U3400 ( .A1(n6909), .A2(n6329), .B(n5640), .C(n5639), .Z(n5641) );
  AOI211D1BWP12T U3401 ( .A1(n6201), .A2(n6870), .B(n5642), .C(n5641), .ZN(
        n5643) );
  OAI21D1BWP12T U3402 ( .A1(n5948), .A2(n6894), .B(n5643), .ZN(n5644) );
  AOI211D1BWP12T U3403 ( .A1(n6898), .A2(n6144), .B(n5645), .C(n5644), .ZN(
        n5646) );
  TPND2D0BWP12T U3404 ( .A1(n5649), .A2(n5652), .ZN(n6159) );
  AOI211D0BWP12T U3405 ( .A1(a[26]), .A2(n5654), .B(n5653), .C(n6862), .ZN(
        n5692) );
  CKND2D0BWP12T U3406 ( .A1(n5660), .A2(n5674), .ZN(n5657) );
  AOI22D0BWP12T U3407 ( .A1(n5661), .A2(n5675), .B1(n5655), .B2(n5673), .ZN(
        n5656) );
  OAI211D1BWP12T U3408 ( .A1(n5658), .A2(n6409), .B(n5657), .C(n5656), .ZN(
        n6378) );
  CKND2D1BWP12T U3409 ( .A1(n5668), .A2(n5667), .ZN(n6340) );
  MUX2ND0BWP12T U3410 ( .I0(n6844), .I1(n6874), .S(a[26]), .ZN(n5670) );
  OAI22D0BWP12T U3411 ( .A1(n6470), .A2(n6751), .B1(n6116), .B2(n6880), .ZN(
        n5669) );
  AOI211D0BWP12T U3412 ( .A1(n6503), .A2(n6745), .B(n5670), .C(n5669), .ZN(
        n5671) );
  OAI211D1BWP12T U3413 ( .A1(n6289), .A2(n6840), .B(n5671), .C(n6686), .ZN(
        n5672) );
  AOI21D1BWP12T U3414 ( .A1(n6688), .A2(n6340), .B(n5672), .ZN(n5690) );
  OAI22D0BWP12T U3415 ( .A1(n6534), .A2(n5674), .B1(n5673), .B2(n6533), .ZN(
        n5679) );
  OAI22D0BWP12T U3416 ( .A1(n5677), .A2(n5676), .B1(n5675), .B2(n6530), .ZN(
        n5678) );
  NR2D1BWP12T U3417 ( .A1(n5679), .A2(n5678), .ZN(n6525) );
  AOI22D0BWP12T U3418 ( .A1(n6552), .A2(n5681), .B1(n5680), .B2(n6553), .ZN(
        n5685) );
  AOI22D0BWP12T U3419 ( .A1(n6556), .A2(n5683), .B1(n5682), .B2(n6549), .ZN(
        n5684) );
  AOI21D1BWP12T U3420 ( .A1(n5685), .A2(n5684), .B(n6557), .ZN(n5686) );
  RCAOI211D0BWP12T U3421 ( .A1(n6562), .A2(n6525), .B(n5686), .C(n6560), .ZN(
        n5687) );
  OA21D1BWP12T U3422 ( .A1(n6565), .A2(n5688), .B(n5687), .Z(n6543) );
  ND2D1BWP12T U3423 ( .A1(n6543), .A2(n6855), .ZN(n5689) );
  OAI211D1BWP12T U3424 ( .A1(n6716), .A2(n6434), .B(n5690), .C(n5689), .ZN(
        n5691) );
  AOI211D1BWP12T U3425 ( .A1(n6214), .A2(n6870), .B(n5692), .C(n5691), .ZN(
        n5699) );
  CKND0BWP12T U3426 ( .I(n5693), .ZN(n6469) );
  TPNR2D0BWP12T U3427 ( .A1(n5694), .A2(n6469), .ZN(n5696) );
  INVD1BWP12T U3428 ( .I(n5999), .ZN(n5695) );
  OAI211D1BWP12T U3429 ( .A1(n5697), .A2(n5696), .B(n5695), .C(n6728), .ZN(
        n5698) );
  OAI211D1BWP12T U3430 ( .A1(n6894), .A2(n5961), .B(n5699), .C(n5698), .ZN(
        n5700) );
  AOI31D1BWP12T U3431 ( .A1(n6898), .A2(n6160), .A3(n6159), .B(n5700), .ZN(
        n5701) );
  XOR2XD0BWP12T U3432 ( .A1(n5702), .A2(n5705), .Z(n5991) );
  XOR2XD0BWP12T U3433 ( .A1(n5703), .A2(n5705), .Z(n6148) );
  CKND1BWP12T U3434 ( .I(n6678), .ZN(n6647) );
  OAI21D1BWP12T U3435 ( .A1(n6647), .A2(n6862), .B(n6844), .ZN(n6679) );
  XOR2XD0BWP12T U3436 ( .A1(n5706), .A2(n5705), .Z(n6205) );
  NR2D1BWP12T U3437 ( .A1(n6205), .A2(n6794), .ZN(n5727) );
  CKND0BWP12T U3438 ( .I(n6518), .ZN(n5709) );
  ND2D1BWP12T U3439 ( .A1(n5707), .A2(n6334), .ZN(n5708) );
  OAI211D1BWP12T U3440 ( .A1(n5709), .A2(n6565), .B(n5708), .C(n6575), .ZN(
        n5710) );
  RCAOI21D0BWP12T U3441 ( .A1(n6578), .A2(n5711), .B(n5710), .ZN(n6579) );
  CKND2D1BWP12T U3442 ( .A1(n6579), .A2(n6855), .ZN(n5718) );
  NR2D0BWP12T U3443 ( .A1(n6399), .A2(n6892), .ZN(n5716) );
  AOI211D1BWP12T U3444 ( .A1(a[17]), .A2(n6874), .B(n5712), .C(n6751), .ZN(
        n5715) );
  OAI22D0BWP12T U3445 ( .A1(n5713), .A2(n6882), .B1(n6115), .B2(n6880), .ZN(
        n5714) );
  NR4D0BWP12T U3446 ( .A1(n5716), .A2(n6661), .A3(n5715), .A4(n5714), .ZN(
        n5717) );
  OAI211D1BWP12T U3447 ( .A1(n6840), .A2(n6317), .B(n5718), .C(n5717), .ZN(
        n5722) );
  OAI22D1BWP12T U3448 ( .A1(n5720), .A2(n6380), .B1(n6395), .B2(n5719), .ZN(
        n5721) );
  AOI211D1BWP12T U3449 ( .A1(n6688), .A2(n6341), .B(n5722), .C(n5721), .ZN(
        n5723) );
  OAI31D1BWP12T U3450 ( .A1(n6647), .A2(n5725), .A3(n5724), .B(n5723), .ZN(
        n5726) );
  NR2D1BWP12T U3451 ( .A1(n6343), .A2(n6565), .ZN(n6387) );
  OAI22D1BWP12T U3452 ( .A1(n5730), .A2(n6334), .B1(n5729), .B2(n6297), .ZN(
        n5734) );
  CKND2D1BWP12T U3453 ( .A1(n5731), .A2(n6479), .ZN(n5732) );
  OAI211D1BWP12T U3454 ( .A1(n6305), .A2(n6308), .B(n6519), .C(n5732), .ZN(
        n5733) );
  AOI211D1BWP12T U3455 ( .A1(n6254), .A2(n6312), .B(n5734), .C(n5733), .ZN(
        n6396) );
  OA21XD1BWP12T U3456 ( .A1(c_in), .A2(n6606), .B(n5735), .Z(n6183) );
  NR2D0BWP12T U3457 ( .A1(n6183), .A2(n6836), .ZN(n5745) );
  CKND0BWP12T U3458 ( .I(n6606), .ZN(n5743) );
  AOI22D0BWP12T U3459 ( .A1(n6488), .A2(n6745), .B1(n5736), .B2(op[1]), .ZN(
        n5742) );
  CKND2D0BWP12T U3460 ( .A1(n6902), .A2(n6880), .ZN(n5737) );
  AOI22D1BWP12T U3461 ( .A1(n6457), .A2(n6621), .B1(n5738), .B2(n5737), .ZN(
        n5741) );
  CKND2D0BWP12T U3462 ( .A1(n6862), .A2(n6874), .ZN(n5739) );
  MUX2ND0BWP12T U3463 ( .I0(n6783), .I1(n5739), .S(a[0]), .ZN(n5740) );
  OAI211D1BWP12T U3464 ( .A1(n5743), .A2(n5742), .B(n5741), .C(n5740), .ZN(
        n5744) );
  AOI211XD0BWP12T U3465 ( .A1(n6870), .A2(n6183), .B(n5745), .C(n5744), .ZN(
        n5746) );
  NR2D1BWP12T U3466 ( .A1(n6396), .A2(n6840), .ZN(n5747) );
  AOI211D1BWP12T U3467 ( .A1(n6387), .A2(n6905), .B(n5748), .C(n5747), .ZN(
        n5749) );
  OAI21D1BWP12T U3468 ( .A1(n6593), .A2(n6852), .B(n5749), .ZN(result[0]) );
  FA1D0BWP12T U3469 ( .A(n5757), .B(n5756), .CI(n5755), .CO(n5898), .S(n5754)
         );
  MAOI222D0BWP12T U3470 ( .A(n5785), .B(n5784), .C(n5783), .ZN(n5796) );
  CKND1BWP12T U3471 ( .I(n5786), .ZN(n5790) );
  INVD1BWP12T U3472 ( .I(n5787), .ZN(n5789) );
  INVD1BWP12T U3473 ( .I(n5791), .ZN(n5793) );
  MAOI222D1BWP12T U3474 ( .A(n5794), .B(n5793), .C(n5792), .ZN(n5795) );
  MAOI222D0BWP12T U3475 ( .A(n5801), .B(n5800), .C(n5799), .ZN(n5835) );
  MUX2ND0BWP12T U3476 ( .I0(n5811), .I1(n5810), .S(b[30]), .ZN(n5815) );
  MUX2ND0BWP12T U3477 ( .I0(n5813), .I1(n5812), .S(b[29]), .ZN(n5814) );
  NR2D1BWP12T U3478 ( .A1(n5815), .A2(n5814), .ZN(n5823) );
  MUX2ND0BWP12T U3479 ( .I0(n5817), .I1(n5816), .S(b[20]), .ZN(n5821) );
  MUX2NXD0BWP12T U3480 ( .I0(n5819), .I1(n5818), .S(b[19]), .ZN(n5820) );
  NR2D1BWP12T U3481 ( .A1(n5821), .A2(n5820), .ZN(n5822) );
  XOR4D1BWP12T U3482 ( .A1(n5825), .A2(n5824), .A3(n5823), .A4(n5822), .Z(
        n5834) );
  MAOI222D0BWP12T U3483 ( .A(n5828), .B(n5827), .C(n5826), .ZN(n5833) );
  MAOI222D0BWP12T U3484 ( .A(n5831), .B(n5830), .C(n5829), .ZN(n5832) );
  XNR4D1BWP12T U3485 ( .A1(n5835), .A2(n5834), .A3(n5833), .A4(n5832), .ZN(
        n5891) );
  MUX2ND0BWP12T U3486 ( .I0(n5837), .I1(n5836), .S(b[24]), .ZN(n5841) );
  MUX2ND0BWP12T U3487 ( .I0(n5839), .I1(n5838), .S(b[23]), .ZN(n5840) );
  NR2D1BWP12T U3488 ( .A1(n5841), .A2(n5840), .ZN(n5857) );
  CKND0BWP12T U3489 ( .I(n5842), .ZN(n5846) );
  XOR2XD0BWP12T U3490 ( .A1(a[25]), .A2(n5843), .Z(n5844) );
  AOI22D0BWP12T U3491 ( .A1(n5847), .A2(n5846), .B1(n5845), .B2(n5844), .ZN(
        n5856) );
  XOR2XD0BWP12T U3492 ( .A1(a[29]), .A2(n6573), .Z(n5848) );
  AOI22D0BWP12T U3493 ( .A1(n5851), .A2(n5850), .B1(n5849), .B2(n5848), .ZN(
        n5855) );
  CKND2D0BWP12T U3494 ( .A1(n5853), .A2(n5852), .ZN(n5854) );
  XNR4D1BWP12T U3495 ( .A1(n5857), .A2(n5856), .A3(n5855), .A4(n5854), .ZN(
        n5890) );
  MUX2ND0BWP12T U3496 ( .I0(n5859), .I1(n5858), .S(b[28]), .ZN(n5863) );
  MUX2ND0BWP12T U3497 ( .I0(n5861), .I1(n5860), .S(b[27]), .ZN(n5862) );
  NR2D1BWP12T U3498 ( .A1(n5863), .A2(n5862), .ZN(n5884) );
  XOR2XD0BWP12T U3499 ( .A1(a[27]), .A2(n5864), .Z(n5865) );
  AOI22D0BWP12T U3500 ( .A1(n5868), .A2(n5867), .B1(n5866), .B2(n5865), .ZN(
        n5883) );
  MUX2NXD0BWP12T U3501 ( .I0(n5872), .I1(n5871), .S(b[17]), .ZN(n5873) );
  NR2D1BWP12T U3502 ( .A1(n5874), .A2(n5873), .ZN(n5882) );
  MUX2ND0BWP12T U3503 ( .I0(n5878), .I1(n5877), .S(b[25]), .ZN(n5879) );
  NR2D1BWP12T U3504 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  XOR4D1BWP12T U3505 ( .A1(n5884), .A2(n5883), .A3(n5882), .A4(n5881), .Z(
        n5889) );
  MAOI222D0BWP12T U3506 ( .A(n5887), .B(n5886), .C(n5885), .ZN(n5888) );
  XNR4D1BWP12T U3507 ( .A1(n5891), .A2(n5890), .A3(n5889), .A4(n5888), .ZN(
        n5896) );
  FA1D0BWP12T U3508 ( .A(n5894), .B(n5893), .CI(n5892), .CO(n5895), .S(n5752)
         );
  TPND2D0BWP12T U3509 ( .A1(n6609), .A2(n6834), .ZN(n5921) );
  OA21D0BWP12T U3510 ( .A1(n5904), .A2(n6505), .B(n5903), .Z(n5905) );
  TPOAI22D0BWP12T U3511 ( .A1(n5906), .A2(n6890), .B1(n5905), .B2(n6836), .ZN(
        n5916) );
  AOI21D0BWP12T U3512 ( .A1(n5922), .A2(n5908), .B(n5907), .ZN(n5909) );
  OAI21D0BWP12T U3513 ( .A1(n5909), .A2(n5910), .B(n6833), .ZN(n5913) );
  AO211D1BWP12T U3514 ( .A1(n5911), .A2(n6110), .B(n5910), .C(n6794), .Z(n5912) );
  ND2D1BWP12T U3515 ( .A1(n5913), .A2(n5912), .ZN(n5915) );
  MUX2NXD0BWP12T U3516 ( .I0(n5916), .I1(n5915), .S(b[31]), .ZN(n5920) );
  NR2D0BWP12T U3517 ( .A1(n6728), .A2(n6898), .ZN(n6611) );
  NR2D0BWP12T U3518 ( .A1(n6833), .A2(n6870), .ZN(n5914) );
  MUX2ND0BWP12T U3519 ( .I0(n6611), .I1(n5914), .S(b[31]), .ZN(n5917) );
  TPOAI31D0BWP12T U3520 ( .A1(n5917), .A2(n5916), .A3(n5915), .B(a[31]), .ZN(
        n5919) );
  ND4D1BWP12T U3521 ( .A1(n5921), .A2(n5920), .A3(n5919), .A4(n5918), .ZN(
        c_out) );
  ND2D1BWP12T U3522 ( .A1(n6841), .A2(n6845), .ZN(n6166) );
  XOR2XD1BWP12T U3523 ( .A1(n5922), .A2(n6166), .Z(n6832) );
  XOR2XD0BWP12T U3524 ( .A1(n5923), .A2(n6168), .Z(n6640) );
  ND2D1BWP12T U3525 ( .A1(n5926), .A2(n5925), .ZN(n6682) );
  XOR2XD0BWP12T U3526 ( .A1(n5927), .A2(n6682), .Z(n6691) );
  AOI21D1BWP12T U3527 ( .A1(n5928), .A2(n5929), .B(n6133), .ZN(n5944) );
  AO31D1BWP12T U3528 ( .A1(n5929), .A2(n6133), .A3(n5928), .B(n5944), .Z(n6806) );
  OAI21D0BWP12T U3529 ( .A1(n5979), .A2(n5931), .B(n5930), .ZN(n6895) );
  ND4D0BWP12T U3530 ( .A1(n5933), .A2(n6833), .A3(n6895), .A4(n5932), .ZN(
        n5934) );
  NR4D0BWP12T U3531 ( .A1(n5937), .A2(n5936), .A3(n5935), .A4(n5934), .ZN(
        n5943) );
  INVD1BWP12T U3532 ( .I(n5938), .ZN(n5939) );
  ND2D1BWP12T U3533 ( .A1(n5939), .A2(n6097), .ZN(n5940) );
  XOR2XD1BWP12T U3534 ( .A1(n5940), .A2(n6134), .Z(n6800) );
  XNR2XD0BWP12T U3535 ( .A1(n5942), .A2(n5941), .ZN(n6724) );
  ND4D0BWP12T U3536 ( .A1(n6806), .A2(n5943), .A3(n6800), .A4(n6724), .ZN(
        n5947) );
  NR4D0BWP12T U3537 ( .A1(n5947), .A2(n5946), .A3(n6772), .A4(n5945), .ZN(
        n5949) );
  ND4D0BWP12T U3538 ( .A1(n5951), .A2(n5950), .A3(n5949), .A4(n5948), .ZN(
        n5952) );
  NR4D0BWP12T U3539 ( .A1(n6691), .A2(n5954), .A3(n5953), .A4(n5952), .ZN(
        n5956) );
  ND4D0BWP12T U3540 ( .A1(n6640), .A2(n6671), .A3(n5956), .A4(n5955), .ZN(
        n5957) );
  NR4D0BWP12T U3541 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(
        n5962) );
  ND4D0BWP12T U3542 ( .A1(n5964), .A2(n5963), .A3(n5962), .A4(n5961), .ZN(
        n5965) );
  NR4D0BWP12T U3543 ( .A1(n6832), .A2(n5967), .A3(n5966), .A4(n5965), .ZN(
        n6005) );
  XOR2XD1BWP12T U3544 ( .A1(n5969), .A2(n6170), .Z(n6674) );
  INVD1BWP12T U3545 ( .I(n5970), .ZN(n6127) );
  XNR2XD0BWP12T U3546 ( .A1(n5973), .A2(n6707), .ZN(n6729) );
  XNR2XD1BWP12T U3547 ( .A1(n5974), .A2(n6175), .ZN(n6775) );
  XOR2XD1BWP12T U3548 ( .A1(n5984), .A2(n6133), .Z(n6830) );
  AOI22D0BWP12T U3549 ( .A1(n6005), .A2(n6004), .B1(n6003), .B2(n6002), .ZN(
        n6607) );
  INVD1BWP12T U3550 ( .I(n6006), .ZN(n6008) );
  ND2D1BWP12T U3551 ( .A1(n6008), .A2(n6007), .ZN(n6010) );
  XNR2D1BWP12T U3552 ( .A1(n6010), .A2(n6009), .ZN(n6645) );
  OAI21D1BWP12T U3553 ( .A1(n6013), .A2(n6012), .B(n6011), .ZN(n6018) );
  INVD1BWP12T U3554 ( .I(n6014), .ZN(n6016) );
  ND2D1BWP12T U3555 ( .A1(n6016), .A2(n6015), .ZN(n6017) );
  XNR2D1BWP12T U3556 ( .A1(n6018), .A2(n6017), .ZN(n6732) );
  INVD1BWP12T U3557 ( .I(n6019), .ZN(n6021) );
  ND2D1BWP12T U3558 ( .A1(n6021), .A2(n6020), .ZN(n6023) );
  XNR2D1BWP12T U3559 ( .A1(n6023), .A2(n6022), .ZN(n6805) );
  ND2D1BWP12T U3560 ( .A1(n6025), .A2(n6024), .ZN(n6027) );
  XNR2D1BWP12T U3561 ( .A1(n6027), .A2(n6026), .ZN(n6733) );
  INVD1BWP12T U3562 ( .I(n6028), .ZN(n6030) );
  ND2D1BWP12T U3563 ( .A1(n6030), .A2(n6029), .ZN(n6032) );
  XOR2XD1BWP12T U3564 ( .A1(n6032), .A2(n6031), .Z(n6804) );
  NR4D0BWP12T U3565 ( .A1(n6037), .A2(n6869), .A3(n6902), .A4(n6036), .ZN(
        n6039) );
  ND4D0BWP12T U3566 ( .A1(n6804), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(
        n6041) );
  NR3D0BWP12T U3567 ( .A1(n6805), .A2(n6733), .A3(n6041), .ZN(n6042) );
  AN4XD1BWP12T U3568 ( .A1(n6732), .A2(n6044), .A3(n6043), .A4(n6042), .Z(
        n6047) );
  AN4XD1BWP12T U3569 ( .A1(n6048), .A2(n6047), .A3(n6046), .A4(n6045), .Z(
        n6051) );
  ND4D1BWP12T U3570 ( .A1(n6052), .A2(n6051), .A3(n6050), .A4(n6049), .ZN(
        n6065) );
  INVD1BWP12T U3571 ( .I(n6056), .ZN(n6058) );
  CKND2D1BWP12T U3572 ( .A1(n6058), .A2(n6057), .ZN(n6059) );
  XNR2D1BWP12T U3573 ( .A1(n6060), .A2(n6059), .ZN(n6697) );
  IND4D1BWP12T U3574 ( .A1(n6065), .B1(n6064), .B2(n6697), .B3(n6675), .ZN(
        n6067) );
  OR4D0BWP12T U3575 ( .A1(n6645), .A2(n6068), .A3(n6067), .A4(n6066), .Z(n6070) );
  OR4XD1BWP12T U3576 ( .A1(n6072), .A2(n6071), .A3(n6070), .A4(n6069), .Z(
        n6088) );
  TPNR2D0BWP12T U3577 ( .A1(n6073), .A2(n6075), .ZN(n6079) );
  TPOAI21D0BWP12T U3578 ( .A1(n6076), .A2(n6075), .B(n6074), .ZN(n6077) );
  AOI21D1BWP12T U3579 ( .A1(n6079), .A2(n6078), .B(n6077), .ZN(n6083) );
  ND2D1BWP12T U3580 ( .A1(n6081), .A2(n6080), .ZN(n6082) );
  XOR2XD1BWP12T U3581 ( .A1(n6083), .A2(n6082), .Z(n6835) );
  OR3XD1BWP12T U3582 ( .A1(n6085), .A2(n6084), .A3(n6608), .Z(n6087) );
  NR4D0BWP12T U3583 ( .A1(n6088), .A2(n6835), .A3(n6087), .A4(n6086), .ZN(
        n6123) );
  OR4D0BWP12T U3584 ( .A1(n6092), .A2(n6091), .A3(n6090), .A4(n6089), .Z(n6120) );
  ND4D0BWP12T U3585 ( .A1(n6095), .A2(n6094), .A3(n6706), .A4(n6093), .ZN(
        n6100) );
  ND4D0BWP12T U3586 ( .A1(n6098), .A2(n6097), .A3(n6811), .A4(n6096), .ZN(
        n6099) );
  NR2XD0BWP12T U3587 ( .A1(n6100), .A2(n6099), .ZN(n6109) );
  CKND2D0BWP12T U3588 ( .A1(b[27]), .A2(a[27]), .ZN(n6103) );
  CKND2D0BWP12T U3589 ( .A1(b[22]), .A2(a[22]), .ZN(n6102) );
  ND4D0BWP12T U3590 ( .A1(n6104), .A2(n6103), .A3(n6102), .A4(n6101), .ZN(
        n6105) );
  AOI211D0BWP12T U3591 ( .A1(a[31]), .A2(b[31]), .B(n6106), .C(n6105), .ZN(
        n6108) );
  ND4D0BWP12T U3592 ( .A1(n6110), .A2(n6109), .A3(n6108), .A4(n6107), .ZN(
        n6119) );
  ND4D0BWP12T U3593 ( .A1(n6113), .A2(n6112), .A3(n6197), .A4(n6111), .ZN(
        n6118) );
  ND4D0BWP12T U3594 ( .A1(n6116), .A2(n6627), .A3(n6115), .A4(n6114), .ZN(
        n6117) );
  NR4D0BWP12T U3595 ( .A1(n6120), .A2(n6119), .A3(n6118), .A4(n6117), .ZN(
        n6122) );
  OAI21D1BWP12T U3596 ( .A1(n6123), .A2(n6122), .B(n6121), .ZN(n6605) );
  INVD0BWP12T U3597 ( .I(n6124), .ZN(n6673) );
  CKND2D0BWP12T U3598 ( .A1(n6125), .A2(n6170), .ZN(n6672) );
  INVD0BWP12T U3599 ( .I(n6130), .ZN(n6131) );
  XOR2XD1BWP12T U3600 ( .A1(n6131), .A2(n6175), .Z(n6734) );
  CKXOR2D1BWP12T U3601 ( .A1(n6135), .A2(n6134), .Z(n6796) );
  OAI21D0BWP12T U3602 ( .A1(n6618), .A2(n6150), .B(n6149), .ZN(n6643) );
  AOI211D0BWP12T U3603 ( .A1(n6160), .A2(n6159), .B(n6158), .C(n6157), .ZN(
        n6603) );
  AN3D0BWP12T U3604 ( .A1(n6163), .A2(n6162), .A3(n6161), .Z(n6602) );
  XOR2XD1BWP12T U3605 ( .A1(n6167), .A2(n6166), .Z(n6865) );
  XNR2XD0BWP12T U3606 ( .A1(n6169), .A2(n6168), .ZN(n6638) );
  CKXOR2D0BWP12T U3607 ( .A1(n6171), .A2(n6170), .Z(n6670) );
  XNR2XD0BWP12T U3608 ( .A1(n6172), .A2(n6682), .ZN(n6690) );
  AOI21D0BWP12T U3609 ( .A1(n6175), .A2(n6174), .B(n6173), .ZN(n6767) );
  OAI21D1BWP12T U3610 ( .A1(n6178), .A2(n6177), .B(n6176), .ZN(n6795) );
  TPAOI21D0BWP12T U3611 ( .A1(n6181), .A2(n6180), .B(n6179), .ZN(n6871) );
  NR4D0BWP12T U3612 ( .A1(n6871), .A2(n6183), .A3(n6182), .A4(n6794), .ZN(
        n6184) );
  ND4D0BWP12T U3613 ( .A1(n6795), .A2(n6186), .A3(n6185), .A4(n6184), .ZN(
        n6192) );
  TPOAI31D0BWP12T U3614 ( .A1(n6190), .A2(n6189), .A3(n6188), .B(n6187), .ZN(
        n6809) );
  NR4D0BWP12T U3615 ( .A1(n6767), .A2(n6192), .A3(n6191), .A4(n6809), .ZN(
        n6194) );
  ND4D0BWP12T U3616 ( .A1(n6196), .A2(n6195), .A3(n6194), .A4(n6193), .ZN(
        n6200) );
  NR4D0BWP12T U3617 ( .A1(n6201), .A2(n6200), .A3(n6199), .A4(n6727), .ZN(
        n6204) );
  ND4D0BWP12T U3618 ( .A1(n6205), .A2(n6204), .A3(n6203), .A4(n6202), .ZN(
        n6206) );
  NR4D0BWP12T U3619 ( .A1(n6207), .A2(n6670), .A3(n6690), .A4(n6206), .ZN(
        n6208) );
  ND4D0BWP12T U3620 ( .A1(n6210), .A2(n6209), .A3(n6638), .A4(n6208), .ZN(
        n6211) );
  NR4D0BWP12T U3621 ( .A1(n6214), .A2(n6213), .A3(n6212), .A4(n6211), .ZN(
        n6216) );
  ND4D0BWP12T U3622 ( .A1(n6218), .A2(n6217), .A3(n6216), .A4(n6215), .ZN(
        n6599) );
  NR4D0BWP12T U3623 ( .A1(n6560), .A2(n6219), .A3(a[31]), .A4(n6874), .ZN(
        n6596) );
  NR3D0BWP12T U3624 ( .A1(n6221), .A2(n6220), .A3(n6862), .ZN(n6225) );
  TPND2D0BWP12T U3625 ( .A1(n6597), .A2(a[31]), .ZN(n6613) );
  OAI21D0BWP12T U3626 ( .A1(n6224), .A2(n6223), .B(n6222), .ZN(n6861) );
  ND4D0BWP12T U3627 ( .A1(n6226), .A2(n6225), .A3(n6613), .A4(n6861), .ZN(
        n6244) );
  ND4D0BWP12T U3628 ( .A1(a[25]), .A2(a[24]), .A3(a[22]), .A4(a[20]), .ZN(
        n6235) );
  ND4D1BWP12T U3629 ( .A1(n6230), .A2(n6249), .A3(n6715), .A4(n6229), .ZN(
        n6234) );
  ND4D1BWP12T U3630 ( .A1(a[19]), .A2(a[18]), .A3(n6232), .A4(n6231), .ZN(
        n6233) );
  NR4D0BWP12T U3631 ( .A1(n6236), .A2(n6235), .A3(n6234), .A4(n6233), .ZN(
        n6242) );
  NR4D0BWP12T U3632 ( .A1(n6240), .A2(n6239), .A3(n6238), .A4(n6237), .ZN(
        n6241) );
  CKND2D1BWP12T U3633 ( .A1(n6242), .A2(n6241), .ZN(n6243) );
  MUX2ND0BWP12T U3634 ( .I0(n6244), .I1(n6243), .S(a[2]), .ZN(n6595) );
  MUX2ND0BWP12T U3635 ( .I0(n6325), .I1(n6321), .S(n6334), .ZN(n6379) );
  AOI21D1BWP12T U3636 ( .A1(n6573), .A2(n6379), .B(n6333), .ZN(n6906) );
  ND2D1BWP12T U3637 ( .A1(n6356), .A2(n6253), .ZN(n6316) );
  CKND2D0BWP12T U3638 ( .A1(n6255), .A2(n6254), .ZN(n6258) );
  AOI21D0BWP12T U3639 ( .A1(n6256), .A2(n6278), .B(n6573), .ZN(n6257) );
  OAI211D1BWP12T U3640 ( .A1(n6259), .A2(n6297), .B(n6258), .C(n6257), .ZN(
        n6261) );
  NR2D1BWP12T U3641 ( .A1(n6298), .A2(n6304), .ZN(n6260) );
  NR2D1BWP12T U3642 ( .A1(n6261), .A2(n6260), .ZN(n6360) );
  AOI21D0BWP12T U3643 ( .A1(n6573), .A2(n6316), .B(n6360), .ZN(n6721) );
  AOI22D1BWP12T U3644 ( .A1(n6264), .A2(n6263), .B1(a[8]), .B2(n6262), .ZN(
        n6265) );
  OAI22D1BWP12T U3645 ( .A1(n6266), .A2(n6308), .B1(n6265), .B2(n6304), .ZN(
        n6272) );
  AOI21D1BWP12T U3646 ( .A1(n6268), .A2(n6267), .B(n6573), .ZN(n6269) );
  OAI21D0BWP12T U3647 ( .A1(n6270), .A2(n6306), .B(n6269), .ZN(n6271) );
  AOI211D1BWP12T U3648 ( .A1(n6313), .A2(n6273), .B(n6272), .C(n6271), .ZN(
        n6776) );
  TPNR2D0BWP12T U3649 ( .A1(n6274), .A2(n6297), .ZN(n6277) );
  NR2D1BWP12T U3650 ( .A1(n6275), .A2(n6304), .ZN(n6276) );
  NR2D1BWP12T U3651 ( .A1(n6277), .A2(n6276), .ZN(n6335) );
  NR2D0BWP12T U3652 ( .A1(n6620), .A2(n6357), .ZN(n6285) );
  AOI211D0BWP12T U3653 ( .A1(n6282), .A2(n6281), .B(n6280), .C(n6279), .ZN(
        n6284) );
  OAI211D0BWP12T U3654 ( .A1(n6776), .A2(n6285), .B(n6284), .C(n6283), .ZN(
        n6286) );
  OR4D0BWP12T U3655 ( .A1(n6287), .A2(n6906), .A3(n6721), .A4(n6286), .Z(n6446) );
  CKND0BWP12T U3656 ( .I(n6446), .ZN(n6296) );
  NR2XD0BWP12T U3657 ( .A1(n6345), .A2(n6288), .ZN(n6808) );
  CKND2D0BWP12T U3658 ( .A1(n6808), .A2(n6289), .ZN(n6402) );
  CKND0BWP12T U3659 ( .I(n6402), .ZN(n6295) );
  INR2D0BWP12T U3660 ( .A1(n6735), .B1(n6290), .ZN(n6320) );
  CKND0BWP12T U3661 ( .I(n6320), .ZN(n6291) );
  NR4D0BWP12T U3662 ( .A1(n6293), .A2(n6292), .A3(n6384), .A4(n6291), .ZN(
        n6294) );
  OAI21D1BWP12T U3663 ( .A1(n6298), .A2(n6297), .B(n6565), .ZN(n6301) );
  NR2D1BWP12T U3664 ( .A1(n6299), .A2(n6304), .ZN(n6300) );
  NR2D1BWP12T U3665 ( .A1(n6301), .A2(n6300), .ZN(n6302) );
  OAI21D0BWP12T U3666 ( .A1(n6303), .A2(n6576), .B(n6302), .ZN(n6346) );
  OAI22D1BWP12T U3667 ( .A1(n6307), .A2(n6306), .B1(n6305), .B2(n6304), .ZN(
        n6311) );
  OAI21D1BWP12T U3668 ( .A1(n6309), .A2(n6308), .B(n6565), .ZN(n6310) );
  AOI211D1BWP12T U3669 ( .A1(n6313), .A2(n6312), .B(n6311), .C(n6310), .ZN(
        n6740) );
  CKND2D0BWP12T U3670 ( .A1(n6320), .A2(n6319), .ZN(n6385) );
  NR4D0BWP12T U3671 ( .A1(n6385), .A2(n6325), .A3(n6324), .A4(n6386), .ZN(
        n6326) );
  AOI21D1BWP12T U3672 ( .A1(n6377), .A2(n6326), .B(n6584), .ZN(n6374) );
  NR4D0BWP12T U3673 ( .A1(n6330), .A2(n6329), .A3(n6328), .A4(n6327), .ZN(
        n6338) );
  AOI211D1BWP12T U3674 ( .A1(n6339), .A2(n6573), .B(n6333), .C(n6560), .ZN(
        n6908) );
  AOI21D1BWP12T U3675 ( .A1(n6629), .A2(n6355), .B(n6350), .ZN(n6337) );
  OAI21D1BWP12T U3676 ( .A1(n6337), .A2(n6776), .B(n6336), .ZN(n6793) );
  INR3XD0BWP12T U3677 ( .A1(n6338), .B1(n6908), .B2(n6793), .ZN(n6371) );
  INVD1BWP12T U3678 ( .I(n6339), .ZN(n6687) );
  CKND0BWP12T U3679 ( .I(n6345), .ZN(n6347) );
  INVD1BWP12T U3680 ( .I(n6346), .ZN(n6824) );
  AOI211D1BWP12T U3681 ( .A1(n6364), .A2(n6347), .B(n6824), .C(n6560), .ZN(
        n6823) );
  AOI211D1BWP12T U3682 ( .A1(n6350), .A2(n6349), .B(n6823), .C(n6348), .ZN(
        n6370) );
  ND4D0BWP12T U3683 ( .A1(n6354), .A2(n6909), .A3(n6353), .A4(n6851), .ZN(
        n6361) );
  OAI31D1BWP12T U3684 ( .A1(n6358), .A2(n6357), .A3(n6356), .B(n6355), .ZN(
        n6359) );
  NR2D1BWP12T U3685 ( .A1(n6360), .A2(n6359), .ZN(n6700) );
  NR4D0BWP12T U3686 ( .A1(n6363), .A2(n6362), .A3(n6361), .A4(n6700), .ZN(
        n6369) );
  AOI211XD0BWP12T U3687 ( .A1(n6735), .A2(n6364), .B(n6740), .C(n6560), .ZN(
        n6766) );
  NR4D0BWP12T U3688 ( .A1(n6367), .A2(n6766), .A3(n6366), .A4(n6365), .ZN(
        n6368) );
  ND4D1BWP12T U3689 ( .A1(n6371), .A2(n6370), .A3(n6369), .A4(n6368), .ZN(
        n6372) );
  TPOAI31D0BWP12T U3690 ( .A1(n6375), .A2(n6374), .A3(n6373), .B(n6372), .ZN(
        n6592) );
  AOI22D0BWP12T U3691 ( .A1(n6377), .A2(n6376), .B1(n6573), .B2(n6742), .ZN(
        n6430) );
  NR2D1BWP12T U3692 ( .A1(n6379), .A2(n6573), .ZN(n6677) );
  ND3D0BWP12T U3693 ( .A1(n6421), .A2(n6857), .A3(n6380), .ZN(n6381) );
  NR4D0BWP12T U3694 ( .A1(n6384), .A2(n6383), .A3(n6382), .A4(n6381), .ZN(
        n6390) );
  NR4D0BWP12T U3695 ( .A1(n6388), .A2(n6387), .A3(n6386), .A4(n6385), .ZN(
        n6389) );
  AN4D0BWP12T U3696 ( .A1(n6689), .A2(n6718), .A3(n6390), .A4(n6389), .Z(n6429) );
  NR2D1BWP12T U3697 ( .A1(n6409), .A2(n6403), .ZN(n6406) );
  OAI22D1BWP12T U3698 ( .A1(n6408), .A2(n6531), .B1(n6407), .B2(n6532), .ZN(
        n6405) );
  TPNR2D0BWP12T U3699 ( .A1(n6410), .A2(n6535), .ZN(n6404) );
  NR3D1BWP12T U3700 ( .A1(n6406), .A2(n6405), .A3(n6404), .ZN(n6440) );
  CKND2D1BWP12T U3701 ( .A1(n6792), .A2(n6717), .ZN(n6435) );
  OAI211D0BWP12T U3702 ( .A1(n6440), .A2(n6565), .B(n6435), .C(n6436), .ZN(
        n6416) );
  OAI22D1BWP12T U3703 ( .A1(n6408), .A2(n6550), .B1(n6407), .B2(n6551), .ZN(
        n6414) );
  NR2D1BWP12T U3704 ( .A1(n6409), .A2(n6555), .ZN(n6413) );
  NR2D0BWP12T U3705 ( .A1(n6410), .A2(n6554), .ZN(n6412) );
  TPOAI31D0BWP12T U3706 ( .A1(n6414), .A2(n6413), .A3(n6412), .B(n6411), .ZN(
        n6415) );
  OAI211D1BWP12T U3707 ( .A1(n6437), .A2(n6417), .B(n6416), .C(n6415), .ZN(
        n6858) );
  OAI22D1BWP12T U3708 ( .A1(n6420), .A2(n6419), .B1(n6418), .B2(n6439), .ZN(
        n6424) );
  CKND0BWP12T U3709 ( .I(n6421), .ZN(n6422) );
  TPOAI21D0BWP12T U3710 ( .A1(n6422), .A2(n6426), .B(n6438), .ZN(n6423) );
  NR2D1BWP12T U3711 ( .A1(n6424), .A2(n6423), .ZN(n6669) );
  AOI211D0BWP12T U3712 ( .A1(n6426), .A2(n6425), .B(n6858), .C(n6669), .ZN(
        n6427) );
  IND4D1BWP12T U3713 ( .A1(n6430), .B1(n6429), .B2(n6428), .B3(n6427), .ZN(
        n6447) );
  ND4D0BWP12T U3714 ( .A1(n6434), .A2(n6433), .A3(n6432), .A4(n6431), .ZN(
        n6445) );
  ND4D0BWP12T U3715 ( .A1(n6443), .A2(n6619), .A3(n6442), .A4(n6441), .ZN(
        n6444) );
  NR4D0BWP12T U3716 ( .A1(n6447), .A2(n6446), .A3(n6445), .A4(n6444), .ZN(
        n6591) );
  INVD0BWP12T U3717 ( .I(n6466), .ZN(n6878) );
  MAOI22D0BWP12T U3718 ( .A1(n6655), .A2(n6476), .B1(n6475), .B2(n6474), .ZN(
        n6589) );
  NR4D0BWP12T U3719 ( .A1(n6486), .A2(n6485), .A3(n6746), .A4(n6484), .ZN(
        n6491) );
  ND4D1BWP12T U3720 ( .A1(n6493), .A2(n6492), .A3(n6491), .A4(n6490), .ZN(
        n6588) );
  NR4D0BWP12T U3721 ( .A1(n6500), .A2(n6499), .A3(n6498), .A4(n6497), .ZN(
        n6508) );
  ND4D1BWP12T U3722 ( .A1(n6509), .A2(n6508), .A3(n6507), .A4(n6506), .ZN(
        n6587) );
  INVD1BWP12T U3723 ( .I(n6511), .ZN(n6738) );
  INVD1BWP12T U3724 ( .I(n6516), .ZN(n6821) );
  INVD1BWP12T U3725 ( .I(n6517), .ZN(n6574) );
  NR2D1BWP12T U3726 ( .A1(n6521), .A2(n6520), .ZN(n6872) );
  TPAOI21D0BWP12T U3727 ( .A1(n6562), .A2(n6524), .B(n6540), .ZN(n6527) );
  CKND2D0BWP12T U3728 ( .A1(n6525), .A2(n6578), .ZN(n6526) );
  OAI211D1BWP12T U3729 ( .A1(n6872), .A2(n6565), .B(n6527), .C(n6526), .ZN(
        n6681) );
  ND3D0BWP12T U3730 ( .A1(n6529), .A2(n6681), .A3(n6528), .ZN(n6544) );
  OAI22D0BWP12T U3731 ( .A1(n6533), .A2(n6532), .B1(n6531), .B2(n6530), .ZN(
        n6537) );
  NR2D0BWP12T U3732 ( .A1(n6535), .A2(n6534), .ZN(n6536) );
  AOI211D0BWP12T U3733 ( .A1(n6556), .A2(n6538), .B(n6537), .C(n6536), .ZN(
        n6548) );
  OAI22D1BWP12T U3734 ( .A1(n6539), .A2(n6576), .B1(n6548), .B2(n6557), .ZN(
        n6541) );
  RCAOI211D0BWP12T U3735 ( .A1(n6573), .A2(n6778), .B(n6541), .C(n6540), .ZN(
        n6633) );
  NR4D0BWP12T U3736 ( .A1(n6544), .A2(n6633), .A3(n6543), .A4(n6542), .ZN(
        n6569) );
  NR4D0BWP12T U3737 ( .A1(n6547), .A2(n6546), .A3(n6545), .A4(n6680), .ZN(
        n6568) );
  CKND0BWP12T U3738 ( .I(n6548), .ZN(n6563) );
  AOI22D0BWP12T U3739 ( .A1(n6552), .A2(n6551), .B1(n6550), .B2(n6549), .ZN(
        n6559) );
  AOI22D0BWP12T U3740 ( .A1(n6556), .A2(n6555), .B1(n6554), .B2(n6553), .ZN(
        n6558) );
  RCAOI21D0BWP12T U3741 ( .A1(n6559), .A2(n6558), .B(n6557), .ZN(n6561) );
  AOI211D0BWP12T U3742 ( .A1(n6563), .A2(n6562), .B(n6561), .C(n6560), .ZN(
        n6564) );
  OAI21D1BWP12T U3743 ( .A1(n6566), .A2(n6565), .B(n6564), .ZN(n6838) );
  AN4D0BWP12T U3744 ( .A1(n6569), .A2(n6568), .A3(n6838), .A4(n6567), .Z(n6583) );
  CKND2D0BWP12T U3745 ( .A1(n6571), .A2(n6570), .ZN(n6580) );
  NR4D0BWP12T U3746 ( .A1(n6581), .A2(n6580), .A3(n6579), .A4(n6650), .ZN(
        n6582) );
  OAI211D1BWP12T U3747 ( .A1(n6585), .A2(n6584), .B(n6583), .C(n6582), .ZN(
        n6586) );
  OAI31D1BWP12T U3748 ( .A1(n6589), .A2(n6588), .A3(n6587), .B(n6586), .ZN(
        n6590) );
  AO211D0BWP12T U3749 ( .A1(n6593), .A2(n6592), .B(n6591), .C(n6590), .Z(n6594) );
  AOI211D0BWP12T U3750 ( .A1(n6597), .A2(n6596), .B(n6595), .C(n6594), .ZN(
        n6598) );
  TPOAI31D0BWP12T U3751 ( .A1(n6865), .A2(n6600), .A3(n6599), .B(n6598), .ZN(
        n6601) );
  TPAOI31D0BWP12T U3752 ( .A1(n6603), .A2(n6602), .A3(n6837), .B(n6601), .ZN(
        n6604) );
  OAI211D1BWP12T U3753 ( .A1(n6607), .A2(n6606), .B(n6605), .C(n6604), .ZN(z)
         );
  XNR2XD1BWP12T U3754 ( .A1(n6609), .A2(n6608), .ZN(n6610) );
  OAI222D1BWP12T U3755 ( .A1(n6613), .A2(n6862), .B1(n6612), .B2(n6611), .C1(
        n6902), .C2(n6610), .ZN(v) );
  TPNR2D0BWP12T U3756 ( .A1(n6615), .A2(n6614), .ZN(n6617) );
  OAI211D1BWP12T U3757 ( .A1(n6618), .A2(n6617), .B(n6616), .C(n6728), .ZN(
        n6642) );
  NR2D1BWP12T U3758 ( .A1(n6619), .A2(n6716), .ZN(n6632) );
  INVD1BWP12T U3759 ( .I(n6620), .ZN(n6777) );
  OAI211D0BWP12T U3760 ( .A1(n6744), .A2(n6627), .B(n6622), .C(n6621), .ZN(
        n6626) );
  AOI22D0BWP12T U3761 ( .A1(n6624), .A2(n6655), .B1(n6783), .B2(n6623), .ZN(
        n6625) );
  OAI211D0BWP12T U3762 ( .A1(n6880), .A2(n6627), .B(n6626), .C(n6625), .ZN(
        n6628) );
  AOI211D1BWP12T U3763 ( .A1(n6688), .A2(n6629), .B(n6661), .C(n6628), .ZN(
        n6630) );
  OAI21D1BWP12T U3764 ( .A1(n6777), .A2(n6840), .B(n6630), .ZN(n6631) );
  AOI211D1BWP12T U3765 ( .A1(n6855), .A2(n6633), .B(n6632), .C(n6631), .ZN(
        n6637) );
  AO211D0BWP12T U3766 ( .A1(a[21]), .A2(n6635), .B(n6634), .C(n6862), .Z(n6636) );
  OAI211D1BWP12T U3767 ( .A1(n6794), .A2(n6638), .B(n6637), .C(n6636), .ZN(
        n6639) );
  RCIAO21D0BWP12T U3768 ( .A1(n6640), .A2(n6894), .B(n6639), .ZN(n6641) );
  OAI211D1BWP12T U3769 ( .A1(n6836), .A2(n6643), .B(n6642), .C(n6641), .ZN(
        n6644) );
  AO21D1BWP12T U3770 ( .A1(n6645), .A2(n6834), .B(n6644), .Z(result[21]) );
  CKND2D0BWP12T U3771 ( .A1(n6647), .A2(n6646), .ZN(n6649) );
  AOI211D1BWP12T U3772 ( .A1(n6649), .A2(a[19]), .B(n6648), .C(n6862), .ZN(
        n6668) );
  CKND2D1BWP12T U3773 ( .A1(n6650), .A2(n6855), .ZN(n6664) );
  CKND0BWP12T U3774 ( .I(n6651), .ZN(n6653) );
  AOI22D0BWP12T U3775 ( .A1(n6653), .A2(n6747), .B1(n6652), .B2(n6744), .ZN(
        n6658) );
  AOI22D1BWP12T U3776 ( .A1(n6656), .A2(n6655), .B1(n6783), .B2(n6654), .ZN(
        n6657) );
  OAI211D0BWP12T U3777 ( .A1(n6659), .A2(n6813), .B(n6658), .C(n6657), .ZN(
        n6660) );
  RCAOI211D0BWP12T U3778 ( .A1(n6688), .A2(n6662), .B(n6661), .C(n6660), .ZN(
        n6663) );
  OAI211D1BWP12T U3779 ( .A1(n6666), .A2(n6665), .B(n6664), .C(n6663), .ZN(
        n6667) );
  AOI21D1BWP12T U3780 ( .A1(n6693), .A2(n6898), .B(n6692), .ZN(n6696) );
  ND2D1BWP12T U3781 ( .A1(n6694), .A2(n6728), .ZN(n6695) );
  OAI211D1BWP12T U3782 ( .A1(n6902), .A2(n6697), .B(n6696), .C(n6695), .ZN(
        result[18]) );
  NR2D1BWP12T U3783 ( .A1(n6698), .A2(n6836), .ZN(n6726) );
  AOI22D1BWP12T U3784 ( .A1(n6700), .A2(n6909), .B1(n6708), .B2(n6699), .ZN(
        n6723) );
  CKND0BWP12T U3785 ( .I(n6703), .ZN(n6705) );
  AOI211D0BWP12T U3786 ( .A1(n6706), .A2(n6810), .B(n6705), .C(n6704), .ZN(
        n6710) );
  AOI211D0BWP12T U3787 ( .A1(n6708), .A2(n6813), .B(n6707), .C(n6882), .ZN(
        n6709) );
  NR4D0BWP12T U3788 ( .A1(n6711), .A2(n6753), .A3(n6710), .A4(n6709), .ZN(
        n6712) );
  OAI31D0BWP12T U3789 ( .A1(n6715), .A2(n6714), .A3(n6713), .B(n6712), .ZN(
        n6720) );
  NR3D1BWP12T U3790 ( .A1(n6718), .A2(n6717), .A3(n6716), .ZN(n6719) );
  RCAOI211D0BWP12T U3791 ( .A1(n6721), .A2(n6905), .B(n6720), .C(n6719), .ZN(
        n6722) );
  OAI211D1BWP12T U3792 ( .A1(n6894), .A2(n6724), .B(n6723), .C(n6722), .ZN(
        n6725) );
  AOI211D1BWP12T U3793 ( .A1(n6870), .A2(n6727), .B(n6726), .C(n6725), .ZN(
        n6731) );
  CKND2D1BWP12T U3794 ( .A1(n6729), .A2(n6728), .ZN(n6730) );
  ND2D1BWP12T U3795 ( .A1(n6733), .A2(n6834), .ZN(n6774) );
  INVD1BWP12T U3796 ( .I(n6734), .ZN(n6770) );
  INVD0BWP12T U3797 ( .I(n6735), .ZN(n6737) );
  AOI21D0BWP12T U3798 ( .A1(n6737), .A2(n6905), .B(n6736), .ZN(n6741) );
  OAI22D1BWP12T U3799 ( .A1(n6741), .A2(n6740), .B1(n6739), .B2(n6738), .ZN(
        n6765) );
  INVD0BWP12T U3800 ( .I(n6742), .ZN(n6754) );
  AOI21D1BWP12T U3801 ( .A1(a[8]), .A2(n6744), .B(n6743), .ZN(n6750) );
  AOI22D0BWP12T U3802 ( .A1(n6748), .A2(n6747), .B1(n6746), .B2(n6745), .ZN(
        n6749) );
  OAI21D1BWP12T U3803 ( .A1(n6751), .A2(n6750), .B(n6749), .ZN(n6752) );
  AOI211D1BWP12T U3804 ( .A1(n6755), .A2(n6754), .B(n6753), .C(n6752), .ZN(
        n6762) );
  INVD1BWP12T U3805 ( .I(n6756), .ZN(n6757) );
  NR2D0BWP12T U3806 ( .A1(n6757), .A2(n6862), .ZN(n6759) );
  OAI21D1BWP12T U3807 ( .A1(n6818), .A2(n6819), .B(a[8]), .ZN(n6758) );
  AOI22D1BWP12T U3808 ( .A1(n6820), .A2(n6760), .B1(n6759), .B2(n6758), .ZN(
        n6761) );
  OAI211D1BWP12T U3809 ( .A1(n6763), .A2(n6892), .B(n6762), .C(n6761), .ZN(
        n6764) );
  AOI211D1BWP12T U3810 ( .A1(n6909), .A2(n6766), .B(n6765), .C(n6764), .ZN(
        n6769) );
  CKND2D1BWP12T U3811 ( .A1(n6767), .A2(n6870), .ZN(n6768) );
  OAI211D1BWP12T U3812 ( .A1(n6836), .A2(n6770), .B(n6769), .C(n6768), .ZN(
        n6771) );
  AOI21D1BWP12T U3813 ( .A1(n6833), .A2(n6772), .B(n6771), .ZN(n6773) );
  OAI211D1BWP12T U3814 ( .A1(n6775), .A2(n6890), .B(n6774), .C(n6773), .ZN(
        result[8]) );
  TPOAI21D0BWP12T U3815 ( .A1(n6779), .A2(op[2]), .B(n6816), .ZN(n6781) );
  CKND2D0BWP12T U3816 ( .A1(n6788), .A2(n6879), .ZN(n6780) );
  OAI211D1BWP12T U3817 ( .A1(n6782), .A2(n6882), .B(n6781), .C(n6780), .ZN(
        n6785) );
  AOI22D0BWP12T U3818 ( .A1(n6785), .A2(n6784), .B1(n6783), .B2(n6788), .ZN(
        n6791) );
  OAI211D1BWP12T U3819 ( .A1(n6789), .A2(n6788), .B(n6787), .C(n6786), .ZN(
        n6790) );
  NR2D1BWP12T U3820 ( .A1(n6796), .A2(n6836), .ZN(n6797) );
  AOI211D1BWP12T U3821 ( .A1(n6728), .A2(n6799), .B(n6798), .C(n6797), .ZN(
        n6803) );
  INVD1BWP12T U3822 ( .I(n6800), .ZN(n6801) );
  ND2D1BWP12T U3823 ( .A1(n6801), .A2(n6833), .ZN(n6802) );
  OAI211D1BWP12T U3824 ( .A1(n6902), .A2(n6804), .B(n6803), .C(n6802), .ZN(
        result[5]) );
  ND2D1BWP12T U3825 ( .A1(n6805), .A2(n6834), .ZN(n6829) );
  NR2D1BWP12T U3826 ( .A1(n6806), .A2(n6894), .ZN(n6826) );
  AOI211D1BWP12T U3827 ( .A1(n6898), .A2(n6827), .B(n6826), .C(n6825), .ZN(
        n6828) );
  OAI211D1BWP12T U3828 ( .A1(n6890), .A2(n6830), .B(n6829), .C(n6828), .ZN(
        result[7]) );
  INVD1BWP12T U3829 ( .I(n6831), .ZN(n6868) );
  AOI22D1BWP12T U3830 ( .A1(n6835), .A2(n6834), .B1(n6833), .B2(n6832), .ZN(
        n6867) );
  NR2D1BWP12T U3831 ( .A1(n6837), .A2(n6836), .ZN(n6864) );
  INVD1BWP12T U3832 ( .I(n6838), .ZN(n6856) );
  NR2D1BWP12T U3833 ( .A1(n6840), .A2(n6839), .ZN(n6854) );
  CKND0BWP12T U3834 ( .I(n6841), .ZN(n6848) );
  OAI22D0BWP12T U3835 ( .A1(n6880), .A2(n6843), .B1(n6842), .B2(n6874), .ZN(
        n6847) );
  OAI22D0BWP12T U3836 ( .A1(n6845), .A2(n6882), .B1(a[29]), .B2(n6844), .ZN(
        n6846) );
  AOI211XD0BWP12T U3837 ( .A1(n6848), .A2(n6879), .B(n6847), .C(n6846), .ZN(
        n6849) );
  OAI211D1BWP12T U3838 ( .A1(n6852), .A2(n6851), .B(n6850), .C(n6849), .ZN(
        n6853) );
  AOI211D1BWP12T U3839 ( .A1(n6856), .A2(n6855), .B(n6854), .C(n6853), .ZN(
        n6860) );
  CKND2D1BWP12T U3840 ( .A1(n6858), .A2(n6857), .ZN(n6859) );
  OAI211D1BWP12T U3841 ( .A1(n6862), .A2(n6861), .B(n6860), .C(n6859), .ZN(
        n6863) );
  AOI211D1BWP12T U3842 ( .A1(n6870), .A2(n6865), .B(n6864), .C(n6863), .ZN(
        n6866) );
  OAI211D1BWP12T U3843 ( .A1(n6868), .A2(n6890), .B(n6867), .C(n6866), .ZN(
        result[29]) );
  INVD1BWP12T U3844 ( .I(n6869), .ZN(n6903) );
  TPNR2D0BWP12T U3845 ( .A1(n6875), .A2(n6874), .ZN(n6876) );
  AO211D1BWP12T U3846 ( .A1(n6879), .A2(n6878), .B(n6877), .C(n6876), .Z(n6885) );
  OAI22D0BWP12T U3847 ( .A1(n6883), .A2(n6882), .B1(n6881), .B2(n6880), .ZN(
        n6884) );
  RCAOI211D0BWP12T U3848 ( .A1(n6887), .A2(n6886), .B(n6885), .C(n6884), .ZN(
        n6889) );
  OAI22D1BWP12T U3849 ( .A1(n6895), .A2(n6894), .B1(n6893), .B2(n6892), .ZN(
        n6896) );
  AOI211D1BWP12T U3850 ( .A1(n6899), .A2(n6898), .B(n6897), .C(n6896), .ZN(
        n6900) );
  OAI211D1BWP12T U3851 ( .A1(n6903), .A2(n6902), .B(n6901), .C(n6900), .ZN(
        n6904) );
  AOI21D1BWP12T U3852 ( .A1(n6906), .A2(n6905), .B(n6904), .ZN(n6907) );
endmodule


module top7 ( clock, reset, MEM_MEMCTRL_from_mem_data, 
        MEMCTRL_MEM_to_mem_read_enable, MEMCTRL_MEM_to_mem_write_enable, 
        MEMCTRL_MEM_to_mem_mem_enable, MEMCTRL_MEM_to_mem_address, 
        MEMCTRL_MEM_to_mem_data );
  input [15:0] MEM_MEMCTRL_from_mem_data;
  output [11:0] MEMCTRL_MEM_to_mem_address;
  output [15:0] MEMCTRL_MEM_to_mem_data;
  input clock, reset;
  output MEMCTRL_MEM_to_mem_read_enable, MEMCTRL_MEM_to_mem_write_enable,
         MEMCTRL_MEM_to_mem_mem_enable;
  wire   ALU_OUT_n, ALU_OUT_c, ALU_OUT_z, ALU_OUT_v, ALU_IN_c,
         memory_interface_inst1_fsm_state_3_,
         memory_interface_inst1_fsm_state_2_,
         memory_interface_inst1_fsm_state_1_,
         memory_interface_inst1_fsm_state_0_, memory_interface_inst1_fsm_N32,
         memory_interface_inst1_fsm_N33, memory_interface_inst1_fsm_N34,
         memory_interface_inst1_fsm_N35,
         memory_interface_inst1_delayed_is_signed,
         memory_interface_inst1_delay_addr_for_adder_0_,
         memory_interface_inst1_delay_addr_for_adder_1_,
         memory_interface_inst1_delay_addr_for_adder_2_,
         memory_interface_inst1_delay_addr_for_adder_3_,
         memory_interface_inst1_delay_addr_for_adder_4_,
         memory_interface_inst1_delay_addr_for_adder_5_,
         memory_interface_inst1_delay_addr_for_adder_6_,
         memory_interface_inst1_delay_addr_for_adder_7_,
         memory_interface_inst1_delay_addr_for_adder_8_,
         memory_interface_inst1_delay_addr_for_adder_9_,
         memory_interface_inst1_delay_addr_for_adder_10_,
         memory_interface_inst1_delay_addr_for_adder_11_,
         register_file_inst1_n2648, register_file_inst1_n2647,
         register_file_inst1_n2646, register_file_inst1_n2645,
         register_file_inst1_n2644, register_file_inst1_n2643,
         register_file_inst1_n2642, register_file_inst1_n2641,
         register_file_inst1_n2640, register_file_inst1_n2639,
         register_file_inst1_n2638, register_file_inst1_n2637,
         register_file_inst1_n2636, register_file_inst1_n2635,
         register_file_inst1_n2634, register_file_inst1_n2633,
         register_file_inst1_n2632, register_file_inst1_n2631,
         register_file_inst1_n2630, register_file_inst1_n2629,
         register_file_inst1_n2628, register_file_inst1_n2627,
         register_file_inst1_n2626, register_file_inst1_n2625,
         register_file_inst1_n2624, register_file_inst1_n2623,
         register_file_inst1_n2622, register_file_inst1_n2621,
         register_file_inst1_n2620, register_file_inst1_n2619,
         register_file_inst1_n2618, register_file_inst1_n2617,
         register_file_inst1_n2616, register_file_inst1_n2615,
         register_file_inst1_n2614, register_file_inst1_n2613,
         register_file_inst1_n2612, register_file_inst1_n2611,
         register_file_inst1_n2610, register_file_inst1_n2609,
         register_file_inst1_n2608, register_file_inst1_n2607,
         register_file_inst1_n2606, register_file_inst1_n2605,
         register_file_inst1_n2604, register_file_inst1_n2603,
         register_file_inst1_n2602, register_file_inst1_n2601,
         register_file_inst1_n2600, register_file_inst1_n2599,
         register_file_inst1_n2598, register_file_inst1_n2597,
         register_file_inst1_n2596, register_file_inst1_n2595,
         register_file_inst1_n2594, register_file_inst1_n2593,
         register_file_inst1_n2592, register_file_inst1_n2591,
         register_file_inst1_n2590, register_file_inst1_n2589,
         register_file_inst1_n2588, register_file_inst1_n2587,
         register_file_inst1_n2586, register_file_inst1_n2585,
         register_file_inst1_n2584, register_file_inst1_n2583,
         register_file_inst1_n2582, register_file_inst1_n2581,
         register_file_inst1_n2580, register_file_inst1_n2579,
         register_file_inst1_n2578, register_file_inst1_n2577,
         register_file_inst1_n2576, register_file_inst1_n2575,
         register_file_inst1_n2574, register_file_inst1_n2573,
         register_file_inst1_n2572, register_file_inst1_n2571,
         register_file_inst1_n2570, register_file_inst1_n2569,
         register_file_inst1_n2568, register_file_inst1_n2567,
         register_file_inst1_n2566, register_file_inst1_n2565,
         register_file_inst1_n2564, register_file_inst1_n2563,
         register_file_inst1_n2562, register_file_inst1_n2561,
         register_file_inst1_n2560, register_file_inst1_n2559,
         register_file_inst1_n2558, register_file_inst1_n2557,
         register_file_inst1_n2556, register_file_inst1_n2555,
         register_file_inst1_n2554, register_file_inst1_n2553,
         register_file_inst1_n2552, register_file_inst1_n2551,
         register_file_inst1_n2550, register_file_inst1_n2549,
         register_file_inst1_n2548, register_file_inst1_n2547,
         register_file_inst1_n2546, register_file_inst1_n2545,
         register_file_inst1_n2544, register_file_inst1_n2543,
         register_file_inst1_n2542, register_file_inst1_n2541,
         register_file_inst1_n2540, register_file_inst1_n2539,
         register_file_inst1_n2538, register_file_inst1_n2537,
         register_file_inst1_n2536, register_file_inst1_n2535,
         register_file_inst1_n2534, register_file_inst1_n2533,
         register_file_inst1_n2532, register_file_inst1_n2531,
         register_file_inst1_n2530, register_file_inst1_n2529,
         register_file_inst1_n2528, register_file_inst1_n2527,
         register_file_inst1_n2526, register_file_inst1_n2525,
         register_file_inst1_n2524, register_file_inst1_n2523,
         register_file_inst1_n2522, register_file_inst1_n2521,
         register_file_inst1_n2520, register_file_inst1_n2519,
         register_file_inst1_n2518, register_file_inst1_n2517,
         register_file_inst1_n2516, register_file_inst1_n2515,
         register_file_inst1_n2514, register_file_inst1_n2513,
         register_file_inst1_n2512, register_file_inst1_n2511,
         register_file_inst1_n2510, register_file_inst1_n2509,
         register_file_inst1_n2508, register_file_inst1_n2507,
         register_file_inst1_n2506, register_file_inst1_n2505,
         register_file_inst1_n2504, register_file_inst1_n2503,
         register_file_inst1_n2502, register_file_inst1_n2501,
         register_file_inst1_n2500, register_file_inst1_n2499,
         register_file_inst1_n2498, register_file_inst1_n2497,
         register_file_inst1_n2496, register_file_inst1_n2495,
         register_file_inst1_n2494, register_file_inst1_n2493,
         register_file_inst1_n2492, register_file_inst1_n2491,
         register_file_inst1_n2490, register_file_inst1_n2489,
         register_file_inst1_n2488, register_file_inst1_n2487,
         register_file_inst1_n2486, register_file_inst1_n2485,
         register_file_inst1_n2484, register_file_inst1_n2483,
         register_file_inst1_n2482, register_file_inst1_n2481,
         register_file_inst1_n2480, register_file_inst1_n2479,
         register_file_inst1_n2478, register_file_inst1_n2477,
         register_file_inst1_n2476, register_file_inst1_n2475,
         register_file_inst1_n2474, register_file_inst1_n2473,
         register_file_inst1_n2472, register_file_inst1_n2471,
         register_file_inst1_n2470, register_file_inst1_n2469,
         register_file_inst1_n2468, register_file_inst1_n2467,
         register_file_inst1_n2466, register_file_inst1_n2465,
         register_file_inst1_n2464, register_file_inst1_n2463,
         register_file_inst1_n2462, register_file_inst1_n2461,
         register_file_inst1_n2460, register_file_inst1_n2459,
         register_file_inst1_n2458, register_file_inst1_n2457,
         register_file_inst1_n2456, register_file_inst1_n2455,
         register_file_inst1_n2454, register_file_inst1_n2453,
         register_file_inst1_n2452, register_file_inst1_n2451,
         register_file_inst1_n2450, register_file_inst1_n2449,
         register_file_inst1_n2448, register_file_inst1_n2447,
         register_file_inst1_n2446, register_file_inst1_n2445,
         register_file_inst1_n2444, register_file_inst1_n2443,
         register_file_inst1_n2442, register_file_inst1_n2441,
         register_file_inst1_n2440, register_file_inst1_n2439,
         register_file_inst1_n2438, register_file_inst1_n2437,
         register_file_inst1_n2436, register_file_inst1_n2435,
         register_file_inst1_n2434, register_file_inst1_n2433,
         register_file_inst1_n2432, register_file_inst1_n2431,
         register_file_inst1_n2430, register_file_inst1_n2429,
         register_file_inst1_n2428, register_file_inst1_n2427,
         register_file_inst1_n2426, register_file_inst1_n2425,
         register_file_inst1_n2424, register_file_inst1_n2423,
         register_file_inst1_n2422, register_file_inst1_n2421,
         register_file_inst1_n2420, register_file_inst1_n2419,
         register_file_inst1_n2418, register_file_inst1_n2417,
         register_file_inst1_n2416, register_file_inst1_n2415,
         register_file_inst1_n2414, register_file_inst1_n2413,
         register_file_inst1_n2412, register_file_inst1_n2411,
         register_file_inst1_n2410, register_file_inst1_n2409,
         register_file_inst1_n2408, register_file_inst1_n2407,
         register_file_inst1_n2406, register_file_inst1_n2405,
         register_file_inst1_n2404, register_file_inst1_n2403,
         register_file_inst1_n2402, register_file_inst1_n2401,
         register_file_inst1_n2400, register_file_inst1_n2399,
         register_file_inst1_n2398, register_file_inst1_n2397,
         register_file_inst1_n2396, register_file_inst1_n2395,
         register_file_inst1_n2394, register_file_inst1_n2393,
         register_file_inst1_n2392, register_file_inst1_n2391,
         register_file_inst1_n2390, register_file_inst1_n2389,
         register_file_inst1_n2388, register_file_inst1_n2387,
         register_file_inst1_n2386, register_file_inst1_n2385,
         register_file_inst1_n2384, register_file_inst1_n2383,
         register_file_inst1_n2382, register_file_inst1_n2381,
         register_file_inst1_n2380, register_file_inst1_n2379,
         register_file_inst1_n2378, register_file_inst1_n2377,
         register_file_inst1_n2376, register_file_inst1_n2375,
         register_file_inst1_n2374, register_file_inst1_n2373,
         register_file_inst1_n2372, register_file_inst1_n2371,
         register_file_inst1_n2370, register_file_inst1_n2369,
         register_file_inst1_n2368, register_file_inst1_n2367,
         register_file_inst1_n2366, register_file_inst1_n2365,
         register_file_inst1_n2364, register_file_inst1_n2363,
         register_file_inst1_n2362, register_file_inst1_n2361,
         register_file_inst1_n2360, register_file_inst1_n2359,
         register_file_inst1_n2358, register_file_inst1_n2357,
         register_file_inst1_n2356, register_file_inst1_n2355,
         register_file_inst1_n2354, register_file_inst1_n2353,
         register_file_inst1_n2352, register_file_inst1_n2351,
         register_file_inst1_n2350, register_file_inst1_n2349,
         register_file_inst1_n2348, register_file_inst1_n2347,
         register_file_inst1_n2346, register_file_inst1_n2345,
         register_file_inst1_n2344, register_file_inst1_n2343,
         register_file_inst1_n2342, register_file_inst1_n2341,
         register_file_inst1_n2340, register_file_inst1_n2339,
         register_file_inst1_n2338, register_file_inst1_n2337,
         register_file_inst1_n2336, register_file_inst1_n2335,
         register_file_inst1_n2334, register_file_inst1_n2333,
         register_file_inst1_n2332, register_file_inst1_n2331,
         register_file_inst1_n2330, register_file_inst1_n2329,
         register_file_inst1_n2328, register_file_inst1_n2327,
         register_file_inst1_n2326, register_file_inst1_n2325,
         register_file_inst1_n2324, register_file_inst1_n2323,
         register_file_inst1_n2322, register_file_inst1_n2321,
         register_file_inst1_n2320, register_file_inst1_n2319,
         register_file_inst1_n2318, register_file_inst1_n2317,
         register_file_inst1_n2316, register_file_inst1_n2315,
         register_file_inst1_n2314, register_file_inst1_n2313,
         register_file_inst1_n2312, register_file_inst1_n2311,
         register_file_inst1_n2310, register_file_inst1_n2309,
         register_file_inst1_n2308, register_file_inst1_n2307,
         register_file_inst1_n2306, register_file_inst1_n2305,
         register_file_inst1_n2304, register_file_inst1_n2303,
         register_file_inst1_n2302, register_file_inst1_n2301,
         register_file_inst1_n2300, register_file_inst1_n2299,
         register_file_inst1_n2298, register_file_inst1_n2297,
         register_file_inst1_n2296, register_file_inst1_n2295,
         register_file_inst1_n2294, register_file_inst1_n2293,
         register_file_inst1_n2292, register_file_inst1_n2291,
         register_file_inst1_n2290, register_file_inst1_n2289,
         register_file_inst1_n2288, register_file_inst1_n2287,
         register_file_inst1_n2286, register_file_inst1_n2285,
         register_file_inst1_n2284, register_file_inst1_n2283,
         register_file_inst1_n2282, register_file_inst1_n2281,
         register_file_inst1_n2280, register_file_inst1_n2279,
         register_file_inst1_n2278, register_file_inst1_n2277,
         register_file_inst1_n2276, register_file_inst1_n2275,
         register_file_inst1_n2274, register_file_inst1_n2273,
         register_file_inst1_n2272, register_file_inst1_n2271,
         register_file_inst1_n2270, register_file_inst1_n2269,
         register_file_inst1_n2268, register_file_inst1_n2267,
         register_file_inst1_n2266, register_file_inst1_n2265,
         register_file_inst1_n2264, register_file_inst1_n2263,
         register_file_inst1_n2262, register_file_inst1_n2261,
         register_file_inst1_n2260, register_file_inst1_n2259,
         register_file_inst1_n2258, register_file_inst1_n2257,
         register_file_inst1_n2256, register_file_inst1_n2255,
         register_file_inst1_n2254, register_file_inst1_n2253,
         register_file_inst1_n2252, register_file_inst1_n2251,
         register_file_inst1_n2250, register_file_inst1_n2249,
         register_file_inst1_n2248, register_file_inst1_n2247,
         register_file_inst1_n2246, register_file_inst1_n2245,
         register_file_inst1_n2244, register_file_inst1_n2243,
         register_file_inst1_n2242, register_file_inst1_n2241,
         register_file_inst1_n2240, register_file_inst1_n2239,
         register_file_inst1_n2238, register_file_inst1_n2237,
         register_file_inst1_n2236, register_file_inst1_n2235,
         register_file_inst1_n2234, register_file_inst1_n2233,
         register_file_inst1_n2232, register_file_inst1_n2231,
         register_file_inst1_n2230, register_file_inst1_n2229,
         register_file_inst1_n2228, register_file_inst1_n2227,
         register_file_inst1_n2226, register_file_inst1_n2225,
         register_file_inst1_n2224, register_file_inst1_n2223,
         register_file_inst1_n2222, register_file_inst1_n2221,
         register_file_inst1_n2220, register_file_inst1_n2219,
         register_file_inst1_n2218, register_file_inst1_n2217,
         register_file_inst1_n2216, register_file_inst1_n2215,
         register_file_inst1_n2214, register_file_inst1_n2213,
         register_file_inst1_n2212, register_file_inst1_n2211,
         register_file_inst1_n2210, register_file_inst1_n2209,
         register_file_inst1_n2208, register_file_inst1_n2207,
         register_file_inst1_n2206, register_file_inst1_n2205,
         register_file_inst1_n2204, register_file_inst1_n2203,
         register_file_inst1_n2202, register_file_inst1_n2201,
         register_file_inst1_n2200, register_file_inst1_n2199,
         register_file_inst1_n2198, register_file_inst1_n2197,
         register_file_inst1_n2196, register_file_inst1_n2195,
         register_file_inst1_n2194, register_file_inst1_n2193,
         register_file_inst1_n2192, register_file_inst1_n2191,
         register_file_inst1_n2190, register_file_inst1_n2189,
         register_file_inst1_n2188, register_file_inst1_n2187,
         register_file_inst1_n2186, register_file_inst1_n2185,
         register_file_inst1_n2184, register_file_inst1_n2183,
         register_file_inst1_n2182, register_file_inst1_n2181,
         register_file_inst1_n2180, register_file_inst1_n2179,
         register_file_inst1_n2178, register_file_inst1_n2177,
         register_file_inst1_n2176, register_file_inst1_n2175,
         register_file_inst1_n2174, register_file_inst1_n2173,
         register_file_inst1_n2172, register_file_inst1_n2171,
         register_file_inst1_n2170, register_file_inst1_n2169,
         register_file_inst1_n2168, register_file_inst1_n2167,
         register_file_inst1_n2166, register_file_inst1_n2165,
         register_file_inst1_n2164, register_file_inst1_n2163,
         register_file_inst1_n2162, register_file_inst1_n2161,
         register_file_inst1_n2160, register_file_inst1_n2159,
         register_file_inst1_n2158, register_file_inst1_n2157,
         register_file_inst1_n2156, register_file_inst1_n2155,
         register_file_inst1_n2154, register_file_inst1_n2153,
         register_file_inst1_n2152, register_file_inst1_n2151,
         register_file_inst1_n2150, register_file_inst1_n2149,
         register_file_inst1_n2148, register_file_inst1_n2147,
         register_file_inst1_n2146, register_file_inst1_n2145,
         register_file_inst1_n2144, register_file_inst1_n2143,
         register_file_inst1_n2142, register_file_inst1_n2141,
         register_file_inst1_n2140, register_file_inst1_n2139,
         register_file_inst1_n2138, register_file_inst1_n2136,
         register_file_inst1_tmp1_0_, register_file_inst1_tmp1_1_,
         register_file_inst1_tmp1_2_, register_file_inst1_tmp1_3_,
         register_file_inst1_tmp1_4_, register_file_inst1_tmp1_5_,
         register_file_inst1_tmp1_6_, register_file_inst1_tmp1_7_,
         register_file_inst1_tmp1_8_, register_file_inst1_tmp1_9_,
         register_file_inst1_tmp1_10_, register_file_inst1_tmp1_11_,
         register_file_inst1_tmp1_12_, register_file_inst1_tmp1_13_,
         register_file_inst1_tmp1_14_, register_file_inst1_tmp1_15_,
         register_file_inst1_tmp1_16_, register_file_inst1_tmp1_17_,
         register_file_inst1_tmp1_18_, register_file_inst1_tmp1_19_,
         register_file_inst1_tmp1_20_, register_file_inst1_tmp1_21_,
         register_file_inst1_tmp1_22_, register_file_inst1_tmp1_23_,
         register_file_inst1_tmp1_24_, register_file_inst1_tmp1_25_,
         register_file_inst1_tmp1_26_, register_file_inst1_tmp1_27_,
         register_file_inst1_tmp1_28_, register_file_inst1_tmp1_29_,
         register_file_inst1_tmp1_30_, register_file_inst1_tmp1_31_,
         register_file_inst1_lr_0_, register_file_inst1_lr_1_,
         register_file_inst1_lr_2_, register_file_inst1_lr_3_,
         register_file_inst1_lr_4_, register_file_inst1_lr_5_,
         register_file_inst1_lr_6_, register_file_inst1_lr_7_,
         register_file_inst1_lr_8_, register_file_inst1_lr_9_,
         register_file_inst1_lr_10_, register_file_inst1_lr_11_,
         register_file_inst1_lr_12_, register_file_inst1_lr_13_,
         register_file_inst1_lr_14_, register_file_inst1_lr_15_,
         register_file_inst1_lr_16_, register_file_inst1_lr_17_,
         register_file_inst1_lr_18_, register_file_inst1_lr_19_,
         register_file_inst1_lr_20_, register_file_inst1_lr_21_,
         register_file_inst1_lr_22_, register_file_inst1_lr_23_,
         register_file_inst1_lr_24_, register_file_inst1_lr_25_,
         register_file_inst1_lr_26_, register_file_inst1_lr_27_,
         register_file_inst1_lr_28_, register_file_inst1_lr_29_,
         register_file_inst1_lr_30_, register_file_inst1_lr_31_,
         register_file_inst1_r12_0_, register_file_inst1_r12_1_,
         register_file_inst1_r12_2_, register_file_inst1_r12_3_,
         register_file_inst1_r12_4_, register_file_inst1_r12_5_,
         register_file_inst1_r12_6_, register_file_inst1_r12_7_,
         register_file_inst1_r12_8_, register_file_inst1_r12_9_,
         register_file_inst1_r12_10_, register_file_inst1_r12_11_,
         register_file_inst1_r12_12_, register_file_inst1_r12_13_,
         register_file_inst1_r12_14_, register_file_inst1_r12_15_,
         register_file_inst1_r12_16_, register_file_inst1_r12_17_,
         register_file_inst1_r12_18_, register_file_inst1_r12_19_,
         register_file_inst1_r12_20_, register_file_inst1_r12_21_,
         register_file_inst1_r12_22_, register_file_inst1_r12_23_,
         register_file_inst1_r12_24_, register_file_inst1_r12_25_,
         register_file_inst1_r12_26_, register_file_inst1_r12_27_,
         register_file_inst1_r12_28_, register_file_inst1_r12_29_,
         register_file_inst1_r12_30_, register_file_inst1_r12_31_,
         register_file_inst1_r11_0_, register_file_inst1_r11_1_,
         register_file_inst1_r11_2_, register_file_inst1_r11_3_,
         register_file_inst1_r11_4_, register_file_inst1_r11_5_,
         register_file_inst1_r11_6_, register_file_inst1_r11_7_,
         register_file_inst1_r11_8_, register_file_inst1_r11_9_,
         register_file_inst1_r11_10_, register_file_inst1_r11_11_,
         register_file_inst1_r11_12_, register_file_inst1_r11_13_,
         register_file_inst1_r11_14_, register_file_inst1_r11_15_,
         register_file_inst1_r11_16_, register_file_inst1_r11_17_,
         register_file_inst1_r11_18_, register_file_inst1_r11_19_,
         register_file_inst1_r11_20_, register_file_inst1_r11_21_,
         register_file_inst1_r11_22_, register_file_inst1_r11_23_,
         register_file_inst1_r11_24_, register_file_inst1_r11_25_,
         register_file_inst1_r11_26_, register_file_inst1_r11_27_,
         register_file_inst1_r11_28_, register_file_inst1_r11_29_,
         register_file_inst1_r11_30_, register_file_inst1_r11_31_,
         register_file_inst1_r10_0_, register_file_inst1_r10_1_,
         register_file_inst1_r10_2_, register_file_inst1_r10_3_,
         register_file_inst1_r10_4_, register_file_inst1_r10_5_,
         register_file_inst1_r10_6_, register_file_inst1_r10_7_,
         register_file_inst1_r10_8_, register_file_inst1_r10_9_,
         register_file_inst1_r10_10_, register_file_inst1_r10_11_,
         register_file_inst1_r10_12_, register_file_inst1_r10_13_,
         register_file_inst1_r10_14_, register_file_inst1_r10_15_,
         register_file_inst1_r10_16_, register_file_inst1_r10_17_,
         register_file_inst1_r10_18_, register_file_inst1_r10_19_,
         register_file_inst1_r10_20_, register_file_inst1_r10_21_,
         register_file_inst1_r10_22_, register_file_inst1_r10_23_,
         register_file_inst1_r10_24_, register_file_inst1_r10_25_,
         register_file_inst1_r10_26_, register_file_inst1_r10_27_,
         register_file_inst1_r10_28_, register_file_inst1_r10_29_,
         register_file_inst1_r10_30_, register_file_inst1_r10_31_,
         register_file_inst1_r9_0_, register_file_inst1_r9_1_,
         register_file_inst1_r9_2_, register_file_inst1_r9_3_,
         register_file_inst1_r9_4_, register_file_inst1_r9_5_,
         register_file_inst1_r9_6_, register_file_inst1_r9_7_,
         register_file_inst1_r9_8_, register_file_inst1_r9_9_,
         register_file_inst1_r9_10_, register_file_inst1_r9_11_,
         register_file_inst1_r9_12_, register_file_inst1_r9_13_,
         register_file_inst1_r9_14_, register_file_inst1_r9_15_,
         register_file_inst1_r9_16_, register_file_inst1_r9_17_,
         register_file_inst1_r9_18_, register_file_inst1_r9_19_,
         register_file_inst1_r9_20_, register_file_inst1_r9_21_,
         register_file_inst1_r9_22_, register_file_inst1_r9_23_,
         register_file_inst1_r9_24_, register_file_inst1_r9_25_,
         register_file_inst1_r9_26_, register_file_inst1_r9_27_,
         register_file_inst1_r9_28_, register_file_inst1_r9_29_,
         register_file_inst1_r9_30_, register_file_inst1_r9_31_,
         register_file_inst1_r8_0_, register_file_inst1_r8_1_,
         register_file_inst1_r8_2_, register_file_inst1_r8_3_,
         register_file_inst1_r8_4_, register_file_inst1_r8_5_,
         register_file_inst1_r8_6_, register_file_inst1_r8_7_,
         register_file_inst1_r8_8_, register_file_inst1_r8_9_,
         register_file_inst1_r8_10_, register_file_inst1_r8_11_,
         register_file_inst1_r8_12_, register_file_inst1_r8_13_,
         register_file_inst1_r8_14_, register_file_inst1_r8_15_,
         register_file_inst1_r8_16_, register_file_inst1_r8_17_,
         register_file_inst1_r8_18_, register_file_inst1_r8_19_,
         register_file_inst1_r8_20_, register_file_inst1_r8_21_,
         register_file_inst1_r8_22_, register_file_inst1_r8_23_,
         register_file_inst1_r8_24_, register_file_inst1_r8_25_,
         register_file_inst1_r8_26_, register_file_inst1_r8_27_,
         register_file_inst1_r8_28_, register_file_inst1_r8_29_,
         register_file_inst1_r8_30_, register_file_inst1_r8_31_,
         register_file_inst1_r7_0_, register_file_inst1_r7_1_,
         register_file_inst1_r7_2_, register_file_inst1_r7_3_,
         register_file_inst1_r7_4_, register_file_inst1_r7_5_,
         register_file_inst1_r7_6_, register_file_inst1_r7_7_,
         register_file_inst1_r7_8_, register_file_inst1_r7_9_,
         register_file_inst1_r7_10_, register_file_inst1_r7_11_,
         register_file_inst1_r7_12_, register_file_inst1_r7_13_,
         register_file_inst1_r7_14_, register_file_inst1_r7_15_,
         register_file_inst1_r7_16_, register_file_inst1_r7_17_,
         register_file_inst1_r7_18_, register_file_inst1_r7_19_,
         register_file_inst1_r7_20_, register_file_inst1_r7_21_,
         register_file_inst1_r7_22_, register_file_inst1_r7_23_,
         register_file_inst1_r7_24_, register_file_inst1_r7_25_,
         register_file_inst1_r7_26_, register_file_inst1_r7_27_,
         register_file_inst1_r7_28_, register_file_inst1_r7_29_,
         register_file_inst1_r7_30_, register_file_inst1_r7_31_,
         register_file_inst1_r6_0_, register_file_inst1_r6_1_,
         register_file_inst1_r6_2_, register_file_inst1_r6_3_,
         register_file_inst1_r6_4_, register_file_inst1_r6_5_,
         register_file_inst1_r6_6_, register_file_inst1_r6_7_,
         register_file_inst1_r6_8_, register_file_inst1_r6_9_,
         register_file_inst1_r6_10_, register_file_inst1_r6_11_,
         register_file_inst1_r6_12_, register_file_inst1_r6_13_,
         register_file_inst1_r6_14_, register_file_inst1_r6_15_,
         register_file_inst1_r6_16_, register_file_inst1_r6_17_,
         register_file_inst1_r6_18_, register_file_inst1_r6_19_,
         register_file_inst1_r6_20_, register_file_inst1_r6_21_,
         register_file_inst1_r6_22_, register_file_inst1_r6_23_,
         register_file_inst1_r6_24_, register_file_inst1_r6_25_,
         register_file_inst1_r6_26_, register_file_inst1_r6_27_,
         register_file_inst1_r6_28_, register_file_inst1_r6_29_,
         register_file_inst1_r6_30_, register_file_inst1_r6_31_,
         register_file_inst1_r5_0_, register_file_inst1_r5_1_,
         register_file_inst1_r5_2_, register_file_inst1_r5_3_,
         register_file_inst1_r5_4_, register_file_inst1_r5_5_,
         register_file_inst1_r5_6_, register_file_inst1_r5_7_,
         register_file_inst1_r5_8_, register_file_inst1_r5_9_,
         register_file_inst1_r5_10_, register_file_inst1_r5_11_,
         register_file_inst1_r5_12_, register_file_inst1_r5_13_,
         register_file_inst1_r5_14_, register_file_inst1_r5_15_,
         register_file_inst1_r5_16_, register_file_inst1_r5_17_,
         register_file_inst1_r5_18_, register_file_inst1_r5_19_,
         register_file_inst1_r5_20_, register_file_inst1_r5_21_,
         register_file_inst1_r5_22_, register_file_inst1_r5_23_,
         register_file_inst1_r5_24_, register_file_inst1_r5_25_,
         register_file_inst1_r5_26_, register_file_inst1_r5_27_,
         register_file_inst1_r5_28_, register_file_inst1_r5_29_,
         register_file_inst1_r5_30_, register_file_inst1_r5_31_,
         register_file_inst1_r4_0_, register_file_inst1_r4_1_,
         register_file_inst1_r4_2_, register_file_inst1_r4_3_,
         register_file_inst1_r4_4_, register_file_inst1_r4_5_,
         register_file_inst1_r4_6_, register_file_inst1_r4_7_,
         register_file_inst1_r4_8_, register_file_inst1_r4_9_,
         register_file_inst1_r4_10_, register_file_inst1_r4_11_,
         register_file_inst1_r4_12_, register_file_inst1_r4_13_,
         register_file_inst1_r4_14_, register_file_inst1_r4_15_,
         register_file_inst1_r4_16_, register_file_inst1_r4_17_,
         register_file_inst1_r4_18_, register_file_inst1_r4_19_,
         register_file_inst1_r4_20_, register_file_inst1_r4_21_,
         register_file_inst1_r4_22_, register_file_inst1_r4_23_,
         register_file_inst1_r4_24_, register_file_inst1_r4_25_,
         register_file_inst1_r4_26_, register_file_inst1_r4_27_,
         register_file_inst1_r4_28_, register_file_inst1_r4_29_,
         register_file_inst1_r4_30_, register_file_inst1_r4_31_,
         register_file_inst1_r3_0_, register_file_inst1_r3_1_,
         register_file_inst1_r3_2_, register_file_inst1_r3_3_,
         register_file_inst1_r3_4_, register_file_inst1_r3_5_,
         register_file_inst1_r3_6_, register_file_inst1_r3_7_,
         register_file_inst1_r3_8_, register_file_inst1_r3_9_,
         register_file_inst1_r3_10_, register_file_inst1_r3_11_,
         register_file_inst1_r3_12_, register_file_inst1_r3_13_,
         register_file_inst1_r3_14_, register_file_inst1_r3_15_,
         register_file_inst1_r3_16_, register_file_inst1_r3_17_,
         register_file_inst1_r3_18_, register_file_inst1_r3_19_,
         register_file_inst1_r3_20_, register_file_inst1_r3_21_,
         register_file_inst1_r3_22_, register_file_inst1_r3_23_,
         register_file_inst1_r3_24_, register_file_inst1_r3_25_,
         register_file_inst1_r3_26_, register_file_inst1_r3_27_,
         register_file_inst1_r3_28_, register_file_inst1_r3_29_,
         register_file_inst1_r3_30_, register_file_inst1_r3_31_,
         register_file_inst1_r2_0_, register_file_inst1_r2_1_,
         register_file_inst1_r2_2_, register_file_inst1_r2_3_,
         register_file_inst1_r2_4_, register_file_inst1_r2_5_,
         register_file_inst1_r2_6_, register_file_inst1_r2_7_,
         register_file_inst1_r2_8_, register_file_inst1_r2_9_,
         register_file_inst1_r2_10_, register_file_inst1_r2_11_,
         register_file_inst1_r2_12_, register_file_inst1_r2_13_,
         register_file_inst1_r2_14_, register_file_inst1_r2_15_,
         register_file_inst1_r2_16_, register_file_inst1_r2_17_,
         register_file_inst1_r2_18_, register_file_inst1_r2_19_,
         register_file_inst1_r2_20_, register_file_inst1_r2_21_,
         register_file_inst1_r2_22_, register_file_inst1_r2_23_,
         register_file_inst1_r2_24_, register_file_inst1_r2_25_,
         register_file_inst1_r2_26_, register_file_inst1_r2_27_,
         register_file_inst1_r2_28_, register_file_inst1_r2_29_,
         register_file_inst1_r2_30_, register_file_inst1_r2_31_,
         register_file_inst1_r1_0_, register_file_inst1_r1_1_,
         register_file_inst1_r1_2_, register_file_inst1_r1_3_,
         register_file_inst1_r1_4_, register_file_inst1_r1_5_,
         register_file_inst1_r1_6_, register_file_inst1_r1_7_,
         register_file_inst1_r1_8_, register_file_inst1_r1_9_,
         register_file_inst1_r1_10_, register_file_inst1_r1_11_,
         register_file_inst1_r1_12_, register_file_inst1_r1_13_,
         register_file_inst1_r1_14_, register_file_inst1_r1_15_,
         register_file_inst1_r1_16_, register_file_inst1_r1_17_,
         register_file_inst1_r1_18_, register_file_inst1_r1_19_,
         register_file_inst1_r1_20_, register_file_inst1_r1_21_,
         register_file_inst1_r1_22_, register_file_inst1_r1_23_,
         register_file_inst1_r1_24_, register_file_inst1_r1_25_,
         register_file_inst1_r1_26_, register_file_inst1_r1_27_,
         register_file_inst1_r1_28_, register_file_inst1_r1_29_,
         register_file_inst1_r1_30_, register_file_inst1_r1_31_,
         register_file_inst1_r0_0_, register_file_inst1_r0_1_,
         register_file_inst1_r0_2_, register_file_inst1_r0_3_,
         register_file_inst1_r0_4_, register_file_inst1_r0_5_,
         register_file_inst1_r0_6_, register_file_inst1_r0_7_,
         register_file_inst1_r0_8_, register_file_inst1_r0_9_,
         register_file_inst1_r0_10_, register_file_inst1_r0_11_,
         register_file_inst1_r0_12_, register_file_inst1_r0_13_,
         register_file_inst1_r0_14_, register_file_inst1_r0_15_,
         register_file_inst1_r0_16_, register_file_inst1_r0_17_,
         register_file_inst1_r0_18_, register_file_inst1_r0_19_,
         register_file_inst1_r0_20_, register_file_inst1_r0_21_,
         register_file_inst1_r0_22_, register_file_inst1_r0_23_,
         register_file_inst1_r0_24_, register_file_inst1_r0_25_,
         register_file_inst1_r0_26_, register_file_inst1_r0_27_,
         register_file_inst1_r0_28_, register_file_inst1_r0_29_,
         register_file_inst1_r0_30_, register_file_inst1_r0_31_, n2243, n2244,
         n2247, n2249, n2251, n2253, n2255, n2257, n2259, n2261, n2262, n2264,
         n2265, n2266, n2267, n2268, n2269, n2342, n2343, n2348, n2396, n2469,
         n2470, n2471, n2515, n2516, n2871, n2874, n2876, n2878, n2880, n2905,
         n2906, n2907, n2908, n2909, n2911, n2912, n2917, n2919, n2920, n3017,
         n3018, n3046, n3047, n3048, n3049, n3054, n3055, n3056, n3059, n3060,
         n3061, n3068, n3095, n3165, n3202, n3217, n3286, n3335, n3420, n3467,
         n3502, n3510, n3519, n3521, n3718, n4090, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407;
  wire   [31:0] ALU_MISC_OUT_result;
  wire   [31:0] RF_next_sp;
  wire   [31:0] RF_ALU_operand_a;
  wire   [31:0] RF_ALU_operand_b;
  wire   [31:0] RF_MEMCTRL_data_reg;
  wire   [11:0] MEMCTRL_IN_address;
  wire   [15:0] memory_interface_inst1_delay_first_two_bytes_out;
  wire   [31:0] memory_interface_inst1_delay_data_in32;
  wire   [11:0] memory_interface_inst1_delay_addr_single;
  wire   [3:0] register_file_inst1_cpsrin;
  wire   [31:0] register_file_inst1_spin;
  tri   clock;
  tri   reset;
  tri   DEC_CPSR_update_flag_n;
  tri   RF_OUT_n;
  tri   DEC_CPSR_update_flag_c;
  tri   RF_OUT_c;
  tri   DEC_CPSR_update_flag_z;
  tri   RF_OUT_z;
  tri   DEC_CPSR_update_flag_v;
  tri   RF_OUT_v;
  tri   [31:0] IF_DEC_instruction;
  tri   IF_DEC_instruction_valid;
  tri   MEMCTRL_write_finished;
  tri   MEMCTRL_read_finished;
  tri   [4:0] DEC_RF_operand_a;
  tri   [4:0] DEC_RF_operand_b;
  tri   [31:0] DEC_RF_offset_a;
  tri   [31:0] DEC_RF_offset_b;
  tri   [4:0] DEC_ALU_alu_opcode;
  tri   [4:0] DEC_RF_alu_write_to_reg;
  tri   DEC_RF_alu_write_to_reg_enable;
  tri   [4:0] DEC_RF_memory_write_to_reg;
  tri   DEC_RF_memory_write_to_reg_enable;
  tri   [4:0] DEC_RF_memory_store_data_reg;
  tri   [4:0] DEC_RF_memory_store_address_reg;
  tri   DEC_MISC_OUT_memory_address_source_is_reg;
  tri   [1:0] DEC_MEMCTRL_load_store_width;
  tri   DEC_MEMCTRL_memorycontroller_sign_extend;
  tri   DEC_MEMCTRL_memory_load_request;
  tri   DEC_MEMCTRL_memory_store_request;
  tri   DEC_IF_stall_to_instructionfetch;
  tri   [15:0] MEMCTRL_RF_IF_data_in;
  tri   [31:0] IF_RF_incremented_pc_out;
  tri   IF_RF_incremented_pc_write_enable;
  tri   [31:0] RF_pc_out;
  tri   IF_memory_load_req;
  tri   [11:0] IF_instruction_memory_address;

  irdecode irdecode_inst1 ( .clock(clock), .reset(reset), .instruction(
        IF_DEC_instruction), .flag_n(RF_OUT_n), .flag_z(RF_OUT_z), .flag_c(
        RF_OUT_c), .flag_v(RF_OUT_v), .instruction_valid(
        IF_DEC_instruction_valid), .memory_write_finished(
        MEMCTRL_write_finished), .memory_read_finished(MEMCTRL_read_finished), 
        .operand_a(DEC_RF_operand_a), .operand_b(DEC_RF_operand_b), .offset_a(
        DEC_RF_offset_a), .offset_b(DEC_RF_offset_b), .alu_opcode(
        DEC_ALU_alu_opcode), .update_flag_n(DEC_CPSR_update_flag_n), 
        .update_flag_z(DEC_CPSR_update_flag_z), .update_flag_c(
        DEC_CPSR_update_flag_c), .update_flag_v(DEC_CPSR_update_flag_v), 
        .alu_write_to_reg(DEC_RF_alu_write_to_reg), .alu_write_to_reg_enable(
        DEC_RF_alu_write_to_reg_enable), .memory_write_to_reg(
        DEC_RF_memory_write_to_reg), .memory_write_to_reg_enable(
        DEC_RF_memory_write_to_reg_enable), .memory_store_data_reg(
        DEC_RF_memory_store_data_reg), .memory_store_address_reg(
        DEC_RF_memory_store_address_reg), .memory_address_source_is_reg(
        DEC_MISC_OUT_memory_address_source_is_reg), .load_store_width(
        DEC_MEMCTRL_load_store_width), .memorycontroller_sign_extend(
        DEC_MEMCTRL_memorycontroller_sign_extend), .memory_load_request(
        DEC_MEMCTRL_memory_load_request), .memory_store_request(
        DEC_MEMCTRL_memory_store_request), .stall_to_instructionfetch(
        DEC_IF_stall_to_instructionfetch) );
  ALU_VARIABLE ALU_VARIABLE_inst1 ( .a(RF_ALU_operand_a), .b(RF_ALU_operand_b), 
        .op(DEC_ALU_alu_opcode[3:0]), .c_in(ALU_IN_c), .result(
        ALU_MISC_OUT_result), .c_out(ALU_OUT_c), .z(ALU_OUT_z), .n(ALU_OUT_n), 
        .v(ALU_OUT_v) );
  Instruction_Fetch Instruction_Fetch_inst1 ( .clk(clock), .reset(reset), 
        .stall_decoder_in(DEC_IF_stall_to_instructionfetch), 
        .memory_output_valid(MEMCTRL_read_finished), .current_pc_in(RF_pc_out), 
        .instruction_in(MEMCTRL_RF_IF_data_in), .memory_load_request(
        IF_memory_load_req), .incremented_pc_write_enable(
        IF_RF_incremented_pc_write_enable), .memory_address(
        IF_instruction_memory_address), .incremented_pc_out(
        IF_RF_incremented_pc_out), .instruction_out(IF_DEC_instruction), 
        .instruction_valid(IF_DEC_instruction_valid) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_1_ ( .D(
        memory_interface_inst1_fsm_N33), .CP(clock), .Q(
        memory_interface_inst1_fsm_state_1_) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_2_ ( .D(
        memory_interface_inst1_fsm_N34), .CP(clock), .Q(
        memory_interface_inst1_fsm_state_2_) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_3_ ( .D(
        memory_interface_inst1_fsm_N35), .CP(clock), .Q(
        memory_interface_inst1_fsm_state_3_) );
  DFQD1BWP12T memory_interface_inst1_delayed_is_signed_reg ( .D(
        DEC_MEMCTRL_memorycontroller_sign_extend), .CP(clock), .Q(
        memory_interface_inst1_delayed_is_signed) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_0_ ( .D(
        MEMCTRL_IN_address[0]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[0]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_1_ ( .D(
        MEMCTRL_IN_address[1]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[1]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_2_ ( .D(
        MEMCTRL_IN_address[2]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_3_ ( .D(
        MEMCTRL_IN_address[3]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_4_ ( .D(
        MEMCTRL_IN_address[4]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[4]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_5_ ( .D(
        MEMCTRL_IN_address[5]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[5]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_6_ ( .D(
        MEMCTRL_IN_address[6]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_7_ ( .D(
        MEMCTRL_IN_address[7]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_8_ ( .D(
        MEMCTRL_IN_address[8]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_9_ ( .D(
        MEMCTRL_IN_address[9]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_10_ ( .D(
        MEMCTRL_IN_address[10]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_11_ ( .D(
        MEMCTRL_IN_address[11]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[11]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_0_ ( .D(
        MEMCTRL_IN_address[0]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_0_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_1_ ( .D(
        MEMCTRL_IN_address[1]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_1_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_2_ ( .D(
        MEMCTRL_IN_address[2]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_2_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_3_ ( .D(
        MEMCTRL_IN_address[3]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_3_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_4_ ( .D(
        MEMCTRL_IN_address[4]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_4_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_5_ ( .D(
        MEMCTRL_IN_address[5]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_5_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_6_ ( .D(
        MEMCTRL_IN_address[6]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_6_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_7_ ( .D(
        MEMCTRL_IN_address[7]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_7_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_8_ ( .D(
        MEMCTRL_IN_address[8]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_8_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_9_ ( .D(
        MEMCTRL_IN_address[9]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_9_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_10_ ( .D(
        MEMCTRL_IN_address[10]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_10_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_11_ ( .D(
        MEMCTRL_IN_address[11]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_11_) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_0_ ( .D(
        RF_MEMCTRL_data_reg[0]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[0]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_1_ ( .D(
        RF_MEMCTRL_data_reg[1]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[1]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_2_ ( .D(
        RF_MEMCTRL_data_reg[2]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_3_ ( .D(
        RF_MEMCTRL_data_reg[3]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_4_ ( .D(
        RF_MEMCTRL_data_reg[4]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[4]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_5_ ( .D(
        RF_MEMCTRL_data_reg[5]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[5]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_6_ ( .D(
        RF_MEMCTRL_data_reg[6]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_7_ ( .D(
        RF_MEMCTRL_data_reg[7]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_8_ ( .D(
        RF_MEMCTRL_data_reg[8]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_9_ ( .D(
        RF_MEMCTRL_data_reg[9]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_10_ ( .D(
        RF_MEMCTRL_data_reg[10]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_11_ ( .D(
        RF_MEMCTRL_data_reg[11]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[11]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_12_ ( .D(
        RF_MEMCTRL_data_reg[12]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[12]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_13_ ( .D(
        RF_MEMCTRL_data_reg[13]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[13]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_14_ ( .D(
        RF_MEMCTRL_data_reg[14]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[14]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_15_ ( .D(
        RF_MEMCTRL_data_reg[15]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[15]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_16_ ( .D(
        RF_MEMCTRL_data_reg[16]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[16]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_17_ ( .D(
        RF_MEMCTRL_data_reg[17]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[17]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_18_ ( .D(
        RF_MEMCTRL_data_reg[18]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[18]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_19_ ( .D(
        RF_MEMCTRL_data_reg[19]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[19]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_20_ ( .D(
        RF_MEMCTRL_data_reg[20]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[20]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_21_ ( .D(
        RF_MEMCTRL_data_reg[21]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[21]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_22_ ( .D(
        RF_MEMCTRL_data_reg[22]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[22]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_23_ ( .D(
        RF_MEMCTRL_data_reg[23]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[23]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_24_ ( .D(
        RF_MEMCTRL_data_reg[24]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[24]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_25_ ( .D(
        RF_MEMCTRL_data_reg[25]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[25]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_26_ ( .D(
        RF_MEMCTRL_data_reg[26]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[26]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_27_ ( .D(
        RF_MEMCTRL_data_reg[27]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[27]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_28_ ( .D(
        RF_MEMCTRL_data_reg[28]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[28]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_29_ ( .D(
        RF_MEMCTRL_data_reg[29]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[29]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_30_ ( .D(
        RF_MEMCTRL_data_reg[30]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[30]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_31_ ( .D(
        RF_MEMCTRL_data_reg[31]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[31]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_0_ ( .D(
        MEM_MEMCTRL_from_mem_data[8]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[0]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_1_ ( .D(
        MEM_MEMCTRL_from_mem_data[9]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[1]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_2_ ( .D(
        MEM_MEMCTRL_from_mem_data[10]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_3_ ( .D(
        MEM_MEMCTRL_from_mem_data[11]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_4_ ( .D(
        MEM_MEMCTRL_from_mem_data[12]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[4]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_5_ ( .D(
        MEM_MEMCTRL_from_mem_data[13]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[5]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_6_ ( .D(
        MEM_MEMCTRL_from_mem_data[14]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_7_ ( .D(
        MEM_MEMCTRL_from_mem_data[15]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_8_ ( .D(
        MEM_MEMCTRL_from_mem_data[0]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_9_ ( .D(
        MEM_MEMCTRL_from_mem_data[1]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_10_ ( .D(
        MEM_MEMCTRL_from_mem_data[2]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_11_ ( .D(
        MEM_MEMCTRL_from_mem_data[3]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[11]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_12_ ( .D(
        MEM_MEMCTRL_from_mem_data[4]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[12]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_13_ ( .D(
        MEM_MEMCTRL_from_mem_data[5]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[13]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_14_ ( .D(
        MEM_MEMCTRL_from_mem_data[6]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[14]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_15_ ( .D(
        MEM_MEMCTRL_from_mem_data[7]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[15]) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_0_ ( .D(register_file_inst1_n2136), 
        .CP(clock), .Q(register_file_inst1_tmp1_0_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_1_ ( .D(register_file_inst1_n2138), 
        .CP(clock), .Q(register_file_inst1_tmp1_1_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_2_ ( .D(register_file_inst1_n2139), 
        .CP(clock), .Q(register_file_inst1_tmp1_2_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_3_ ( .D(register_file_inst1_n2140), 
        .CP(clock), .Q(register_file_inst1_tmp1_3_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_4_ ( .D(register_file_inst1_n2141), 
        .CP(clock), .Q(register_file_inst1_tmp1_4_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_5_ ( .D(register_file_inst1_n2142), 
        .CP(clock), .Q(register_file_inst1_tmp1_5_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_6_ ( .D(register_file_inst1_n2143), 
        .CP(clock), .Q(register_file_inst1_tmp1_6_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_7_ ( .D(register_file_inst1_n2144), 
        .CP(clock), .Q(register_file_inst1_tmp1_7_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_8_ ( .D(register_file_inst1_n2145), 
        .CP(clock), .Q(register_file_inst1_tmp1_8_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_9_ ( .D(register_file_inst1_n2146), 
        .CP(clock), .Q(register_file_inst1_tmp1_9_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_10_ ( .D(register_file_inst1_n2147), 
        .CP(clock), .Q(register_file_inst1_tmp1_10_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_11_ ( .D(register_file_inst1_n2148), 
        .CP(clock), .Q(register_file_inst1_tmp1_11_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_12_ ( .D(register_file_inst1_n2149), 
        .CP(clock), .Q(register_file_inst1_tmp1_12_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_13_ ( .D(register_file_inst1_n2150), 
        .CP(clock), .Q(register_file_inst1_tmp1_13_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_14_ ( .D(register_file_inst1_n2151), 
        .CP(clock), .Q(register_file_inst1_tmp1_14_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_15_ ( .D(register_file_inst1_n2152), 
        .CP(clock), .Q(register_file_inst1_tmp1_15_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_16_ ( .D(register_file_inst1_n2153), 
        .CP(clock), .Q(register_file_inst1_tmp1_16_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_17_ ( .D(register_file_inst1_n2154), 
        .CP(clock), .Q(register_file_inst1_tmp1_17_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_18_ ( .D(register_file_inst1_n2155), 
        .CP(clock), .Q(register_file_inst1_tmp1_18_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_19_ ( .D(register_file_inst1_n2156), 
        .CP(clock), .Q(register_file_inst1_tmp1_19_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_20_ ( .D(register_file_inst1_n2157), 
        .CP(clock), .Q(register_file_inst1_tmp1_20_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_21_ ( .D(register_file_inst1_n2158), 
        .CP(clock), .Q(register_file_inst1_tmp1_21_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_22_ ( .D(register_file_inst1_n2159), 
        .CP(clock), .Q(register_file_inst1_tmp1_22_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_23_ ( .D(register_file_inst1_n2160), 
        .CP(clock), .Q(register_file_inst1_tmp1_23_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_24_ ( .D(register_file_inst1_n2161), 
        .CP(clock), .Q(register_file_inst1_tmp1_24_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_25_ ( .D(register_file_inst1_n2162), 
        .CP(clock), .Q(register_file_inst1_tmp1_25_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_26_ ( .D(register_file_inst1_n2163), 
        .CP(clock), .Q(register_file_inst1_tmp1_26_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_27_ ( .D(register_file_inst1_n2164), 
        .CP(clock), .Q(register_file_inst1_tmp1_27_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_28_ ( .D(register_file_inst1_n2165), 
        .CP(clock), .Q(register_file_inst1_tmp1_28_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_29_ ( .D(register_file_inst1_n2166), 
        .CP(clock), .Q(register_file_inst1_tmp1_29_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_30_ ( .D(register_file_inst1_n2167), 
        .CP(clock), .Q(register_file_inst1_tmp1_30_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_31_ ( .D(register_file_inst1_n2168), 
        .CP(clock), .Q(register_file_inst1_tmp1_31_) );
  DFQD1BWP12T register_file_inst1_cpsr_reg_0_ ( .D(
        register_file_inst1_cpsrin[0]), .CP(clock), .Q(RF_OUT_v) );
  DFQD1BWP12T register_file_inst1_cpsr_reg_1_ ( .D(
        register_file_inst1_cpsrin[1]), .CP(clock), .Q(RF_OUT_z) );
  DFQD1BWP12T register_file_inst1_cpsr_reg_2_ ( .D(
        register_file_inst1_cpsrin[2]), .CP(clock), .Q(RF_OUT_c) );
  DFQD1BWP12T register_file_inst1_cpsr_reg_3_ ( .D(
        register_file_inst1_cpsrin[3]), .CP(clock), .Q(RF_OUT_n) );
  DFQD1BWP12T register_file_inst1_pc_reg_0_ ( .D(register_file_inst1_n2169), 
        .CP(clock), .Q(RF_pc_out[0]) );
  DFQD1BWP12T register_file_inst1_pc_reg_1_ ( .D(register_file_inst1_n2170), 
        .CP(clock), .Q(RF_pc_out[1]) );
  DFQD1BWP12T register_file_inst1_pc_reg_2_ ( .D(register_file_inst1_n2171), 
        .CP(clock), .Q(RF_pc_out[2]) );
  DFQD1BWP12T register_file_inst1_pc_reg_3_ ( .D(register_file_inst1_n2172), 
        .CP(clock), .Q(RF_pc_out[3]) );
  DFQD1BWP12T register_file_inst1_pc_reg_4_ ( .D(register_file_inst1_n2173), 
        .CP(clock), .Q(RF_pc_out[4]) );
  DFQD1BWP12T register_file_inst1_pc_reg_5_ ( .D(register_file_inst1_n2174), 
        .CP(clock), .Q(RF_pc_out[5]) );
  DFQD1BWP12T register_file_inst1_pc_reg_6_ ( .D(register_file_inst1_n2175), 
        .CP(clock), .Q(RF_pc_out[6]) );
  DFQD1BWP12T register_file_inst1_pc_reg_7_ ( .D(register_file_inst1_n2176), 
        .CP(clock), .Q(RF_pc_out[7]) );
  DFQD1BWP12T register_file_inst1_pc_reg_8_ ( .D(register_file_inst1_n2177), 
        .CP(clock), .Q(RF_pc_out[8]) );
  DFQD1BWP12T register_file_inst1_pc_reg_9_ ( .D(register_file_inst1_n2178), 
        .CP(clock), .Q(RF_pc_out[9]) );
  DFQD1BWP12T register_file_inst1_pc_reg_10_ ( .D(register_file_inst1_n2179), 
        .CP(clock), .Q(RF_pc_out[10]) );
  DFQD1BWP12T register_file_inst1_pc_reg_11_ ( .D(register_file_inst1_n2180), 
        .CP(clock), .Q(RF_pc_out[11]) );
  DFQD1BWP12T register_file_inst1_pc_reg_12_ ( .D(register_file_inst1_n2181), 
        .CP(clock), .Q(RF_pc_out[12]) );
  DFQD1BWP12T register_file_inst1_pc_reg_13_ ( .D(register_file_inst1_n2182), 
        .CP(clock), .Q(RF_pc_out[13]) );
  DFQD1BWP12T register_file_inst1_pc_reg_14_ ( .D(register_file_inst1_n2183), 
        .CP(clock), .Q(RF_pc_out[14]) );
  DFQD1BWP12T register_file_inst1_pc_reg_15_ ( .D(register_file_inst1_n2184), 
        .CP(clock), .Q(RF_pc_out[15]) );
  DFQD1BWP12T register_file_inst1_pc_reg_16_ ( .D(register_file_inst1_n2185), 
        .CP(clock), .Q(RF_pc_out[16]) );
  DFQD1BWP12T register_file_inst1_pc_reg_17_ ( .D(register_file_inst1_n2186), 
        .CP(clock), .Q(RF_pc_out[17]) );
  DFQD1BWP12T register_file_inst1_pc_reg_18_ ( .D(register_file_inst1_n2187), 
        .CP(clock), .Q(RF_pc_out[18]) );
  DFQD1BWP12T register_file_inst1_pc_reg_19_ ( .D(register_file_inst1_n2188), 
        .CP(clock), .Q(RF_pc_out[19]) );
  DFQD1BWP12T register_file_inst1_pc_reg_20_ ( .D(register_file_inst1_n2189), 
        .CP(clock), .Q(RF_pc_out[20]) );
  DFQD1BWP12T register_file_inst1_pc_reg_21_ ( .D(register_file_inst1_n2190), 
        .CP(clock), .Q(RF_pc_out[21]) );
  DFQD1BWP12T register_file_inst1_pc_reg_22_ ( .D(register_file_inst1_n2191), 
        .CP(clock), .Q(RF_pc_out[22]) );
  DFQD1BWP12T register_file_inst1_pc_reg_23_ ( .D(register_file_inst1_n2192), 
        .CP(clock), .Q(RF_pc_out[23]) );
  DFQD1BWP12T register_file_inst1_pc_reg_24_ ( .D(register_file_inst1_n2193), 
        .CP(clock), .Q(RF_pc_out[24]) );
  DFQD1BWP12T register_file_inst1_pc_reg_25_ ( .D(register_file_inst1_n2194), 
        .CP(clock), .Q(RF_pc_out[25]) );
  DFQD1BWP12T register_file_inst1_pc_reg_26_ ( .D(register_file_inst1_n2195), 
        .CP(clock), .Q(RF_pc_out[26]) );
  DFQD1BWP12T register_file_inst1_pc_reg_27_ ( .D(register_file_inst1_n2196), 
        .CP(clock), .Q(RF_pc_out[27]) );
  DFQD1BWP12T register_file_inst1_pc_reg_28_ ( .D(register_file_inst1_n2197), 
        .CP(clock), .Q(RF_pc_out[28]) );
  DFQD1BWP12T register_file_inst1_pc_reg_29_ ( .D(register_file_inst1_n2198), 
        .CP(clock), .Q(RF_pc_out[29]) );
  DFQD1BWP12T register_file_inst1_pc_reg_30_ ( .D(register_file_inst1_n2199), 
        .CP(clock), .Q(RF_pc_out[30]) );
  DFQD1BWP12T register_file_inst1_pc_reg_31_ ( .D(register_file_inst1_n2200), 
        .CP(clock), .Q(RF_pc_out[31]) );
  DFQD1BWP12T register_file_inst1_sp_reg_0_ ( .D(register_file_inst1_spin[0]), 
        .CP(clock), .Q(RF_next_sp[0]) );
  DFQD1BWP12T register_file_inst1_sp_reg_1_ ( .D(register_file_inst1_spin[1]), 
        .CP(clock), .Q(RF_next_sp[1]) );
  DFQD1BWP12T register_file_inst1_sp_reg_2_ ( .D(register_file_inst1_spin[2]), 
        .CP(clock), .Q(RF_next_sp[2]) );
  DFQD1BWP12T register_file_inst1_sp_reg_3_ ( .D(register_file_inst1_spin[3]), 
        .CP(clock), .Q(RF_next_sp[3]) );
  DFQD1BWP12T register_file_inst1_sp_reg_4_ ( .D(register_file_inst1_spin[4]), 
        .CP(clock), .Q(RF_next_sp[4]) );
  DFQD1BWP12T register_file_inst1_sp_reg_5_ ( .D(register_file_inst1_spin[5]), 
        .CP(clock), .Q(RF_next_sp[5]) );
  DFQD1BWP12T register_file_inst1_sp_reg_6_ ( .D(register_file_inst1_spin[6]), 
        .CP(clock), .Q(RF_next_sp[6]) );
  DFQD1BWP12T register_file_inst1_sp_reg_7_ ( .D(register_file_inst1_spin[7]), 
        .CP(clock), .Q(RF_next_sp[7]) );
  DFQD1BWP12T register_file_inst1_sp_reg_8_ ( .D(register_file_inst1_spin[8]), 
        .CP(clock), .Q(RF_next_sp[8]) );
  DFQD1BWP12T register_file_inst1_sp_reg_9_ ( .D(register_file_inst1_spin[9]), 
        .CP(clock), .Q(RF_next_sp[9]) );
  DFQD1BWP12T register_file_inst1_sp_reg_10_ ( .D(register_file_inst1_spin[10]), .CP(clock), .Q(RF_next_sp[10]) );
  DFQD1BWP12T register_file_inst1_sp_reg_11_ ( .D(register_file_inst1_spin[11]), .CP(clock), .Q(RF_next_sp[11]) );
  DFQD1BWP12T register_file_inst1_sp_reg_12_ ( .D(register_file_inst1_spin[12]), .CP(clock), .Q(RF_next_sp[12]) );
  DFQD1BWP12T register_file_inst1_sp_reg_13_ ( .D(register_file_inst1_spin[13]), .CP(clock), .Q(RF_next_sp[13]) );
  DFQD1BWP12T register_file_inst1_sp_reg_14_ ( .D(register_file_inst1_spin[14]), .CP(clock), .Q(RF_next_sp[14]) );
  DFQD1BWP12T register_file_inst1_sp_reg_15_ ( .D(register_file_inst1_spin[15]), .CP(clock), .Q(RF_next_sp[15]) );
  DFQD1BWP12T register_file_inst1_sp_reg_16_ ( .D(register_file_inst1_spin[16]), .CP(clock), .Q(RF_next_sp[16]) );
  DFQD1BWP12T register_file_inst1_sp_reg_17_ ( .D(register_file_inst1_spin[17]), .CP(clock), .Q(RF_next_sp[17]) );
  DFQD1BWP12T register_file_inst1_sp_reg_18_ ( .D(register_file_inst1_spin[18]), .CP(clock), .Q(RF_next_sp[18]) );
  DFQD1BWP12T register_file_inst1_sp_reg_19_ ( .D(register_file_inst1_spin[19]), .CP(clock), .Q(RF_next_sp[19]) );
  DFQD1BWP12T register_file_inst1_sp_reg_20_ ( .D(register_file_inst1_spin[20]), .CP(clock), .Q(RF_next_sp[20]) );
  DFQD1BWP12T register_file_inst1_sp_reg_21_ ( .D(register_file_inst1_spin[21]), .CP(clock), .Q(RF_next_sp[21]) );
  DFQD1BWP12T register_file_inst1_sp_reg_22_ ( .D(register_file_inst1_spin[22]), .CP(clock), .Q(RF_next_sp[22]) );
  DFQD1BWP12T register_file_inst1_sp_reg_23_ ( .D(register_file_inst1_spin[23]), .CP(clock), .Q(RF_next_sp[23]) );
  DFQD1BWP12T register_file_inst1_sp_reg_24_ ( .D(register_file_inst1_spin[24]), .CP(clock), .Q(RF_next_sp[24]) );
  DFQD1BWP12T register_file_inst1_sp_reg_25_ ( .D(register_file_inst1_spin[25]), .CP(clock), .Q(RF_next_sp[25]) );
  DFQD1BWP12T register_file_inst1_sp_reg_26_ ( .D(register_file_inst1_spin[26]), .CP(clock), .Q(RF_next_sp[26]) );
  DFQD1BWP12T register_file_inst1_sp_reg_27_ ( .D(register_file_inst1_spin[27]), .CP(clock), .Q(RF_next_sp[27]) );
  DFQD1BWP12T register_file_inst1_sp_reg_28_ ( .D(register_file_inst1_spin[28]), .CP(clock), .Q(RF_next_sp[28]) );
  DFQD1BWP12T register_file_inst1_sp_reg_29_ ( .D(register_file_inst1_spin[29]), .CP(clock), .Q(RF_next_sp[29]) );
  DFQD1BWP12T register_file_inst1_sp_reg_30_ ( .D(register_file_inst1_spin[30]), .CP(clock), .Q(RF_next_sp[30]) );
  DFQD1BWP12T register_file_inst1_sp_reg_31_ ( .D(register_file_inst1_spin[31]), .CP(clock), .Q(RF_next_sp[31]) );
  DFQD1BWP12T register_file_inst1_lr_reg_0_ ( .D(register_file_inst1_n2201), 
        .CP(clock), .Q(register_file_inst1_lr_0_) );
  DFQD1BWP12T register_file_inst1_lr_reg_1_ ( .D(register_file_inst1_n2202), 
        .CP(clock), .Q(register_file_inst1_lr_1_) );
  DFQD1BWP12T register_file_inst1_lr_reg_2_ ( .D(register_file_inst1_n2203), 
        .CP(clock), .Q(register_file_inst1_lr_2_) );
  DFQD1BWP12T register_file_inst1_lr_reg_3_ ( .D(register_file_inst1_n2204), 
        .CP(clock), .Q(register_file_inst1_lr_3_) );
  DFQD1BWP12T register_file_inst1_lr_reg_4_ ( .D(register_file_inst1_n2205), 
        .CP(clock), .Q(register_file_inst1_lr_4_) );
  DFQD1BWP12T register_file_inst1_lr_reg_5_ ( .D(register_file_inst1_n2206), 
        .CP(clock), .Q(register_file_inst1_lr_5_) );
  DFQD1BWP12T register_file_inst1_lr_reg_7_ ( .D(register_file_inst1_n2208), 
        .CP(clock), .Q(register_file_inst1_lr_7_) );
  DFQD1BWP12T register_file_inst1_lr_reg_8_ ( .D(register_file_inst1_n2209), 
        .CP(clock), .Q(register_file_inst1_lr_8_) );
  DFQD1BWP12T register_file_inst1_lr_reg_9_ ( .D(register_file_inst1_n2210), 
        .CP(clock), .Q(register_file_inst1_lr_9_) );
  DFQD1BWP12T register_file_inst1_lr_reg_10_ ( .D(register_file_inst1_n2211), 
        .CP(clock), .Q(register_file_inst1_lr_10_) );
  DFQD1BWP12T register_file_inst1_lr_reg_11_ ( .D(register_file_inst1_n2212), 
        .CP(clock), .Q(register_file_inst1_lr_11_) );
  DFQD1BWP12T register_file_inst1_lr_reg_13_ ( .D(register_file_inst1_n2214), 
        .CP(clock), .Q(register_file_inst1_lr_13_) );
  DFQD1BWP12T register_file_inst1_lr_reg_14_ ( .D(register_file_inst1_n2215), 
        .CP(clock), .Q(register_file_inst1_lr_14_) );
  DFQD1BWP12T register_file_inst1_lr_reg_15_ ( .D(register_file_inst1_n2216), 
        .CP(clock), .Q(register_file_inst1_lr_15_) );
  DFQD1BWP12T register_file_inst1_lr_reg_16_ ( .D(register_file_inst1_n2217), 
        .CP(clock), .Q(register_file_inst1_lr_16_) );
  DFQD1BWP12T register_file_inst1_lr_reg_17_ ( .D(register_file_inst1_n2218), 
        .CP(clock), .Q(register_file_inst1_lr_17_) );
  DFQD1BWP12T register_file_inst1_lr_reg_18_ ( .D(register_file_inst1_n2219), 
        .CP(clock), .Q(register_file_inst1_lr_18_) );
  DFQD1BWP12T register_file_inst1_lr_reg_19_ ( .D(register_file_inst1_n2220), 
        .CP(clock), .Q(register_file_inst1_lr_19_) );
  DFQD1BWP12T register_file_inst1_lr_reg_20_ ( .D(register_file_inst1_n2221), 
        .CP(clock), .Q(register_file_inst1_lr_20_) );
  DFQD1BWP12T register_file_inst1_lr_reg_21_ ( .D(register_file_inst1_n2222), 
        .CP(clock), .Q(register_file_inst1_lr_21_) );
  DFQD1BWP12T register_file_inst1_lr_reg_22_ ( .D(register_file_inst1_n2223), 
        .CP(clock), .Q(register_file_inst1_lr_22_) );
  DFQD1BWP12T register_file_inst1_lr_reg_23_ ( .D(register_file_inst1_n2224), 
        .CP(clock), .Q(register_file_inst1_lr_23_) );
  DFQD1BWP12T register_file_inst1_lr_reg_24_ ( .D(register_file_inst1_n2225), 
        .CP(clock), .Q(register_file_inst1_lr_24_) );
  DFQD1BWP12T register_file_inst1_lr_reg_25_ ( .D(register_file_inst1_n2226), 
        .CP(clock), .Q(register_file_inst1_lr_25_) );
  DFQD1BWP12T register_file_inst1_lr_reg_26_ ( .D(register_file_inst1_n2227), 
        .CP(clock), .Q(register_file_inst1_lr_26_) );
  DFQD1BWP12T register_file_inst1_lr_reg_27_ ( .D(register_file_inst1_n2228), 
        .CP(clock), .Q(register_file_inst1_lr_27_) );
  DFQD1BWP12T register_file_inst1_lr_reg_28_ ( .D(register_file_inst1_n2229), 
        .CP(clock), .Q(register_file_inst1_lr_28_) );
  DFQD1BWP12T register_file_inst1_lr_reg_29_ ( .D(register_file_inst1_n2230), 
        .CP(clock), .Q(register_file_inst1_lr_29_) );
  DFQD1BWP12T register_file_inst1_lr_reg_30_ ( .D(register_file_inst1_n2231), 
        .CP(clock), .Q(register_file_inst1_lr_30_) );
  DFQD1BWP12T register_file_inst1_lr_reg_31_ ( .D(register_file_inst1_n2232), 
        .CP(clock), .Q(register_file_inst1_lr_31_) );
  DFQD1BWP12T register_file_inst1_r12_reg_0_ ( .D(register_file_inst1_n2233), 
        .CP(clock), .Q(register_file_inst1_r12_0_) );
  DFQD1BWP12T register_file_inst1_r12_reg_1_ ( .D(register_file_inst1_n2234), 
        .CP(clock), .Q(register_file_inst1_r12_1_) );
  DFQD1BWP12T register_file_inst1_r12_reg_3_ ( .D(register_file_inst1_n2236), 
        .CP(clock), .Q(register_file_inst1_r12_3_) );
  DFQD1BWP12T register_file_inst1_r12_reg_4_ ( .D(register_file_inst1_n2237), 
        .CP(clock), .Q(register_file_inst1_r12_4_) );
  DFQD1BWP12T register_file_inst1_r12_reg_5_ ( .D(register_file_inst1_n2238), 
        .CP(clock), .Q(register_file_inst1_r12_5_) );
  DFQD1BWP12T register_file_inst1_r12_reg_6_ ( .D(register_file_inst1_n2239), 
        .CP(clock), .Q(register_file_inst1_r12_6_) );
  DFQD1BWP12T register_file_inst1_r12_reg_7_ ( .D(register_file_inst1_n2240), 
        .CP(clock), .Q(register_file_inst1_r12_7_) );
  DFQD1BWP12T register_file_inst1_r12_reg_8_ ( .D(register_file_inst1_n2241), 
        .CP(clock), .Q(register_file_inst1_r12_8_) );
  DFQD1BWP12T register_file_inst1_r12_reg_9_ ( .D(register_file_inst1_n2242), 
        .CP(clock), .Q(register_file_inst1_r12_9_) );
  DFQD1BWP12T register_file_inst1_r12_reg_10_ ( .D(register_file_inst1_n2243), 
        .CP(clock), .Q(register_file_inst1_r12_10_) );
  DFQD1BWP12T register_file_inst1_r12_reg_11_ ( .D(register_file_inst1_n2244), 
        .CP(clock), .Q(register_file_inst1_r12_11_) );
  DFQD1BWP12T register_file_inst1_r12_reg_12_ ( .D(register_file_inst1_n2245), 
        .CP(clock), .Q(register_file_inst1_r12_12_) );
  DFQD1BWP12T register_file_inst1_r12_reg_13_ ( .D(register_file_inst1_n2246), 
        .CP(clock), .Q(register_file_inst1_r12_13_) );
  DFQD1BWP12T register_file_inst1_r12_reg_14_ ( .D(register_file_inst1_n2247), 
        .CP(clock), .Q(register_file_inst1_r12_14_) );
  DFQD1BWP12T register_file_inst1_r12_reg_15_ ( .D(register_file_inst1_n2248), 
        .CP(clock), .Q(register_file_inst1_r12_15_) );
  DFQD1BWP12T register_file_inst1_r12_reg_16_ ( .D(register_file_inst1_n2249), 
        .CP(clock), .Q(register_file_inst1_r12_16_) );
  DFQD1BWP12T register_file_inst1_r12_reg_17_ ( .D(register_file_inst1_n2250), 
        .CP(clock), .Q(register_file_inst1_r12_17_) );
  DFQD1BWP12T register_file_inst1_r12_reg_18_ ( .D(register_file_inst1_n2251), 
        .CP(clock), .Q(register_file_inst1_r12_18_) );
  DFQD1BWP12T register_file_inst1_r12_reg_19_ ( .D(register_file_inst1_n2252), 
        .CP(clock), .Q(register_file_inst1_r12_19_) );
  DFQD1BWP12T register_file_inst1_r12_reg_20_ ( .D(register_file_inst1_n2253), 
        .CP(clock), .Q(register_file_inst1_r12_20_) );
  DFQD1BWP12T register_file_inst1_r12_reg_21_ ( .D(register_file_inst1_n2254), 
        .CP(clock), .Q(register_file_inst1_r12_21_) );
  DFQD1BWP12T register_file_inst1_r12_reg_22_ ( .D(register_file_inst1_n2255), 
        .CP(clock), .Q(register_file_inst1_r12_22_) );
  DFQD1BWP12T register_file_inst1_r12_reg_23_ ( .D(register_file_inst1_n2256), 
        .CP(clock), .Q(register_file_inst1_r12_23_) );
  DFQD1BWP12T register_file_inst1_r12_reg_24_ ( .D(register_file_inst1_n2257), 
        .CP(clock), .Q(register_file_inst1_r12_24_) );
  DFQD1BWP12T register_file_inst1_r12_reg_25_ ( .D(register_file_inst1_n2258), 
        .CP(clock), .Q(register_file_inst1_r12_25_) );
  DFQD1BWP12T register_file_inst1_r12_reg_26_ ( .D(register_file_inst1_n2259), 
        .CP(clock), .Q(register_file_inst1_r12_26_) );
  DFQD1BWP12T register_file_inst1_r12_reg_27_ ( .D(register_file_inst1_n2260), 
        .CP(clock), .Q(register_file_inst1_r12_27_) );
  DFQD1BWP12T register_file_inst1_r12_reg_28_ ( .D(register_file_inst1_n2261), 
        .CP(clock), .Q(register_file_inst1_r12_28_) );
  DFQD1BWP12T register_file_inst1_r12_reg_29_ ( .D(register_file_inst1_n2262), 
        .CP(clock), .Q(register_file_inst1_r12_29_) );
  DFQD1BWP12T register_file_inst1_r12_reg_30_ ( .D(register_file_inst1_n2263), 
        .CP(clock), .Q(register_file_inst1_r12_30_) );
  DFQD1BWP12T register_file_inst1_r12_reg_31_ ( .D(register_file_inst1_n2264), 
        .CP(clock), .Q(register_file_inst1_r12_31_) );
  DFQD1BWP12T register_file_inst1_r11_reg_0_ ( .D(register_file_inst1_n2265), 
        .CP(clock), .Q(register_file_inst1_r11_0_) );
  DFQD1BWP12T register_file_inst1_r11_reg_1_ ( .D(register_file_inst1_n2266), 
        .CP(clock), .Q(register_file_inst1_r11_1_) );
  DFQD1BWP12T register_file_inst1_r11_reg_2_ ( .D(register_file_inst1_n2267), 
        .CP(clock), .Q(register_file_inst1_r11_2_) );
  DFQD1BWP12T register_file_inst1_r11_reg_3_ ( .D(register_file_inst1_n2268), 
        .CP(clock), .Q(register_file_inst1_r11_3_) );
  DFQD1BWP12T register_file_inst1_r11_reg_4_ ( .D(register_file_inst1_n2269), 
        .CP(clock), .Q(register_file_inst1_r11_4_) );
  DFQD1BWP12T register_file_inst1_r11_reg_5_ ( .D(register_file_inst1_n2270), 
        .CP(clock), .Q(register_file_inst1_r11_5_) );
  DFQD1BWP12T register_file_inst1_r11_reg_6_ ( .D(register_file_inst1_n2271), 
        .CP(clock), .Q(register_file_inst1_r11_6_) );
  DFQD1BWP12T register_file_inst1_r11_reg_8_ ( .D(register_file_inst1_n2273), 
        .CP(clock), .Q(register_file_inst1_r11_8_) );
  DFQD1BWP12T register_file_inst1_r11_reg_10_ ( .D(register_file_inst1_n2275), 
        .CP(clock), .Q(register_file_inst1_r11_10_) );
  DFQD1BWP12T register_file_inst1_r11_reg_11_ ( .D(register_file_inst1_n2276), 
        .CP(clock), .Q(register_file_inst1_r11_11_) );
  DFQD1BWP12T register_file_inst1_r11_reg_12_ ( .D(register_file_inst1_n2277), 
        .CP(clock), .Q(register_file_inst1_r11_12_) );
  DFQD1BWP12T register_file_inst1_r11_reg_13_ ( .D(register_file_inst1_n2278), 
        .CP(clock), .Q(register_file_inst1_r11_13_) );
  DFQD1BWP12T register_file_inst1_r11_reg_14_ ( .D(register_file_inst1_n2279), 
        .CP(clock), .Q(register_file_inst1_r11_14_) );
  DFQD1BWP12T register_file_inst1_r11_reg_15_ ( .D(register_file_inst1_n2280), 
        .CP(clock), .Q(register_file_inst1_r11_15_) );
  DFQD1BWP12T register_file_inst1_r11_reg_16_ ( .D(register_file_inst1_n2281), 
        .CP(clock), .Q(register_file_inst1_r11_16_) );
  DFQD1BWP12T register_file_inst1_r11_reg_17_ ( .D(register_file_inst1_n2282), 
        .CP(clock), .Q(register_file_inst1_r11_17_) );
  DFQD1BWP12T register_file_inst1_r11_reg_18_ ( .D(register_file_inst1_n2283), 
        .CP(clock), .Q(register_file_inst1_r11_18_) );
  DFQD1BWP12T register_file_inst1_r11_reg_19_ ( .D(register_file_inst1_n2284), 
        .CP(clock), .Q(register_file_inst1_r11_19_) );
  DFQD1BWP12T register_file_inst1_r11_reg_20_ ( .D(register_file_inst1_n2285), 
        .CP(clock), .Q(register_file_inst1_r11_20_) );
  DFQD1BWP12T register_file_inst1_r11_reg_21_ ( .D(register_file_inst1_n2286), 
        .CP(clock), .Q(register_file_inst1_r11_21_) );
  DFQD1BWP12T register_file_inst1_r11_reg_22_ ( .D(register_file_inst1_n2287), 
        .CP(clock), .Q(register_file_inst1_r11_22_) );
  DFQD1BWP12T register_file_inst1_r11_reg_23_ ( .D(register_file_inst1_n2288), 
        .CP(clock), .Q(register_file_inst1_r11_23_) );
  DFQD1BWP12T register_file_inst1_r11_reg_24_ ( .D(register_file_inst1_n2289), 
        .CP(clock), .Q(register_file_inst1_r11_24_) );
  DFQD1BWP12T register_file_inst1_r11_reg_25_ ( .D(register_file_inst1_n2290), 
        .CP(clock), .Q(register_file_inst1_r11_25_) );
  DFQD1BWP12T register_file_inst1_r11_reg_26_ ( .D(register_file_inst1_n2291), 
        .CP(clock), .Q(register_file_inst1_r11_26_) );
  DFQD1BWP12T register_file_inst1_r11_reg_27_ ( .D(register_file_inst1_n2292), 
        .CP(clock), .Q(register_file_inst1_r11_27_) );
  DFQD1BWP12T register_file_inst1_r11_reg_28_ ( .D(register_file_inst1_n2293), 
        .CP(clock), .Q(register_file_inst1_r11_28_) );
  DFQD1BWP12T register_file_inst1_r11_reg_29_ ( .D(register_file_inst1_n2294), 
        .CP(clock), .Q(register_file_inst1_r11_29_) );
  DFQD1BWP12T register_file_inst1_r11_reg_30_ ( .D(register_file_inst1_n2295), 
        .CP(clock), .Q(register_file_inst1_r11_30_) );
  DFQD1BWP12T register_file_inst1_r11_reg_31_ ( .D(register_file_inst1_n2296), 
        .CP(clock), .Q(register_file_inst1_r11_31_) );
  DFQD1BWP12T register_file_inst1_r10_reg_0_ ( .D(register_file_inst1_n2297), 
        .CP(clock), .Q(register_file_inst1_r10_0_) );
  DFQD1BWP12T register_file_inst1_r10_reg_1_ ( .D(register_file_inst1_n2298), 
        .CP(clock), .Q(register_file_inst1_r10_1_) );
  DFQD1BWP12T register_file_inst1_r10_reg_2_ ( .D(register_file_inst1_n2299), 
        .CP(clock), .Q(register_file_inst1_r10_2_) );
  DFQD1BWP12T register_file_inst1_r10_reg_3_ ( .D(register_file_inst1_n2300), 
        .CP(clock), .Q(register_file_inst1_r10_3_) );
  DFQD1BWP12T register_file_inst1_r10_reg_4_ ( .D(register_file_inst1_n2301), 
        .CP(clock), .Q(register_file_inst1_r10_4_) );
  DFQD1BWP12T register_file_inst1_r10_reg_5_ ( .D(register_file_inst1_n2302), 
        .CP(clock), .Q(register_file_inst1_r10_5_) );
  DFQD1BWP12T register_file_inst1_r10_reg_6_ ( .D(register_file_inst1_n2303), 
        .CP(clock), .Q(register_file_inst1_r10_6_) );
  DFQD1BWP12T register_file_inst1_r10_reg_8_ ( .D(register_file_inst1_n2305), 
        .CP(clock), .Q(register_file_inst1_r10_8_) );
  DFQD1BWP12T register_file_inst1_r10_reg_9_ ( .D(register_file_inst1_n2306), 
        .CP(clock), .Q(register_file_inst1_r10_9_) );
  DFQD1BWP12T register_file_inst1_r10_reg_10_ ( .D(register_file_inst1_n2307), 
        .CP(clock), .Q(register_file_inst1_r10_10_) );
  DFQD1BWP12T register_file_inst1_r10_reg_11_ ( .D(register_file_inst1_n2308), 
        .CP(clock), .Q(register_file_inst1_r10_11_) );
  DFQD1BWP12T register_file_inst1_r10_reg_12_ ( .D(register_file_inst1_n2309), 
        .CP(clock), .Q(register_file_inst1_r10_12_) );
  DFQD1BWP12T register_file_inst1_r10_reg_13_ ( .D(register_file_inst1_n2310), 
        .CP(clock), .Q(register_file_inst1_r10_13_) );
  DFQD1BWP12T register_file_inst1_r10_reg_14_ ( .D(register_file_inst1_n2311), 
        .CP(clock), .Q(register_file_inst1_r10_14_) );
  DFQD1BWP12T register_file_inst1_r10_reg_15_ ( .D(register_file_inst1_n2312), 
        .CP(clock), .Q(register_file_inst1_r10_15_) );
  DFQD1BWP12T register_file_inst1_r10_reg_16_ ( .D(register_file_inst1_n2313), 
        .CP(clock), .Q(register_file_inst1_r10_16_) );
  DFQD1BWP12T register_file_inst1_r10_reg_17_ ( .D(register_file_inst1_n2314), 
        .CP(clock), .Q(register_file_inst1_r10_17_) );
  DFQD1BWP12T register_file_inst1_r10_reg_18_ ( .D(register_file_inst1_n2315), 
        .CP(clock), .Q(register_file_inst1_r10_18_) );
  DFQD1BWP12T register_file_inst1_r10_reg_19_ ( .D(register_file_inst1_n2316), 
        .CP(clock), .Q(register_file_inst1_r10_19_) );
  DFQD1BWP12T register_file_inst1_r10_reg_20_ ( .D(register_file_inst1_n2317), 
        .CP(clock), .Q(register_file_inst1_r10_20_) );
  DFQD1BWP12T register_file_inst1_r10_reg_21_ ( .D(register_file_inst1_n2318), 
        .CP(clock), .Q(register_file_inst1_r10_21_) );
  DFQD1BWP12T register_file_inst1_r10_reg_22_ ( .D(register_file_inst1_n2319), 
        .CP(clock), .Q(register_file_inst1_r10_22_) );
  DFQD1BWP12T register_file_inst1_r10_reg_23_ ( .D(register_file_inst1_n2320), 
        .CP(clock), .Q(register_file_inst1_r10_23_) );
  DFQD1BWP12T register_file_inst1_r10_reg_24_ ( .D(register_file_inst1_n2321), 
        .CP(clock), .Q(register_file_inst1_r10_24_) );
  DFQD1BWP12T register_file_inst1_r10_reg_25_ ( .D(register_file_inst1_n2322), 
        .CP(clock), .Q(register_file_inst1_r10_25_) );
  DFQD1BWP12T register_file_inst1_r10_reg_26_ ( .D(register_file_inst1_n2323), 
        .CP(clock), .Q(register_file_inst1_r10_26_) );
  DFQD1BWP12T register_file_inst1_r10_reg_27_ ( .D(register_file_inst1_n2324), 
        .CP(clock), .Q(register_file_inst1_r10_27_) );
  DFQD1BWP12T register_file_inst1_r10_reg_28_ ( .D(register_file_inst1_n2325), 
        .CP(clock), .Q(register_file_inst1_r10_28_) );
  DFQD1BWP12T register_file_inst1_r10_reg_29_ ( .D(register_file_inst1_n2326), 
        .CP(clock), .Q(register_file_inst1_r10_29_) );
  DFQD1BWP12T register_file_inst1_r10_reg_30_ ( .D(register_file_inst1_n2327), 
        .CP(clock), .Q(register_file_inst1_r10_30_) );
  DFQD1BWP12T register_file_inst1_r10_reg_31_ ( .D(register_file_inst1_n2328), 
        .CP(clock), .Q(register_file_inst1_r10_31_) );
  DFQD1BWP12T register_file_inst1_r9_reg_0_ ( .D(register_file_inst1_n2329), 
        .CP(clock), .Q(register_file_inst1_r9_0_) );
  DFQD1BWP12T register_file_inst1_r9_reg_1_ ( .D(register_file_inst1_n2330), 
        .CP(clock), .Q(register_file_inst1_r9_1_) );
  DFQD1BWP12T register_file_inst1_r9_reg_2_ ( .D(register_file_inst1_n2331), 
        .CP(clock), .Q(register_file_inst1_r9_2_) );
  DFQD1BWP12T register_file_inst1_r9_reg_3_ ( .D(register_file_inst1_n2332), 
        .CP(clock), .Q(register_file_inst1_r9_3_) );
  DFQD1BWP12T register_file_inst1_r9_reg_4_ ( .D(register_file_inst1_n2333), 
        .CP(clock), .Q(register_file_inst1_r9_4_) );
  DFQD1BWP12T register_file_inst1_r9_reg_5_ ( .D(register_file_inst1_n2334), 
        .CP(clock), .Q(register_file_inst1_r9_5_) );
  DFQD1BWP12T register_file_inst1_r9_reg_6_ ( .D(register_file_inst1_n2335), 
        .CP(clock), .Q(register_file_inst1_r9_6_) );
  DFQD1BWP12T register_file_inst1_r9_reg_7_ ( .D(register_file_inst1_n2336), 
        .CP(clock), .Q(register_file_inst1_r9_7_) );
  DFQD1BWP12T register_file_inst1_r9_reg_8_ ( .D(register_file_inst1_n2337), 
        .CP(clock), .Q(register_file_inst1_r9_8_) );
  DFQD1BWP12T register_file_inst1_r9_reg_9_ ( .D(register_file_inst1_n2338), 
        .CP(clock), .Q(register_file_inst1_r9_9_) );
  DFQD1BWP12T register_file_inst1_r9_reg_10_ ( .D(register_file_inst1_n2339), 
        .CP(clock), .Q(register_file_inst1_r9_10_) );
  DFQD1BWP12T register_file_inst1_r9_reg_11_ ( .D(register_file_inst1_n2340), 
        .CP(clock), .Q(register_file_inst1_r9_11_) );
  DFQD1BWP12T register_file_inst1_r9_reg_12_ ( .D(register_file_inst1_n2341), 
        .CP(clock), .Q(register_file_inst1_r9_12_) );
  DFQD1BWP12T register_file_inst1_r9_reg_13_ ( .D(register_file_inst1_n2342), 
        .CP(clock), .Q(register_file_inst1_r9_13_) );
  DFQD1BWP12T register_file_inst1_r9_reg_14_ ( .D(register_file_inst1_n2343), 
        .CP(clock), .Q(register_file_inst1_r9_14_) );
  DFQD1BWP12T register_file_inst1_r9_reg_15_ ( .D(register_file_inst1_n2344), 
        .CP(clock), .Q(register_file_inst1_r9_15_) );
  DFQD1BWP12T register_file_inst1_r9_reg_16_ ( .D(register_file_inst1_n2345), 
        .CP(clock), .Q(register_file_inst1_r9_16_) );
  DFQD1BWP12T register_file_inst1_r9_reg_17_ ( .D(register_file_inst1_n2346), 
        .CP(clock), .Q(register_file_inst1_r9_17_) );
  DFQD1BWP12T register_file_inst1_r9_reg_18_ ( .D(register_file_inst1_n2347), 
        .CP(clock), .Q(register_file_inst1_r9_18_) );
  DFQD1BWP12T register_file_inst1_r9_reg_19_ ( .D(register_file_inst1_n2348), 
        .CP(clock), .Q(register_file_inst1_r9_19_) );
  DFQD1BWP12T register_file_inst1_r9_reg_20_ ( .D(register_file_inst1_n2349), 
        .CP(clock), .Q(register_file_inst1_r9_20_) );
  DFQD1BWP12T register_file_inst1_r9_reg_21_ ( .D(register_file_inst1_n2350), 
        .CP(clock), .Q(register_file_inst1_r9_21_) );
  DFQD1BWP12T register_file_inst1_r9_reg_22_ ( .D(register_file_inst1_n2351), 
        .CP(clock), .Q(register_file_inst1_r9_22_) );
  DFQD1BWP12T register_file_inst1_r9_reg_23_ ( .D(register_file_inst1_n2352), 
        .CP(clock), .Q(register_file_inst1_r9_23_) );
  DFQD1BWP12T register_file_inst1_r9_reg_24_ ( .D(register_file_inst1_n2353), 
        .CP(clock), .Q(register_file_inst1_r9_24_) );
  DFQD1BWP12T register_file_inst1_r9_reg_25_ ( .D(register_file_inst1_n2354), 
        .CP(clock), .Q(register_file_inst1_r9_25_) );
  DFQD1BWP12T register_file_inst1_r9_reg_26_ ( .D(register_file_inst1_n2355), 
        .CP(clock), .Q(register_file_inst1_r9_26_) );
  DFQD1BWP12T register_file_inst1_r9_reg_27_ ( .D(register_file_inst1_n2356), 
        .CP(clock), .Q(register_file_inst1_r9_27_) );
  DFQD1BWP12T register_file_inst1_r9_reg_28_ ( .D(register_file_inst1_n2357), 
        .CP(clock), .Q(register_file_inst1_r9_28_) );
  DFQD1BWP12T register_file_inst1_r9_reg_29_ ( .D(register_file_inst1_n2358), 
        .CP(clock), .Q(register_file_inst1_r9_29_) );
  DFQD1BWP12T register_file_inst1_r9_reg_30_ ( .D(register_file_inst1_n2359), 
        .CP(clock), .Q(register_file_inst1_r9_30_) );
  DFQD1BWP12T register_file_inst1_r9_reg_31_ ( .D(register_file_inst1_n2360), 
        .CP(clock), .Q(register_file_inst1_r9_31_) );
  DFQD1BWP12T register_file_inst1_r8_reg_0_ ( .D(register_file_inst1_n2361), 
        .CP(clock), .Q(register_file_inst1_r8_0_) );
  DFQD1BWP12T register_file_inst1_r8_reg_1_ ( .D(register_file_inst1_n2362), 
        .CP(clock), .Q(register_file_inst1_r8_1_) );
  DFQD1BWP12T register_file_inst1_r8_reg_3_ ( .D(register_file_inst1_n2364), 
        .CP(clock), .Q(register_file_inst1_r8_3_) );
  DFQD1BWP12T register_file_inst1_r8_reg_4_ ( .D(register_file_inst1_n2365), 
        .CP(clock), .Q(register_file_inst1_r8_4_) );
  DFQD1BWP12T register_file_inst1_r8_reg_5_ ( .D(register_file_inst1_n2366), 
        .CP(clock), .Q(register_file_inst1_r8_5_) );
  DFQD1BWP12T register_file_inst1_r8_reg_6_ ( .D(register_file_inst1_n2367), 
        .CP(clock), .Q(register_file_inst1_r8_6_) );
  DFQD1BWP12T register_file_inst1_r8_reg_7_ ( .D(register_file_inst1_n2368), 
        .CP(clock), .Q(register_file_inst1_r8_7_) );
  DFQD1BWP12T register_file_inst1_r8_reg_9_ ( .D(register_file_inst1_n2370), 
        .CP(clock), .Q(register_file_inst1_r8_9_) );
  DFQD1BWP12T register_file_inst1_r8_reg_10_ ( .D(register_file_inst1_n2371), 
        .CP(clock), .Q(register_file_inst1_r8_10_) );
  DFQD1BWP12T register_file_inst1_r8_reg_12_ ( .D(register_file_inst1_n2373), 
        .CP(clock), .Q(register_file_inst1_r8_12_) );
  DFQD1BWP12T register_file_inst1_r8_reg_13_ ( .D(register_file_inst1_n2374), 
        .CP(clock), .Q(register_file_inst1_r8_13_) );
  DFQD1BWP12T register_file_inst1_r8_reg_14_ ( .D(register_file_inst1_n2375), 
        .CP(clock), .Q(register_file_inst1_r8_14_) );
  DFQD1BWP12T register_file_inst1_r8_reg_16_ ( .D(register_file_inst1_n2377), 
        .CP(clock), .Q(register_file_inst1_r8_16_) );
  DFQD1BWP12T register_file_inst1_r8_reg_17_ ( .D(register_file_inst1_n2378), 
        .CP(clock), .Q(register_file_inst1_r8_17_) );
  DFQD1BWP12T register_file_inst1_r8_reg_18_ ( .D(register_file_inst1_n2379), 
        .CP(clock), .Q(register_file_inst1_r8_18_) );
  DFQD1BWP12T register_file_inst1_r8_reg_19_ ( .D(register_file_inst1_n2380), 
        .CP(clock), .Q(register_file_inst1_r8_19_) );
  DFQD1BWP12T register_file_inst1_r8_reg_20_ ( .D(register_file_inst1_n2381), 
        .CP(clock), .Q(register_file_inst1_r8_20_) );
  DFQD1BWP12T register_file_inst1_r8_reg_21_ ( .D(register_file_inst1_n2382), 
        .CP(clock), .Q(register_file_inst1_r8_21_) );
  DFQD1BWP12T register_file_inst1_r8_reg_22_ ( .D(register_file_inst1_n2383), 
        .CP(clock), .Q(register_file_inst1_r8_22_) );
  DFQD1BWP12T register_file_inst1_r8_reg_23_ ( .D(register_file_inst1_n2384), 
        .CP(clock), .Q(register_file_inst1_r8_23_) );
  DFQD1BWP12T register_file_inst1_r8_reg_24_ ( .D(register_file_inst1_n2385), 
        .CP(clock), .Q(register_file_inst1_r8_24_) );
  DFQD1BWP12T register_file_inst1_r8_reg_25_ ( .D(register_file_inst1_n2386), 
        .CP(clock), .Q(register_file_inst1_r8_25_) );
  DFQD1BWP12T register_file_inst1_r8_reg_26_ ( .D(register_file_inst1_n2387), 
        .CP(clock), .Q(register_file_inst1_r8_26_) );
  DFQD1BWP12T register_file_inst1_r8_reg_27_ ( .D(register_file_inst1_n2388), 
        .CP(clock), .Q(register_file_inst1_r8_27_) );
  DFQD1BWP12T register_file_inst1_r8_reg_28_ ( .D(register_file_inst1_n2389), 
        .CP(clock), .Q(register_file_inst1_r8_28_) );
  DFQD1BWP12T register_file_inst1_r8_reg_29_ ( .D(register_file_inst1_n2390), 
        .CP(clock), .Q(register_file_inst1_r8_29_) );
  DFQD1BWP12T register_file_inst1_r8_reg_30_ ( .D(register_file_inst1_n2391), 
        .CP(clock), .Q(register_file_inst1_r8_30_) );
  DFQD1BWP12T register_file_inst1_r8_reg_31_ ( .D(register_file_inst1_n2392), 
        .CP(clock), .Q(register_file_inst1_r8_31_) );
  DFQD1BWP12T register_file_inst1_r7_reg_0_ ( .D(register_file_inst1_n2393), 
        .CP(clock), .Q(register_file_inst1_r7_0_) );
  DFQD1BWP12T register_file_inst1_r7_reg_1_ ( .D(register_file_inst1_n2394), 
        .CP(clock), .Q(register_file_inst1_r7_1_) );
  DFQD1BWP12T register_file_inst1_r7_reg_2_ ( .D(register_file_inst1_n2395), 
        .CP(clock), .Q(register_file_inst1_r7_2_) );
  DFQD1BWP12T register_file_inst1_r7_reg_4_ ( .D(register_file_inst1_n2397), 
        .CP(clock), .Q(register_file_inst1_r7_4_) );
  DFQD1BWP12T register_file_inst1_r7_reg_5_ ( .D(register_file_inst1_n2398), 
        .CP(clock), .Q(register_file_inst1_r7_5_) );
  DFQD1BWP12T register_file_inst1_r7_reg_6_ ( .D(register_file_inst1_n2399), 
        .CP(clock), .Q(register_file_inst1_r7_6_) );
  DFQD1BWP12T register_file_inst1_r7_reg_7_ ( .D(register_file_inst1_n2400), 
        .CP(clock), .Q(register_file_inst1_r7_7_) );
  DFQD1BWP12T register_file_inst1_r7_reg_8_ ( .D(register_file_inst1_n2401), 
        .CP(clock), .Q(register_file_inst1_r7_8_) );
  DFQD1BWP12T register_file_inst1_r7_reg_10_ ( .D(register_file_inst1_n2403), 
        .CP(clock), .Q(register_file_inst1_r7_10_) );
  DFQD1BWP12T register_file_inst1_r7_reg_11_ ( .D(register_file_inst1_n2404), 
        .CP(clock), .Q(register_file_inst1_r7_11_) );
  DFQD1BWP12T register_file_inst1_r7_reg_12_ ( .D(register_file_inst1_n2405), 
        .CP(clock), .Q(register_file_inst1_r7_12_) );
  DFQD1BWP12T register_file_inst1_r7_reg_13_ ( .D(register_file_inst1_n2406), 
        .CP(clock), .Q(register_file_inst1_r7_13_) );
  DFQD1BWP12T register_file_inst1_r7_reg_14_ ( .D(register_file_inst1_n2407), 
        .CP(clock), .Q(register_file_inst1_r7_14_) );
  DFQD1BWP12T register_file_inst1_r7_reg_15_ ( .D(register_file_inst1_n2408), 
        .CP(clock), .Q(register_file_inst1_r7_15_) );
  DFQD1BWP12T register_file_inst1_r7_reg_16_ ( .D(register_file_inst1_n2409), 
        .CP(clock), .Q(register_file_inst1_r7_16_) );
  DFQD1BWP12T register_file_inst1_r7_reg_17_ ( .D(register_file_inst1_n2410), 
        .CP(clock), .Q(register_file_inst1_r7_17_) );
  DFQD1BWP12T register_file_inst1_r7_reg_18_ ( .D(register_file_inst1_n2411), 
        .CP(clock), .Q(register_file_inst1_r7_18_) );
  DFQD1BWP12T register_file_inst1_r7_reg_19_ ( .D(register_file_inst1_n2412), 
        .CP(clock), .Q(register_file_inst1_r7_19_) );
  DFQD1BWP12T register_file_inst1_r7_reg_20_ ( .D(register_file_inst1_n2413), 
        .CP(clock), .Q(register_file_inst1_r7_20_) );
  DFQD1BWP12T register_file_inst1_r7_reg_21_ ( .D(register_file_inst1_n2414), 
        .CP(clock), .Q(register_file_inst1_r7_21_) );
  DFQD1BWP12T register_file_inst1_r7_reg_22_ ( .D(register_file_inst1_n2415), 
        .CP(clock), .Q(register_file_inst1_r7_22_) );
  DFQD1BWP12T register_file_inst1_r7_reg_23_ ( .D(register_file_inst1_n2416), 
        .CP(clock), .Q(register_file_inst1_r7_23_) );
  DFQD1BWP12T register_file_inst1_r7_reg_24_ ( .D(register_file_inst1_n2417), 
        .CP(clock), .Q(register_file_inst1_r7_24_) );
  DFQD1BWP12T register_file_inst1_r7_reg_25_ ( .D(register_file_inst1_n2418), 
        .CP(clock), .Q(register_file_inst1_r7_25_) );
  DFQD1BWP12T register_file_inst1_r7_reg_26_ ( .D(register_file_inst1_n2419), 
        .CP(clock), .Q(register_file_inst1_r7_26_) );
  DFQD1BWP12T register_file_inst1_r7_reg_27_ ( .D(register_file_inst1_n2420), 
        .CP(clock), .Q(register_file_inst1_r7_27_) );
  DFQD1BWP12T register_file_inst1_r7_reg_28_ ( .D(register_file_inst1_n2421), 
        .CP(clock), .Q(register_file_inst1_r7_28_) );
  DFQD1BWP12T register_file_inst1_r7_reg_29_ ( .D(register_file_inst1_n2422), 
        .CP(clock), .Q(register_file_inst1_r7_29_) );
  DFQD1BWP12T register_file_inst1_r7_reg_30_ ( .D(register_file_inst1_n2423), 
        .CP(clock), .Q(register_file_inst1_r7_30_) );
  DFQD1BWP12T register_file_inst1_r7_reg_31_ ( .D(register_file_inst1_n2424), 
        .CP(clock), .Q(register_file_inst1_r7_31_) );
  DFQD1BWP12T register_file_inst1_r6_reg_0_ ( .D(register_file_inst1_n2425), 
        .CP(clock), .Q(register_file_inst1_r6_0_) );
  DFQD1BWP12T register_file_inst1_r6_reg_1_ ( .D(register_file_inst1_n2426), 
        .CP(clock), .Q(register_file_inst1_r6_1_) );
  DFQD1BWP12T register_file_inst1_r6_reg_2_ ( .D(register_file_inst1_n2427), 
        .CP(clock), .Q(register_file_inst1_r6_2_) );
  DFQD1BWP12T register_file_inst1_r6_reg_3_ ( .D(register_file_inst1_n2428), 
        .CP(clock), .Q(register_file_inst1_r6_3_) );
  DFQD1BWP12T register_file_inst1_r6_reg_4_ ( .D(register_file_inst1_n2429), 
        .CP(clock), .Q(register_file_inst1_r6_4_) );
  DFQD1BWP12T register_file_inst1_r6_reg_5_ ( .D(register_file_inst1_n2430), 
        .CP(clock), .Q(register_file_inst1_r6_5_) );
  DFQD1BWP12T register_file_inst1_r6_reg_6_ ( .D(register_file_inst1_n2431), 
        .CP(clock), .Q(register_file_inst1_r6_6_) );
  DFQD1BWP12T register_file_inst1_r6_reg_7_ ( .D(register_file_inst1_n2432), 
        .CP(clock), .Q(register_file_inst1_r6_7_) );
  DFQD1BWP12T register_file_inst1_r6_reg_8_ ( .D(register_file_inst1_n2433), 
        .CP(clock), .Q(register_file_inst1_r6_8_) );
  DFQD1BWP12T register_file_inst1_r6_reg_10_ ( .D(register_file_inst1_n2435), 
        .CP(clock), .Q(register_file_inst1_r6_10_) );
  DFQD1BWP12T register_file_inst1_r6_reg_11_ ( .D(register_file_inst1_n2436), 
        .CP(clock), .Q(register_file_inst1_r6_11_) );
  DFQD1BWP12T register_file_inst1_r6_reg_12_ ( .D(register_file_inst1_n2437), 
        .CP(clock), .Q(register_file_inst1_r6_12_) );
  DFQD1BWP12T register_file_inst1_r6_reg_13_ ( .D(register_file_inst1_n2438), 
        .CP(clock), .Q(register_file_inst1_r6_13_) );
  DFQD1BWP12T register_file_inst1_r6_reg_14_ ( .D(register_file_inst1_n2439), 
        .CP(clock), .Q(register_file_inst1_r6_14_) );
  DFQD1BWP12T register_file_inst1_r6_reg_15_ ( .D(register_file_inst1_n2440), 
        .CP(clock), .Q(register_file_inst1_r6_15_) );
  DFQD1BWP12T register_file_inst1_r6_reg_16_ ( .D(register_file_inst1_n2441), 
        .CP(clock), .Q(register_file_inst1_r6_16_) );
  DFQD1BWP12T register_file_inst1_r6_reg_17_ ( .D(register_file_inst1_n2442), 
        .CP(clock), .Q(register_file_inst1_r6_17_) );
  DFQD1BWP12T register_file_inst1_r6_reg_18_ ( .D(register_file_inst1_n2443), 
        .CP(clock), .Q(register_file_inst1_r6_18_) );
  DFQD1BWP12T register_file_inst1_r6_reg_19_ ( .D(register_file_inst1_n2444), 
        .CP(clock), .Q(register_file_inst1_r6_19_) );
  DFQD1BWP12T register_file_inst1_r6_reg_20_ ( .D(register_file_inst1_n2445), 
        .CP(clock), .Q(register_file_inst1_r6_20_) );
  DFQD1BWP12T register_file_inst1_r6_reg_21_ ( .D(register_file_inst1_n2446), 
        .CP(clock), .Q(register_file_inst1_r6_21_) );
  DFQD1BWP12T register_file_inst1_r6_reg_22_ ( .D(register_file_inst1_n2447), 
        .CP(clock), .Q(register_file_inst1_r6_22_) );
  DFQD1BWP12T register_file_inst1_r6_reg_23_ ( .D(register_file_inst1_n2448), 
        .CP(clock), .Q(register_file_inst1_r6_23_) );
  DFQD1BWP12T register_file_inst1_r6_reg_24_ ( .D(register_file_inst1_n2449), 
        .CP(clock), .Q(register_file_inst1_r6_24_) );
  DFQD1BWP12T register_file_inst1_r6_reg_25_ ( .D(register_file_inst1_n2450), 
        .CP(clock), .Q(register_file_inst1_r6_25_) );
  DFQD1BWP12T register_file_inst1_r6_reg_26_ ( .D(register_file_inst1_n2451), 
        .CP(clock), .Q(register_file_inst1_r6_26_) );
  DFQD1BWP12T register_file_inst1_r6_reg_27_ ( .D(register_file_inst1_n2452), 
        .CP(clock), .Q(register_file_inst1_r6_27_) );
  DFQD1BWP12T register_file_inst1_r6_reg_28_ ( .D(register_file_inst1_n2453), 
        .CP(clock), .Q(register_file_inst1_r6_28_) );
  DFQD1BWP12T register_file_inst1_r6_reg_29_ ( .D(register_file_inst1_n2454), 
        .CP(clock), .Q(register_file_inst1_r6_29_) );
  DFQD1BWP12T register_file_inst1_r6_reg_30_ ( .D(register_file_inst1_n2455), 
        .CP(clock), .Q(register_file_inst1_r6_30_) );
  DFQD1BWP12T register_file_inst1_r6_reg_31_ ( .D(register_file_inst1_n2456), 
        .CP(clock), .Q(register_file_inst1_r6_31_) );
  DFQD1BWP12T register_file_inst1_r5_reg_0_ ( .D(register_file_inst1_n2457), 
        .CP(clock), .Q(register_file_inst1_r5_0_) );
  DFQD1BWP12T register_file_inst1_r5_reg_1_ ( .D(register_file_inst1_n2458), 
        .CP(clock), .Q(register_file_inst1_r5_1_) );
  DFQD1BWP12T register_file_inst1_r5_reg_2_ ( .D(register_file_inst1_n2459), 
        .CP(clock), .Q(register_file_inst1_r5_2_) );
  DFQD1BWP12T register_file_inst1_r5_reg_3_ ( .D(register_file_inst1_n2460), 
        .CP(clock), .Q(register_file_inst1_r5_3_) );
  DFQD1BWP12T register_file_inst1_r5_reg_4_ ( .D(register_file_inst1_n2461), 
        .CP(clock), .Q(register_file_inst1_r5_4_) );
  DFQD1BWP12T register_file_inst1_r5_reg_5_ ( .D(register_file_inst1_n2462), 
        .CP(clock), .Q(register_file_inst1_r5_5_) );
  DFQD1BWP12T register_file_inst1_r5_reg_6_ ( .D(register_file_inst1_n2463), 
        .CP(clock), .Q(register_file_inst1_r5_6_) );
  DFQD1BWP12T register_file_inst1_r5_reg_8_ ( .D(register_file_inst1_n2465), 
        .CP(clock), .Q(register_file_inst1_r5_8_) );
  DFQD1BWP12T register_file_inst1_r5_reg_9_ ( .D(register_file_inst1_n2466), 
        .CP(clock), .Q(register_file_inst1_r5_9_) );
  DFQD1BWP12T register_file_inst1_r5_reg_10_ ( .D(register_file_inst1_n2467), 
        .CP(clock), .Q(register_file_inst1_r5_10_) );
  DFQD1BWP12T register_file_inst1_r5_reg_11_ ( .D(register_file_inst1_n2468), 
        .CP(clock), .Q(register_file_inst1_r5_11_) );
  DFQD1BWP12T register_file_inst1_r5_reg_12_ ( .D(register_file_inst1_n2469), 
        .CP(clock), .Q(register_file_inst1_r5_12_) );
  DFQD1BWP12T register_file_inst1_r5_reg_13_ ( .D(register_file_inst1_n2470), 
        .CP(clock), .Q(register_file_inst1_r5_13_) );
  DFQD1BWP12T register_file_inst1_r5_reg_14_ ( .D(register_file_inst1_n2471), 
        .CP(clock), .Q(register_file_inst1_r5_14_) );
  DFQD1BWP12T register_file_inst1_r5_reg_15_ ( .D(register_file_inst1_n2472), 
        .CP(clock), .Q(register_file_inst1_r5_15_) );
  DFQD1BWP12T register_file_inst1_r5_reg_16_ ( .D(register_file_inst1_n2473), 
        .CP(clock), .Q(register_file_inst1_r5_16_) );
  DFQD1BWP12T register_file_inst1_r5_reg_17_ ( .D(register_file_inst1_n2474), 
        .CP(clock), .Q(register_file_inst1_r5_17_) );
  DFQD1BWP12T register_file_inst1_r5_reg_18_ ( .D(register_file_inst1_n2475), 
        .CP(clock), .Q(register_file_inst1_r5_18_) );
  DFQD1BWP12T register_file_inst1_r5_reg_19_ ( .D(register_file_inst1_n2476), 
        .CP(clock), .Q(register_file_inst1_r5_19_) );
  DFQD1BWP12T register_file_inst1_r5_reg_20_ ( .D(register_file_inst1_n2477), 
        .CP(clock), .Q(register_file_inst1_r5_20_) );
  DFQD1BWP12T register_file_inst1_r5_reg_21_ ( .D(register_file_inst1_n2478), 
        .CP(clock), .Q(register_file_inst1_r5_21_) );
  DFQD1BWP12T register_file_inst1_r5_reg_22_ ( .D(register_file_inst1_n2479), 
        .CP(clock), .Q(register_file_inst1_r5_22_) );
  DFQD1BWP12T register_file_inst1_r5_reg_23_ ( .D(register_file_inst1_n2480), 
        .CP(clock), .Q(register_file_inst1_r5_23_) );
  DFQD1BWP12T register_file_inst1_r5_reg_24_ ( .D(register_file_inst1_n2481), 
        .CP(clock), .Q(register_file_inst1_r5_24_) );
  DFQD1BWP12T register_file_inst1_r5_reg_25_ ( .D(register_file_inst1_n2482), 
        .CP(clock), .Q(register_file_inst1_r5_25_) );
  DFQD1BWP12T register_file_inst1_r5_reg_26_ ( .D(register_file_inst1_n2483), 
        .CP(clock), .Q(register_file_inst1_r5_26_) );
  DFQD1BWP12T register_file_inst1_r5_reg_27_ ( .D(register_file_inst1_n2484), 
        .CP(clock), .Q(register_file_inst1_r5_27_) );
  DFQD1BWP12T register_file_inst1_r5_reg_28_ ( .D(register_file_inst1_n2485), 
        .CP(clock), .Q(register_file_inst1_r5_28_) );
  DFQD1BWP12T register_file_inst1_r5_reg_29_ ( .D(register_file_inst1_n2486), 
        .CP(clock), .Q(register_file_inst1_r5_29_) );
  DFQD1BWP12T register_file_inst1_r5_reg_30_ ( .D(register_file_inst1_n2487), 
        .CP(clock), .Q(register_file_inst1_r5_30_) );
  DFQD1BWP12T register_file_inst1_r5_reg_31_ ( .D(register_file_inst1_n2488), 
        .CP(clock), .Q(register_file_inst1_r5_31_) );
  DFQD1BWP12T register_file_inst1_r4_reg_0_ ( .D(register_file_inst1_n2489), 
        .CP(clock), .Q(register_file_inst1_r4_0_) );
  DFQD1BWP12T register_file_inst1_r4_reg_1_ ( .D(register_file_inst1_n2490), 
        .CP(clock), .Q(register_file_inst1_r4_1_) );
  DFQD1BWP12T register_file_inst1_r4_reg_2_ ( .D(register_file_inst1_n2491), 
        .CP(clock), .Q(register_file_inst1_r4_2_) );
  DFQD1BWP12T register_file_inst1_r4_reg_3_ ( .D(register_file_inst1_n2492), 
        .CP(clock), .Q(register_file_inst1_r4_3_) );
  DFQD1BWP12T register_file_inst1_r4_reg_4_ ( .D(register_file_inst1_n2493), 
        .CP(clock), .Q(register_file_inst1_r4_4_) );
  DFQD1BWP12T register_file_inst1_r4_reg_5_ ( .D(register_file_inst1_n2494), 
        .CP(clock), .Q(register_file_inst1_r4_5_) );
  DFQD1BWP12T register_file_inst1_r4_reg_6_ ( .D(register_file_inst1_n2495), 
        .CP(clock), .Q(register_file_inst1_r4_6_) );
  DFQD1BWP12T register_file_inst1_r4_reg_7_ ( .D(register_file_inst1_n2496), 
        .CP(clock), .Q(register_file_inst1_r4_7_) );
  DFQD1BWP12T register_file_inst1_r4_reg_8_ ( .D(register_file_inst1_n2497), 
        .CP(clock), .Q(register_file_inst1_r4_8_) );
  DFQD1BWP12T register_file_inst1_r4_reg_9_ ( .D(register_file_inst1_n2498), 
        .CP(clock), .Q(register_file_inst1_r4_9_) );
  DFQD1BWP12T register_file_inst1_r4_reg_10_ ( .D(register_file_inst1_n2499), 
        .CP(clock), .Q(register_file_inst1_r4_10_) );
  DFQD1BWP12T register_file_inst1_r4_reg_11_ ( .D(register_file_inst1_n2500), 
        .CP(clock), .Q(register_file_inst1_r4_11_) );
  DFQD1BWP12T register_file_inst1_r4_reg_12_ ( .D(register_file_inst1_n2501), 
        .CP(clock), .Q(register_file_inst1_r4_12_) );
  DFQD1BWP12T register_file_inst1_r4_reg_13_ ( .D(register_file_inst1_n2502), 
        .CP(clock), .Q(register_file_inst1_r4_13_) );
  DFQD1BWP12T register_file_inst1_r4_reg_14_ ( .D(register_file_inst1_n2503), 
        .CP(clock), .Q(register_file_inst1_r4_14_) );
  DFQD1BWP12T register_file_inst1_r4_reg_15_ ( .D(register_file_inst1_n2504), 
        .CP(clock), .Q(register_file_inst1_r4_15_) );
  DFQD1BWP12T register_file_inst1_r4_reg_16_ ( .D(register_file_inst1_n2505), 
        .CP(clock), .Q(register_file_inst1_r4_16_) );
  DFQD1BWP12T register_file_inst1_r4_reg_17_ ( .D(register_file_inst1_n2506), 
        .CP(clock), .Q(register_file_inst1_r4_17_) );
  DFQD1BWP12T register_file_inst1_r4_reg_18_ ( .D(register_file_inst1_n2507), 
        .CP(clock), .Q(register_file_inst1_r4_18_) );
  DFQD1BWP12T register_file_inst1_r4_reg_19_ ( .D(register_file_inst1_n2508), 
        .CP(clock), .Q(register_file_inst1_r4_19_) );
  DFQD1BWP12T register_file_inst1_r4_reg_20_ ( .D(register_file_inst1_n2509), 
        .CP(clock), .Q(register_file_inst1_r4_20_) );
  DFQD1BWP12T register_file_inst1_r4_reg_21_ ( .D(register_file_inst1_n2510), 
        .CP(clock), .Q(register_file_inst1_r4_21_) );
  DFQD1BWP12T register_file_inst1_r4_reg_22_ ( .D(register_file_inst1_n2511), 
        .CP(clock), .Q(register_file_inst1_r4_22_) );
  DFQD1BWP12T register_file_inst1_r4_reg_23_ ( .D(register_file_inst1_n2512), 
        .CP(clock), .Q(register_file_inst1_r4_23_) );
  DFQD1BWP12T register_file_inst1_r4_reg_24_ ( .D(register_file_inst1_n2513), 
        .CP(clock), .Q(register_file_inst1_r4_24_) );
  DFQD1BWP12T register_file_inst1_r4_reg_25_ ( .D(register_file_inst1_n2514), 
        .CP(clock), .Q(register_file_inst1_r4_25_) );
  DFQD1BWP12T register_file_inst1_r4_reg_26_ ( .D(register_file_inst1_n2515), 
        .CP(clock), .Q(register_file_inst1_r4_26_) );
  DFQD1BWP12T register_file_inst1_r4_reg_27_ ( .D(register_file_inst1_n2516), 
        .CP(clock), .Q(register_file_inst1_r4_27_) );
  DFQD1BWP12T register_file_inst1_r4_reg_28_ ( .D(register_file_inst1_n2517), 
        .CP(clock), .Q(register_file_inst1_r4_28_) );
  DFQD1BWP12T register_file_inst1_r4_reg_29_ ( .D(register_file_inst1_n2518), 
        .CP(clock), .Q(register_file_inst1_r4_29_) );
  DFQD1BWP12T register_file_inst1_r4_reg_30_ ( .D(register_file_inst1_n2519), 
        .CP(clock), .Q(register_file_inst1_r4_30_) );
  DFQD1BWP12T register_file_inst1_r4_reg_31_ ( .D(register_file_inst1_n2520), 
        .CP(clock), .Q(register_file_inst1_r4_31_) );
  DFQD1BWP12T register_file_inst1_r3_reg_0_ ( .D(register_file_inst1_n2521), 
        .CP(clock), .Q(register_file_inst1_r3_0_) );
  DFQD1BWP12T register_file_inst1_r3_reg_1_ ( .D(register_file_inst1_n2522), 
        .CP(clock), .Q(register_file_inst1_r3_1_) );
  DFQD1BWP12T register_file_inst1_r3_reg_2_ ( .D(register_file_inst1_n2523), 
        .CP(clock), .Q(register_file_inst1_r3_2_) );
  DFQD1BWP12T register_file_inst1_r3_reg_3_ ( .D(register_file_inst1_n2524), 
        .CP(clock), .Q(register_file_inst1_r3_3_) );
  DFQD1BWP12T register_file_inst1_r3_reg_4_ ( .D(register_file_inst1_n2525), 
        .CP(clock), .Q(register_file_inst1_r3_4_) );
  DFQD1BWP12T register_file_inst1_r3_reg_5_ ( .D(register_file_inst1_n2526), 
        .CP(clock), .Q(register_file_inst1_r3_5_) );
  DFQD1BWP12T register_file_inst1_r3_reg_6_ ( .D(register_file_inst1_n2527), 
        .CP(clock), .Q(register_file_inst1_r3_6_) );
  DFQD1BWP12T register_file_inst1_r3_reg_7_ ( .D(register_file_inst1_n2528), 
        .CP(clock), .Q(register_file_inst1_r3_7_) );
  DFQD1BWP12T register_file_inst1_r3_reg_8_ ( .D(register_file_inst1_n2529), 
        .CP(clock), .Q(register_file_inst1_r3_8_) );
  DFQD1BWP12T register_file_inst1_r3_reg_10_ ( .D(register_file_inst1_n2531), 
        .CP(clock), .Q(register_file_inst1_r3_10_) );
  DFQD1BWP12T register_file_inst1_r3_reg_11_ ( .D(register_file_inst1_n2532), 
        .CP(clock), .Q(register_file_inst1_r3_11_) );
  DFQD1BWP12T register_file_inst1_r3_reg_12_ ( .D(register_file_inst1_n2533), 
        .CP(clock), .Q(register_file_inst1_r3_12_) );
  DFQD1BWP12T register_file_inst1_r3_reg_13_ ( .D(register_file_inst1_n2534), 
        .CP(clock), .Q(register_file_inst1_r3_13_) );
  DFQD1BWP12T register_file_inst1_r3_reg_14_ ( .D(register_file_inst1_n2535), 
        .CP(clock), .Q(register_file_inst1_r3_14_) );
  DFQD1BWP12T register_file_inst1_r3_reg_15_ ( .D(register_file_inst1_n2536), 
        .CP(clock), .Q(register_file_inst1_r3_15_) );
  DFQD1BWP12T register_file_inst1_r3_reg_16_ ( .D(register_file_inst1_n2537), 
        .CP(clock), .Q(register_file_inst1_r3_16_) );
  DFQD1BWP12T register_file_inst1_r3_reg_17_ ( .D(register_file_inst1_n2538), 
        .CP(clock), .Q(register_file_inst1_r3_17_) );
  DFQD1BWP12T register_file_inst1_r3_reg_18_ ( .D(register_file_inst1_n2539), 
        .CP(clock), .Q(register_file_inst1_r3_18_) );
  DFQD1BWP12T register_file_inst1_r3_reg_19_ ( .D(register_file_inst1_n2540), 
        .CP(clock), .Q(register_file_inst1_r3_19_) );
  DFQD1BWP12T register_file_inst1_r3_reg_20_ ( .D(register_file_inst1_n2541), 
        .CP(clock), .Q(register_file_inst1_r3_20_) );
  DFQD1BWP12T register_file_inst1_r3_reg_21_ ( .D(register_file_inst1_n2542), 
        .CP(clock), .Q(register_file_inst1_r3_21_) );
  DFQD1BWP12T register_file_inst1_r3_reg_22_ ( .D(register_file_inst1_n2543), 
        .CP(clock), .Q(register_file_inst1_r3_22_) );
  DFQD1BWP12T register_file_inst1_r3_reg_23_ ( .D(register_file_inst1_n2544), 
        .CP(clock), .Q(register_file_inst1_r3_23_) );
  DFQD1BWP12T register_file_inst1_r3_reg_24_ ( .D(register_file_inst1_n2545), 
        .CP(clock), .Q(register_file_inst1_r3_24_) );
  DFQD1BWP12T register_file_inst1_r3_reg_25_ ( .D(register_file_inst1_n2546), 
        .CP(clock), .Q(register_file_inst1_r3_25_) );
  DFQD1BWP12T register_file_inst1_r3_reg_26_ ( .D(register_file_inst1_n2547), 
        .CP(clock), .Q(register_file_inst1_r3_26_) );
  DFQD1BWP12T register_file_inst1_r3_reg_27_ ( .D(register_file_inst1_n2548), 
        .CP(clock), .Q(register_file_inst1_r3_27_) );
  DFQD1BWP12T register_file_inst1_r3_reg_28_ ( .D(register_file_inst1_n2549), 
        .CP(clock), .Q(register_file_inst1_r3_28_) );
  DFQD1BWP12T register_file_inst1_r3_reg_29_ ( .D(register_file_inst1_n2550), 
        .CP(clock), .Q(register_file_inst1_r3_29_) );
  DFQD1BWP12T register_file_inst1_r3_reg_30_ ( .D(register_file_inst1_n2551), 
        .CP(clock), .Q(register_file_inst1_r3_30_) );
  DFQD1BWP12T register_file_inst1_r3_reg_31_ ( .D(register_file_inst1_n2552), 
        .CP(clock), .Q(register_file_inst1_r3_31_) );
  DFQD1BWP12T register_file_inst1_r2_reg_1_ ( .D(register_file_inst1_n2554), 
        .CP(clock), .Q(register_file_inst1_r2_1_) );
  DFQD1BWP12T register_file_inst1_r2_reg_2_ ( .D(register_file_inst1_n2555), 
        .CP(clock), .Q(register_file_inst1_r2_2_) );
  DFQD1BWP12T register_file_inst1_r2_reg_3_ ( .D(register_file_inst1_n2556), 
        .CP(clock), .Q(register_file_inst1_r2_3_) );
  DFQD1BWP12T register_file_inst1_r2_reg_4_ ( .D(register_file_inst1_n2557), 
        .CP(clock), .Q(register_file_inst1_r2_4_) );
  DFQD1BWP12T register_file_inst1_r2_reg_5_ ( .D(register_file_inst1_n2558), 
        .CP(clock), .Q(register_file_inst1_r2_5_) );
  DFQD1BWP12T register_file_inst1_r2_reg_6_ ( .D(register_file_inst1_n2559), 
        .CP(clock), .Q(register_file_inst1_r2_6_) );
  DFQD1BWP12T register_file_inst1_r2_reg_7_ ( .D(register_file_inst1_n2560), 
        .CP(clock), .Q(register_file_inst1_r2_7_) );
  DFQD1BWP12T register_file_inst1_r2_reg_8_ ( .D(register_file_inst1_n2561), 
        .CP(clock), .Q(register_file_inst1_r2_8_) );
  DFQD1BWP12T register_file_inst1_r2_reg_9_ ( .D(register_file_inst1_n2562), 
        .CP(clock), .Q(register_file_inst1_r2_9_) );
  DFQD1BWP12T register_file_inst1_r2_reg_10_ ( .D(register_file_inst1_n2563), 
        .CP(clock), .Q(register_file_inst1_r2_10_) );
  DFQD1BWP12T register_file_inst1_r2_reg_11_ ( .D(register_file_inst1_n2564), 
        .CP(clock), .Q(register_file_inst1_r2_11_) );
  DFQD1BWP12T register_file_inst1_r2_reg_12_ ( .D(register_file_inst1_n2565), 
        .CP(clock), .Q(register_file_inst1_r2_12_) );
  DFQD1BWP12T register_file_inst1_r2_reg_13_ ( .D(register_file_inst1_n2566), 
        .CP(clock), .Q(register_file_inst1_r2_13_) );
  DFQD1BWP12T register_file_inst1_r2_reg_14_ ( .D(register_file_inst1_n2567), 
        .CP(clock), .Q(register_file_inst1_r2_14_) );
  DFQD1BWP12T register_file_inst1_r2_reg_15_ ( .D(register_file_inst1_n2568), 
        .CP(clock), .Q(register_file_inst1_r2_15_) );
  DFQD1BWP12T register_file_inst1_r2_reg_16_ ( .D(register_file_inst1_n2569), 
        .CP(clock), .Q(register_file_inst1_r2_16_) );
  DFQD1BWP12T register_file_inst1_r2_reg_17_ ( .D(register_file_inst1_n2570), 
        .CP(clock), .Q(register_file_inst1_r2_17_) );
  DFQD1BWP12T register_file_inst1_r2_reg_18_ ( .D(register_file_inst1_n2571), 
        .CP(clock), .Q(register_file_inst1_r2_18_) );
  DFQD1BWP12T register_file_inst1_r2_reg_19_ ( .D(register_file_inst1_n2572), 
        .CP(clock), .Q(register_file_inst1_r2_19_) );
  DFQD1BWP12T register_file_inst1_r2_reg_20_ ( .D(register_file_inst1_n2573), 
        .CP(clock), .Q(register_file_inst1_r2_20_) );
  DFQD1BWP12T register_file_inst1_r2_reg_21_ ( .D(register_file_inst1_n2574), 
        .CP(clock), .Q(register_file_inst1_r2_21_) );
  DFQD1BWP12T register_file_inst1_r2_reg_22_ ( .D(register_file_inst1_n2575), 
        .CP(clock), .Q(register_file_inst1_r2_22_) );
  DFQD1BWP12T register_file_inst1_r2_reg_23_ ( .D(register_file_inst1_n2576), 
        .CP(clock), .Q(register_file_inst1_r2_23_) );
  DFQD1BWP12T register_file_inst1_r2_reg_24_ ( .D(register_file_inst1_n2577), 
        .CP(clock), .Q(register_file_inst1_r2_24_) );
  DFQD1BWP12T register_file_inst1_r2_reg_25_ ( .D(register_file_inst1_n2578), 
        .CP(clock), .Q(register_file_inst1_r2_25_) );
  DFQD1BWP12T register_file_inst1_r2_reg_26_ ( .D(register_file_inst1_n2579), 
        .CP(clock), .Q(register_file_inst1_r2_26_) );
  DFQD1BWP12T register_file_inst1_r2_reg_27_ ( .D(register_file_inst1_n2580), 
        .CP(clock), .Q(register_file_inst1_r2_27_) );
  DFQD1BWP12T register_file_inst1_r2_reg_28_ ( .D(register_file_inst1_n2581), 
        .CP(clock), .Q(register_file_inst1_r2_28_) );
  DFQD1BWP12T register_file_inst1_r2_reg_29_ ( .D(register_file_inst1_n2582), 
        .CP(clock), .Q(register_file_inst1_r2_29_) );
  DFQD1BWP12T register_file_inst1_r2_reg_30_ ( .D(register_file_inst1_n2583), 
        .CP(clock), .Q(register_file_inst1_r2_30_) );
  DFQD1BWP12T register_file_inst1_r2_reg_31_ ( .D(register_file_inst1_n2584), 
        .CP(clock), .Q(register_file_inst1_r2_31_) );
  DFQD1BWP12T register_file_inst1_r1_reg_0_ ( .D(register_file_inst1_n2585), 
        .CP(clock), .Q(register_file_inst1_r1_0_) );
  DFQD1BWP12T register_file_inst1_r1_reg_1_ ( .D(register_file_inst1_n2586), 
        .CP(clock), .Q(register_file_inst1_r1_1_) );
  DFQD1BWP12T register_file_inst1_r1_reg_2_ ( .D(register_file_inst1_n2587), 
        .CP(clock), .Q(register_file_inst1_r1_2_) );
  DFQD1BWP12T register_file_inst1_r1_reg_3_ ( .D(register_file_inst1_n2588), 
        .CP(clock), .Q(register_file_inst1_r1_3_) );
  DFQD1BWP12T register_file_inst1_r1_reg_4_ ( .D(register_file_inst1_n2589), 
        .CP(clock), .Q(register_file_inst1_r1_4_) );
  DFQD1BWP12T register_file_inst1_r1_reg_5_ ( .D(register_file_inst1_n2590), 
        .CP(clock), .Q(register_file_inst1_r1_5_) );
  DFQD1BWP12T register_file_inst1_r1_reg_6_ ( .D(register_file_inst1_n2591), 
        .CP(clock), .Q(register_file_inst1_r1_6_) );
  DFQD1BWP12T register_file_inst1_r1_reg_7_ ( .D(register_file_inst1_n2592), 
        .CP(clock), .Q(register_file_inst1_r1_7_) );
  DFQD1BWP12T register_file_inst1_r1_reg_8_ ( .D(register_file_inst1_n2593), 
        .CP(clock), .Q(register_file_inst1_r1_8_) );
  DFQD1BWP12T register_file_inst1_r1_reg_9_ ( .D(register_file_inst1_n2594), 
        .CP(clock), .Q(register_file_inst1_r1_9_) );
  DFQD1BWP12T register_file_inst1_r1_reg_10_ ( .D(register_file_inst1_n2595), 
        .CP(clock), .Q(register_file_inst1_r1_10_) );
  DFQD1BWP12T register_file_inst1_r1_reg_11_ ( .D(register_file_inst1_n2596), 
        .CP(clock), .Q(register_file_inst1_r1_11_) );
  DFQD1BWP12T register_file_inst1_r1_reg_12_ ( .D(register_file_inst1_n2597), 
        .CP(clock), .Q(register_file_inst1_r1_12_) );
  DFQD1BWP12T register_file_inst1_r1_reg_13_ ( .D(register_file_inst1_n2598), 
        .CP(clock), .Q(register_file_inst1_r1_13_) );
  DFQD1BWP12T register_file_inst1_r1_reg_14_ ( .D(register_file_inst1_n2599), 
        .CP(clock), .Q(register_file_inst1_r1_14_) );
  DFQD1BWP12T register_file_inst1_r1_reg_15_ ( .D(register_file_inst1_n2600), 
        .CP(clock), .Q(register_file_inst1_r1_15_) );
  DFQD1BWP12T register_file_inst1_r1_reg_16_ ( .D(register_file_inst1_n2601), 
        .CP(clock), .Q(register_file_inst1_r1_16_) );
  DFQD1BWP12T register_file_inst1_r1_reg_17_ ( .D(register_file_inst1_n2602), 
        .CP(clock), .Q(register_file_inst1_r1_17_) );
  DFQD1BWP12T register_file_inst1_r1_reg_18_ ( .D(register_file_inst1_n2603), 
        .CP(clock), .Q(register_file_inst1_r1_18_) );
  DFQD1BWP12T register_file_inst1_r1_reg_19_ ( .D(register_file_inst1_n2604), 
        .CP(clock), .Q(register_file_inst1_r1_19_) );
  DFQD1BWP12T register_file_inst1_r1_reg_20_ ( .D(register_file_inst1_n2605), 
        .CP(clock), .Q(register_file_inst1_r1_20_) );
  DFQD1BWP12T register_file_inst1_r1_reg_21_ ( .D(register_file_inst1_n2606), 
        .CP(clock), .Q(register_file_inst1_r1_21_) );
  DFQD1BWP12T register_file_inst1_r1_reg_22_ ( .D(register_file_inst1_n2607), 
        .CP(clock), .Q(register_file_inst1_r1_22_) );
  DFQD1BWP12T register_file_inst1_r1_reg_23_ ( .D(register_file_inst1_n2608), 
        .CP(clock), .Q(register_file_inst1_r1_23_) );
  DFQD1BWP12T register_file_inst1_r1_reg_24_ ( .D(register_file_inst1_n2609), 
        .CP(clock), .Q(register_file_inst1_r1_24_) );
  DFQD1BWP12T register_file_inst1_r1_reg_25_ ( .D(register_file_inst1_n2610), 
        .CP(clock), .Q(register_file_inst1_r1_25_) );
  DFQD1BWP12T register_file_inst1_r1_reg_26_ ( .D(register_file_inst1_n2611), 
        .CP(clock), .Q(register_file_inst1_r1_26_) );
  DFQD1BWP12T register_file_inst1_r1_reg_27_ ( .D(register_file_inst1_n2612), 
        .CP(clock), .Q(register_file_inst1_r1_27_) );
  DFQD1BWP12T register_file_inst1_r1_reg_28_ ( .D(register_file_inst1_n2613), 
        .CP(clock), .Q(register_file_inst1_r1_28_) );
  DFQD1BWP12T register_file_inst1_r1_reg_29_ ( .D(register_file_inst1_n2614), 
        .CP(clock), .Q(register_file_inst1_r1_29_) );
  DFQD1BWP12T register_file_inst1_r1_reg_30_ ( .D(register_file_inst1_n2615), 
        .CP(clock), .Q(register_file_inst1_r1_30_) );
  DFQD1BWP12T register_file_inst1_r1_reg_31_ ( .D(register_file_inst1_n2616), 
        .CP(clock), .Q(register_file_inst1_r1_31_) );
  DFQD1BWP12T register_file_inst1_r0_reg_0_ ( .D(register_file_inst1_n2617), 
        .CP(clock), .Q(register_file_inst1_r0_0_) );
  DFQD1BWP12T register_file_inst1_r0_reg_1_ ( .D(register_file_inst1_n2618), 
        .CP(clock), .Q(register_file_inst1_r0_1_) );
  DFQD1BWP12T register_file_inst1_r0_reg_2_ ( .D(register_file_inst1_n2619), 
        .CP(clock), .Q(register_file_inst1_r0_2_) );
  DFQD1BWP12T register_file_inst1_r0_reg_3_ ( .D(register_file_inst1_n2620), 
        .CP(clock), .Q(register_file_inst1_r0_3_) );
  DFQD1BWP12T register_file_inst1_r0_reg_4_ ( .D(register_file_inst1_n2621), 
        .CP(clock), .Q(register_file_inst1_r0_4_) );
  DFQD1BWP12T register_file_inst1_r0_reg_5_ ( .D(register_file_inst1_n2622), 
        .CP(clock), .Q(register_file_inst1_r0_5_) );
  DFQD1BWP12T register_file_inst1_r0_reg_6_ ( .D(register_file_inst1_n2623), 
        .CP(clock), .Q(register_file_inst1_r0_6_) );
  DFQD1BWP12T register_file_inst1_r0_reg_7_ ( .D(register_file_inst1_n2624), 
        .CP(clock), .Q(register_file_inst1_r0_7_) );
  DFQD1BWP12T register_file_inst1_r0_reg_8_ ( .D(register_file_inst1_n2625), 
        .CP(clock), .Q(register_file_inst1_r0_8_) );
  DFQD1BWP12T register_file_inst1_r0_reg_9_ ( .D(register_file_inst1_n2626), 
        .CP(clock), .Q(register_file_inst1_r0_9_) );
  DFQD1BWP12T register_file_inst1_r0_reg_10_ ( .D(register_file_inst1_n2627), 
        .CP(clock), .Q(register_file_inst1_r0_10_) );
  DFQD1BWP12T register_file_inst1_r0_reg_11_ ( .D(register_file_inst1_n2628), 
        .CP(clock), .Q(register_file_inst1_r0_11_) );
  DFQD1BWP12T register_file_inst1_r0_reg_12_ ( .D(register_file_inst1_n2629), 
        .CP(clock), .Q(register_file_inst1_r0_12_) );
  DFQD1BWP12T register_file_inst1_r0_reg_13_ ( .D(register_file_inst1_n2630), 
        .CP(clock), .Q(register_file_inst1_r0_13_) );
  DFQD1BWP12T register_file_inst1_r0_reg_14_ ( .D(register_file_inst1_n2631), 
        .CP(clock), .Q(register_file_inst1_r0_14_) );
  DFQD1BWP12T register_file_inst1_r0_reg_15_ ( .D(register_file_inst1_n2632), 
        .CP(clock), .Q(register_file_inst1_r0_15_) );
  DFQD1BWP12T register_file_inst1_r0_reg_16_ ( .D(register_file_inst1_n2633), 
        .CP(clock), .Q(register_file_inst1_r0_16_) );
  DFQD1BWP12T register_file_inst1_r0_reg_17_ ( .D(register_file_inst1_n2634), 
        .CP(clock), .Q(register_file_inst1_r0_17_) );
  DFQD1BWP12T register_file_inst1_r0_reg_18_ ( .D(register_file_inst1_n2635), 
        .CP(clock), .Q(register_file_inst1_r0_18_) );
  DFQD1BWP12T register_file_inst1_r0_reg_19_ ( .D(register_file_inst1_n2636), 
        .CP(clock), .Q(register_file_inst1_r0_19_) );
  DFQD1BWP12T register_file_inst1_r0_reg_20_ ( .D(register_file_inst1_n2637), 
        .CP(clock), .Q(register_file_inst1_r0_20_) );
  DFQD1BWP12T register_file_inst1_r0_reg_21_ ( .D(register_file_inst1_n2638), 
        .CP(clock), .Q(register_file_inst1_r0_21_) );
  DFQD1BWP12T register_file_inst1_r0_reg_22_ ( .D(register_file_inst1_n2639), 
        .CP(clock), .Q(register_file_inst1_r0_22_) );
  DFQD1BWP12T register_file_inst1_r0_reg_23_ ( .D(register_file_inst1_n2640), 
        .CP(clock), .Q(register_file_inst1_r0_23_) );
  DFQD1BWP12T register_file_inst1_r0_reg_24_ ( .D(register_file_inst1_n2641), 
        .CP(clock), .Q(register_file_inst1_r0_24_) );
  DFQD1BWP12T register_file_inst1_r0_reg_25_ ( .D(register_file_inst1_n2642), 
        .CP(clock), .Q(register_file_inst1_r0_25_) );
  DFQD1BWP12T register_file_inst1_r0_reg_26_ ( .D(register_file_inst1_n2643), 
        .CP(clock), .Q(register_file_inst1_r0_26_) );
  DFQD1BWP12T register_file_inst1_r0_reg_27_ ( .D(register_file_inst1_n2644), 
        .CP(clock), .Q(register_file_inst1_r0_27_) );
  DFQD1BWP12T register_file_inst1_r0_reg_28_ ( .D(register_file_inst1_n2645), 
        .CP(clock), .Q(register_file_inst1_r0_28_) );
  DFQD1BWP12T register_file_inst1_r0_reg_29_ ( .D(register_file_inst1_n2646), 
        .CP(clock), .Q(register_file_inst1_r0_29_) );
  DFQD1BWP12T register_file_inst1_r0_reg_30_ ( .D(register_file_inst1_n2647), 
        .CP(clock), .Q(register_file_inst1_r0_30_) );
  DFQD1BWP12T register_file_inst1_r0_reg_31_ ( .D(register_file_inst1_n2648), 
        .CP(clock), .Q(register_file_inst1_r0_31_) );
  DFQD1BWP12T register_file_inst1_r2_reg_0_ ( .D(register_file_inst1_n2553), 
        .CP(clock), .Q(register_file_inst1_r2_0_) );
  DFQD1BWP12T register_file_inst1_r7_reg_3_ ( .D(register_file_inst1_n2396), 
        .CP(clock), .Q(register_file_inst1_r7_3_) );
  DFQD1BWP12T register_file_inst1_r3_reg_9_ ( .D(register_file_inst1_n2530), 
        .CP(clock), .Q(register_file_inst1_r3_9_) );
  AO211D0BWP12T U2778 ( .A1(memory_interface_inst1_fsm_state_0_), .A2(n6400), 
        .B(n6399), .C(n5985), .Z(MEMCTRL_read_finished) );
  OAI21D1BWP12T U2975 ( .A1(n6407), .A2(n5985), .B(n2265), .ZN(
        MEMCTRL_RF_IF_data_in[7]) );
  AOI211D1BWP12T U2993 ( .A1(n4090), .A2(n2244), .B(n2243), .C(n6401), .ZN(
        MEMCTRL_write_finished) );
  OAI211D1BWP12T U3003 ( .A1(n2264), .A2(n4101), .B(n2262), .C(n2255), .ZN(
        MEMCTRL_RF_IF_data_in[11]) );
  OAI211D1BWP12T U3004 ( .A1(n2264), .A2(n4100), .B(n2262), .C(n2253), .ZN(
        MEMCTRL_RF_IF_data_in[12]) );
  OAI211D1BWP12T U3005 ( .A1(n2264), .A2(n4099), .B(n2262), .C(n2251), .ZN(
        MEMCTRL_RF_IF_data_in[13]) );
  OAI211D1BWP12T U3006 ( .A1(n2264), .A2(n4098), .B(n2262), .C(n2249), .ZN(
        MEMCTRL_RF_IF_data_in[14]) );
  OAI211D1BWP12T U3007 ( .A1(n2264), .A2(n4097), .B(n2262), .C(n2247), .ZN(
        MEMCTRL_RF_IF_data_in[15]) );
  OAI211D1BWP12T U3008 ( .A1(n2264), .A2(n4104), .B(n2262), .C(n2261), .ZN(
        MEMCTRL_RF_IF_data_in[8]) );
  OAI211D1BWP12T U3009 ( .A1(n2264), .A2(n4103), .B(n2262), .C(n2259), .ZN(
        MEMCTRL_RF_IF_data_in[9]) );
  OAI211D1BWP12T U3010 ( .A1(n2264), .A2(n4102), .B(n2262), .C(n2257), .ZN(
        MEMCTRL_RF_IF_data_in[10]) );
  DFQD4BWP12T register_file_inst1_r8_reg_15_ ( .D(register_file_inst1_n2376), 
        .CP(clock), .Q(register_file_inst1_r8_15_) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_0_ ( .D(
        memory_interface_inst1_fsm_N32), .CP(clock), .Q(
        memory_interface_inst1_fsm_state_0_) );
  INR2D1BWP12T U370 ( .A1(DEC_RF_operand_b[3]), .B1(DEC_RF_operand_b[4]), .ZN(
        n2515) );
  NR2D1BWP12T U818 ( .A1(DEC_RF_memory_write_to_reg[3]), .A2(n2880), .ZN(n2876) );
  NR2D1BWP12T U366 ( .A1(DEC_RF_operand_b[4]), .A2(DEC_RF_operand_b[3]), .ZN(
        n2516) );
  NR2D1BWP12T U297 ( .A1(DEC_RF_operand_a[3]), .A2(DEC_RF_operand_a[4]), .ZN(
        n2470) );
  NR2D1BWP12T U315 ( .A1(DEC_RF_operand_a[4]), .A2(n6402), .ZN(n2471) );
  NR2D1BWP12T U305 ( .A1(DEC_RF_operand_a[0]), .A2(DEC_RF_operand_a[4]), .ZN(
        n2469) );
  AOI22D1BWP12T U1530 ( .A1(ALU_MISC_OUT_result[10]), .A2(n6396), .B1(
        IF_memory_load_req), .B2(IF_instruction_memory_address[9]), .ZN(n3420)
         );
  ND2D1BWP12T U1085 ( .A1(DEC_RF_memory_store_address_reg[0]), .A2(
        DEC_RF_memory_store_address_reg[1]), .ZN(n3054) );
  INVD1BWP12T U1086 ( .I(DEC_RF_memory_store_address_reg[2]), .ZN(n3046) );
  INVD1BWP12T U1097 ( .I(DEC_RF_memory_store_address_reg[3]), .ZN(n3047) );
  ND2D1BWP12T U1093 ( .A1(DEC_RF_memory_store_address_reg[3]), .A2(
        DEC_RF_memory_store_address_reg[2]), .ZN(n3059) );
  INVD1BWP12T U1095 ( .I(DEC_RF_memory_store_address_reg[1]), .ZN(n3048) );
  INVD1BWP12T U1089 ( .I(DEC_RF_memory_store_address_reg[0]), .ZN(n3049) );
  ND2D1BWP12T U1098 ( .A1(DEC_RF_memory_store_address_reg[2]), .A2(n3047), 
        .ZN(n3060) );
  ND2D1BWP12T U1087 ( .A1(DEC_RF_memory_store_address_reg[3]), .A2(n3046), 
        .ZN(n3055) );
  ND2D1BWP12T U1096 ( .A1(DEC_RF_memory_store_address_reg[0]), .A2(n3048), 
        .ZN(n3056) );
  ND2D1BWP12T U1090 ( .A1(DEC_RF_memory_store_address_reg[1]), .A2(n3049), 
        .ZN(n3061) );
  AOI22D1BWP12T U1248 ( .A1(ALU_MISC_OUT_result[6]), .A2(n6396), .B1(
        IF_memory_load_req), .B2(IF_instruction_memory_address[5]), .ZN(n3165)
         );
  AOI22D1BWP12T U1560 ( .A1(ALU_MISC_OUT_result[4]), .A2(n6396), .B1(
        IF_memory_load_req), .B2(IF_instruction_memory_address[3]), .ZN(n3467)
         );
  AOI22D1BWP12T U1167 ( .A1(ALU_MISC_OUT_result[2]), .A2(n6396), .B1(
        IF_memory_load_req), .B2(IF_instruction_memory_address[1]), .ZN(n3095)
         );
  AOI22D1BWP12T U1289 ( .A1(ALU_MISC_OUT_result[3]), .A2(n6396), .B1(
        IF_memory_load_req), .B2(IF_instruction_memory_address[2]), .ZN(n3202)
         );
  NR2D1BWP12T U184 ( .A1(IF_memory_load_req), .A2(
        DEC_MEMCTRL_memory_load_request), .ZN(n2342) );
  INVD1BWP12T U190 ( .I(DEC_MEMCTRL_memory_store_request), .ZN(n3017) );
  OAI32D1BWP12T U191 ( .A1(n6406), .A2(DEC_MEMCTRL_load_store_width[1]), .A3(
        n3017), .B1(n2342), .B2(DEC_MEMCTRL_load_store_width[0]), .ZN(n2343)
         );
  INVD1BWP12T U906 ( .I(DEC_RF_memory_store_data_reg[1]), .ZN(n2905) );
  ND2D1BWP12T U907 ( .A1(DEC_RF_memory_store_data_reg[0]), .A2(n2905), .ZN(
        n2909) );
  INVD1BWP12T U921 ( .I(DEC_RF_memory_store_data_reg[3]), .ZN(n2907) );
  INVD1BWP12T U908 ( .I(DEC_RF_memory_store_data_reg[2]), .ZN(n2908) );
  ND2D1BWP12T U902 ( .A1(DEC_RF_memory_store_data_reg[1]), .A2(
        DEC_RF_memory_store_data_reg[0]), .ZN(n2911) );
  INVD1BWP12T U913 ( .I(DEC_RF_memory_store_data_reg[0]), .ZN(n2906) );
  ND2D1BWP12T U918 ( .A1(DEC_RF_memory_store_data_reg[1]), .A2(n2906), .ZN(
        n2920) );
  ND2D1BWP12T U922 ( .A1(DEC_RF_memory_store_data_reg[2]), .A2(n2907), .ZN(
        n2912) );
  ND3D1BWP12T U904 ( .A1(DEC_RF_memory_store_data_reg[2]), .A2(
        DEC_RF_memory_store_data_reg[3]), .A3(n3502), .ZN(n2919) );
  ND3D1BWP12T U909 ( .A1(DEC_RF_memory_store_data_reg[3]), .A2(n3502), .A3(
        n2908), .ZN(n2917) );
  OAI21D1BWP12T U1050 ( .A1(DEC_MEMCTRL_load_store_width[0]), .A2(
        DEC_MEMCTRL_load_store_width[1]), .B(n6398), .ZN(n3018) );
  NR2D1BWP12T U58 ( .A1(DEC_RF_alu_write_to_reg[4]), .A2(n3519), .ZN(n2878) );
  IND2D1BWP12T U845 ( .A1(DEC_RF_alu_write_to_reg[2]), .B1(
        DEC_RF_alu_write_to_reg[1]), .ZN(n3510) );
  IND2D1BWP12T U52 ( .A1(DEC_RF_memory_write_to_reg[4]), .B1(
        DEC_RF_memory_write_to_reg_enable), .ZN(n2880) );
  MAOI22D0BWP12T U183 ( .A1(DEC_MEMCTRL_load_store_width[0]), .A2(
        DEC_MEMCTRL_load_store_width[1]), .B1(DEC_MEMCTRL_load_store_width[0]), 
        .B2(DEC_MEMCTRL_load_store_width[1]), .ZN(n2348) );
  AN2D1BWP12T U1080 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[0]), .Z(MEMCTRL_IN_address[0]) );
  NR2D1BWP12T U795 ( .A1(reset), .A2(DEC_RF_alu_write_to_reg[1]), .ZN(n2874)
         );
  NR2D0BWP12T U1588 ( .A1(DEC_RF_memory_write_to_reg[0]), .A2(n6403), .ZN(
        n3521) );
  MUX2D0BWP12T U3017 ( .I0(MEM_MEMCTRL_from_mem_data[11]), .I1(
        memory_interface_inst1_delay_first_two_bytes_out[3]), .S(n5985), .Z(
        MEMCTRL_RF_IF_data_in[3]) );
  MUX2D0BWP12T U3018 ( .I0(MEM_MEMCTRL_from_mem_data[10]), .I1(
        memory_interface_inst1_delay_first_two_bytes_out[2]), .S(n5985), .Z(
        MEMCTRL_RF_IF_data_in[2]) );
  MUX2D0BWP12T U3016 ( .I0(MEM_MEMCTRL_from_mem_data[9]), .I1(
        memory_interface_inst1_delay_first_two_bytes_out[1]), .S(n5985), .Z(
        MEMCTRL_RF_IF_data_in[1]) );
  TPOAI21D0BWP12T U2977 ( .A1(n5985), .A2(n4095), .B(n2268), .ZN(
        MEMCTRL_RF_IF_data_in[4]) );
  TPOAI21D0BWP12T U2978 ( .A1(n5985), .A2(n4094), .B(n2267), .ZN(
        MEMCTRL_RF_IF_data_in[5]) );
  OAI21D0BWP12T U2976 ( .A1(n5985), .A2(n4096), .B(n2269), .ZN(
        MEMCTRL_RF_IF_data_in[0]) );
  TPOAI21D0BWP12T U2979 ( .A1(n5985), .A2(n4093), .B(n2266), .ZN(
        MEMCTRL_RF_IF_data_in[6]) );
  AO222D1BWP12T U244 ( .A1(n2396), .A2(n6395), .B1(n6007), .B2(RF_pc_out[0]), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[0]), .Z(
        register_file_inst1_n2169) );
  AOI22D0BWP12T U1384 ( .A1(ALU_MISC_OUT_result[5]), .A2(n6396), .B1(
        IF_memory_load_req), .B2(IF_instruction_memory_address[4]), .ZN(n3286)
         );
  AOI22D0BWP12T U1305 ( .A1(ALU_MISC_OUT_result[8]), .A2(n6396), .B1(
        IF_memory_load_req), .B2(IF_instruction_memory_address[7]), .ZN(n3217)
         );
  AOI22D0BWP12T U1439 ( .A1(ALU_MISC_OUT_result[7]), .A2(n6396), .B1(
        IF_memory_load_req), .B2(IF_instruction_memory_address[6]), .ZN(n3335)
         );
  AOI22D0BWP12T U1126 ( .A1(ALU_MISC_OUT_result[9]), .A2(n6396), .B1(
        IF_memory_load_req), .B2(IF_instruction_memory_address[8]), .ZN(n3068)
         );
  DFQD1BWP12T register_file_inst1_r7_reg_9_ ( .D(register_file_inst1_n2402), 
        .CP(clock), .Q(register_file_inst1_r7_9_) );
  DFQD1BWP12T register_file_inst1_r6_reg_9_ ( .D(register_file_inst1_n2434), 
        .CP(clock), .Q(register_file_inst1_r6_9_) );
  DFQD1BWP12T register_file_inst1_r8_reg_8_ ( .D(register_file_inst1_n2369), 
        .CP(clock), .Q(register_file_inst1_r8_8_) );
  DFQD2BWP12T register_file_inst1_r10_reg_7_ ( .D(register_file_inst1_n2304), 
        .CP(clock), .Q(register_file_inst1_r10_7_) );
  DFQD1BWP12T register_file_inst1_r11_reg_9_ ( .D(register_file_inst1_n2274), 
        .CP(clock), .Q(register_file_inst1_r11_9_) );
  DFQD1BWP12T register_file_inst1_r8_reg_2_ ( .D(register_file_inst1_n2363), 
        .CP(clock), .Q(register_file_inst1_r8_2_) );
  DFQD1BWP12T register_file_inst1_lr_reg_6_ ( .D(register_file_inst1_n2207), 
        .CP(clock), .Q(register_file_inst1_lr_6_) );
  DFQD1BWP12T register_file_inst1_r8_reg_11_ ( .D(register_file_inst1_n2372), 
        .CP(clock), .Q(register_file_inst1_r8_11_) );
  DFQD1BWP12T register_file_inst1_r5_reg_7_ ( .D(register_file_inst1_n2464), 
        .CP(clock), .Q(register_file_inst1_r5_7_) );
  DFQD1BWP12T register_file_inst1_r12_reg_2_ ( .D(register_file_inst1_n2235), 
        .CP(clock), .Q(register_file_inst1_r12_2_) );
  DFQD1BWP12T register_file_inst1_lr_reg_12_ ( .D(register_file_inst1_n2213), 
        .CP(clock), .Q(register_file_inst1_lr_12_) );
  DFQD1BWP12T register_file_inst1_r11_reg_7_ ( .D(register_file_inst1_n2272), 
        .CP(clock), .Q(register_file_inst1_r11_7_) );
  TIELBWP12T U2511 ( .ZN(n4106) );
  INVD1BWP12T U2512 ( .I(n4106), .ZN(MEMCTRL_MEM_to_mem_mem_enable) );
  NR2D1BWP12T U2513 ( .A1(ALU_MISC_OUT_result[10]), .A2(n5984), .ZN(n4124) );
  OAI22D1BWP12T U2514 ( .A1(n5804), .A2(n5959), .B1(n5803), .B2(n5912), .ZN(
        n5809) );
  AOI22D1BWP12T U2515 ( .A1(register_file_inst1_r5_13_), .A2(n5948), .B1(
        register_file_inst1_r8_13_), .B2(n6230), .ZN(n5593) );
  AOI22D1BWP12T U2516 ( .A1(RF_pc_out[13]), .A2(n6006), .B1(
        register_file_inst1_r12_13_), .B2(n6228), .ZN(n6187) );
  AOI22D1BWP12T U2517 ( .A1(RF_pc_out[1]), .A2(n5996), .B1(
        register_file_inst1_r10_1_), .B2(n5995), .ZN(n6055) );
  OR4XD1BWP12T U2518 ( .A1(n5548), .A2(n5547), .A3(n5546), .A4(n5545), .Z(
        RF_ALU_operand_a[16]) );
  ND4D1BWP12T U2519 ( .A1(n5841), .A2(n5840), .A3(n5839), .A4(n5838), .ZN(
        RF_ALU_operand_a[1]) );
  AOI22D1BWP12T U2520 ( .A1(RF_pc_out[16]), .A2(n5996), .B1(
        register_file_inst1_r10_16_), .B2(n5995), .ZN(n6115) );
  AOI22D1BWP12T U2521 ( .A1(RF_pc_out[20]), .A2(n5996), .B1(
        register_file_inst1_r10_20_), .B2(n5995), .ZN(n6123) );
  NR2D1BWP12T U2522 ( .A1(ALU_MISC_OUT_result[3]), .A2(n5984), .ZN(n4125) );
  OR4XD1BWP12T U2523 ( .A1(n5856), .A2(n5855), .A3(n5854), .A4(n5853), .Z(
        RF_ALU_operand_a[0]) );
  AOI22D1BWP12T U2524 ( .A1(RF_pc_out[9]), .A2(n5996), .B1(
        register_file_inst1_r5_9_), .B2(n6002), .ZN(n6088) );
  AOI22D1BWP12T U2525 ( .A1(RF_pc_out[25]), .A2(n5996), .B1(
        register_file_inst1_r10_25_), .B2(n5995), .ZN(n6133) );
  AOI22D1BWP12T U2526 ( .A1(RF_pc_out[27]), .A2(n5996), .B1(
        register_file_inst1_r10_27_), .B2(n5995), .ZN(n6137) );
  AOI22D1BWP12T U2527 ( .A1(RF_pc_out[23]), .A2(n5996), .B1(
        register_file_inst1_r10_23_), .B2(n5995), .ZN(n6129) );
  AOI22D1BWP12T U2528 ( .A1(RF_pc_out[15]), .A2(n5996), .B1(
        register_file_inst1_r10_15_), .B2(n5995), .ZN(n6106) );
  AOI22D1BWP12T U2529 ( .A1(RF_pc_out[6]), .A2(n5996), .B1(
        register_file_inst1_r10_6_), .B2(n5995), .ZN(n6077) );
  AOI22D1BWP12T U2530 ( .A1(register_file_inst1_r5_13_), .A2(n6002), .B1(
        register_file_inst1_lr_13_), .B2(n5970), .ZN(n4709) );
  AOI22D1BWP12T U2531 ( .A1(RF_pc_out[13]), .A2(n5996), .B1(
        register_file_inst1_r10_13_), .B2(n5995), .ZN(n6102) );
  AOI22D1BWP12T U2532 ( .A1(RF_pc_out[28]), .A2(n5996), .B1(
        register_file_inst1_r10_28_), .B2(n5995), .ZN(n6139) );
  AOI22D1BWP12T U2533 ( .A1(RF_pc_out[26]), .A2(n5996), .B1(
        register_file_inst1_r10_26_), .B2(n5995), .ZN(n6135) );
  AOI22D1BWP12T U2534 ( .A1(RF_pc_out[19]), .A2(n5996), .B1(
        register_file_inst1_r10_19_), .B2(n5995), .ZN(n6121) );
  AOI22D1BWP12T U2535 ( .A1(RF_pc_out[17]), .A2(n5996), .B1(
        register_file_inst1_r10_17_), .B2(n5995), .ZN(n6117) );
  ND2D1BWP12T U2536 ( .A1(n4217), .A2(n6030), .ZN(n5231) );
  ND2D1BWP12T U2537 ( .A1(n4181), .A2(n6017), .ZN(n5240) );
  ND2D1BWP12T U2538 ( .A1(n4183), .A2(n4185), .ZN(n5256) );
  ND2D1BWP12T U2539 ( .A1(n4187), .A2(n4189), .ZN(n5203) );
  ND2D1BWP12T U2540 ( .A1(n4217), .A2(n6034), .ZN(n5226) );
  ND2D1BWP12T U2541 ( .A1(n4208), .A2(n6018), .ZN(n5249) );
  ND2D1BWP12T U2542 ( .A1(n4217), .A2(n6027), .ZN(n5229) );
  ND2D1BWP12T U2543 ( .A1(n6027), .A2(n6026), .ZN(n5227) );
  ND2D1BWP12T U2544 ( .A1(n4205), .A2(n6031), .ZN(n5246) );
  ND2D1BWP12T U2545 ( .A1(n4212), .A2(n6029), .ZN(n5237) );
  ND2D1BWP12T U2546 ( .A1(n6287), .A2(n6030), .ZN(n5238) );
  ND2D1BWP12T U2547 ( .A1(n4194), .A2(n4195), .ZN(n5252) );
  ND2D1BWP12T U2548 ( .A1(n6024), .A2(n6023), .ZN(n5219) );
  ND2D1BWP12T U2549 ( .A1(n4222), .A2(n6035), .ZN(n5243) );
  ND2D1BWP12T U2550 ( .A1(n6027), .A2(n4221), .ZN(n5223) );
  ND2D1BWP12T U2551 ( .A1(n4198), .A2(n6028), .ZN(n5233) );
  AN3XD1BWP12T U2552 ( .A1(n6386), .A2(IF_RF_incremented_pc_write_enable), 
        .A3(n6391), .Z(n6393) );
  INVD1BWP12T U2553 ( .I(ALU_MISC_OUT_result[31]), .ZN(n5258) );
  INVD1BWP12T U2554 ( .I(ALU_MISC_OUT_result[27]), .ZN(n5177) );
  INVD1BWP12T U2555 ( .I(ALU_MISC_OUT_result[26]), .ZN(n5167) );
  INVD1BWP12T U2556 ( .I(ALU_MISC_OUT_result[25]), .ZN(n5262) );
  INVD2BWP12T U2557 ( .I(ALU_MISC_OUT_result[24]), .ZN(n5260) );
  INVD1BWP12T U2558 ( .I(ALU_MISC_OUT_result[23]), .ZN(n5136) );
  INVD1BWP12T U2559 ( .I(ALU_MISC_OUT_result[21]), .ZN(n5119) );
  INVD1BWP12T U2560 ( .I(ALU_MISC_OUT_result[19]), .ZN(n5114) );
  INVD1BWP12T U2561 ( .I(ALU_MISC_OUT_result[17]), .ZN(n5098) );
  INVD1BWP12T U2562 ( .I(MEMCTRL_RF_IF_data_in[15]), .ZN(n6340) );
  INVD1BWP12T U2563 ( .I(MEMCTRL_RF_IF_data_in[14]), .ZN(n6343) );
  INVD1BWP12T U2564 ( .I(MEMCTRL_RF_IF_data_in[13]), .ZN(n6346) );
  INVD1BWP12T U2565 ( .I(MEMCTRL_RF_IF_data_in[12]), .ZN(n6349) );
  INVD1BWP12T U2566 ( .I(MEMCTRL_RF_IF_data_in[11]), .ZN(n6352) );
  INVD1BWP12T U2567 ( .I(MEMCTRL_RF_IF_data_in[10]), .ZN(n6355) );
  INVD1BWP12T U2568 ( .I(MEMCTRL_RF_IF_data_in[9]), .ZN(n6308) );
  INVD1BWP12T U2569 ( .I(MEMCTRL_RF_IF_data_in[8]), .ZN(n6307) );
  INVD1BWP12T U2570 ( .I(MEMCTRL_RF_IF_data_in[6]), .ZN(n6367) );
  INVD1BWP12T U2571 ( .I(MEMCTRL_RF_IF_data_in[5]), .ZN(n6304) );
  INVD1BWP12T U2572 ( .I(MEMCTRL_RF_IF_data_in[4]), .ZN(n6303) );
  INVD1BWP12T U2573 ( .I(MEMCTRL_RF_IF_data_in[3]), .ZN(n6063) );
  INVD1BWP12T U2574 ( .I(MEMCTRL_RF_IF_data_in[2]), .ZN(n6302) );
  INVD1BWP12T U2575 ( .I(MEMCTRL_RF_IF_data_in[1]), .ZN(n6054) );
  INVD1BWP12T U2576 ( .I(MEMCTRL_RF_IF_data_in[0]), .ZN(n3718) );
  INVD1BWP12T U2577 ( .I(n4672), .ZN(n5009) );
  INVD1BWP12T U2578 ( .I(n4674), .ZN(n5980) );
  NR2D1BWP12T U2579 ( .A1(n2920), .A2(n2912), .ZN(n5004) );
  NR2D1BWP12T U2580 ( .A1(n2912), .A2(n4547), .ZN(n5003) );
  NR2D1BWP12T U2581 ( .A1(n2909), .A2(n4396), .ZN(n5001) );
  NR2D1BWP12T U2582 ( .A1(n2909), .A2(n2917), .ZN(n6005) );
  NR2D1BWP12T U2583 ( .A1(n2909), .A2(n2919), .ZN(n5010) );
  INVD1BWP12T U2584 ( .I(DEC_RF_memory_store_data_reg[4]), .ZN(n3502) );
  INVD1BWP12T U2585 ( .I(reset), .ZN(n6391) );
  INR2D1BWP12T U2586 ( .A1(n4120), .B1(n4670), .ZN(n5985) );
  INVD1BWP12T U2587 ( .I(register_file_inst1_r1_0_), .ZN(n5843) );
  NR2D1BWP12T U2588 ( .A1(n6156), .A2(n6157), .ZN(n5946) );
  AN3XD1BWP12T U2589 ( .A1(DEC_RF_operand_a[1]), .A2(n2471), .A3(n6158), .Z(
        n6229) );
  CKBD1BWP12T U2590 ( .I(n6230), .Z(n5947) );
  INVD1BWP12T U2591 ( .I(n5981), .ZN(n5962) );
  NR2D1BWP12T U2592 ( .A1(n6038), .A2(n6047), .ZN(n5964) );
  NR2D1BWP12T U2593 ( .A1(n4678), .A2(n6046), .ZN(n5968) );
  NR2D1BWP12T U2594 ( .A1(n6046), .A2(n6045), .ZN(n5967) );
  NR2D1BWP12T U2595 ( .A1(n6051), .A2(n6048), .ZN(n6001) );
  NR2D1BWP12T U2596 ( .A1(n6046), .A2(n6049), .ZN(n5969) );
  NR2D1BWP12T U2597 ( .A1(n4676), .A2(n4640), .ZN(n6004) );
  NR2D1BWP12T U2598 ( .A1(n4676), .A2(n6154), .ZN(n6003) );
  NR2D1BWP12T U2599 ( .A1(n4678), .A2(n4677), .ZN(n5994) );
  NR2D1BWP12T U2600 ( .A1(n6044), .A2(n6039), .ZN(n5993) );
  NR2D1BWP12T U2601 ( .A1(n4676), .A2(n6156), .ZN(n5998) );
  NR2D2BWP12T U2602 ( .A1(n6049), .A2(n4677), .ZN(n5995) );
  AN3XD1BWP12T U2603 ( .A1(DEC_RF_operand_a[3]), .A2(n6155), .A3(n2469), .Z(
        n6228) );
  OAI22D1BWP12T U2604 ( .A1(n4618), .A2(n5912), .B1(n5843), .B2(n5857), .ZN(
        n4623) );
  OAI22D1BWP12T U2605 ( .A1(n4621), .A2(n5959), .B1(n4743), .B2(n5805), .ZN(
        n4622) );
  AOI22D1BWP12T U2606 ( .A1(register_file_inst1_r5_3_), .A2(n5948), .B1(
        register_file_inst1_r8_3_), .B2(n5947), .ZN(n5782) );
  AOI22D1BWP12T U2607 ( .A1(RF_pc_out[11]), .A2(n6006), .B1(
        register_file_inst1_r12_11_), .B2(n6228), .ZN(n6182) );
  AOI22D1BWP12T U2608 ( .A1(RF_pc_out[15]), .A2(n6006), .B1(
        register_file_inst1_r12_15_), .B2(n6228), .ZN(n6191) );
  AOI22D1BWP12T U2609 ( .A1(RF_pc_out[7]), .A2(n6006), .B1(
        register_file_inst1_r12_7_), .B2(n6228), .ZN(n6175) );
  AOI22D1BWP12T U2610 ( .A1(RF_pc_out[29]), .A2(n5996), .B1(
        register_file_inst1_r10_29_), .B2(n5995), .ZN(n6141) );
  AOI22D1BWP12T U2611 ( .A1(RF_pc_out[30]), .A2(n5996), .B1(
        register_file_inst1_r10_30_), .B2(n5995), .ZN(n6143) );
  AOI22D1BWP12T U2612 ( .A1(RF_pc_out[31]), .A2(n5996), .B1(
        register_file_inst1_r10_31_), .B2(n5995), .ZN(n6146) );
  AOI22D1BWP12T U2613 ( .A1(RF_pc_out[1]), .A2(n6006), .B1(
        register_file_inst1_r12_1_), .B2(n6228), .ZN(n6162) );
  AOI22D1BWP12T U2614 ( .A1(RF_pc_out[3]), .A2(n6006), .B1(
        register_file_inst1_r12_3_), .B2(n6228), .ZN(n6166) );
  AOI22D1BWP12T U2615 ( .A1(RF_pc_out[4]), .A2(n6006), .B1(
        register_file_inst1_r12_4_), .B2(n6228), .ZN(n6168) );
  ND3D1BWP12T U2616 ( .A1(n5566), .A2(n5565), .A3(n6190), .ZN(n5571) );
  INVD1BWP12T U2617 ( .I(RF_pc_out[0]), .ZN(n6040) );
  IAO21D0BWP12T U2618 ( .A1(MEM_MEMCTRL_from_mem_data[7]), .A2(n4173), .B(
        n4163), .ZN(n4122) );
  ND4D0BWP12T U2619 ( .A1(n6400), .A2(MEM_MEMCTRL_from_mem_data[7]), .A3(
        memory_interface_inst1_delayed_is_signed), .A4(n4119), .ZN(n4164) );
  CKND0BWP12T U2620 ( .I(memory_interface_inst1_delayed_is_signed), .ZN(n4107)
         );
  OAI21D0BWP12T U2621 ( .A1(n5157), .A2(n4107), .B(n4119), .ZN(n4108) );
  IOA21D0BWP12T U2622 ( .A1(MEM_MEMCTRL_from_mem_data[15]), .A2(n4108), .B(
        n4164), .ZN(n4173) );
  MUX2ND0BWP12T U2623 ( .I0(n5259), .I1(n5260), .S(n6008), .ZN(n4109) );
  CKND2D0BWP12T U2624 ( .A1(n5215), .A2(n4109), .ZN(n6323) );
  IOA21D0BWP12T U2625 ( .A1(MEM_MEMCTRL_from_mem_data[14]), .A2(n5985), .B(
        n4160), .ZN(n4749) );
  AN4XD1BWP12T U2626 ( .A1(n5730), .A2(n5731), .A3(n6172), .A4(n5732), .Z(
        n4110) );
  AOI22D0BWP12T U2627 ( .A1(n5836), .A2(register_file_inst1_lr_6_), .B1(n5837), 
        .B2(register_file_inst1_r1_6_), .ZN(n4111) );
  AOI22D1BWP12T U2628 ( .A1(n5835), .A2(RF_next_sp[6]), .B1(n5848), .B2(
        register_file_inst1_r7_6_), .ZN(n4112) );
  AN4XD1BWP12T U2629 ( .A1(n5734), .A2(n6173), .A3(n5733), .A4(n4112), .Z(
        n4113) );
  ND3D1BWP12T U2630 ( .A1(n4110), .A2(n4111), .A3(n4113), .ZN(
        RF_ALU_operand_a[6]) );
  IND2D0BWP12T U2631 ( .A1(n4198), .B1(n6028), .ZN(n5232) );
  IOA21D0BWP12T U2632 ( .A1(MEM_MEMCTRL_from_mem_data[12]), .A2(n5985), .B(
        n4160), .ZN(n4761) );
  IAO21D0BWP12T U2633 ( .A1(MEM_MEMCTRL_from_mem_data[10]), .A2(n4173), .B(
        n4163), .ZN(n4754) );
  IOA21D0BWP12T U2634 ( .A1(MEM_MEMCTRL_from_mem_data[8]), .A2(n5985), .B(
        n4160), .ZN(n4753) );
  AOI21D0BWP12T U2635 ( .A1(n5985), .A2(MEM_MEMCTRL_from_mem_data[3]), .B(
        n4173), .ZN(n5178) );
  AOI21D0BWP12T U2636 ( .A1(n5985), .A2(MEM_MEMCTRL_from_mem_data[2]), .B(
        n4173), .ZN(n5263) );
  AOI21D0BWP12T U2637 ( .A1(n5985), .A2(MEM_MEMCTRL_from_mem_data[1]), .B(
        n4173), .ZN(n5261) );
  AOI21D0BWP12T U2638 ( .A1(n5985), .A2(MEM_MEMCTRL_from_mem_data[0]), .B(
        n4173), .ZN(n5259) );
  IND2D0BWP12T U2639 ( .A1(n4181), .B1(n6017), .ZN(n5239) );
  AO21D0BWP12T U2640 ( .A1(n4164), .A2(n6407), .B(n4163), .Z(n5135) );
  NR4D0BWP12T U2641 ( .A1(n5985), .A2(n6234), .A3(n6400), .A4(
        MEM_MEMCTRL_from_mem_data[15]), .ZN(n4114) );
  OAI21D0BWP12T U2642 ( .A1(memory_interface_inst1_delayed_is_signed), .A2(
        n5157), .B(n4114), .ZN(n2262) );
  INR2D0BWP12T U2643 ( .A1(n4221), .B1(n3510), .ZN(n4193) );
  ND3D1BWP12T U2644 ( .A1(n5553), .A2(n5552), .A3(n6105), .ZN(n5558) );
  IND3D1BWP12T U2645 ( .A1(n4219), .B1(n6391), .B2(n5226), .ZN(n5225) );
  IND2D0BWP12T U2646 ( .A1(n4205), .B1(n6031), .ZN(n5244) );
  AOI21D0BWP12T U2647 ( .A1(n5985), .A2(MEM_MEMCTRL_from_mem_data[13]), .B(
        n4173), .ZN(n5120) );
  IND2D0BWP12T U2648 ( .A1(memory_interface_inst1_fsm_state_1_), .B1(
        memory_interface_inst1_fsm_state_2_), .ZN(n4670) );
  AOI22D1BWP12T U2649 ( .A1(RF_pc_out[2]), .A2(n6006), .B1(
        register_file_inst1_r12_2_), .B2(n6228), .ZN(n6164) );
  INR2D0BWP12T U2650 ( .A1(n4197), .B1(n6403), .ZN(n6297) );
  AOI22D1BWP12T U2651 ( .A1(RF_pc_out[21]), .A2(n5996), .B1(
        register_file_inst1_r10_21_), .B2(n5995), .ZN(n6125) );
  IND3D1BWP12T U2652 ( .A1(n4199), .B1(n6391), .B2(n5231), .ZN(n5096) );
  IND2D0BWP12T U2653 ( .A1(n4208), .B1(n6018), .ZN(n5247) );
  IND3D1BWP12T U2654 ( .A1(n4194), .B1(n6391), .B2(n4195), .ZN(n5250) );
  AOI21D0BWP12T U2655 ( .A1(n5985), .A2(MEM_MEMCTRL_from_mem_data[11]), .B(
        n4173), .ZN(n5115) );
  MAOI22D0BWP12T U2656 ( .A1(n4927), .A2(
        memory_interface_inst1_delay_addr_for_adder_10_), .B1(n4927), .B2(
        memory_interface_inst1_delay_addr_for_adder_10_), .ZN(n4115) );
  AO222D0BWP12T U2657 ( .A1(MEMCTRL_IN_address[10]), .A2(n6295), .B1(n6294), 
        .B2(memory_interface_inst1_delay_addr_single[10]), .C1(n4928), .C2(
        n4115), .Z(MEMCTRL_MEM_to_mem_address[10]) );
  IND2D0BWP12T U2658 ( .A1(n6151), .B1(n2469), .ZN(n5940) );
  AOI22D1BWP12T U2659 ( .A1(RF_pc_out[5]), .A2(n5996), .B1(
        register_file_inst1_r10_5_), .B2(n5995), .ZN(n6073) );
  INR2D0BWP12T U2660 ( .A1(n6026), .B1(n3510), .ZN(n4186) );
  INR2D0BWP12T U2661 ( .A1(n2878), .B1(n6019), .ZN(n4221) );
  IND2D0BWP12T U2662 ( .A1(n4212), .B1(n6029), .ZN(n5235) );
  IND2D0BWP12T U2663 ( .A1(n6023), .B1(n6024), .ZN(n5217) );
  IND2D0BWP12T U2664 ( .A1(n4222), .B1(n6035), .ZN(n5242) );
  AOI21D1BWP12T U2665 ( .A1(ALU_MISC_OUT_result[1]), .A2(n6008), .B(n5982), 
        .ZN(n5021) );
  AOI21D0BWP12T U2666 ( .A1(n5985), .A2(MEM_MEMCTRL_from_mem_data[9]), .B(
        n4173), .ZN(n5099) );
  IND2D0BWP12T U2667 ( .A1(n4838), .B1(n4822), .ZN(n5017) );
  CKND2D0BWP12T U2668 ( .A1(n4927), .A2(
        memory_interface_inst1_delay_addr_for_adder_10_), .ZN(n4116) );
  MOAI22D0BWP12T U2669 ( .A1(memory_interface_inst1_delay_addr_for_adder_11_), 
        .A2(n4116), .B1(memory_interface_inst1_delay_addr_for_adder_11_), .B2(
        n4116), .ZN(n4117) );
  AO222D0BWP12T U2670 ( .A1(MEMCTRL_IN_address[11]), .A2(n6295), .B1(n6294), 
        .B2(memory_interface_inst1_delay_addr_single[11]), .C1(n4117), .C2(
        n4928), .Z(MEMCTRL_MEM_to_mem_address[11]) );
  CKND0BWP12T U2671 ( .I(n6398), .ZN(n4118) );
  MAOI22D0BWP12T U2672 ( .A1(n4841), .A2(n4118), .B1(n6406), .B2(n3018), .ZN(
        MEMCTRL_MEM_to_mem_read_enable) );
  IND2D0BWP12T U2673 ( .A1(n4626), .B1(n6050), .ZN(n5910) );
  ND2D1BWP12T U2674 ( .A1(n4180), .A2(n6310), .ZN(register_file_inst1_n2200)
         );
  TPOAI21D1BWP12T U2675 ( .A1(ALU_MISC_OUT_result[11]), .A2(n5984), .B(n4140), 
        .ZN(n4141) );
  TPNR2D1BWP12T U2676 ( .A1(n4125), .A2(n6301), .ZN(n4128) );
  AOI22D1BWP12T U2677 ( .A1(RF_pc_out[17]), .A2(n6006), .B1(
        register_file_inst1_r12_17_), .B2(n6228), .ZN(n6195) );
  CKND0BWP12T U2678 ( .I(register_file_inst1_r12_6_), .ZN(n5030) );
  AOI22D1BWP12T U2679 ( .A1(RF_pc_out[6]), .A2(n6006), .B1(
        register_file_inst1_r12_6_), .B2(n6228), .ZN(n6172) );
  TPAOI21D8BWP12T U2680 ( .A1(ALU_MISC_OUT_result[24]), .A2(n6008), .B(n4168), 
        .ZN(n4169) );
  AOI22D2BWP12T U2681 ( .A1(register_file_inst1_r4_3_), .A2(n5900), .B1(
        register_file_inst1_r9_3_), .B2(n6225), .ZN(n5785) );
  OR4D2BWP12T U2682 ( .A1(n5666), .A2(n5665), .A3(n5664), .A4(n5663), .Z(
        RF_ALU_operand_b[9]) );
  AOI22D1BWP12T U2683 ( .A1(RF_pc_out[5]), .A2(n6006), .B1(
        register_file_inst1_r12_5_), .B2(n6228), .ZN(n6170) );
  TPAOI21D8BWP12T U2684 ( .A1(n5102), .A2(n6008), .B(n4148), .ZN(n4149) );
  TPAOI21D2BWP12T U2685 ( .A1(n5082), .A2(n6008), .B(n6309), .ZN(n4142) );
  ND4D4BWP12T U2686 ( .A1(n4667), .A2(n4666), .A3(n4665), .A4(n4664), .ZN(
        RF_ALU_operand_a[2]) );
  OAI222D0BWP12T U2687 ( .A1(n5127), .A2(n5235), .B1(n5237), .B2(n5132), .C1(
        n5131), .C2(n5238), .ZN(register_file_inst1_n2351) );
  OAI222D0BWP12T U2688 ( .A1(n5461), .A2(n5094), .B1(n5158), .B2(n5132), .C1(
        n5131), .C2(n5227), .ZN(register_file_inst1_n2415) );
  OAI222D0BWP12T U2689 ( .A1(n5449), .A2(n5096), .B1(n5230), .B2(n5132), .C1(
        n5131), .C2(n5231), .ZN(register_file_inst1_n2639) );
  OAI222D0BWP12T U2690 ( .A1(n5448), .A2(n5095), .B1(n5228), .B2(n5132), .C1(
        n5131), .C2(n5229), .ZN(register_file_inst1_n2447) );
  OAI222D0BWP12T U2691 ( .A1(n5462), .A2(n5222), .B1(n5160), .B2(n5132), .C1(
        n5131), .C2(n5223), .ZN(register_file_inst1_n2223) );
  OAI222D0BWP12T U2692 ( .A1(n5129), .A2(n5225), .B1(n5205), .B2(n5132), .C1(
        n5131), .C2(n5226), .ZN(register_file_inst1_n2511) );
  OAI222D0BWP12T U2693 ( .A1(n5133), .A2(n5250), .B1(n5252), .B2(n5132), .C1(
        n5131), .C2(n5253), .ZN(register_file_inst1_n2319) );
  OAI222D0BWP12T U2694 ( .A1(n5450), .A2(n5254), .B1(n5256), .B2(n5132), .C1(
        n5131), .C2(n5257), .ZN(register_file_inst1_n2575) );
  OAI222D0BWP12T U2695 ( .A1(n4750), .A2(n4758), .B1(n5203), .B2(n5132), .C1(
        n5131), .C2(n5200), .ZN(register_file_inst1_n2543) );
  OAI222D0BWP12T U2696 ( .A1(n5126), .A2(n5247), .B1(n5249), .B2(n5132), .C1(
        n5131), .C2(n5143), .ZN(register_file_inst1_n2479) );
  OAI222D0BWP12T U2697 ( .A1(n5128), .A2(n5242), .B1(n5243), .B2(n5132), .C1(
        n5131), .C2(n5140), .ZN(register_file_inst1_n2255) );
  OAI222D0BWP12T U2698 ( .A1(n5460), .A2(n5232), .B1(n5233), .B2(n5132), .C1(
        n5131), .C2(n5234), .ZN(register_file_inst1_spin[22]) );
  OAI222D0BWP12T U2699 ( .A1(n5463), .A2(n5239), .B1(n5240), .B2(n5132), .C1(
        n5131), .C2(n5074), .ZN(register_file_inst1_n2607) );
  OAI222D0BWP12T U2700 ( .A1(n5125), .A2(n5244), .B1(n5246), .B2(n5132), .C1(
        n5131), .C2(n5145), .ZN(register_file_inst1_n2383) );
  OAI222D0BWP12T U2701 ( .A1(n5130), .A2(n5217), .B1(n5219), .B2(n5132), .C1(
        n5131), .C2(n5220), .ZN(register_file_inst1_n2287) );
  OAI222D0BWP12T U2702 ( .A1(n5124), .A2(n4683), .B1(n5212), .B2(n5132), .C1(
        n5131), .C2(n6144), .ZN(register_file_inst1_n2159) );
  INVD2BWP12T U2703 ( .I(register_file_inst1_r4_0_), .ZN(n4743) );
  OA222D0BWP12T U2704 ( .A1(n5270), .A2(n6313), .B1(n5269), .B2(n5268), .C1(
        n5267), .C2(n5266), .Z(n5272) );
  INVD8BWP12T U2705 ( .I(ALU_MISC_OUT_result[6]), .ZN(n5034) );
  ND4D2BWP12T U2706 ( .A1(n5790), .A2(n5789), .A3(n5788), .A4(n5787), .ZN(
        RF_ALU_operand_a[3]) );
  ND4D4BWP12T U2707 ( .A1(n5829), .A2(n5828), .A3(n5827), .A4(n5826), .ZN(
        RF_ALU_operand_b[1]) );
  TPNR2D3BWP12T U2708 ( .A1(n4132), .A2(n4131), .ZN(n5046) );
  TPNR2D2BWP12T U2709 ( .A1(n4124), .A2(n6300), .ZN(n4139) );
  AOI222D0BWP12T U2710 ( .A1(ALU_MISC_OUT_result[9]), .A2(n6376), .B1(n6395), 
        .B2(n6362), .C1(n6379), .C2(MEMCTRL_RF_IF_data_in[9]), .ZN(n6359) );
  TPND2D3BWP12T U2711 ( .A1(n4145), .A2(n5137), .ZN(n6345) );
  TPNR2D3BWP12T U2712 ( .A1(n6366), .A2(n4136), .ZN(n6362) );
  OR4D2BWP12T U2713 ( .A1(n4729), .A2(n4728), .A3(n4727), .A4(n4726), .Z(
        RF_ALU_operand_b[14]) );
  NR2D1BWP12T U2714 ( .A1(n4547), .A2(n4396), .ZN(n5002) );
  NR2D1BWP12T U2715 ( .A1(n2920), .A2(n2917), .ZN(n5011) );
  NR2D1BWP12T U2716 ( .A1(n2911), .A2(n4396), .ZN(n4989) );
  NR2D1BWP12T U2717 ( .A1(n2912), .A2(n2909), .ZN(n4990) );
  NR2D1BWP12T U2718 ( .A1(n2920), .A2(n4396), .ZN(n4962) );
  NR2D1BWP12T U2719 ( .A1(n2912), .A2(n2911), .ZN(n4991) );
  ND2D1BWP12T U2720 ( .A1(n6287), .A2(n6286), .ZN(n5984) );
  INVD1BWP12T U2721 ( .I(n5984), .ZN(n6008) );
  ND2D1BWP12T U2722 ( .A1(n6008), .A2(n6391), .ZN(n5269) );
  INVD1BWP12T U2723 ( .I(n5269), .ZN(n6376) );
  NR2D1BWP12T U2724 ( .A1(memory_interface_inst1_fsm_state_0_), .A2(
        memory_interface_inst1_fsm_state_3_), .ZN(n4120) );
  INVD1BWP12T U2725 ( .I(n5985), .ZN(n5182) );
  NR3D1BWP12T U2726 ( .A1(memory_interface_inst1_fsm_state_1_), .A2(
        memory_interface_inst1_fsm_state_2_), .A3(
        memory_interface_inst1_fsm_state_3_), .ZN(n6400) );
  INR2D1BWP12T U2727 ( .A1(n6400), .B1(memory_interface_inst1_fsm_state_0_), 
        .ZN(n6282) );
  NR2D1BWP12T U2728 ( .A1(n6234), .A2(n6282), .ZN(n4119) );
  CKND1BWP12T U2729 ( .I(memory_interface_inst1_fsm_state_2_), .ZN(n4765) );
  ND2D1BWP12T U2730 ( .A1(n4765), .A2(memory_interface_inst1_fsm_state_1_), 
        .ZN(n4090) );
  INR2D1BWP12T U2731 ( .A1(n4120), .B1(n4090), .ZN(n6399) );
  INVD1BWP12T U2732 ( .I(n6399), .ZN(n5157) );
  INR2D1BWP12T U2733 ( .A1(n5182), .B1(n4173), .ZN(n4163) );
  INVD1BWP12T U2734 ( .I(n4122), .ZN(n5255) );
  ND2D1BWP12T U2735 ( .A1(n6395), .A2(n5984), .ZN(n5267) );
  TPNR2D0BWP12T U2736 ( .A1(n5255), .A2(n5267), .ZN(n4121) );
  AOI21D0BWP12T U2737 ( .A1(n6376), .A2(ALU_MISC_OUT_result[31]), .B(n4121), 
        .ZN(n4179) );
  OA22XD0BWP12T U2738 ( .A1(ALU_MISC_OUT_result[31]), .A2(n5269), .B1(n4122), 
        .B2(n5267), .Z(n4178) );
  AOI21D1BWP12T U2739 ( .A1(n5985), .A2(MEM_MEMCTRL_from_mem_data[6]), .B(
        n4173), .ZN(n5266) );
  NR2D1BWP12T U2740 ( .A1(ALU_MISC_OUT_result[29]), .A2(n5984), .ZN(n4176) );
  INVD1BWP12T U2741 ( .I(MEM_MEMCTRL_from_mem_data[5]), .ZN(n4099) );
  INVD1BWP12T U2742 ( .I(n4173), .ZN(n4160) );
  OAI21D1BWP12T U2743 ( .A1(n5182), .A2(n4099), .B(n4160), .ZN(n4764) );
  NR2D0BWP12T U2744 ( .A1(n4764), .A2(n6008), .ZN(n4175) );
  NR2D1BWP12T U2745 ( .A1(ALU_MISC_OUT_result[14]), .A2(n5984), .ZN(n4123) );
  NR2D1BWP12T U2746 ( .A1(n4123), .A2(n6299), .ZN(n4145) );
  NR2D1BWP12T U2747 ( .A1(ALU_MISC_OUT_result[9]), .A2(n5984), .ZN(n4138) );
  NR2D1BWP12T U2748 ( .A1(ALU_MISC_OUT_result[5]), .A2(n5984), .ZN(n4132) );
  CKND2D1BWP12T U2749 ( .A1(n6302), .A2(n5984), .ZN(n4126) );
  TPOAI21D1BWP12T U2750 ( .A1(ALU_MISC_OUT_result[2]), .A2(n5984), .B(n4126), 
        .ZN(n4127) );
  NR2XD1BWP12T U2751 ( .A1(n5021), .A2(n4127), .ZN(n6382) );
  TPND2D1BWP12T U2752 ( .A1(n4128), .A2(n6382), .ZN(n6378) );
  CKND2D1BWP12T U2753 ( .A1(n6303), .A2(n5984), .ZN(n4129) );
  OAI21D1BWP12T U2754 ( .A1(ALU_MISC_OUT_result[4]), .A2(n5984), .B(n4129), 
        .ZN(n4130) );
  NR2XD1BWP12T U2755 ( .A1(n6378), .A2(n4130), .ZN(n6374) );
  IOA21D2BWP12T U2756 ( .A1(n5984), .A2(n6304), .B(n6374), .ZN(n4131) );
  AOI21D1BWP12T U2757 ( .A1(n5034), .A2(n6008), .B(n6305), .ZN(n4133) );
  TPND2D2BWP12T U2758 ( .A1(n5046), .A2(n4133), .ZN(n6369) );
  TPNR2D2BWP12T U2759 ( .A1(n6369), .A2(n6306), .ZN(n4134) );
  TPOAI21D1BWP12T U2760 ( .A1(ALU_MISC_OUT_result[7]), .A2(n5984), .B(n4134), 
        .ZN(n6366) );
  ND2D1BWP12T U2761 ( .A1(n6307), .A2(n5984), .ZN(n4135) );
  OAI21D1BWP12T U2762 ( .A1(ALU_MISC_OUT_result[8]), .A2(n5984), .B(n4135), 
        .ZN(n4136) );
  IOA21D2BWP12T U2763 ( .A1(n5984), .A2(n6308), .B(n6362), .ZN(n4137) );
  TPNR2D2BWP12T U2764 ( .A1(n4138), .A2(n4137), .ZN(n5117) );
  TPND2D2BWP12T U2765 ( .A1(n4139), .A2(n5117), .ZN(n6357) );
  CKND2D1BWP12T U2766 ( .A1(n6352), .A2(n5984), .ZN(n4140) );
  TPNR2D2BWP12T U2767 ( .A1(n6357), .A2(n4141), .ZN(n5122) );
  INVD3BWP12T U2768 ( .I(ALU_MISC_OUT_result[12]), .ZN(n5082) );
  TPND2D2BWP12T U2769 ( .A1(n5122), .A2(n4142), .ZN(n6351) );
  ND2D1BWP12T U2770 ( .A1(n6346), .A2(n5984), .ZN(n4143) );
  OAI21D1BWP12T U2771 ( .A1(ALU_MISC_OUT_result[13]), .A2(n5984), .B(n4143), 
        .ZN(n4144) );
  TPNR2D2BWP12T U2772 ( .A1(n6351), .A2(n4144), .ZN(n5137) );
  CKND2D1BWP12T U2773 ( .A1(n6340), .A2(n5984), .ZN(n4146) );
  OAI21D1BWP12T U2774 ( .A1(ALU_MISC_OUT_result[15]), .A2(n5984), .B(n4146), 
        .ZN(n4147) );
  NR2XD3BWP12T U2775 ( .A1(n6345), .A2(n4147), .ZN(n4752) );
  INVD8BWP12T U2776 ( .I(ALU_MISC_OUT_result[16]), .ZN(n5102) );
  NR2D1BWP12T U2777 ( .A1(n4753), .A2(n6008), .ZN(n4148) );
  TPND2D2BWP12T U2779 ( .A1(n4752), .A2(n4149), .ZN(n6339) );
  ND2D1BWP12T U2780 ( .A1(n5099), .A2(n5984), .ZN(n4150) );
  OAI21D1BWP12T U2781 ( .A1(ALU_MISC_OUT_result[17]), .A2(n5984), .B(n4150), 
        .ZN(n4151) );
  TPNR2D2BWP12T U2782 ( .A1(n6339), .A2(n4151), .ZN(n4755) );
  INVD3BWP12T U2783 ( .I(ALU_MISC_OUT_result[18]), .ZN(n4690) );
  NR2D1BWP12T U2784 ( .A1(n4754), .A2(n6008), .ZN(n4152) );
  TPAOI21D2BWP12T U2785 ( .A1(n4690), .A2(n6008), .B(n4152), .ZN(n4153) );
  TPND2D2BWP12T U2786 ( .A1(n4755), .A2(n4153), .ZN(n6335) );
  TPND2D0BWP12T U2787 ( .A1(n5115), .A2(n5984), .ZN(n4154) );
  OAI21D1BWP12T U2788 ( .A1(ALU_MISC_OUT_result[19]), .A2(n5984), .B(n4154), 
        .ZN(n4155) );
  TPNR2D2BWP12T U2789 ( .A1(n6335), .A2(n4155), .ZN(n4760) );
  INVD3BWP12T U2790 ( .I(ALU_MISC_OUT_result[20]), .ZN(n5111) );
  NR2D1BWP12T U2791 ( .A1(n4761), .A2(n6008), .ZN(n4156) );
  TPAOI21D4BWP12T U2792 ( .A1(n5111), .A2(n6008), .B(n4156), .ZN(n4157) );
  TPND2D2BWP12T U2793 ( .A1(n4760), .A2(n4157), .ZN(n6331) );
  ND2D1BWP12T U2794 ( .A1(n5120), .A2(n5984), .ZN(n4158) );
  OAI21D1BWP12T U2795 ( .A1(ALU_MISC_OUT_result[21]), .A2(n5984), .B(n4158), 
        .ZN(n4159) );
  TPNR2D3BWP12T U2796 ( .A1(n6331), .A2(n4159), .ZN(n4730) );
  INVD4BWP12T U2797 ( .I(ALU_MISC_OUT_result[22]), .ZN(n5131) );
  NR2D1BWP12T U2798 ( .A1(n4749), .A2(n6008), .ZN(n4161) );
  TPAOI21D2BWP12T U2799 ( .A1(n5131), .A2(n6008), .B(n4161), .ZN(n4162) );
  TPND2D2BWP12T U2800 ( .A1(n4730), .A2(n4162), .ZN(n6327) );
  INVD1BWP12T U2801 ( .I(MEM_MEMCTRL_from_mem_data[15]), .ZN(n6407) );
  ND2D1BWP12T U2802 ( .A1(n5135), .A2(n5984), .ZN(n4165) );
  TPOAI21D2BWP12T U2803 ( .A1(ALU_MISC_OUT_result[23]), .A2(n5984), .B(n4165), 
        .ZN(n4166) );
  TPNR2D3BWP12T U2804 ( .A1(n6327), .A2(n4166), .ZN(n5215) );
  ND2D1BWP12T U2805 ( .A1(n5261), .A2(n5984), .ZN(n4167) );
  TPOAI21D2BWP12T U2806 ( .A1(ALU_MISC_OUT_result[25]), .A2(n5984), .B(n4167), 
        .ZN(n5216) );
  NR3D1BWP12T U2807 ( .A1(n5259), .A2(n5263), .A3(n6008), .ZN(n4168) );
  NR2XD3BWP12T U2808 ( .A1(n5216), .A2(n4169), .ZN(n4170) );
  OAI211D4BWP12T U2809 ( .A1(n5984), .A2(ALU_MISC_OUT_result[26]), .B(n5215), 
        .C(n4170), .ZN(n6319) );
  TPND2D0BWP12T U2810 ( .A1(n5178), .A2(n5984), .ZN(n4171) );
  OAI21D1BWP12T U2811 ( .A1(ALU_MISC_OUT_result[27]), .A2(n5984), .B(n4171), 
        .ZN(n4172) );
  NR2XD3BWP12T U2812 ( .A1(n6319), .A2(n4172), .ZN(n4763) );
  AOI21D1BWP12T U2813 ( .A1(n5985), .A2(MEM_MEMCTRL_from_mem_data[4]), .B(
        n4173), .ZN(n5190) );
  ND2D1BWP12T U2814 ( .A1(n5190), .A2(n5984), .ZN(n4174) );
  OAI211D4BWP12T U2815 ( .A1(n5984), .A2(ALU_MISC_OUT_result[28]), .B(n4763), 
        .C(n4174), .ZN(n6315) );
  OR3XD4BWP12T U2816 ( .A1(n4176), .A2(n4175), .A3(n6315), .Z(n6313) );
  TPNR2D1BWP12T U2817 ( .A1(ALU_MISC_OUT_result[30]), .A2(n5984), .ZN(n4177)
         );
  RCAOI211D4BWP12T U2818 ( .A1(n5266), .A2(n5984), .B(n6313), .C(n4177), .ZN(
        n5271) );
  MUX2D1BWP12T U2819 ( .I0(n4179), .I1(n4178), .S(n5271), .Z(n4180) );
  ND2D1BWP12T U2820 ( .A1(n6030), .A2(n6026), .ZN(n5074) );
  ND2D1BWP12T U2821 ( .A1(n6014), .A2(n6021), .ZN(n4210) );
  NR2D1BWP12T U2822 ( .A1(n2880), .A2(n6404), .ZN(n4197) );
  ND2D1BWP12T U2823 ( .A1(n4197), .A2(n6403), .ZN(n4207) );
  NR2D1BWP12T U2824 ( .A1(n4210), .A2(n4207), .ZN(n4181) );
  INVD1BWP12T U2825 ( .I(register_file_inst1_r1_24_), .ZN(n5410) );
  OAI222D0BWP12T U2826 ( .A1(n5074), .A2(n5260), .B1(n5240), .B2(n5259), .C1(
        n5239), .C2(n5410), .ZN(register_file_inst1_n2609) );
  NR2D1BWP12T U2827 ( .A1(n3510), .A2(n6012), .ZN(n4182) );
  ND2D1BWP12T U2828 ( .A1(n4182), .A2(n6391), .ZN(n5257) );
  ND2D1BWP12T U2829 ( .A1(n2876), .A2(n6404), .ZN(n4218) );
  NR2D1BWP12T U2830 ( .A1(n6025), .A2(n4218), .ZN(n4183) );
  INVD1BWP12T U2831 ( .I(n4182), .ZN(n4185) );
  INVD0BWP12T U2832 ( .I(n4183), .ZN(n4184) );
  ND3D1BWP12T U2833 ( .A1(n6391), .A2(n4185), .A3(n4184), .ZN(n5254) );
  INVD1BWP12T U2834 ( .I(register_file_inst1_r2_24_), .ZN(n5413) );
  OAI222D0BWP12T U2835 ( .A1(n5257), .A2(n5260), .B1(n5256), .B2(n5259), .C1(
        n5254), .C2(n5413), .ZN(register_file_inst1_n2577) );
  ND2D1BWP12T U2836 ( .A1(n4186), .A2(n6391), .ZN(n5200) );
  NR2D1BWP12T U2837 ( .A1(n6025), .A2(n4207), .ZN(n4187) );
  INVD1BWP12T U2838 ( .I(n4186), .ZN(n4189) );
  INVD0BWP12T U2839 ( .I(n4187), .ZN(n4188) );
  ND3D1BWP12T U2840 ( .A1(n6391), .A2(n4189), .A3(n4188), .ZN(n4758) );
  CKND0BWP12T U2841 ( .I(register_file_inst1_r3_24_), .ZN(n4190) );
  OAI222D0BWP12T U2842 ( .A1(n5200), .A2(n5260), .B1(n5203), .B2(n5259), .C1(
        n4758), .C2(n4190), .ZN(register_file_inst1_n2545) );
  INVD1BWP12T U2843 ( .I(n6296), .ZN(n4202) );
  NR2D1BWP12T U2844 ( .A1(n4202), .A2(n4207), .ZN(n4191) );
  ND3D1BWP12T U2845 ( .A1(n4191), .A2(n6391), .A3(n5227), .ZN(n5158) );
  INVD0BWP12T U2846 ( .I(n4191), .ZN(n4192) );
  ND3D1BWP12T U2847 ( .A1(n6391), .A2(n5227), .A3(n4192), .ZN(n5094) );
  INVD1BWP12T U2848 ( .I(register_file_inst1_r7_24_), .ZN(n5399) );
  OAI222D0BWP12T U2849 ( .A1(n5227), .A2(n5260), .B1(n5158), .B2(n5259), .C1(
        n5094), .C2(n5399), .ZN(register_file_inst1_n2417) );
  ND2D1BWP12T U2850 ( .A1(n4193), .A2(n6391), .ZN(n5253) );
  NR2D1BWP12T U2851 ( .A1(n6025), .A2(n6032), .ZN(n4194) );
  INVD1BWP12T U2852 ( .I(n4193), .ZN(n4195) );
  CKND0BWP12T U2853 ( .I(register_file_inst1_r10_24_), .ZN(n4196) );
  OAI222D0BWP12T U2854 ( .A1(n5253), .A2(n5260), .B1(n5252), .B2(n5259), .C1(
        n5250), .C2(n4196), .ZN(register_file_inst1_n2321) );
  ND2D1BWP12T U2855 ( .A1(n6287), .A2(n6034), .ZN(n5234) );
  INVD1BWP12T U2856 ( .I(n6297), .ZN(n4211) );
  NR2D1BWP12T U2857 ( .A1(n4211), .A2(n6033), .ZN(n4198) );
  INVD1BWP12T U2858 ( .I(RF_next_sp[24]), .ZN(n5398) );
  OAI222D0BWP12T U2859 ( .A1(n5234), .A2(n5260), .B1(n5233), .B2(n5259), .C1(
        n5232), .C2(n5398), .ZN(register_file_inst1_spin[24]) );
  INVD1BWP12T U2860 ( .I(n6012), .ZN(n4217) );
  NR2D1BWP12T U2861 ( .A1(n4218), .A2(n4210), .ZN(n4199) );
  ND3D1BWP12T U2862 ( .A1(n4199), .A2(n6391), .A3(n5231), .ZN(n5230) );
  INVD1BWP12T U2863 ( .I(register_file_inst1_r0_24_), .ZN(n5412) );
  OAI222D0BWP12T U2864 ( .A1(n5231), .A2(n5260), .B1(n5230), .B2(n5259), .C1(
        n5096), .C2(n5412), .ZN(register_file_inst1_n2641) );
  CKND0BWP12T U2865 ( .I(n3510), .ZN(n6022) );
  ND3D1BWP12T U2866 ( .A1(n6287), .A2(n6391), .A3(n6022), .ZN(n5220) );
  INVD0BWP12T U2867 ( .I(register_file_inst1_r11_24_), .ZN(n4668) );
  OAI222D0BWP12T U2868 ( .A1(n5220), .A2(n5260), .B1(n5219), .B2(n5259), .C1(
        n5217), .C2(n4668), .ZN(register_file_inst1_n2289) );
  NR2D1BWP12T U2869 ( .A1(n4202), .A2(n4218), .ZN(n4200) );
  ND3D1BWP12T U2870 ( .A1(n4200), .A2(n6391), .A3(n5229), .ZN(n5228) );
  INVD0BWP12T U2871 ( .I(n4200), .ZN(n4201) );
  ND3D1BWP12T U2872 ( .A1(n6391), .A2(n5229), .A3(n4201), .ZN(n5095) );
  INVD1BWP12T U2873 ( .I(register_file_inst1_r6_24_), .ZN(n5411) );
  OAI222D0BWP12T U2874 ( .A1(n5229), .A2(n5260), .B1(n5228), .B2(n5259), .C1(
        n5095), .C2(n5411), .ZN(register_file_inst1_n2449) );
  NR2D1BWP12T U2875 ( .A1(n4202), .A2(n6032), .ZN(n4203) );
  ND3D1BWP12T U2876 ( .A1(n4203), .A2(n6391), .A3(n5223), .ZN(n5160) );
  INVD0BWP12T U2877 ( .I(n4203), .ZN(n4204) );
  ND3D1BWP12T U2878 ( .A1(n6391), .A2(n5223), .A3(n4204), .ZN(n5222) );
  INVD1BWP12T U2879 ( .I(register_file_inst1_lr_24_), .ZN(n5400) );
  OAI222D0BWP12T U2880 ( .A1(n5223), .A2(n5260), .B1(n5160), .B2(n5259), .C1(
        n5222), .C2(n5400), .ZN(register_file_inst1_n2225) );
  INVD1BWP12T U2881 ( .I(register_file_inst1_r1_23_), .ZN(n5438) );
  OAI222D0BWP12T U2882 ( .A1(n5136), .A2(n5074), .B1(n5240), .B2(n5135), .C1(
        n5239), .C2(n5438), .ZN(register_file_inst1_n2608) );
  ND2D1BWP12T U2883 ( .A1(n6030), .A2(n4221), .ZN(n5145) );
  NR2D1BWP12T U2884 ( .A1(n4210), .A2(n6032), .ZN(n4205) );
  CKND0BWP12T U2885 ( .I(register_file_inst1_r8_23_), .ZN(n4206) );
  OAI222D0BWP12T U2886 ( .A1(n5136), .A2(n5145), .B1(n5246), .B2(n5135), .C1(
        n5244), .C2(n4206), .ZN(register_file_inst1_n2384) );
  INVD1BWP12T U2887 ( .I(register_file_inst1_r2_23_), .ZN(n5425) );
  OAI222D0BWP12T U2888 ( .A1(n5136), .A2(n5257), .B1(n5256), .B2(n5135), .C1(
        n5254), .C2(n5425), .ZN(register_file_inst1_n2576) );
  ND2D1BWP12T U2889 ( .A1(n6034), .A2(n6026), .ZN(n5143) );
  NR2D1BWP12T U2890 ( .A1(n6033), .A2(n4207), .ZN(n4208) );
  CKND0BWP12T U2891 ( .I(register_file_inst1_r5_23_), .ZN(n4209) );
  OAI222D0BWP12T U2892 ( .A1(n5136), .A2(n5143), .B1(n5249), .B2(n5135), .C1(
        n5247), .C2(n4209), .ZN(register_file_inst1_n2480) );
  NR2D1BWP12T U2893 ( .A1(n4211), .A2(n4210), .ZN(n4212) );
  CKND0BWP12T U2894 ( .I(register_file_inst1_r9_23_), .ZN(n4213) );
  OAI222D0BWP12T U2895 ( .A1(n5136), .A2(n5238), .B1(n5237), .B2(n5135), .C1(
        n5235), .C2(n4213), .ZN(register_file_inst1_n2352) );
  CKND0BWP12T U2896 ( .I(register_file_inst1_r10_23_), .ZN(n4214) );
  OAI222D0BWP12T U2897 ( .A1(n5136), .A2(n5253), .B1(n5252), .B2(n5135), .C1(
        n5250), .C2(n4214), .ZN(register_file_inst1_n2320) );
  INVD1BWP12T U2898 ( .I(register_file_inst1_lr_23_), .ZN(n5437) );
  OAI222D0BWP12T U2899 ( .A1(n5136), .A2(n5223), .B1(n5160), .B2(n5135), .C1(
        n5222), .C2(n5437), .ZN(register_file_inst1_n2224) );
  INVD1BWP12T U2900 ( .I(register_file_inst1_r6_23_), .ZN(n5423) );
  OAI222D0BWP12T U2901 ( .A1(n5136), .A2(n5229), .B1(n5228), .B2(n5135), .C1(
        n5095), .C2(n5423), .ZN(register_file_inst1_n2448) );
  INVD1BWP12T U2902 ( .I(RF_next_sp[23]), .ZN(n5435) );
  OAI222D0BWP12T U2903 ( .A1(n5136), .A2(n5234), .B1(n5233), .B2(n5135), .C1(
        n5232), .C2(n5435), .ZN(register_file_inst1_spin[23]) );
  CKND0BWP12T U2904 ( .I(register_file_inst1_r3_23_), .ZN(n4215) );
  OAI222D0BWP12T U2905 ( .A1(n5136), .A2(n5200), .B1(n5203), .B2(n5135), .C1(
        n4758), .C2(n4215), .ZN(register_file_inst1_n2544) );
  CKND0BWP12T U2906 ( .I(register_file_inst1_r11_23_), .ZN(n4216) );
  OAI222D0BWP12T U2907 ( .A1(n5136), .A2(n5220), .B1(n5219), .B2(n5135), .C1(
        n5217), .C2(n4216), .ZN(register_file_inst1_n2288) );
  INVD1BWP12T U2908 ( .I(register_file_inst1_r7_23_), .ZN(n5436) );
  OAI222D0BWP12T U2909 ( .A1(n5136), .A2(n5227), .B1(n5158), .B2(n5135), .C1(
        n5094), .C2(n5436), .ZN(register_file_inst1_n2416) );
  NR2D1BWP12T U2910 ( .A1(n4218), .A2(n6033), .ZN(n4219) );
  ND3D1BWP12T U2911 ( .A1(n4219), .A2(n6391), .A3(n5226), .ZN(n5205) );
  CKND0BWP12T U2912 ( .I(register_file_inst1_r4_23_), .ZN(n4220) );
  OAI222D0BWP12T U2913 ( .A1(n5136), .A2(n5226), .B1(n5205), .B2(n5135), .C1(
        n5225), .C2(n4220), .ZN(register_file_inst1_n2512) );
  ND2D1BWP12T U2914 ( .A1(n6034), .A2(n4221), .ZN(n5140) );
  NR2D1BWP12T U2915 ( .A1(n6033), .A2(n6032), .ZN(n4222) );
  CKND0BWP12T U2916 ( .I(register_file_inst1_r12_23_), .ZN(n4223) );
  OAI222D0BWP12T U2917 ( .A1(n5136), .A2(n5140), .B1(n5243), .B2(n5135), .C1(
        n5242), .C2(n4223), .ZN(register_file_inst1_n2256) );
  INVD1BWP12T U2918 ( .I(register_file_inst1_r0_23_), .ZN(n5424) );
  OAI222D0BWP12T U2919 ( .A1(n5136), .A2(n5231), .B1(n5230), .B2(n5135), .C1(
        n5096), .C2(n5424), .ZN(register_file_inst1_n2640) );
  INVD1BWP12T U2920 ( .I(register_file_inst1_lr_21_), .ZN(n5873) );
  OAI222D0BWP12T U2921 ( .A1(n5873), .A2(n5222), .B1(n5160), .B2(n5120), .C1(
        n5119), .C2(n5223), .ZN(register_file_inst1_n2222) );
  CKND0BWP12T U2922 ( .I(register_file_inst1_r4_21_), .ZN(n4224) );
  OAI222D0BWP12T U2923 ( .A1(n4224), .A2(n5225), .B1(n5205), .B2(n5120), .C1(
        n5119), .C2(n5226), .ZN(register_file_inst1_n2510) );
  CKND0BWP12T U2924 ( .I(register_file_inst1_r9_21_), .ZN(n4225) );
  OAI222D0BWP12T U2925 ( .A1(n4225), .A2(n5235), .B1(n5237), .B2(n5120), .C1(
        n5119), .C2(n5238), .ZN(register_file_inst1_n2350) );
  INVD1BWP12T U2926 ( .I(register_file_inst1_r0_21_), .ZN(n4732) );
  OAI222D0BWP12T U2927 ( .A1(n4732), .A2(n5096), .B1(n5230), .B2(n5120), .C1(
        n5119), .C2(n5231), .ZN(register_file_inst1_n2638) );
  INVD1BWP12T U2928 ( .I(RF_next_sp[21]), .ZN(n5871) );
  OAI222D0BWP12T U2929 ( .A1(n5871), .A2(n5232), .B1(n5233), .B2(n5120), .C1(
        n5119), .C2(n5234), .ZN(register_file_inst1_spin[21]) );
  INVD1BWP12T U2930 ( .I(register_file_inst1_r7_21_), .ZN(n5872) );
  OAI222D0BWP12T U2931 ( .A1(n5872), .A2(n5094), .B1(n5158), .B2(n5120), .C1(
        n5119), .C2(n5227), .ZN(register_file_inst1_n2414) );
  CKND0BWP12T U2932 ( .I(register_file_inst1_r5_21_), .ZN(n4226) );
  OAI222D0BWP12T U2933 ( .A1(n4226), .A2(n5247), .B1(n5249), .B2(n5120), .C1(
        n5119), .C2(n5143), .ZN(register_file_inst1_n2478) );
  CKND0BWP12T U2934 ( .I(register_file_inst1_r12_21_), .ZN(n4227) );
  OAI222D0BWP12T U2935 ( .A1(n4227), .A2(n5242), .B1(n5243), .B2(n5120), .C1(
        n5119), .C2(n5140), .ZN(register_file_inst1_n2254) );
  INVD1BWP12T U2936 ( .I(register_file_inst1_r1_21_), .ZN(n5874) );
  OAI222D0BWP12T U2937 ( .A1(n5874), .A2(n5239), .B1(n5240), .B2(n5120), .C1(
        n5119), .C2(n5074), .ZN(register_file_inst1_n2606) );
  CKND0BWP12T U2938 ( .I(register_file_inst1_r10_21_), .ZN(n4228) );
  OAI222D0BWP12T U2939 ( .A1(n4228), .A2(n5250), .B1(n5252), .B2(n5120), .C1(
        n5119), .C2(n5253), .ZN(register_file_inst1_n2318) );
  INVD1BWP12T U2940 ( .I(register_file_inst1_r6_21_), .ZN(n4731) );
  OAI222D0BWP12T U2941 ( .A1(n4731), .A2(n5095), .B1(n5228), .B2(n5120), .C1(
        n5119), .C2(n5229), .ZN(register_file_inst1_n2446) );
  INVD1BWP12T U2942 ( .I(register_file_inst1_r2_21_), .ZN(n4733) );
  OAI222D0BWP12T U2943 ( .A1(n4733), .A2(n5254), .B1(n5256), .B2(n5120), .C1(
        n5119), .C2(n5257), .ZN(register_file_inst1_n2574) );
  CKND0BWP12T U2944 ( .I(register_file_inst1_r3_21_), .ZN(n4229) );
  OAI222D0BWP12T U2945 ( .A1(n4229), .A2(n4758), .B1(n5203), .B2(n5120), .C1(
        n5119), .C2(n5200), .ZN(register_file_inst1_n2542) );
  CKND0BWP12T U2946 ( .I(register_file_inst1_r8_21_), .ZN(n4230) );
  OAI222D0BWP12T U2947 ( .A1(n4230), .A2(n5244), .B1(n5246), .B2(n5120), .C1(
        n5119), .C2(n5145), .ZN(register_file_inst1_n2382) );
  CKND0BWP12T U2948 ( .I(register_file_inst1_r11_21_), .ZN(n4231) );
  OAI222D0BWP12T U2949 ( .A1(n4231), .A2(n5217), .B1(n5219), .B2(n5120), .C1(
        n5119), .C2(n5220), .ZN(register_file_inst1_n2286) );
  INVD1BWP12T U2950 ( .I(register_file_inst1_r12_19_), .ZN(n4232) );
  OAI222D0BWP12T U2951 ( .A1(n4232), .A2(n5242), .B1(n5243), .B2(n5115), .C1(
        n5114), .C2(n5140), .ZN(register_file_inst1_n2252) );
  INVD1BWP12T U2952 ( .I(register_file_inst1_lr_19_), .ZN(n5475) );
  OAI222D0BWP12T U2953 ( .A1(n5475), .A2(n5222), .B1(n5160), .B2(n5115), .C1(
        n5114), .C2(n5223), .ZN(register_file_inst1_n2220) );
  INVD1BWP12T U2954 ( .I(register_file_inst1_r1_19_), .ZN(n5476) );
  OAI222D0BWP12T U2955 ( .A1(n5476), .A2(n5239), .B1(n5240), .B2(n5115), .C1(
        n5114), .C2(n5074), .ZN(register_file_inst1_n2604) );
  INVD1BWP12T U2956 ( .I(register_file_inst1_r3_19_), .ZN(n4233) );
  OAI222D0BWP12T U2957 ( .A1(n4233), .A2(n4758), .B1(n5203), .B2(n5115), .C1(
        n5114), .C2(n5200), .ZN(register_file_inst1_n2540) );
  INVD1BWP12T U2958 ( .I(register_file_inst1_r9_19_), .ZN(n4234) );
  OAI222D0BWP12T U2959 ( .A1(n4234), .A2(n5235), .B1(n5237), .B2(n5115), .C1(
        n5114), .C2(n5238), .ZN(register_file_inst1_n2348) );
  CKND0BWP12T U2960 ( .I(register_file_inst1_r4_19_), .ZN(n4235) );
  OAI222D0BWP12T U2961 ( .A1(n4235), .A2(n5225), .B1(n5205), .B2(n5115), .C1(
        n5114), .C2(n5226), .ZN(register_file_inst1_n2508) );
  INVD1BWP12T U2962 ( .I(register_file_inst1_r8_19_), .ZN(n4236) );
  OAI222D0BWP12T U2963 ( .A1(n4236), .A2(n5244), .B1(n5246), .B2(n5115), .C1(
        n5114), .C2(n5145), .ZN(register_file_inst1_n2380) );
  INVD1BWP12T U2964 ( .I(RF_next_sp[19]), .ZN(n5473) );
  OAI222D0BWP12T U2965 ( .A1(n5473), .A2(n5232), .B1(n5233), .B2(n5115), .C1(
        n5114), .C2(n5234), .ZN(register_file_inst1_spin[19]) );
  INVD1BWP12T U2966 ( .I(register_file_inst1_r7_19_), .ZN(n5474) );
  OAI222D0BWP12T U2967 ( .A1(n5474), .A2(n5094), .B1(n5158), .B2(n5115), .C1(
        n5114), .C2(n5227), .ZN(register_file_inst1_n2412) );
  CKND0BWP12T U2968 ( .I(register_file_inst1_r5_19_), .ZN(n4237) );
  OAI222D0BWP12T U2969 ( .A1(n4237), .A2(n5247), .B1(n5249), .B2(n5115), .C1(
        n5114), .C2(n5143), .ZN(register_file_inst1_n2476) );
  INVD1BWP12T U2970 ( .I(register_file_inst1_r10_19_), .ZN(n4238) );
  OAI222D0BWP12T U2971 ( .A1(n4238), .A2(n5250), .B1(n5252), .B2(n5115), .C1(
        n5114), .C2(n5253), .ZN(register_file_inst1_n2316) );
  INVD1BWP12T U2972 ( .I(register_file_inst1_r6_19_), .ZN(n4692) );
  OAI222D0BWP12T U2973 ( .A1(n4692), .A2(n5095), .B1(n5228), .B2(n5115), .C1(
        n5114), .C2(n5229), .ZN(register_file_inst1_n2444) );
  INVD1BWP12T U2974 ( .I(register_file_inst1_r0_19_), .ZN(n4693) );
  OAI222D0BWP12T U2980 ( .A1(n4693), .A2(n5096), .B1(n5230), .B2(n5115), .C1(
        n5114), .C2(n5231), .ZN(register_file_inst1_n2636) );
  CKND0BWP12T U2981 ( .I(register_file_inst1_r11_19_), .ZN(n4239) );
  OAI222D0BWP12T U2982 ( .A1(n4239), .A2(n5217), .B1(n5219), .B2(n5115), .C1(
        n5114), .C2(n5220), .ZN(register_file_inst1_n2284) );
  INVD1BWP12T U2983 ( .I(register_file_inst1_r2_19_), .ZN(n4694) );
  OAI222D0BWP12T U2984 ( .A1(n4694), .A2(n5254), .B1(n5256), .B2(n5115), .C1(
        n5114), .C2(n5257), .ZN(register_file_inst1_n2572) );
  INVD1BWP12T U2985 ( .I(ALU_MISC_OUT_result[15]), .ZN(n5088) );
  INVD1BWP12T U2986 ( .I(register_file_inst1_r2_15_), .ZN(n5551) );
  OAI222D0BWP12T U2987 ( .A1(n5088), .A2(n5257), .B1(n5256), .B2(n6340), .C1(
        n5254), .C2(n5551), .ZN(register_file_inst1_n2568) );
  INVD1BWP12T U2988 ( .I(register_file_inst1_r7_17_), .ZN(n5512) );
  OAI222D0BWP12T U2989 ( .A1(n5512), .A2(n5094), .B1(n5158), .B2(n5099), .C1(
        n5098), .C2(n5227), .ZN(register_file_inst1_n2410) );
  INVD1BWP12T U2990 ( .I(register_file_inst1_r10_15_), .ZN(n4240) );
  OAI222D0BWP12T U2991 ( .A1(n5088), .A2(n5253), .B1(n5252), .B2(n6340), .C1(
        n5250), .C2(n4240), .ZN(register_file_inst1_n2312) );
  INVD1BWP12T U2992 ( .I(RF_next_sp[15]), .ZN(n5561) );
  OAI222D0BWP12T U2994 ( .A1(n5088), .A2(n5234), .B1(n5233), .B2(n6340), .C1(
        n5232), .C2(n5561), .ZN(register_file_inst1_spin[15]) );
  INVD1BWP12T U2995 ( .I(register_file_inst1_r2_17_), .ZN(n4649) );
  OAI222D0BWP12T U2996 ( .A1(n4649), .A2(n5254), .B1(n5256), .B2(n5099), .C1(
        n5098), .C2(n5257), .ZN(register_file_inst1_n2570) );
  INVD1BWP12T U2997 ( .I(register_file_inst1_lr_15_), .ZN(n5563) );
  OAI222D0BWP12T U2998 ( .A1(n5088), .A2(n5223), .B1(n5160), .B2(n6340), .C1(
        n5222), .C2(n5563), .ZN(register_file_inst1_n2216) );
  CKND0BWP12T U2999 ( .I(register_file_inst1_r9_17_), .ZN(n4241) );
  OAI222D0BWP12T U3000 ( .A1(n4241), .A2(n5235), .B1(n5237), .B2(n5099), .C1(
        n5098), .C2(n5238), .ZN(register_file_inst1_n2346) );
  INVD1BWP12T U3001 ( .I(RF_next_sp[17]), .ZN(n5511) );
  OAI222D0BWP12T U3002 ( .A1(n5511), .A2(n5232), .B1(n5233), .B2(n5099), .C1(
        n5098), .C2(n5234), .ZN(register_file_inst1_spin[17]) );
  INVD1BWP12T U3011 ( .I(register_file_inst1_r7_15_), .ZN(n5562) );
  OAI222D0BWP12T U3012 ( .A1(n5088), .A2(n5227), .B1(n5158), .B2(n6340), .C1(
        n5094), .C2(n5562), .ZN(register_file_inst1_n2408) );
  INVD1BWP12T U3013 ( .I(register_file_inst1_lr_17_), .ZN(n5513) );
  OAI222D0BWP12T U3014 ( .A1(n5513), .A2(n5222), .B1(n5160), .B2(n5099), .C1(
        n5098), .C2(n5223), .ZN(register_file_inst1_n2218) );
  INVD1BWP12T U3015 ( .I(register_file_inst1_r6_15_), .ZN(n5549) );
  OAI222D0BWP12T U3019 ( .A1(n5088), .A2(n5229), .B1(n5228), .B2(n6340), .C1(
        n5095), .C2(n5549), .ZN(register_file_inst1_n2440) );
  INVD1BWP12T U3020 ( .I(register_file_inst1_r9_15_), .ZN(n4242) );
  OAI222D0BWP12T U3021 ( .A1(n5088), .A2(n5238), .B1(n5237), .B2(n6340), .C1(
        n5235), .C2(n4242), .ZN(register_file_inst1_n2344) );
  CKND0BWP12T U3022 ( .I(register_file_inst1_r5_17_), .ZN(n4243) );
  OAI222D0BWP12T U3023 ( .A1(n4243), .A2(n5247), .B1(n5249), .B2(n5099), .C1(
        n5098), .C2(n5143), .ZN(register_file_inst1_n2474) );
  CKND0BWP12T U3024 ( .I(register_file_inst1_r10_17_), .ZN(n4244) );
  OAI222D0BWP12T U3025 ( .A1(n4244), .A2(n5250), .B1(n5252), .B2(n5099), .C1(
        n5098), .C2(n5253), .ZN(register_file_inst1_n2314) );
  INVD1BWP12T U3026 ( .I(register_file_inst1_r12_15_), .ZN(n4245) );
  OAI222D0BWP12T U3027 ( .A1(n5088), .A2(n5140), .B1(n5243), .B2(n6340), .C1(
        n5242), .C2(n4245), .ZN(register_file_inst1_n2248) );
  INVD1BWP12T U3028 ( .I(register_file_inst1_r12_17_), .ZN(n4246) );
  OAI222D0BWP12T U3029 ( .A1(n4246), .A2(n5242), .B1(n5243), .B2(n5099), .C1(
        n5098), .C2(n5140), .ZN(register_file_inst1_n2250) );
  INVD1BWP12T U3030 ( .I(register_file_inst1_r6_17_), .ZN(n4647) );
  OAI222D0BWP12T U3031 ( .A1(n4647), .A2(n5095), .B1(n5228), .B2(n5099), .C1(
        n5098), .C2(n5229), .ZN(register_file_inst1_n2442) );
  CKND0BWP12T U3032 ( .I(register_file_inst1_r11_15_), .ZN(n4247) );
  OAI222D0BWP12T U3033 ( .A1(n5088), .A2(n5220), .B1(n5219), .B2(n6340), .C1(
        n5217), .C2(n4247), .ZN(register_file_inst1_n2280) );
  CKND0BWP12T U3034 ( .I(register_file_inst1_r11_17_), .ZN(n4248) );
  OAI222D0BWP12T U3035 ( .A1(n4248), .A2(n5217), .B1(n5219), .B2(n5099), .C1(
        n5098), .C2(n5220), .ZN(register_file_inst1_n2282) );
  INVD1BWP12T U3036 ( .I(register_file_inst1_r5_15_), .ZN(n4249) );
  OAI222D0BWP12T U3037 ( .A1(n5088), .A2(n5143), .B1(n5249), .B2(n6340), .C1(
        n5247), .C2(n4249), .ZN(register_file_inst1_n2472) );
  INVD1BWP12T U3038 ( .I(register_file_inst1_r1_15_), .ZN(n5564) );
  OAI222D0BWP12T U3039 ( .A1(n5088), .A2(n5074), .B1(n5240), .B2(n6340), .C1(
        n5239), .C2(n5564), .ZN(register_file_inst1_n2600) );
  CKND0BWP12T U3040 ( .I(register_file_inst1_r8_17_), .ZN(n4250) );
  OAI222D0BWP12T U3041 ( .A1(n4250), .A2(n5244), .B1(n5246), .B2(n5099), .C1(
        n5098), .C2(n5145), .ZN(register_file_inst1_n2378) );
  INVD1BWP12T U3042 ( .I(register_file_inst1_r0_15_), .ZN(n5550) );
  OAI222D0BWP12T U3043 ( .A1(n5088), .A2(n5231), .B1(n5230), .B2(n6340), .C1(
        n5096), .C2(n5550), .ZN(register_file_inst1_n2632) );
  CKND0BWP12T U3044 ( .I(register_file_inst1_r4_17_), .ZN(n4251) );
  OAI222D0BWP12T U3045 ( .A1(n4251), .A2(n5225), .B1(n5205), .B2(n5099), .C1(
        n5098), .C2(n5226), .ZN(register_file_inst1_n2506) );
  CKND0BWP12T U3046 ( .I(register_file_inst1_r4_15_), .ZN(n4252) );
  OAI222D0BWP12T U3047 ( .A1(n5088), .A2(n5226), .B1(n5205), .B2(n6340), .C1(
        n5225), .C2(n4252), .ZN(register_file_inst1_n2504) );
  INVD1BWP12T U3048 ( .I(register_file_inst1_r3_15_), .ZN(n4253) );
  OAI222D0BWP12T U3049 ( .A1(n5088), .A2(n5200), .B1(n5203), .B2(n6340), .C1(
        n4758), .C2(n4253), .ZN(register_file_inst1_n2536) );
  INVD1BWP12T U3050 ( .I(register_file_inst1_r0_17_), .ZN(n4648) );
  OAI222D0BWP12T U3051 ( .A1(n4648), .A2(n5096), .B1(n5230), .B2(n5099), .C1(
        n5098), .C2(n5231), .ZN(register_file_inst1_n2634) );
  INVD1BWP12T U3052 ( .I(register_file_inst1_r1_17_), .ZN(n5514) );
  OAI222D0BWP12T U3053 ( .A1(n5514), .A2(n5239), .B1(n5240), .B2(n5099), .C1(
        n5098), .C2(n5074), .ZN(register_file_inst1_n2602) );
  CKND0BWP12T U3054 ( .I(register_file_inst1_r3_17_), .ZN(n4254) );
  OAI222D0BWP12T U3055 ( .A1(n4254), .A2(n4758), .B1(n5203), .B2(n5099), .C1(
        n5098), .C2(n5200), .ZN(register_file_inst1_n2538) );
  INVD0BWP12T U3056 ( .I(register_file_inst1_r8_15_), .ZN(n4255) );
  OAI222D0BWP12T U3057 ( .A1(n5088), .A2(n5145), .B1(n5246), .B2(n6340), .C1(
        n5244), .C2(n4255), .ZN(register_file_inst1_n2376) );
  INVD1BWP12T U3058 ( .I(ALU_MISC_OUT_result[13]), .ZN(n5084) );
  CKND0BWP12T U3059 ( .I(register_file_inst1_r3_13_), .ZN(n4256) );
  OAI222D0BWP12T U3060 ( .A1(n5084), .A2(n5200), .B1(n5203), .B2(n6346), .C1(
        n4758), .C2(n4256), .ZN(register_file_inst1_n2534) );
  INVD1BWP12T U3061 ( .I(ALU_MISC_OUT_result[11]), .ZN(n4717) );
  INVD1BWP12T U3062 ( .I(register_file_inst1_r5_11_), .ZN(n4257) );
  OAI222D0BWP12T U3063 ( .A1(n4717), .A2(n5143), .B1(n5249), .B2(n6352), .C1(
        n5247), .C2(n4257), .ZN(register_file_inst1_n2468) );
  INVD1BWP12T U3064 ( .I(register_file_inst1_r0_13_), .ZN(n4705) );
  OAI222D0BWP12T U3065 ( .A1(n5084), .A2(n5231), .B1(n5230), .B2(n6346), .C1(
        n5096), .C2(n4705), .ZN(register_file_inst1_n2630) );
  CKND0BWP12T U3066 ( .I(register_file_inst1_r9_11_), .ZN(n4258) );
  OAI222D0BWP12T U3067 ( .A1(n4717), .A2(n5238), .B1(n5237), .B2(n6352), .C1(
        n5235), .C2(n4258), .ZN(register_file_inst1_n2340) );
  INVD1BWP12T U3068 ( .I(register_file_inst1_r0_11_), .ZN(n5633) );
  OAI222D0BWP12T U3069 ( .A1(n4717), .A2(n5231), .B1(n5230), .B2(n6352), .C1(
        n5096), .C2(n5633), .ZN(register_file_inst1_n2628) );
  INVD1BWP12T U3070 ( .I(register_file_inst1_r12_13_), .ZN(n4259) );
  OAI222D0BWP12T U3071 ( .A1(n5084), .A2(n5140), .B1(n5243), .B2(n6346), .C1(
        n5242), .C2(n4259), .ZN(register_file_inst1_n2246) );
  INVD1BWP12T U3072 ( .I(register_file_inst1_r4_11_), .ZN(n4260) );
  OAI222D0BWP12T U3073 ( .A1(n4717), .A2(n5226), .B1(n5205), .B2(n6352), .C1(
        n5225), .C2(n4260), .ZN(register_file_inst1_n2500) );
  CKND0BWP12T U3074 ( .I(register_file_inst1_r9_13_), .ZN(n4261) );
  OAI222D0BWP12T U3075 ( .A1(n5084), .A2(n5238), .B1(n5237), .B2(n6346), .C1(
        n5235), .C2(n4261), .ZN(register_file_inst1_n2342) );
  CKND0BWP12T U3076 ( .I(register_file_inst1_r7_11_), .ZN(n4262) );
  OAI222D0BWP12T U3077 ( .A1(n4717), .A2(n5227), .B1(n5158), .B2(n6352), .C1(
        n5094), .C2(n4262), .ZN(register_file_inst1_n2404) );
  INVD1BWP12T U3078 ( .I(register_file_inst1_r1_13_), .ZN(n5590) );
  OAI222D0BWP12T U3079 ( .A1(n5084), .A2(n5074), .B1(n5240), .B2(n6346), .C1(
        n5239), .C2(n5590), .ZN(register_file_inst1_n2598) );
  INVD1BWP12T U3080 ( .I(register_file_inst1_r12_11_), .ZN(n4263) );
  OAI222D0BWP12T U3081 ( .A1(n4717), .A2(n5140), .B1(n5243), .B2(n6352), .C1(
        n5242), .C2(n4263), .ZN(register_file_inst1_n2244) );
  INVD1BWP12T U3082 ( .I(register_file_inst1_r3_11_), .ZN(n4264) );
  OAI222D0BWP12T U3083 ( .A1(n4717), .A2(n5200), .B1(n5203), .B2(n6352), .C1(
        n4758), .C2(n4264), .ZN(register_file_inst1_n2532) );
  INVD1BWP12T U3084 ( .I(register_file_inst1_r1_11_), .ZN(n5631) );
  OAI222D0BWP12T U3085 ( .A1(n4717), .A2(n5074), .B1(n5240), .B2(n6352), .C1(
        n5239), .C2(n5631), .ZN(register_file_inst1_n2596) );
  CKND0BWP12T U3086 ( .I(register_file_inst1_r4_13_), .ZN(n4265) );
  OAI222D0BWP12T U3087 ( .A1(n5084), .A2(n5226), .B1(n5205), .B2(n6346), .C1(
        n5225), .C2(n4265), .ZN(register_file_inst1_n2502) );
  INVD0BWP12T U3088 ( .I(register_file_inst1_r8_11_), .ZN(n4266) );
  OAI222D0BWP12T U3089 ( .A1(n4717), .A2(n5145), .B1(n5246), .B2(n6352), .C1(
        n5244), .C2(n4266), .ZN(register_file_inst1_n2372) );
  INVD1BWP12T U3090 ( .I(register_file_inst1_r7_13_), .ZN(n5588) );
  OAI222D0BWP12T U3091 ( .A1(n5084), .A2(n5227), .B1(n5158), .B2(n6346), .C1(
        n5094), .C2(n5588), .ZN(register_file_inst1_n2406) );
  CKND0BWP12T U3092 ( .I(register_file_inst1_r5_13_), .ZN(n4267) );
  OAI222D0BWP12T U3093 ( .A1(n5084), .A2(n5143), .B1(n5249), .B2(n6346), .C1(
        n5247), .C2(n4267), .ZN(register_file_inst1_n2470) );
  INVD1BWP12T U3094 ( .I(register_file_inst1_r2_13_), .ZN(n4706) );
  OAI222D0BWP12T U3095 ( .A1(n5084), .A2(n5257), .B1(n5256), .B2(n6346), .C1(
        n5254), .C2(n4706), .ZN(register_file_inst1_n2566) );
  INVD1BWP12T U3096 ( .I(register_file_inst1_r10_11_), .ZN(n4268) );
  OAI222D0BWP12T U3097 ( .A1(n4717), .A2(n5253), .B1(n5252), .B2(n6352), .C1(
        n5250), .C2(n4268), .ZN(register_file_inst1_n2308) );
  CKND0BWP12T U3098 ( .I(register_file_inst1_r11_13_), .ZN(n4269) );
  OAI222D0BWP12T U3099 ( .A1(n5084), .A2(n5220), .B1(n5219), .B2(n6346), .C1(
        n5217), .C2(n4269), .ZN(register_file_inst1_n2278) );
  CKND0BWP12T U3100 ( .I(register_file_inst1_r8_13_), .ZN(n4270) );
  OAI222D0BWP12T U3101 ( .A1(n5084), .A2(n5145), .B1(n5246), .B2(n6346), .C1(
        n5244), .C2(n4270), .ZN(register_file_inst1_n2374) );
  INVD1BWP12T U3102 ( .I(register_file_inst1_r11_11_), .ZN(n4271) );
  OAI222D0BWP12T U3103 ( .A1(n4717), .A2(n5220), .B1(n5219), .B2(n6352), .C1(
        n5217), .C2(n4271), .ZN(register_file_inst1_n2276) );
  INVD1BWP12T U3104 ( .I(register_file_inst1_lr_13_), .ZN(n5589) );
  OAI222D0BWP12T U3105 ( .A1(n5084), .A2(n5223), .B1(n5160), .B2(n6346), .C1(
        n5222), .C2(n5589), .ZN(register_file_inst1_n2214) );
  INVD1BWP12T U3106 ( .I(register_file_inst1_lr_11_), .ZN(n4272) );
  OAI222D0BWP12T U3107 ( .A1(n4717), .A2(n5223), .B1(n5160), .B2(n6352), .C1(
        n5222), .C2(n4272), .ZN(register_file_inst1_n2212) );
  INVD1BWP12T U3108 ( .I(register_file_inst1_r2_11_), .ZN(n5634) );
  OAI222D0BWP12T U3109 ( .A1(n4717), .A2(n5257), .B1(n5256), .B2(n6352), .C1(
        n5254), .C2(n5634), .ZN(register_file_inst1_n2564) );
  CKND0BWP12T U3110 ( .I(register_file_inst1_r10_13_), .ZN(n4273) );
  OAI222D0BWP12T U3111 ( .A1(n5084), .A2(n5253), .B1(n5252), .B2(n6346), .C1(
        n5250), .C2(n4273), .ZN(register_file_inst1_n2310) );
  INVD1BWP12T U3112 ( .I(RF_next_sp[13]), .ZN(n5587) );
  OAI222D0BWP12T U3113 ( .A1(n5084), .A2(n5234), .B1(n5233), .B2(n6346), .C1(
        n5232), .C2(n5587), .ZN(register_file_inst1_spin[13]) );
  ND3D1BWP12T U3114 ( .A1(n6020), .A2(n6391), .A3(n6144), .ZN(n5212) );
  CKND0BWP12T U3115 ( .I(n6020), .ZN(n4274) );
  ND3D1BWP12T U3116 ( .A1(n6391), .A2(n6144), .A3(n4274), .ZN(n4683) );
  CKND0BWP12T U3117 ( .I(register_file_inst1_tmp1_11_), .ZN(n4275) );
  OAI222D0BWP12T U3118 ( .A1(n4717), .A2(n6144), .B1(n5212), .B2(n6352), .C1(
        n4683), .C2(n4275), .ZN(register_file_inst1_n2148) );
  INVD1BWP12T U3119 ( .I(register_file_inst1_r6_11_), .ZN(n5632) );
  OAI222D0BWP12T U3120 ( .A1(n4717), .A2(n5229), .B1(n5228), .B2(n6352), .C1(
        n5095), .C2(n5632), .ZN(register_file_inst1_n2436) );
  INVD1BWP12T U3121 ( .I(register_file_inst1_r6_13_), .ZN(n4704) );
  OAI222D0BWP12T U3122 ( .A1(n5084), .A2(n5229), .B1(n5228), .B2(n6346), .C1(
        n5095), .C2(n4704), .ZN(register_file_inst1_n2438) );
  TPOAI21D0BWP12T U3123 ( .A1(n4717), .A2(n5234), .B(n6093), .ZN(
        register_file_inst1_spin[11]) );
  INVD1BWP12T U3124 ( .I(ALU_MISC_OUT_result[9]), .ZN(n4307) );
  INVD1BWP12T U3125 ( .I(register_file_inst1_lr_9_), .ZN(n5654) );
  OAI222D0BWP12T U3126 ( .A1(n5160), .A2(n6308), .B1(n5223), .B2(n4307), .C1(
        n5222), .C2(n5654), .ZN(register_file_inst1_n2210) );
  INVD1BWP12T U3127 ( .I(ALU_MISC_OUT_result[14]), .ZN(n5086) );
  INVD1BWP12T U3128 ( .I(register_file_inst1_r6_14_), .ZN(n4718) );
  OAI222D0BWP12T U3129 ( .A1(n5086), .A2(n5229), .B1(n5228), .B2(n6343), .C1(
        n5095), .C2(n4718), .ZN(register_file_inst1_n2439) );
  CKND0BWP12T U3130 ( .I(register_file_inst1_r5_14_), .ZN(n4276) );
  OAI222D0BWP12T U3131 ( .A1(n5086), .A2(n5143), .B1(n5249), .B2(n6343), .C1(
        n5247), .C2(n4276), .ZN(register_file_inst1_n2471) );
  CKND0BWP12T U3132 ( .I(register_file_inst1_r9_14_), .ZN(n4277) );
  OAI222D0BWP12T U3133 ( .A1(n5086), .A2(n5238), .B1(n5237), .B2(n6343), .C1(
        n5235), .C2(n4277), .ZN(register_file_inst1_n2343) );
  INVD1BWP12T U3134 ( .I(register_file_inst1_lr_14_), .ZN(n5576) );
  OAI222D0BWP12T U3135 ( .A1(n5086), .A2(n5223), .B1(n5160), .B2(n6343), .C1(
        n5222), .C2(n5576), .ZN(register_file_inst1_n2215) );
  INVD1BWP12T U3136 ( .I(ALU_MISC_OUT_result[10]), .ZN(n4304) );
  CKND0BWP12T U3137 ( .I(register_file_inst1_lr_10_), .ZN(n4278) );
  OAI222D0BWP12T U3138 ( .A1(n4304), .A2(n5223), .B1(n5160), .B2(n6355), .C1(
        n5222), .C2(n4278), .ZN(register_file_inst1_n2211) );
  CKND0BWP12T U3139 ( .I(register_file_inst1_r10_10_), .ZN(n4279) );
  OAI222D0BWP12T U3140 ( .A1(n4304), .A2(n5253), .B1(n5252), .B2(n6355), .C1(
        n5250), .C2(n4279), .ZN(register_file_inst1_n2307) );
  INVD1BWP12T U3141 ( .I(RF_next_sp[14]), .ZN(n5574) );
  OAI222D0BWP12T U3142 ( .A1(n5086), .A2(n5234), .B1(n5233), .B2(n6343), .C1(
        n5232), .C2(n5574), .ZN(register_file_inst1_spin[14]) );
  INVD1BWP12T U3143 ( .I(register_file_inst1_r0_9_), .ZN(n5656) );
  OAI222D0BWP12T U3144 ( .A1(n5230), .A2(n6308), .B1(n5231), .B2(n4307), .C1(
        n5096), .C2(n5656), .ZN(register_file_inst1_n2626) );
  CKND0BWP12T U3145 ( .I(register_file_inst1_tmp1_10_), .ZN(n4280) );
  OAI222D0BWP12T U3146 ( .A1(n4304), .A2(n6144), .B1(n5212), .B2(n6355), .C1(
        n4683), .C2(n4280), .ZN(register_file_inst1_n2147) );
  INVD0BWP12T U3147 ( .I(register_file_inst1_r7_9_), .ZN(n4281) );
  OAI222D0BWP12T U3148 ( .A1(n5158), .A2(n6308), .B1(n5227), .B2(n4307), .C1(
        n5094), .C2(n4281), .ZN(register_file_inst1_n2402) );
  CKND0BWP12T U3149 ( .I(register_file_inst1_r6_9_), .ZN(n4282) );
  OAI222D0BWP12T U3150 ( .A1(n5228), .A2(n6308), .B1(n5229), .B2(n4307), .C1(
        n5095), .C2(n4282), .ZN(register_file_inst1_n2434) );
  INVD1BWP12T U3151 ( .I(register_file_inst1_r0_10_), .ZN(n5860) );
  OAI222D0BWP12T U3152 ( .A1(n4304), .A2(n5231), .B1(n5230), .B2(n6355), .C1(
        n5096), .C2(n5860), .ZN(register_file_inst1_n2627) );
  INVD1BWP12T U3153 ( .I(register_file_inst1_r6_10_), .ZN(n5859) );
  OAI222D0BWP12T U3154 ( .A1(n4304), .A2(n5229), .B1(n5228), .B2(n6355), .C1(
        n5095), .C2(n5859), .ZN(register_file_inst1_n2435) );
  INVD1BWP12T U3155 ( .I(register_file_inst1_r12_14_), .ZN(n4283) );
  OAI222D0BWP12T U3156 ( .A1(n5086), .A2(n5140), .B1(n5243), .B2(n6343), .C1(
        n5242), .C2(n4283), .ZN(register_file_inst1_n2247) );
  CKND0BWP12T U3157 ( .I(register_file_inst1_tmp1_9_), .ZN(n4284) );
  OAI222D0BWP12T U3158 ( .A1(n5212), .A2(n6308), .B1(n6144), .B2(n4307), .C1(
        n4683), .C2(n4284), .ZN(register_file_inst1_n2146) );
  INVD1BWP12T U3159 ( .I(register_file_inst1_r10_9_), .ZN(n4285) );
  OAI222D0BWP12T U3160 ( .A1(n5252), .A2(n6308), .B1(n5253), .B2(n4307), .C1(
        n5250), .C2(n4285), .ZN(register_file_inst1_n2306) );
  INVD1BWP12T U3161 ( .I(register_file_inst1_r2_9_), .ZN(n5657) );
  OAI222D0BWP12T U3162 ( .A1(n5256), .A2(n6308), .B1(n5257), .B2(n4307), .C1(
        n5254), .C2(n5657), .ZN(register_file_inst1_n2562) );
  INVD1BWP12T U3163 ( .I(register_file_inst1_r5_9_), .ZN(n4286) );
  OAI222D0BWP12T U3164 ( .A1(n5249), .A2(n6308), .B1(n5143), .B2(n4307), .C1(
        n5247), .C2(n4286), .ZN(register_file_inst1_n2466) );
  INVD1BWP12T U3165 ( .I(register_file_inst1_r10_14_), .ZN(n4287) );
  OAI222D0BWP12T U3166 ( .A1(n5086), .A2(n5253), .B1(n5252), .B2(n6343), .C1(
        n5250), .C2(n4287), .ZN(register_file_inst1_n2311) );
  INVD1BWP12T U3167 ( .I(register_file_inst1_r1_9_), .ZN(n5655) );
  OAI222D0BWP12T U3168 ( .A1(n5240), .A2(n6308), .B1(n5074), .B2(n4307), .C1(
        n5239), .C2(n5655), .ZN(register_file_inst1_n2594) );
  INVD1BWP12T U3169 ( .I(register_file_inst1_r2_10_), .ZN(n5861) );
  OAI222D0BWP12T U3170 ( .A1(n4304), .A2(n5257), .B1(n5256), .B2(n6355), .C1(
        n5254), .C2(n5861), .ZN(register_file_inst1_n2563) );
  CKND0BWP12T U3171 ( .I(register_file_inst1_r3_14_), .ZN(n4288) );
  OAI222D0BWP12T U3172 ( .A1(n5086), .A2(n5200), .B1(n5203), .B2(n6343), .C1(
        n4758), .C2(n4288), .ZN(register_file_inst1_n2535) );
  INVD1BWP12T U3173 ( .I(register_file_inst1_r3_9_), .ZN(n4289) );
  OAI222D0BWP12T U3174 ( .A1(n5203), .A2(n6308), .B1(n5200), .B2(n4307), .C1(
        n4758), .C2(n4289), .ZN(register_file_inst1_n2530) );
  INVD1BWP12T U3175 ( .I(register_file_inst1_r1_10_), .ZN(n5858) );
  OAI222D0BWP12T U3176 ( .A1(n4304), .A2(n5074), .B1(n5240), .B2(n6355), .C1(
        n5239), .C2(n5858), .ZN(register_file_inst1_n2595) );
  CKND0BWP12T U3177 ( .I(register_file_inst1_r5_10_), .ZN(n4290) );
  OAI222D0BWP12T U3178 ( .A1(n4304), .A2(n5143), .B1(n5249), .B2(n6355), .C1(
        n5247), .C2(n4290), .ZN(register_file_inst1_n2467) );
  CKND0BWP12T U3179 ( .I(register_file_inst1_r4_14_), .ZN(n4291) );
  OAI222D0BWP12T U3180 ( .A1(n5086), .A2(n5226), .B1(n5205), .B2(n6343), .C1(
        n5225), .C2(n4291), .ZN(register_file_inst1_n2503) );
  CKND0BWP12T U3181 ( .I(register_file_inst1_r9_10_), .ZN(n4292) );
  OAI222D0BWP12T U3182 ( .A1(n4304), .A2(n5238), .B1(n5237), .B2(n6355), .C1(
        n5235), .C2(n4292), .ZN(register_file_inst1_n2339) );
  INVD1BWP12T U3183 ( .I(register_file_inst1_r2_14_), .ZN(n4720) );
  OAI222D0BWP12T U3184 ( .A1(n5086), .A2(n5257), .B1(n5256), .B2(n6343), .C1(
        n5254), .C2(n4720), .ZN(register_file_inst1_n2567) );
  CKND0BWP12T U3185 ( .I(register_file_inst1_r12_10_), .ZN(n4293) );
  OAI222D0BWP12T U3186 ( .A1(n4304), .A2(n5140), .B1(n5243), .B2(n6355), .C1(
        n5242), .C2(n4293), .ZN(register_file_inst1_n2243) );
  INVD1BWP12T U3187 ( .I(register_file_inst1_r11_9_), .ZN(n4294) );
  OAI222D0BWP12T U3188 ( .A1(n5219), .A2(n6308), .B1(n5220), .B2(n4307), .C1(
        n5217), .C2(n4294), .ZN(register_file_inst1_n2274) );
  CKND0BWP12T U3189 ( .I(register_file_inst1_r8_9_), .ZN(n4295) );
  OAI222D0BWP12T U3190 ( .A1(n5246), .A2(n6308), .B1(n5145), .B2(n4307), .C1(
        n5244), .C2(n4295), .ZN(register_file_inst1_n2370) );
  CKND0BWP12T U3191 ( .I(register_file_inst1_r8_14_), .ZN(n4296) );
  OAI222D0BWP12T U3192 ( .A1(n5086), .A2(n5145), .B1(n5246), .B2(n6343), .C1(
        n5244), .C2(n4296), .ZN(register_file_inst1_n2375) );
  CKND0BWP12T U3193 ( .I(register_file_inst1_r8_10_), .ZN(n4297) );
  OAI222D0BWP12T U3194 ( .A1(n4304), .A2(n5145), .B1(n5246), .B2(n6355), .C1(
        n5244), .C2(n4297), .ZN(register_file_inst1_n2371) );
  INVD1BWP12T U3195 ( .I(register_file_inst1_r1_14_), .ZN(n5577) );
  OAI222D0BWP12T U3196 ( .A1(n5086), .A2(n5074), .B1(n5240), .B2(n6343), .C1(
        n5239), .C2(n5577), .ZN(register_file_inst1_n2599) );
  CKND0BWP12T U3197 ( .I(register_file_inst1_r11_10_), .ZN(n4298) );
  OAI222D0BWP12T U3198 ( .A1(n4304), .A2(n5220), .B1(n5219), .B2(n6355), .C1(
        n5217), .C2(n4298), .ZN(register_file_inst1_n2275) );
  INVD1BWP12T U3199 ( .I(register_file_inst1_r7_14_), .ZN(n5575) );
  OAI222D0BWP12T U3200 ( .A1(n5086), .A2(n5227), .B1(n5158), .B2(n6343), .C1(
        n5094), .C2(n5575), .ZN(register_file_inst1_n2407) );
  INVD1BWP12T U3201 ( .I(register_file_inst1_r12_9_), .ZN(n4299) );
  OAI222D0BWP12T U3202 ( .A1(n5243), .A2(n6308), .B1(n5140), .B2(n4307), .C1(
        n5242), .C2(n4299), .ZN(register_file_inst1_n2242) );
  INVD1BWP12T U3203 ( .I(register_file_inst1_r0_14_), .ZN(n4719) );
  OAI222D0BWP12T U3204 ( .A1(n5086), .A2(n5231), .B1(n5230), .B2(n6343), .C1(
        n5096), .C2(n4719), .ZN(register_file_inst1_n2631) );
  INVD1BWP12T U3205 ( .I(register_file_inst1_r9_9_), .ZN(n4300) );
  OAI222D0BWP12T U3206 ( .A1(n5237), .A2(n6308), .B1(n5238), .B2(n4307), .C1(
        n5235), .C2(n4300), .ZN(register_file_inst1_n2338) );
  CKND0BWP12T U3207 ( .I(register_file_inst1_r7_10_), .ZN(n4301) );
  OAI222D0BWP12T U3208 ( .A1(n4304), .A2(n5227), .B1(n5158), .B2(n6355), .C1(
        n5094), .C2(n4301), .ZN(register_file_inst1_n2403) );
  CKND0BWP12T U3209 ( .I(register_file_inst1_r4_10_), .ZN(n4302) );
  OAI222D0BWP12T U3210 ( .A1(n4304), .A2(n5226), .B1(n5205), .B2(n6355), .C1(
        n5225), .C2(n4302), .ZN(register_file_inst1_n2499) );
  CKND0BWP12T U3211 ( .I(register_file_inst1_r3_10_), .ZN(n4303) );
  OAI222D0BWP12T U3212 ( .A1(n4304), .A2(n5200), .B1(n5203), .B2(n6355), .C1(
        n4758), .C2(n4303), .ZN(register_file_inst1_n2531) );
  INVD1BWP12T U3213 ( .I(register_file_inst1_r11_14_), .ZN(n4305) );
  OAI222D0BWP12T U3214 ( .A1(n5086), .A2(n5220), .B1(n5219), .B2(n6343), .C1(
        n5217), .C2(n4305), .ZN(register_file_inst1_n2279) );
  CKND0BWP12T U3215 ( .I(register_file_inst1_r4_9_), .ZN(n4306) );
  OAI222D0BWP12T U3216 ( .A1(n5205), .A2(n6308), .B1(n5226), .B2(n4307), .C1(
        n5225), .C2(n4306), .ZN(register_file_inst1_n2498) );
  INVD1BWP12T U3217 ( .I(ALU_MISC_OUT_result[7]), .ZN(n4691) );
  INVD1BWP12T U3218 ( .I(register_file_inst1_r8_7_), .ZN(n4308) );
  OAI222D0BWP12T U3219 ( .A1(n5246), .A2(n6364), .B1(n5145), .B2(n4691), .C1(
        n5244), .C2(n4308), .ZN(register_file_inst1_n2368) );
  INVD1BWP12T U3220 ( .I(register_file_inst1_r11_7_), .ZN(n4309) );
  OAI222D0BWP12T U3221 ( .A1(n5219), .A2(n6364), .B1(n5220), .B2(n4691), .C1(
        n5217), .C2(n4309), .ZN(register_file_inst1_n2272) );
  INVD1BWP12T U3222 ( .I(register_file_inst1_r6_7_), .ZN(n5705) );
  OAI222D0BWP12T U3223 ( .A1(n5228), .A2(n6364), .B1(n5229), .B2(n4691), .C1(
        n5095), .C2(n5705), .ZN(register_file_inst1_n2432) );
  TPOAI21D0BWP12T U3224 ( .A1(n4691), .A2(n5234), .B(n6079), .ZN(
        register_file_inst1_spin[7]) );
  INVD1BWP12T U3225 ( .I(register_file_inst1_r1_7_), .ZN(n5704) );
  OAI222D0BWP12T U3226 ( .A1(n5240), .A2(n6364), .B1(n5074), .B2(n4691), .C1(
        n5239), .C2(n5704), .ZN(register_file_inst1_n2592) );
  INVD1BWP12T U3227 ( .I(register_file_inst1_r0_7_), .ZN(n5706) );
  OAI222D0BWP12T U3228 ( .A1(n5230), .A2(n6364), .B1(n5231), .B2(n4691), .C1(
        n5096), .C2(n5706), .ZN(register_file_inst1_n2624) );
  INVD1BWP12T U3229 ( .I(register_file_inst1_r3_7_), .ZN(n4310) );
  OAI222D0BWP12T U3230 ( .A1(n5203), .A2(n6364), .B1(n5200), .B2(n4691), .C1(
        n4758), .C2(n4310), .ZN(register_file_inst1_n2528) );
  CKND0BWP12T U3231 ( .I(register_file_inst1_r4_7_), .ZN(n4311) );
  OAI222D0BWP12T U3232 ( .A1(n5205), .A2(n6364), .B1(n5226), .B2(n4691), .C1(
        n5225), .C2(n4311), .ZN(register_file_inst1_n2496) );
  INVD1BWP12T U3233 ( .I(register_file_inst1_r12_7_), .ZN(n4312) );
  OAI222D0BWP12T U3234 ( .A1(n5243), .A2(n6364), .B1(n5140), .B2(n4691), .C1(
        n5242), .C2(n4312), .ZN(register_file_inst1_n2240) );
  INVD1BWP12T U3235 ( .I(register_file_inst1_r10_7_), .ZN(n4313) );
  OAI222D0BWP12T U3236 ( .A1(n5252), .A2(n6364), .B1(n5253), .B2(n4691), .C1(
        n5250), .C2(n4313), .ZN(register_file_inst1_n2304) );
  INVD1BWP12T U3237 ( .I(register_file_inst1_r2_7_), .ZN(n5707) );
  OAI222D0BWP12T U3238 ( .A1(n5256), .A2(n6364), .B1(n5257), .B2(n4691), .C1(
        n5254), .C2(n5707), .ZN(register_file_inst1_n2560) );
  INVD1BWP12T U3239 ( .I(register_file_inst1_r9_7_), .ZN(n4314) );
  OAI222D0BWP12T U3240 ( .A1(n5237), .A2(n6364), .B1(n5238), .B2(n4691), .C1(
        n5235), .C2(n4314), .ZN(register_file_inst1_n2336) );
  CKND0BWP12T U3241 ( .I(register_file_inst1_tmp1_7_), .ZN(n4315) );
  OAI222D0BWP12T U3242 ( .A1(n5212), .A2(n6364), .B1(n6144), .B2(n4691), .C1(
        n4683), .C2(n4315), .ZN(register_file_inst1_n2144) );
  INVD1BWP12T U3243 ( .I(register_file_inst1_r7_7_), .ZN(n5693) );
  OAI222D0BWP12T U3244 ( .A1(n5158), .A2(n6364), .B1(n5227), .B2(n4691), .C1(
        n5094), .C2(n5693), .ZN(register_file_inst1_n2400) );
  INVD1BWP12T U3245 ( .I(register_file_inst1_lr_7_), .ZN(n5694) );
  OAI222D0BWP12T U3246 ( .A1(n5160), .A2(n6364), .B1(n5223), .B2(n4691), .C1(
        n5222), .C2(n5694), .ZN(register_file_inst1_n2208) );
  INVD1BWP12T U3247 ( .I(register_file_inst1_r5_7_), .ZN(n4316) );
  OAI222D0BWP12T U3248 ( .A1(n5249), .A2(n6364), .B1(n5143), .B2(n4691), .C1(
        n5247), .C2(n4316), .ZN(register_file_inst1_n2464) );
  INVD1BWP12T U3249 ( .I(ALU_MISC_OUT_result[8]), .ZN(n4716) );
  CKND0BWP12T U3250 ( .I(register_file_inst1_r11_8_), .ZN(n4317) );
  OAI222D0BWP12T U3251 ( .A1(n4716), .A2(n5220), .B1(n5219), .B2(n6307), .C1(
        n5217), .C2(n4317), .ZN(register_file_inst1_n2273) );
  INVD1BWP12T U3252 ( .I(register_file_inst1_r1_8_), .ZN(n5682) );
  OAI222D0BWP12T U3253 ( .A1(n4716), .A2(n5074), .B1(n5240), .B2(n6307), .C1(
        n5239), .C2(n5682), .ZN(register_file_inst1_n2593) );
  CKND0BWP12T U3254 ( .I(register_file_inst1_tmp1_8_), .ZN(n4318) );
  OAI222D0BWP12T U3255 ( .A1(n4716), .A2(n6144), .B1(n5212), .B2(n6307), .C1(
        n4683), .C2(n4318), .ZN(register_file_inst1_n2145) );
  CKND0BWP12T U3256 ( .I(register_file_inst1_r9_8_), .ZN(n4319) );
  OAI222D0BWP12T U3257 ( .A1(n4716), .A2(n5238), .B1(n5237), .B2(n6307), .C1(
        n5235), .C2(n4319), .ZN(register_file_inst1_n2337) );
  INVD1BWP12T U3258 ( .I(register_file_inst1_lr_8_), .ZN(n5681) );
  OAI222D0BWP12T U3259 ( .A1(n4716), .A2(n5223), .B1(n5160), .B2(n6307), .C1(
        n5222), .C2(n5681), .ZN(register_file_inst1_n2209) );
  CKND0BWP12T U3260 ( .I(register_file_inst1_r12_8_), .ZN(n4320) );
  OAI222D0BWP12T U3261 ( .A1(n4716), .A2(n5140), .B1(n5243), .B2(n6307), .C1(
        n5242), .C2(n4320), .ZN(register_file_inst1_n2241) );
  INVD1BWP12T U3262 ( .I(register_file_inst1_r6_8_), .ZN(n5667) );
  OAI222D0BWP12T U3263 ( .A1(n4716), .A2(n5229), .B1(n5228), .B2(n6307), .C1(
        n5095), .C2(n5667), .ZN(register_file_inst1_n2433) );
  INVD0BWP12T U3264 ( .I(register_file_inst1_r8_8_), .ZN(n4321) );
  OAI222D0BWP12T U3265 ( .A1(n4716), .A2(n5145), .B1(n5246), .B2(n6307), .C1(
        n5244), .C2(n4321), .ZN(register_file_inst1_n2369) );
  INVD1BWP12T U3266 ( .I(register_file_inst1_r0_8_), .ZN(n5668) );
  OAI222D0BWP12T U3267 ( .A1(n4716), .A2(n5231), .B1(n5230), .B2(n6307), .C1(
        n5096), .C2(n5668), .ZN(register_file_inst1_n2625) );
  CKND0BWP12T U3268 ( .I(register_file_inst1_r4_8_), .ZN(n4322) );
  OAI222D0BWP12T U3269 ( .A1(n4716), .A2(n5226), .B1(n5205), .B2(n6307), .C1(
        n5225), .C2(n4322), .ZN(register_file_inst1_n2497) );
  CKND0BWP12T U3270 ( .I(register_file_inst1_r10_8_), .ZN(n4323) );
  OAI222D0BWP12T U3271 ( .A1(n4716), .A2(n5253), .B1(n5252), .B2(n6307), .C1(
        n5250), .C2(n4323), .ZN(register_file_inst1_n2305) );
  CKND0BWP12T U3272 ( .I(register_file_inst1_r3_8_), .ZN(n4324) );
  OAI222D0BWP12T U3273 ( .A1(n4716), .A2(n5200), .B1(n5203), .B2(n6307), .C1(
        n4758), .C2(n4324), .ZN(register_file_inst1_n2529) );
  TPOAI21D0BWP12T U3274 ( .A1(n4716), .A2(n5234), .B(n6083), .ZN(
        register_file_inst1_spin[8]) );
  INVD1BWP12T U3275 ( .I(register_file_inst1_r7_8_), .ZN(n5680) );
  OAI222D0BWP12T U3276 ( .A1(n4716), .A2(n5227), .B1(n5158), .B2(n6307), .C1(
        n5094), .C2(n5680), .ZN(register_file_inst1_n2401) );
  CKND0BWP12T U3277 ( .I(register_file_inst1_r5_8_), .ZN(n4325) );
  OAI222D0BWP12T U3278 ( .A1(n4716), .A2(n5143), .B1(n5249), .B2(n6307), .C1(
        n5247), .C2(n4325), .ZN(register_file_inst1_n2465) );
  INVD1BWP12T U3279 ( .I(register_file_inst1_r2_8_), .ZN(n5669) );
  OAI222D0BWP12T U3280 ( .A1(n4716), .A2(n5257), .B1(n5256), .B2(n6307), .C1(
        n5254), .C2(n5669), .ZN(register_file_inst1_n2561) );
  INVD1BWP12T U3281 ( .I(ALU_MISC_OUT_result[4]), .ZN(n5023) );
  CKND0BWP12T U3282 ( .I(register_file_inst1_r5_4_), .ZN(n4326) );
  OAI222D0BWP12T U3283 ( .A1(n5023), .A2(n5143), .B1(n5249), .B2(n6303), .C1(
        n5247), .C2(n4326), .ZN(register_file_inst1_n2461) );
  INVD1BWP12T U3284 ( .I(ALU_MISC_OUT_result[5]), .ZN(n4346) );
  CKND0BWP12T U3285 ( .I(register_file_inst1_r3_5_), .ZN(n4327) );
  OAI222D0BWP12T U3286 ( .A1(n5203), .A2(n6304), .B1(n5200), .B2(n4346), .C1(
        n4758), .C2(n4327), .ZN(register_file_inst1_n2526) );
  INVD1BWP12T U3287 ( .I(register_file_inst1_r0_4_), .ZN(n5760) );
  OAI222D0BWP12T U3288 ( .A1(n5023), .A2(n5231), .B1(n5230), .B2(n6303), .C1(
        n5096), .C2(n5760), .ZN(register_file_inst1_n2621) );
  CKND0BWP12T U3289 ( .I(register_file_inst1_tmp1_5_), .ZN(n4328) );
  OAI222D0BWP12T U3290 ( .A1(n5212), .A2(n6304), .B1(n6144), .B2(n4346), .C1(
        n4683), .C2(n4328), .ZN(register_file_inst1_n2142) );
  CKND0BWP12T U3291 ( .I(register_file_inst1_lr_5_), .ZN(n4329) );
  OAI222D0BWP12T U3292 ( .A1(n5160), .A2(n6304), .B1(n5223), .B2(n4346), .C1(
        n5222), .C2(n4329), .ZN(register_file_inst1_n2206) );
  INVD1BWP12T U3293 ( .I(register_file_inst1_r6_5_), .ZN(n5736) );
  OAI222D0BWP12T U3294 ( .A1(n5228), .A2(n6304), .B1(n5229), .B2(n4346), .C1(
        n5095), .C2(n5736), .ZN(register_file_inst1_n2430) );
  INVD1BWP12T U3295 ( .I(register_file_inst1_tmp1_4_), .ZN(n5763) );
  OAI222D0BWP12T U3296 ( .A1(n5023), .A2(n6144), .B1(n5212), .B2(n6303), .C1(
        n4683), .C2(n5763), .ZN(register_file_inst1_n2141) );
  CKND0BWP12T U3297 ( .I(register_file_inst1_r5_5_), .ZN(n4330) );
  OAI222D0BWP12T U3298 ( .A1(n5249), .A2(n6304), .B1(n5143), .B2(n4346), .C1(
        n5247), .C2(n4330), .ZN(register_file_inst1_n2462) );
  INVD1BWP12T U3299 ( .I(register_file_inst1_r0_5_), .ZN(n5737) );
  OAI222D0BWP12T U3300 ( .A1(n5230), .A2(n6304), .B1(n5231), .B2(n4346), .C1(
        n5096), .C2(n5737), .ZN(register_file_inst1_n2622) );
  INVD1BWP12T U3301 ( .I(register_file_inst1_r6_4_), .ZN(n5759) );
  OAI222D0BWP12T U3302 ( .A1(n5023), .A2(n5229), .B1(n5228), .B2(n6303), .C1(
        n5095), .C2(n5759), .ZN(register_file_inst1_n2429) );
  CKND0BWP12T U3303 ( .I(register_file_inst1_r3_4_), .ZN(n4331) );
  OAI222D0BWP12T U3304 ( .A1(n5023), .A2(n5200), .B1(n5203), .B2(n6303), .C1(
        n4758), .C2(n4331), .ZN(register_file_inst1_n2525) );
  CKND0BWP12T U3305 ( .I(register_file_inst1_r9_5_), .ZN(n4332) );
  OAI222D0BWP12T U3306 ( .A1(n5237), .A2(n6304), .B1(n5238), .B2(n4346), .C1(
        n5235), .C2(n4332), .ZN(register_file_inst1_n2334) );
  CKND0BWP12T U3307 ( .I(register_file_inst1_r9_4_), .ZN(n4333) );
  OAI222D0BWP12T U3308 ( .A1(n5023), .A2(n5238), .B1(n5237), .B2(n6303), .C1(
        n5235), .C2(n4333), .ZN(register_file_inst1_n2333) );
  CKND0BWP12T U3309 ( .I(register_file_inst1_r12_4_), .ZN(n4334) );
  OAI222D0BWP12T U3310 ( .A1(n5023), .A2(n5140), .B1(n5243), .B2(n6303), .C1(
        n5242), .C2(n4334), .ZN(register_file_inst1_n2237) );
  CKND0BWP12T U3311 ( .I(register_file_inst1_lr_4_), .ZN(n4335) );
  OAI222D0BWP12T U3312 ( .A1(n5023), .A2(n5223), .B1(n5160), .B2(n6303), .C1(
        n5222), .C2(n4335), .ZN(register_file_inst1_n2205) );
  INVD1BWP12T U3313 ( .I(register_file_inst1_r12_5_), .ZN(n4336) );
  OAI222D0BWP12T U3314 ( .A1(n5243), .A2(n6304), .B1(n5140), .B2(n4346), .C1(
        n5242), .C2(n4336), .ZN(register_file_inst1_n2238) );
  INVD1BWP12T U3315 ( .I(register_file_inst1_r4_4_), .ZN(n5762) );
  OAI222D0BWP12T U3316 ( .A1(n5023), .A2(n5226), .B1(n5205), .B2(n6303), .C1(
        n5225), .C2(n5762), .ZN(register_file_inst1_n2493) );
  CKND0BWP12T U3317 ( .I(register_file_inst1_r8_4_), .ZN(n4337) );
  OAI222D0BWP12T U3318 ( .A1(n5023), .A2(n5145), .B1(n5246), .B2(n6303), .C1(
        n5244), .C2(n4337), .ZN(register_file_inst1_n2365) );
  INVD1BWP12T U3319 ( .I(register_file_inst1_r2_5_), .ZN(n5738) );
  OAI222D0BWP12T U3320 ( .A1(n5256), .A2(n6304), .B1(n5257), .B2(n4346), .C1(
        n5254), .C2(n5738), .ZN(register_file_inst1_n2558) );
  CKND0BWP12T U3321 ( .I(register_file_inst1_r8_5_), .ZN(n4338) );
  OAI222D0BWP12T U3322 ( .A1(n5246), .A2(n6304), .B1(n5145), .B2(n4346), .C1(
        n5244), .C2(n4338), .ZN(register_file_inst1_n2366) );
  INVD1BWP12T U3323 ( .I(register_file_inst1_r2_4_), .ZN(n5761) );
  OAI222D0BWP12T U3324 ( .A1(n5023), .A2(n5257), .B1(n5256), .B2(n6303), .C1(
        n5254), .C2(n5761), .ZN(register_file_inst1_n2557) );
  CKND0BWP12T U3325 ( .I(register_file_inst1_r11_5_), .ZN(n4339) );
  OAI222D0BWP12T U3326 ( .A1(n5219), .A2(n6304), .B1(n5220), .B2(n4346), .C1(
        n5217), .C2(n4339), .ZN(register_file_inst1_n2270) );
  CKND0BWP12T U3327 ( .I(register_file_inst1_r11_4_), .ZN(n4340) );
  OAI222D0BWP12T U3328 ( .A1(n5023), .A2(n5220), .B1(n5219), .B2(n6303), .C1(
        n5217), .C2(n4340), .ZN(register_file_inst1_n2269) );
  CKND0BWP12T U3329 ( .I(register_file_inst1_r7_5_), .ZN(n4341) );
  OAI222D0BWP12T U3330 ( .A1(n5158), .A2(n6304), .B1(n5227), .B2(n4346), .C1(
        n5094), .C2(n4341), .ZN(register_file_inst1_n2398) );
  CKND0BWP12T U3331 ( .I(register_file_inst1_r7_4_), .ZN(n4342) );
  OAI222D0BWP12T U3332 ( .A1(n5023), .A2(n5227), .B1(n5158), .B2(n6303), .C1(
        n5094), .C2(n4342), .ZN(register_file_inst1_n2397) );
  TPOAI21D0BWP12T U3333 ( .A1(n4346), .A2(n5234), .B(n6071), .ZN(
        register_file_inst1_spin[5]) );
  TPOAI21D0BWP12T U3334 ( .A1(n5023), .A2(n5234), .B(n6067), .ZN(
        register_file_inst1_spin[4]) );
  CKND0BWP12T U3335 ( .I(register_file_inst1_r4_5_), .ZN(n4343) );
  OAI222D0BWP12T U3336 ( .A1(n5205), .A2(n6304), .B1(n5226), .B2(n4346), .C1(
        n5225), .C2(n4343), .ZN(register_file_inst1_n2494) );
  CKND0BWP12T U3337 ( .I(register_file_inst1_r10_4_), .ZN(n4344) );
  OAI222D0BWP12T U3338 ( .A1(n5023), .A2(n5253), .B1(n5252), .B2(n6303), .C1(
        n5250), .C2(n4344), .ZN(register_file_inst1_n2301) );
  INVD1BWP12T U3339 ( .I(register_file_inst1_r10_5_), .ZN(n4345) );
  OAI222D0BWP12T U3340 ( .A1(n5252), .A2(n6304), .B1(n5253), .B2(n4346), .C1(
        n5250), .C2(n4345), .ZN(register_file_inst1_n2302) );
  INVD1BWP12T U3341 ( .I(register_file_inst1_r1_4_), .ZN(n5758) );
  OAI222D0BWP12T U3342 ( .A1(n5023), .A2(n5074), .B1(n5240), .B2(n6303), .C1(
        n5239), .C2(n5758), .ZN(register_file_inst1_n2589) );
  INVD1BWP12T U3343 ( .I(register_file_inst1_r1_5_), .ZN(n5735) );
  OAI222D0BWP12T U3344 ( .A1(n5240), .A2(n6304), .B1(n5074), .B2(n4346), .C1(
        n5239), .C2(n5735), .ZN(register_file_inst1_n2590) );
  INVD1BWP12T U3345 ( .I(ALU_MISC_OUT_result[2]), .ZN(n5022) );
  CKND0BWP12T U3346 ( .I(register_file_inst1_r3_2_), .ZN(n4347) );
  OAI222D0BWP12T U3347 ( .A1(n5022), .A2(n5200), .B1(n5203), .B2(n6302), .C1(
        n4758), .C2(n4347), .ZN(register_file_inst1_n2523) );
  CKND0BWP12T U3348 ( .I(register_file_inst1_r5_2_), .ZN(n4348) );
  OAI222D0BWP12T U3349 ( .A1(n5022), .A2(n5143), .B1(n5249), .B2(n6302), .C1(
        n5247), .C2(n4348), .ZN(register_file_inst1_n2459) );
  INVD1BWP12T U3350 ( .I(register_file_inst1_r12_2_), .ZN(n4349) );
  OAI222D0BWP12T U3351 ( .A1(n5022), .A2(n5140), .B1(n5243), .B2(n6302), .C1(
        n5242), .C2(n4349), .ZN(register_file_inst1_n2235) );
  CKND0BWP12T U3352 ( .I(register_file_inst1_r9_2_), .ZN(n4350) );
  OAI222D0BWP12T U3353 ( .A1(n5022), .A2(n5238), .B1(n5237), .B2(n6302), .C1(
        n5235), .C2(n4350), .ZN(register_file_inst1_n2331) );
  INVD1BWP12T U3354 ( .I(register_file_inst1_r1_2_), .ZN(n5801) );
  OAI222D0BWP12T U3355 ( .A1(n5022), .A2(n5074), .B1(n5240), .B2(n6302), .C1(
        n5239), .C2(n5801), .ZN(register_file_inst1_n2587) );
  INVD1BWP12T U3356 ( .I(register_file_inst1_tmp1_2_), .ZN(n5807) );
  OAI222D0BWP12T U3357 ( .A1(n5022), .A2(n6144), .B1(n5212), .B2(n6302), .C1(
        n4683), .C2(n5807), .ZN(register_file_inst1_n2139) );
  CKND0BWP12T U3358 ( .I(register_file_inst1_r7_2_), .ZN(n4351) );
  OAI222D0BWP12T U3359 ( .A1(n5022), .A2(n5227), .B1(n5158), .B2(n6302), .C1(
        n5094), .C2(n4351), .ZN(register_file_inst1_n2395) );
  INVD1BWP12T U3360 ( .I(register_file_inst1_r0_2_), .ZN(n5803) );
  OAI222D0BWP12T U3361 ( .A1(n5022), .A2(n5231), .B1(n5230), .B2(n6302), .C1(
        n5096), .C2(n5803), .ZN(register_file_inst1_n2619) );
  INVD1BWP12T U3362 ( .I(register_file_inst1_r6_2_), .ZN(n5802) );
  OAI222D0BWP12T U3363 ( .A1(n5022), .A2(n5229), .B1(n5228), .B2(n6302), .C1(
        n5095), .C2(n5802), .ZN(register_file_inst1_n2427) );
  INVD1BWP12T U3364 ( .I(register_file_inst1_r4_2_), .ZN(n5806) );
  OAI222D0BWP12T U3365 ( .A1(n5022), .A2(n5226), .B1(n5205), .B2(n6302), .C1(
        n5225), .C2(n5806), .ZN(register_file_inst1_n2491) );
  TPOAI21D0BWP12T U3366 ( .A1(n5022), .A2(n5234), .B(n6058), .ZN(
        register_file_inst1_spin[2]) );
  CKND0BWP12T U3367 ( .I(register_file_inst1_r11_2_), .ZN(n4352) );
  OAI222D0BWP12T U3368 ( .A1(n5022), .A2(n5220), .B1(n5219), .B2(n6302), .C1(
        n5217), .C2(n4352), .ZN(register_file_inst1_n2267) );
  CKND0BWP12T U3369 ( .I(register_file_inst1_lr_2_), .ZN(n4353) );
  OAI222D0BWP12T U3370 ( .A1(n5022), .A2(n5223), .B1(n5160), .B2(n6302), .C1(
        n5222), .C2(n4353), .ZN(register_file_inst1_n2203) );
  INVD0BWP12T U3371 ( .I(register_file_inst1_r8_2_), .ZN(n4354) );
  OAI222D0BWP12T U3372 ( .A1(n5022), .A2(n5145), .B1(n5246), .B2(n6302), .C1(
        n5244), .C2(n4354), .ZN(register_file_inst1_n2363) );
  CKND0BWP12T U3373 ( .I(register_file_inst1_r10_2_), .ZN(n4355) );
  OAI222D0BWP12T U3374 ( .A1(n5022), .A2(n5253), .B1(n5252), .B2(n6302), .C1(
        n5250), .C2(n4355), .ZN(register_file_inst1_n2299) );
  INVD1BWP12T U3375 ( .I(register_file_inst1_r2_2_), .ZN(n5804) );
  OAI222D0BWP12T U3376 ( .A1(n5022), .A2(n5257), .B1(n5256), .B2(n6302), .C1(
        n5254), .C2(n5804), .ZN(register_file_inst1_n2555) );
  INVD1BWP12T U3377 ( .I(ALU_MISC_OUT_result[1]), .ZN(n4386) );
  INVD1BWP12T U3378 ( .I(register_file_inst1_r4_1_), .ZN(n4356) );
  OAI222D0BWP12T U3379 ( .A1(n6054), .A2(n5205), .B1(n4386), .B2(n5226), .C1(
        n5225), .C2(n4356), .ZN(register_file_inst1_n2490) );
  INVD1BWP12T U3380 ( .I(ALU_MISC_OUT_result[3]), .ZN(n4385) );
  INVD1BWP12T U3381 ( .I(register_file_inst1_r11_3_), .ZN(n4357) );
  OAI222D0BWP12T U3382 ( .A1(n4385), .A2(n5220), .B1(n5219), .B2(n6063), .C1(
        n5217), .C2(n4357), .ZN(register_file_inst1_n2268) );
  INVD1BWP12T U3383 ( .I(register_file_inst1_r10_3_), .ZN(n4358) );
  OAI222D0BWP12T U3384 ( .A1(n4385), .A2(n5253), .B1(n5252), .B2(n6063), .C1(
        n5250), .C2(n4358), .ZN(register_file_inst1_n2300) );
  TPOAI21D0BWP12T U3385 ( .A1(n4386), .A2(n5234), .B(n6053), .ZN(
        register_file_inst1_spin[1]) );
  INVD1BWP12T U3386 ( .I(register_file_inst1_r10_1_), .ZN(n4359) );
  OAI222D0BWP12T U3387 ( .A1(n4359), .A2(n5250), .B1(n4386), .B2(n5253), .C1(
        n6054), .C2(n5252), .ZN(register_file_inst1_n2298) );
  CKND0BWP12T U3388 ( .I(register_file_inst1_r2_1_), .ZN(n4360) );
  OAI222D0BWP12T U3389 ( .A1(n4360), .A2(n5254), .B1(n4386), .B2(n5257), .C1(
        n5256), .C2(n6054), .ZN(register_file_inst1_n2554) );
  CKND0BWP12T U3390 ( .I(register_file_inst1_r0_1_), .ZN(n4361) );
  OAI222D0BWP12T U3391 ( .A1(n4361), .A2(n5096), .B1(n4386), .B2(n5231), .C1(
        n6054), .C2(n5230), .ZN(register_file_inst1_n2618) );
  INVD1BWP12T U3392 ( .I(register_file_inst1_r8_3_), .ZN(n4362) );
  OAI222D0BWP12T U3393 ( .A1(n4385), .A2(n5145), .B1(n5246), .B2(n6063), .C1(
        n5244), .C2(n4362), .ZN(register_file_inst1_n2364) );
  CKND0BWP12T U3394 ( .I(register_file_inst1_r2_3_), .ZN(n4363) );
  OAI222D0BWP12T U3395 ( .A1(n4385), .A2(n5257), .B1(n5256), .B2(n6063), .C1(
        n5254), .C2(n4363), .ZN(register_file_inst1_n2556) );
  INVD1BWP12T U3396 ( .I(register_file_inst1_r6_1_), .ZN(n4364) );
  OAI222D0BWP12T U3397 ( .A1(n4364), .A2(n5095), .B1(n4386), .B2(n5229), .C1(
        n6054), .C2(n5228), .ZN(register_file_inst1_n2426) );
  TPOAI21D0BWP12T U3398 ( .A1(n4385), .A2(n5234), .B(n6062), .ZN(
        register_file_inst1_spin[3]) );
  INVD1BWP12T U3399 ( .I(register_file_inst1_r8_1_), .ZN(n4365) );
  OAI222D0BWP12T U3400 ( .A1(n4365), .A2(n5244), .B1(n4386), .B2(n5145), .C1(
        n6054), .C2(n5246), .ZN(register_file_inst1_n2362) );
  INVD1BWP12T U3401 ( .I(register_file_inst1_r11_1_), .ZN(n4366) );
  OAI222D0BWP12T U3402 ( .A1(n4366), .A2(n5217), .B1(n4386), .B2(n5220), .C1(
        n6054), .C2(n5219), .ZN(register_file_inst1_n2266) );
  CKND0BWP12T U3403 ( .I(register_file_inst1_r0_3_), .ZN(n4367) );
  OAI222D0BWP12T U3404 ( .A1(n4385), .A2(n5231), .B1(n5230), .B2(n6063), .C1(
        n5096), .C2(n4367), .ZN(register_file_inst1_n2620) );
  CKND0BWP12T U3405 ( .I(register_file_inst1_r4_3_), .ZN(n4368) );
  OAI222D0BWP12T U3406 ( .A1(n4385), .A2(n5226), .B1(n5205), .B2(n6063), .C1(
        n5225), .C2(n4368), .ZN(register_file_inst1_n2492) );
  INVD1BWP12T U3407 ( .I(register_file_inst1_lr_1_), .ZN(n4369) );
  OAI222D0BWP12T U3408 ( .A1(n6054), .A2(n5160), .B1(n4386), .B2(n5223), .C1(
        n5222), .C2(n4369), .ZN(register_file_inst1_n2202) );
  CKND0BWP12T U3409 ( .I(register_file_inst1_r1_3_), .ZN(n4370) );
  OAI222D0BWP12T U3410 ( .A1(n4385), .A2(n5074), .B1(n5240), .B2(n6063), .C1(
        n5239), .C2(n4370), .ZN(register_file_inst1_n2588) );
  INVD1BWP12T U3411 ( .I(register_file_inst1_lr_3_), .ZN(n4371) );
  OAI222D0BWP12T U3412 ( .A1(n4385), .A2(n5223), .B1(n5160), .B2(n6063), .C1(
        n5222), .C2(n4371), .ZN(register_file_inst1_n2204) );
  INVD1BWP12T U3413 ( .I(register_file_inst1_r6_3_), .ZN(n4372) );
  OAI222D0BWP12T U3414 ( .A1(n4385), .A2(n5229), .B1(n5228), .B2(n6063), .C1(
        n5095), .C2(n4372), .ZN(register_file_inst1_n2428) );
  INVD1BWP12T U3415 ( .I(register_file_inst1_r7_1_), .ZN(n4373) );
  OAI222D0BWP12T U3416 ( .A1(n4373), .A2(n5094), .B1(n4386), .B2(n5227), .C1(
        n6054), .C2(n5158), .ZN(register_file_inst1_n2394) );
  CKND0BWP12T U3417 ( .I(register_file_inst1_tmp1_1_), .ZN(n4374) );
  OAI222D0BWP12T U3418 ( .A1(n6054), .A2(n5212), .B1(n4386), .B2(n6144), .C1(
        n4683), .C2(n4374), .ZN(register_file_inst1_n2138) );
  INVD1BWP12T U3419 ( .I(register_file_inst1_r9_3_), .ZN(n4375) );
  OAI222D0BWP12T U3420 ( .A1(n4385), .A2(n5238), .B1(n5237), .B2(n6063), .C1(
        n5235), .C2(n4375), .ZN(register_file_inst1_n2332) );
  INVD1BWP12T U3421 ( .I(register_file_inst1_r5_3_), .ZN(n4376) );
  OAI222D0BWP12T U3422 ( .A1(n4385), .A2(n5143), .B1(n5249), .B2(n6063), .C1(
        n5247), .C2(n4376), .ZN(register_file_inst1_n2460) );
  INVD1BWP12T U3423 ( .I(register_file_inst1_r12_1_), .ZN(n4377) );
  OAI222D0BWP12T U3424 ( .A1(n6054), .A2(n5243), .B1(n4386), .B2(n5140), .C1(
        n5242), .C2(n4377), .ZN(register_file_inst1_n2234) );
  INVD1BWP12T U3425 ( .I(register_file_inst1_r12_3_), .ZN(n4378) );
  OAI222D0BWP12T U3426 ( .A1(n4385), .A2(n5140), .B1(n5243), .B2(n6063), .C1(
        n5242), .C2(n4378), .ZN(register_file_inst1_n2236) );
  INVD1BWP12T U3427 ( .I(register_file_inst1_r9_1_), .ZN(n4379) );
  OAI222D0BWP12T U3428 ( .A1(n4379), .A2(n5235), .B1(n4386), .B2(n5238), .C1(
        n6054), .C2(n5237), .ZN(register_file_inst1_n2330) );
  CKND0BWP12T U3429 ( .I(register_file_inst1_r7_3_), .ZN(n4380) );
  OAI222D0BWP12T U3430 ( .A1(n4385), .A2(n5227), .B1(n5158), .B2(n6063), .C1(
        n5094), .C2(n4380), .ZN(register_file_inst1_n2396) );
  INVD1BWP12T U3431 ( .I(register_file_inst1_r5_1_), .ZN(n4381) );
  OAI222D0BWP12T U3432 ( .A1(n4381), .A2(n5247), .B1(n4386), .B2(n5143), .C1(
        n6054), .C2(n5249), .ZN(register_file_inst1_n2458) );
  INVD1BWP12T U3433 ( .I(register_file_inst1_r3_3_), .ZN(n4382) );
  OAI222D0BWP12T U3434 ( .A1(n4385), .A2(n5200), .B1(n5203), .B2(n6063), .C1(
        n4758), .C2(n4382), .ZN(register_file_inst1_n2524) );
  INVD1BWP12T U3435 ( .I(register_file_inst1_r3_1_), .ZN(n4383) );
  OAI222D0BWP12T U3436 ( .A1(n6054), .A2(n5203), .B1(n4386), .B2(n5200), .C1(
        n4758), .C2(n4383), .ZN(register_file_inst1_n2522) );
  CKND0BWP12T U3437 ( .I(register_file_inst1_tmp1_3_), .ZN(n4384) );
  OAI222D0BWP12T U3438 ( .A1(n4385), .A2(n6144), .B1(n5212), .B2(n6063), .C1(
        n4683), .C2(n4384), .ZN(register_file_inst1_n2140) );
  CKND0BWP12T U3439 ( .I(register_file_inst1_r1_1_), .ZN(n4387) );
  OAI222D0BWP12T U3440 ( .A1(n4387), .A2(n5239), .B1(n4386), .B2(n5074), .C1(
        n6054), .C2(n5240), .ZN(register_file_inst1_n2586) );
  INVD1BWP12T U3441 ( .I(register_file_inst1_r0_0_), .ZN(n4618) );
  INVD1BWP12T U3442 ( .I(ALU_MISC_OUT_result[0]), .ZN(n5020) );
  OAI222D0BWP12T U3443 ( .A1(n4618), .A2(n5096), .B1(n5020), .B2(n5231), .C1(
        n3718), .C2(n5230), .ZN(register_file_inst1_n2617) );
  INVD1BWP12T U3444 ( .I(register_file_inst1_lr_0_), .ZN(n5846) );
  OAI222D0BWP12T U3445 ( .A1(n3718), .A2(n5160), .B1(n5020), .B2(n5223), .C1(
        n5222), .C2(n5846), .ZN(register_file_inst1_n2201) );
  INVD1BWP12T U3446 ( .I(register_file_inst1_r5_0_), .ZN(n4388) );
  OAI222D0BWP12T U3447 ( .A1(n4388), .A2(n5247), .B1(n5020), .B2(n5143), .C1(
        n3718), .C2(n5249), .ZN(register_file_inst1_n2457) );
  INVD1BWP12T U3448 ( .I(RF_next_sp[0]), .ZN(n5842) );
  OAI222D0BWP12T U3449 ( .A1(n5842), .A2(n5232), .B1(n5020), .B2(n5234), .C1(
        n3718), .C2(n5233), .ZN(register_file_inst1_spin[0]) );
  CKND0BWP12T U3450 ( .I(register_file_inst1_r12_0_), .ZN(n4389) );
  OAI222D0BWP12T U3451 ( .A1(n3718), .A2(n5243), .B1(n5020), .B2(n5140), .C1(
        n5242), .C2(n4389), .ZN(register_file_inst1_n2233) );
  INVD1BWP12T U3452 ( .I(register_file_inst1_r9_0_), .ZN(n4390) );
  OAI222D0BWP12T U3453 ( .A1(n4390), .A2(n5235), .B1(n5020), .B2(n5238), .C1(
        n3718), .C2(n5237), .ZN(register_file_inst1_n2329) );
  INVD1BWP12T U3454 ( .I(register_file_inst1_r6_0_), .ZN(n4391) );
  OAI222D0BWP12T U3455 ( .A1(n4391), .A2(n5095), .B1(n5020), .B2(n5229), .C1(
        n3718), .C2(n5228), .ZN(register_file_inst1_n2425) );
  INVD1BWP12T U3456 ( .I(register_file_inst1_r3_0_), .ZN(n4392) );
  OAI222D0BWP12T U3457 ( .A1(n3718), .A2(n5203), .B1(n5020), .B2(n5200), .C1(
        n4758), .C2(n4392), .ZN(register_file_inst1_n2521) );
  INVD1BWP12T U3458 ( .I(register_file_inst1_r2_0_), .ZN(n4621) );
  OAI222D0BWP12T U3459 ( .A1(n4621), .A2(n5254), .B1(n5020), .B2(n5257), .C1(
        n5256), .C2(n3718), .ZN(register_file_inst1_n2553) );
  OAI222D0BWP12T U3460 ( .A1(n5843), .A2(n5239), .B1(n5020), .B2(n5074), .C1(
        n3718), .C2(n5240), .ZN(register_file_inst1_n2585) );
  INVD1BWP12T U3461 ( .I(register_file_inst1_r7_0_), .ZN(n4393) );
  OAI222D0BWP12T U3462 ( .A1(n4393), .A2(n5094), .B1(n5020), .B2(n5227), .C1(
        n3718), .C2(n5158), .ZN(register_file_inst1_n2393) );
  INVD1BWP12T U3463 ( .I(register_file_inst1_r8_0_), .ZN(n4394) );
  OAI222D0BWP12T U3464 ( .A1(n4394), .A2(n5244), .B1(n5020), .B2(n5145), .C1(
        n3718), .C2(n5246), .ZN(register_file_inst1_n2361) );
  INVD1BWP12T U3465 ( .I(register_file_inst1_r10_0_), .ZN(n5845) );
  OAI222D0BWP12T U3466 ( .A1(n5845), .A2(n5250), .B1(n5020), .B2(n5253), .C1(
        n3718), .C2(n5252), .ZN(register_file_inst1_n2297) );
  INVD1BWP12T U3467 ( .I(register_file_inst1_r11_0_), .ZN(n4395) );
  OAI222D0BWP12T U3468 ( .A1(n4395), .A2(n5217), .B1(n5020), .B2(n5220), .C1(
        n3718), .C2(n5219), .ZN(register_file_inst1_n2265) );
  ND2D1BWP12T U3469 ( .A1(n2907), .A2(n2908), .ZN(n4396) );
  AOI22D0BWP12T U3470 ( .A1(register_file_inst1_r1_13_), .A2(n5001), .B1(
        register_file_inst1_r3_13_), .B2(n4989), .ZN(n4400) );
  ND2D1BWP12T U3471 ( .A1(n2906), .A2(n2905), .ZN(n4547) );
  AOI22D0BWP12T U3472 ( .A1(register_file_inst1_r2_13_), .A2(n4962), .B1(
        register_file_inst1_r0_13_), .B2(n5002), .ZN(n4399) );
  AOI22D0BWP12T U3473 ( .A1(register_file_inst1_r4_13_), .A2(n5003), .B1(
        register_file_inst1_r5_13_), .B2(n4990), .ZN(n4398) );
  AOI22D0BWP12T U3474 ( .A1(register_file_inst1_r6_13_), .A2(n5004), .B1(
        register_file_inst1_r7_13_), .B2(n4991), .ZN(n4397) );
  ND4D1BWP12T U3475 ( .A1(n4400), .A2(n4399), .A3(n4398), .A4(n4397), .ZN(
        n4405) );
  NR2D1BWP12T U3476 ( .A1(n2920), .A2(n2919), .ZN(n4437) );
  NR2D1BWP12T U3477 ( .A1(n2919), .A2(n4547), .ZN(n4510) );
  INVD1BWP12T U3478 ( .I(n4510), .ZN(n4673) );
  AOI22D1BWP12T U3479 ( .A1(register_file_inst1_lr_13_), .A2(n4437), .B1(
        register_file_inst1_r12_13_), .B2(n4510), .ZN(n4403) );
  OR2XD1BWP12T U3480 ( .A1(n2911), .A2(n2917), .Z(n4672) );
  AOI22D1BWP12T U3481 ( .A1(RF_next_sp[13]), .A2(n5010), .B1(
        register_file_inst1_r11_13_), .B2(n5009), .ZN(n4402) );
  AOI22D0BWP12T U3482 ( .A1(register_file_inst1_r9_13_), .A2(n6005), .B1(
        register_file_inst1_r10_13_), .B2(n5011), .ZN(n4401) );
  ND4D1BWP12T U3483 ( .A1(n6238), .A2(n4403), .A3(n4402), .A4(n4401), .ZN(
        n4404) );
  AO21D1BWP12T U3484 ( .A1(n3502), .A2(n4405), .B(n4404), .Z(
        RF_MEMCTRL_data_reg[13]) );
  AOI22D1BWP12T U3485 ( .A1(register_file_inst1_r1_15_), .A2(n5001), .B1(
        register_file_inst1_r3_15_), .B2(n4989), .ZN(n4409) );
  AOI22D0BWP12T U3486 ( .A1(register_file_inst1_r2_15_), .A2(n4962), .B1(
        register_file_inst1_r0_15_), .B2(n5002), .ZN(n4408) );
  AOI22D1BWP12T U3487 ( .A1(register_file_inst1_r4_15_), .A2(n5003), .B1(
        register_file_inst1_r5_15_), .B2(n4990), .ZN(n4407) );
  AOI22D1BWP12T U3488 ( .A1(register_file_inst1_r6_15_), .A2(n5004), .B1(
        register_file_inst1_r7_15_), .B2(n4991), .ZN(n4406) );
  ND4D1BWP12T U3489 ( .A1(n4409), .A2(n4408), .A3(n4407), .A4(n4406), .ZN(
        n4414) );
  AOI22D1BWP12T U3490 ( .A1(register_file_inst1_lr_15_), .A2(n4437), .B1(
        register_file_inst1_r12_15_), .B2(n4510), .ZN(n4412) );
  AOI22D1BWP12T U3491 ( .A1(RF_next_sp[15]), .A2(n5010), .B1(
        register_file_inst1_r11_15_), .B2(n5009), .ZN(n4411) );
  AOI22D1BWP12T U3492 ( .A1(register_file_inst1_r9_15_), .A2(n6005), .B1(
        register_file_inst1_r10_15_), .B2(n5011), .ZN(n4410) );
  ND4D1BWP12T U3493 ( .A1(n6268), .A2(n4412), .A3(n4411), .A4(n4410), .ZN(
        n4413) );
  AO21D1BWP12T U3494 ( .A1(n3502), .A2(n4414), .B(n4413), .Z(
        RF_MEMCTRL_data_reg[15]) );
  AOI22D0BWP12T U3495 ( .A1(register_file_inst1_r1_14_), .A2(n5001), .B1(
        register_file_inst1_r3_14_), .B2(n4989), .ZN(n4418) );
  AOI22D0BWP12T U3496 ( .A1(register_file_inst1_r2_14_), .A2(n4962), .B1(
        register_file_inst1_r0_14_), .B2(n5002), .ZN(n4417) );
  AOI22D0BWP12T U3497 ( .A1(register_file_inst1_r4_14_), .A2(n5003), .B1(
        register_file_inst1_r5_14_), .B2(n4990), .ZN(n4416) );
  AOI22D0BWP12T U3498 ( .A1(register_file_inst1_r6_14_), .A2(n5004), .B1(
        register_file_inst1_r7_14_), .B2(n4991), .ZN(n4415) );
  ND4D1BWP12T U3499 ( .A1(n4418), .A2(n4417), .A3(n4416), .A4(n4415), .ZN(
        n4423) );
  AOI22D1BWP12T U3500 ( .A1(register_file_inst1_lr_14_), .A2(n4437), .B1(
        register_file_inst1_r12_14_), .B2(n4510), .ZN(n4421) );
  AOI22D1BWP12T U3501 ( .A1(RF_next_sp[14]), .A2(n5010), .B1(
        register_file_inst1_r11_14_), .B2(n5009), .ZN(n4420) );
  AOI22D1BWP12T U3502 ( .A1(register_file_inst1_r9_14_), .A2(n6005), .B1(
        register_file_inst1_r10_14_), .B2(n5011), .ZN(n4419) );
  ND4D1BWP12T U3503 ( .A1(n6259), .A2(n4421), .A3(n4420), .A4(n4419), .ZN(
        n4422) );
  AO21D1BWP12T U3504 ( .A1(n3502), .A2(n4423), .B(n4422), .Z(
        RF_MEMCTRL_data_reg[14]) );
  AOI22D0BWP12T U3505 ( .A1(register_file_inst1_r1_8_), .A2(n5001), .B1(
        register_file_inst1_r3_8_), .B2(n4989), .ZN(n4427) );
  AOI22D0BWP12T U3506 ( .A1(register_file_inst1_r2_8_), .A2(n4962), .B1(
        register_file_inst1_r0_8_), .B2(n5002), .ZN(n4426) );
  AOI22D0BWP12T U3507 ( .A1(register_file_inst1_r4_8_), .A2(n5003), .B1(
        register_file_inst1_r5_8_), .B2(n4990), .ZN(n4425) );
  AOI22D0BWP12T U3508 ( .A1(register_file_inst1_r6_8_), .A2(n5004), .B1(
        register_file_inst1_r7_8_), .B2(n4991), .ZN(n4424) );
  ND4D1BWP12T U3509 ( .A1(n4427), .A2(n4426), .A3(n4425), .A4(n4424), .ZN(
        n4432) );
  AOI22D1BWP12T U3510 ( .A1(register_file_inst1_lr_8_), .A2(n4437), .B1(
        register_file_inst1_r12_8_), .B2(n4510), .ZN(n4430) );
  AOI22D1BWP12T U3511 ( .A1(register_file_inst1_r11_8_), .A2(n5009), .B1(
        RF_next_sp[8]), .B2(n5010), .ZN(n4429) );
  AOI22D0BWP12T U3512 ( .A1(register_file_inst1_r9_8_), .A2(n6005), .B1(
        register_file_inst1_r10_8_), .B2(n5011), .ZN(n4428) );
  ND4D1BWP12T U3513 ( .A1(n6277), .A2(n4430), .A3(n4429), .A4(n4428), .ZN(
        n4431) );
  AO21D1BWP12T U3514 ( .A1(n3502), .A2(n4432), .B(n4431), .Z(
        RF_MEMCTRL_data_reg[8]) );
  AOI22D1BWP12T U3515 ( .A1(register_file_inst1_r1_9_), .A2(n5001), .B1(
        register_file_inst1_r3_9_), .B2(n4989), .ZN(n4436) );
  AOI22D1BWP12T U3516 ( .A1(register_file_inst1_r2_9_), .A2(n4962), .B1(
        register_file_inst1_r0_9_), .B2(n5002), .ZN(n4435) );
  AOI22D1BWP12T U3517 ( .A1(register_file_inst1_r4_9_), .A2(n5003), .B1(
        register_file_inst1_r5_9_), .B2(n4990), .ZN(n4434) );
  AOI22D0BWP12T U3518 ( .A1(register_file_inst1_r6_9_), .A2(n5004), .B1(
        register_file_inst1_r7_9_), .B2(n4991), .ZN(n4433) );
  ND4D1BWP12T U3519 ( .A1(n4436), .A2(n4435), .A3(n4434), .A4(n4433), .ZN(
        n4442) );
  AOI22D1BWP12T U3520 ( .A1(register_file_inst1_lr_9_), .A2(n4437), .B1(
        register_file_inst1_r12_9_), .B2(n4510), .ZN(n4440) );
  AOI22D1BWP12T U3521 ( .A1(register_file_inst1_r11_9_), .A2(n5009), .B1(
        RF_next_sp[9]), .B2(n5010), .ZN(n4439) );
  AOI22D1BWP12T U3522 ( .A1(register_file_inst1_r9_9_), .A2(n6005), .B1(
        register_file_inst1_r10_9_), .B2(n5011), .ZN(n4438) );
  ND4D1BWP12T U3523 ( .A1(n6233), .A2(n4440), .A3(n4439), .A4(n4438), .ZN(
        n4441) );
  AO21D1BWP12T U3524 ( .A1(n3502), .A2(n4442), .B(n4441), .Z(
        RF_MEMCTRL_data_reg[9]) );
  AOI22D0BWP12T U3525 ( .A1(register_file_inst1_r1_10_), .A2(n5001), .B1(
        register_file_inst1_r3_10_), .B2(n4989), .ZN(n4446) );
  AOI22D0BWP12T U3526 ( .A1(register_file_inst1_r2_10_), .A2(n4962), .B1(
        register_file_inst1_r0_10_), .B2(n5002), .ZN(n4445) );
  AOI22D0BWP12T U3527 ( .A1(register_file_inst1_r4_10_), .A2(n5003), .B1(
        register_file_inst1_r5_10_), .B2(n4990), .ZN(n4444) );
  AOI22D0BWP12T U3528 ( .A1(register_file_inst1_r6_10_), .A2(n5004), .B1(
        register_file_inst1_r7_10_), .B2(n4991), .ZN(n4443) );
  ND4D1BWP12T U3529 ( .A1(n4446), .A2(n4445), .A3(n4444), .A4(n4443), .ZN(
        n4451) );
  AOI22D1BWP12T U3530 ( .A1(register_file_inst1_lr_10_), .A2(n4437), .B1(
        register_file_inst1_r12_10_), .B2(n4510), .ZN(n4449) );
  AOI22D1BWP12T U3531 ( .A1(register_file_inst1_r11_10_), .A2(n5009), .B1(
        RF_next_sp[10]), .B2(n5010), .ZN(n4448) );
  AOI22D0BWP12T U3532 ( .A1(register_file_inst1_r9_10_), .A2(n6005), .B1(
        register_file_inst1_r10_10_), .B2(n5011), .ZN(n4447) );
  ND4D1BWP12T U3533 ( .A1(n6250), .A2(n4449), .A3(n4448), .A4(n4447), .ZN(
        n4450) );
  AO21D1BWP12T U3534 ( .A1(n3502), .A2(n4451), .B(n4450), .Z(
        RF_MEMCTRL_data_reg[10]) );
  AOI22D1BWP12T U3535 ( .A1(register_file_inst1_r3_11_), .A2(n4989), .B1(
        register_file_inst1_r1_11_), .B2(n5001), .ZN(n4455) );
  AOI22D0BWP12T U3536 ( .A1(register_file_inst1_r2_11_), .A2(n4962), .B1(
        register_file_inst1_r0_11_), .B2(n5002), .ZN(n4454) );
  AOI22D1BWP12T U3537 ( .A1(register_file_inst1_r5_11_), .A2(n4990), .B1(
        register_file_inst1_r4_11_), .B2(n5003), .ZN(n4453) );
  AOI22D0BWP12T U3538 ( .A1(register_file_inst1_r7_11_), .A2(n4991), .B1(
        register_file_inst1_r6_11_), .B2(n5004), .ZN(n4452) );
  ND4D1BWP12T U3539 ( .A1(n4455), .A2(n4454), .A3(n4453), .A4(n4452), .ZN(
        n4460) );
  AOI22D1BWP12T U3540 ( .A1(register_file_inst1_lr_11_), .A2(n4437), .B1(
        register_file_inst1_r12_11_), .B2(n4510), .ZN(n4458) );
  AOI22D1BWP12T U3541 ( .A1(RF_next_sp[11]), .A2(n5010), .B1(
        register_file_inst1_r11_11_), .B2(n5009), .ZN(n4457) );
  AOI22D0BWP12T U3542 ( .A1(register_file_inst1_r9_11_), .A2(n6005), .B1(
        register_file_inst1_r10_11_), .B2(n5011), .ZN(n4456) );
  ND4D1BWP12T U3543 ( .A1(n6281), .A2(n4458), .A3(n4457), .A4(n4456), .ZN(
        n4459) );
  AO21D1BWP12T U3544 ( .A1(n3502), .A2(n4460), .B(n4459), .Z(
        RF_MEMCTRL_data_reg[11]) );
  AOI22D1BWP12T U3545 ( .A1(register_file_inst1_r3_12_), .A2(n4989), .B1(
        register_file_inst1_r1_12_), .B2(n5001), .ZN(n4464) );
  AOI22D0BWP12T U3546 ( .A1(register_file_inst1_r2_12_), .A2(n4962), .B1(
        register_file_inst1_r0_12_), .B2(n5002), .ZN(n4463) );
  AOI22D1BWP12T U3547 ( .A1(register_file_inst1_r5_12_), .A2(n4990), .B1(
        register_file_inst1_r4_12_), .B2(n5003), .ZN(n4462) );
  AOI22D0BWP12T U3548 ( .A1(register_file_inst1_r7_12_), .A2(n4991), .B1(
        register_file_inst1_r6_12_), .B2(n5004), .ZN(n4461) );
  ND4D1BWP12T U3549 ( .A1(n4464), .A2(n4463), .A3(n4462), .A4(n4461), .ZN(
        n4469) );
  AOI22D1BWP12T U3550 ( .A1(register_file_inst1_lr_12_), .A2(n4437), .B1(
        register_file_inst1_r12_12_), .B2(n4510), .ZN(n4467) );
  AOI22D1BWP12T U3551 ( .A1(RF_next_sp[12]), .A2(n5010), .B1(
        register_file_inst1_r11_12_), .B2(n5009), .ZN(n4466) );
  AOI22D1BWP12T U3552 ( .A1(register_file_inst1_r9_12_), .A2(n6005), .B1(
        register_file_inst1_r10_12_), .B2(n5011), .ZN(n4465) );
  ND4D1BWP12T U3553 ( .A1(n6255), .A2(n4467), .A3(n4466), .A4(n4465), .ZN(
        n4468) );
  AO21D1BWP12T U3554 ( .A1(n3502), .A2(n4469), .B(n4468), .Z(
        RF_MEMCTRL_data_reg[12]) );
  AOI22D1BWP12T U3555 ( .A1(register_file_inst1_r1_1_), .A2(n5001), .B1(
        register_file_inst1_r3_1_), .B2(n4989), .ZN(n4473) );
  AOI22D0BWP12T U3556 ( .A1(register_file_inst1_r2_1_), .A2(n4962), .B1(
        register_file_inst1_r0_1_), .B2(n5002), .ZN(n4472) );
  AOI22D1BWP12T U3557 ( .A1(register_file_inst1_r4_1_), .A2(n5003), .B1(
        register_file_inst1_r5_1_), .B2(n4990), .ZN(n4471) );
  AOI22D1BWP12T U3558 ( .A1(register_file_inst1_r6_1_), .A2(n5004), .B1(
        register_file_inst1_r7_1_), .B2(n4991), .ZN(n4470) );
  ND4D1BWP12T U3559 ( .A1(n4473), .A2(n4472), .A3(n4471), .A4(n4470), .ZN(
        n4478) );
  AOI22D1BWP12T U3560 ( .A1(register_file_inst1_lr_1_), .A2(n4437), .B1(
        register_file_inst1_r12_1_), .B2(n4510), .ZN(n4476) );
  AOI22D1BWP12T U3561 ( .A1(register_file_inst1_r11_1_), .A2(n5009), .B1(
        RF_next_sp[1]), .B2(n5010), .ZN(n4475) );
  AOI22D1BWP12T U3562 ( .A1(register_file_inst1_r9_1_), .A2(n6005), .B1(
        register_file_inst1_r10_1_), .B2(n5011), .ZN(n4474) );
  ND4D1BWP12T U3563 ( .A1(n6248), .A2(n4476), .A3(n4475), .A4(n4474), .ZN(
        n4477) );
  AO21D1BWP12T U3564 ( .A1(n3502), .A2(n4478), .B(n4477), .Z(
        RF_MEMCTRL_data_reg[1]) );
  AOI22D0BWP12T U3565 ( .A1(register_file_inst1_r1_17_), .A2(n5001), .B1(
        register_file_inst1_r3_17_), .B2(n4989), .ZN(n4482) );
  AOI22D0BWP12T U3566 ( .A1(register_file_inst1_r2_17_), .A2(n4962), .B1(
        register_file_inst1_r0_17_), .B2(n5002), .ZN(n4481) );
  AOI22D0BWP12T U3567 ( .A1(register_file_inst1_r4_17_), .A2(n5003), .B1(
        register_file_inst1_r5_17_), .B2(n4990), .ZN(n4480) );
  AOI22D0BWP12T U3568 ( .A1(register_file_inst1_r6_17_), .A2(n5004), .B1(
        register_file_inst1_r7_17_), .B2(n4991), .ZN(n4479) );
  ND4D1BWP12T U3569 ( .A1(n4482), .A2(n4481), .A3(n4480), .A4(n4479), .ZN(
        n4487) );
  AOI22D1BWP12T U3570 ( .A1(register_file_inst1_lr_17_), .A2(n4437), .B1(
        register_file_inst1_r12_17_), .B2(n4510), .ZN(n4485) );
  AOI22D1BWP12T U3571 ( .A1(RF_next_sp[17]), .A2(n5010), .B1(
        register_file_inst1_r11_17_), .B2(n5009), .ZN(n4484) );
  AOI22D0BWP12T U3572 ( .A1(register_file_inst1_r9_17_), .A2(n6005), .B1(
        register_file_inst1_r10_17_), .B2(n5011), .ZN(n4483) );
  ND4D1BWP12T U3573 ( .A1(n6247), .A2(n4485), .A3(n4484), .A4(n4483), .ZN(
        n4486) );
  AO21D1BWP12T U3574 ( .A1(n3502), .A2(n4487), .B(n4486), .Z(
        RF_MEMCTRL_data_reg[17]) );
  AOI22D0BWP12T U3575 ( .A1(register_file_inst1_r1_5_), .A2(n5001), .B1(
        register_file_inst1_r3_5_), .B2(n4989), .ZN(n4491) );
  AOI22D0BWP12T U3576 ( .A1(register_file_inst1_r2_5_), .A2(n4962), .B1(
        register_file_inst1_r0_5_), .B2(n5002), .ZN(n4490) );
  AOI22D0BWP12T U3577 ( .A1(register_file_inst1_r4_5_), .A2(n5003), .B1(
        register_file_inst1_r5_5_), .B2(n4990), .ZN(n4489) );
  AOI22D0BWP12T U3578 ( .A1(register_file_inst1_r6_5_), .A2(n5004), .B1(
        register_file_inst1_r7_5_), .B2(n4991), .ZN(n4488) );
  ND4D1BWP12T U3579 ( .A1(n4491), .A2(n4490), .A3(n4489), .A4(n4488), .ZN(
        n4496) );
  AOI22D1BWP12T U3580 ( .A1(register_file_inst1_lr_5_), .A2(n4437), .B1(
        register_file_inst1_r12_5_), .B2(n4510), .ZN(n4494) );
  AOI22D1BWP12T U3581 ( .A1(register_file_inst1_r11_5_), .A2(n5009), .B1(
        RF_next_sp[5]), .B2(n5010), .ZN(n4493) );
  AOI22D1BWP12T U3582 ( .A1(register_file_inst1_r9_5_), .A2(n6005), .B1(
        register_file_inst1_r10_5_), .B2(n5011), .ZN(n4492) );
  ND4D1BWP12T U3583 ( .A1(n6263), .A2(n4494), .A3(n4493), .A4(n4492), .ZN(
        n4495) );
  AO21D1BWP12T U3584 ( .A1(n3502), .A2(n4496), .B(n4495), .Z(
        RF_MEMCTRL_data_reg[5]) );
  AOI22D0BWP12T U3585 ( .A1(register_file_inst1_r1_21_), .A2(n5001), .B1(
        register_file_inst1_r3_21_), .B2(n4989), .ZN(n4500) );
  AOI22D0BWP12T U3586 ( .A1(register_file_inst1_r2_21_), .A2(n4962), .B1(
        register_file_inst1_r0_21_), .B2(n5002), .ZN(n4499) );
  AOI22D0BWP12T U3587 ( .A1(register_file_inst1_r4_21_), .A2(n5003), .B1(
        register_file_inst1_r5_21_), .B2(n4990), .ZN(n4498) );
  AOI22D0BWP12T U3588 ( .A1(register_file_inst1_r6_21_), .A2(n5004), .B1(
        register_file_inst1_r7_21_), .B2(n4991), .ZN(n4497) );
  ND4D1BWP12T U3589 ( .A1(n4500), .A2(n4499), .A3(n4498), .A4(n4497), .ZN(
        n4505) );
  AOI22D0BWP12T U3590 ( .A1(register_file_inst1_lr_21_), .A2(n4437), .B1(
        register_file_inst1_r12_21_), .B2(n4510), .ZN(n4503) );
  AOI22D1BWP12T U3591 ( .A1(RF_next_sp[21]), .A2(n5010), .B1(
        register_file_inst1_r11_21_), .B2(n5009), .ZN(n4502) );
  AOI22D0BWP12T U3592 ( .A1(register_file_inst1_r9_21_), .A2(n6005), .B1(
        register_file_inst1_r10_21_), .B2(n5011), .ZN(n4501) );
  ND4D1BWP12T U3593 ( .A1(n6262), .A2(n4503), .A3(n4502), .A4(n4501), .ZN(
        n4504) );
  AO21D1BWP12T U3594 ( .A1(n3502), .A2(n4505), .B(n4504), .Z(
        RF_MEMCTRL_data_reg[21]) );
  AOI22D1BWP12T U3595 ( .A1(register_file_inst1_r1_7_), .A2(n5001), .B1(
        register_file_inst1_r3_7_), .B2(n4989), .ZN(n4509) );
  AOI22D0BWP12T U3596 ( .A1(register_file_inst1_r2_7_), .A2(n4962), .B1(
        register_file_inst1_r0_7_), .B2(n5002), .ZN(n4508) );
  AOI22D0BWP12T U3597 ( .A1(register_file_inst1_r4_7_), .A2(n5003), .B1(
        register_file_inst1_r5_7_), .B2(n4990), .ZN(n4507) );
  AOI22D0BWP12T U3598 ( .A1(register_file_inst1_r6_7_), .A2(n5004), .B1(
        register_file_inst1_r7_7_), .B2(n4991), .ZN(n4506) );
  ND4D1BWP12T U3599 ( .A1(n4509), .A2(n4508), .A3(n4507), .A4(n4506), .ZN(
        n4515) );
  AOI22D1BWP12T U3600 ( .A1(register_file_inst1_lr_7_), .A2(n4437), .B1(
        register_file_inst1_r12_7_), .B2(n4510), .ZN(n4513) );
  AOI22D1BWP12T U3601 ( .A1(register_file_inst1_r11_7_), .A2(n5009), .B1(
        RF_next_sp[7]), .B2(n5010), .ZN(n4512) );
  AOI22D1BWP12T U3602 ( .A1(register_file_inst1_r9_7_), .A2(n6005), .B1(
        register_file_inst1_r10_7_), .B2(n5011), .ZN(n4511) );
  ND4D1BWP12T U3603 ( .A1(n6280), .A2(n4513), .A3(n4512), .A4(n4511), .ZN(
        n4514) );
  AO21D1BWP12T U3604 ( .A1(n3502), .A2(n4515), .B(n4514), .Z(
        RF_MEMCTRL_data_reg[7]) );
  AOI22D0BWP12T U3605 ( .A1(register_file_inst1_r1_23_), .A2(n5001), .B1(
        register_file_inst1_r3_23_), .B2(n4989), .ZN(n4519) );
  AOI22D0BWP12T U3606 ( .A1(register_file_inst1_r2_23_), .A2(n4962), .B1(
        register_file_inst1_r0_23_), .B2(n5002), .ZN(n4518) );
  AOI22D0BWP12T U3607 ( .A1(register_file_inst1_r4_23_), .A2(n5003), .B1(
        register_file_inst1_r5_23_), .B2(n4990), .ZN(n4517) );
  AOI22D0BWP12T U3608 ( .A1(register_file_inst1_r6_23_), .A2(n5004), .B1(
        register_file_inst1_r7_23_), .B2(n4991), .ZN(n4516) );
  ND4D1BWP12T U3609 ( .A1(n4519), .A2(n4518), .A3(n4517), .A4(n4516), .ZN(
        n4524) );
  AOI22D1BWP12T U3610 ( .A1(register_file_inst1_lr_23_), .A2(n4437), .B1(
        register_file_inst1_r12_23_), .B2(n4510), .ZN(n4522) );
  AOI22D1BWP12T U3611 ( .A1(RF_next_sp[23]), .A2(n5010), .B1(
        register_file_inst1_r11_23_), .B2(n5009), .ZN(n4521) );
  AOI22D0BWP12T U3612 ( .A1(register_file_inst1_r9_23_), .A2(n6005), .B1(
        register_file_inst1_r10_23_), .B2(n5011), .ZN(n4520) );
  ND4D1BWP12T U3613 ( .A1(n6279), .A2(n4522), .A3(n4521), .A4(n4520), .ZN(
        n4523) );
  AO21D1BWP12T U3614 ( .A1(n3502), .A2(n4524), .B(n4523), .Z(
        RF_MEMCTRL_data_reg[23]) );
  AOI22D0BWP12T U3615 ( .A1(register_file_inst1_r1_2_), .A2(n5001), .B1(
        register_file_inst1_r3_2_), .B2(n4989), .ZN(n4528) );
  AOI22D0BWP12T U3616 ( .A1(register_file_inst1_r2_2_), .A2(n4962), .B1(
        register_file_inst1_r0_2_), .B2(n5002), .ZN(n4527) );
  AOI22D0BWP12T U3617 ( .A1(register_file_inst1_r4_2_), .A2(n5003), .B1(
        register_file_inst1_r5_2_), .B2(n4990), .ZN(n4526) );
  AOI22D0BWP12T U3618 ( .A1(register_file_inst1_r6_2_), .A2(n5004), .B1(
        register_file_inst1_r7_2_), .B2(n4991), .ZN(n4525) );
  ND4D1BWP12T U3619 ( .A1(n4528), .A2(n4527), .A3(n4526), .A4(n4525), .ZN(
        n4533) );
  AOI22D1BWP12T U3620 ( .A1(register_file_inst1_lr_2_), .A2(n4437), .B1(
        register_file_inst1_r12_2_), .B2(n4510), .ZN(n4531) );
  AOI22D1BWP12T U3621 ( .A1(register_file_inst1_r11_2_), .A2(n5009), .B1(
        RF_next_sp[2]), .B2(n5010), .ZN(n4530) );
  AOI22D0BWP12T U3622 ( .A1(register_file_inst1_r9_2_), .A2(n6005), .B1(
        register_file_inst1_r10_2_), .B2(n5011), .ZN(n4529) );
  ND4D1BWP12T U3623 ( .A1(n6272), .A2(n4531), .A3(n4530), .A4(n4529), .ZN(
        n4532) );
  AO21D1BWP12T U3624 ( .A1(n3502), .A2(n4533), .B(n4532), .Z(
        RF_MEMCTRL_data_reg[2]) );
  AOI22D0BWP12T U3625 ( .A1(register_file_inst1_r1_18_), .A2(n5001), .B1(
        register_file_inst1_r3_18_), .B2(n4989), .ZN(n4537) );
  AOI22D0BWP12T U3626 ( .A1(register_file_inst1_r2_18_), .A2(n4962), .B1(
        register_file_inst1_r0_18_), .B2(n5002), .ZN(n4536) );
  AOI22D0BWP12T U3627 ( .A1(register_file_inst1_r4_18_), .A2(n5003), .B1(
        register_file_inst1_r5_18_), .B2(n4990), .ZN(n4535) );
  AOI22D0BWP12T U3628 ( .A1(register_file_inst1_r6_18_), .A2(n5004), .B1(
        register_file_inst1_r7_18_), .B2(n4991), .ZN(n4534) );
  ND4D1BWP12T U3629 ( .A1(n4537), .A2(n4536), .A3(n4535), .A4(n4534), .ZN(
        n4542) );
  AOI22D1BWP12T U3630 ( .A1(register_file_inst1_lr_18_), .A2(n4437), .B1(
        register_file_inst1_r12_18_), .B2(n4510), .ZN(n4540) );
  AOI22D1BWP12T U3631 ( .A1(RF_next_sp[18]), .A2(n5010), .B1(
        register_file_inst1_r11_18_), .B2(n5009), .ZN(n4539) );
  AOI22D1BWP12T U3632 ( .A1(register_file_inst1_r9_18_), .A2(n6005), .B1(
        register_file_inst1_r10_18_), .B2(n5011), .ZN(n4538) );
  ND4D1BWP12T U3633 ( .A1(n6271), .A2(n4540), .A3(n4539), .A4(n4538), .ZN(
        n4541) );
  AO21D1BWP12T U3634 ( .A1(n3502), .A2(n4542), .B(n4541), .Z(
        RF_MEMCTRL_data_reg[18]) );
  AOI22D1BWP12T U3635 ( .A1(register_file_inst1_r1_0_), .A2(n5001), .B1(
        register_file_inst1_r3_0_), .B2(n4989), .ZN(n4546) );
  AOI22D1BWP12T U3636 ( .A1(register_file_inst1_r2_0_), .A2(n4962), .B1(
        register_file_inst1_r0_0_), .B2(n5002), .ZN(n4545) );
  AOI22D1BWP12T U3637 ( .A1(register_file_inst1_r4_0_), .A2(n5003), .B1(
        register_file_inst1_r5_0_), .B2(n4990), .ZN(n4544) );
  AOI22D1BWP12T U3638 ( .A1(register_file_inst1_r6_0_), .A2(n5004), .B1(
        register_file_inst1_r7_0_), .B2(n4991), .ZN(n4543) );
  ND4D1BWP12T U3639 ( .A1(n4546), .A2(n4545), .A3(n4544), .A4(n4543), .ZN(
        n4552) );
  OR2XD1BWP12T U3640 ( .A1(n2917), .A2(n4547), .Z(n4674) );
  AOI22D1BWP12T U3641 ( .A1(register_file_inst1_lr_0_), .A2(n4437), .B1(
        register_file_inst1_r8_0_), .B2(n5980), .ZN(n4550) );
  AOI22D1BWP12T U3642 ( .A1(RF_next_sp[0]), .A2(n5010), .B1(
        register_file_inst1_r12_0_), .B2(n4510), .ZN(n4549) );
  AOI22D1BWP12T U3643 ( .A1(register_file_inst1_r10_0_), .A2(n5011), .B1(
        register_file_inst1_r11_0_), .B2(n5009), .ZN(n4548) );
  ND4D1BWP12T U3644 ( .A1(n4550), .A2(n6243), .A3(n4549), .A4(n4548), .ZN(
        n4551) );
  AO21D1BWP12T U3645 ( .A1(n3502), .A2(n4552), .B(n4551), .Z(
        RF_MEMCTRL_data_reg[0]) );
  AOI22D1BWP12T U3646 ( .A1(register_file_inst1_r1_16_), .A2(n5001), .B1(
        register_file_inst1_r3_16_), .B2(n4989), .ZN(n4556) );
  AOI22D0BWP12T U3647 ( .A1(register_file_inst1_r2_16_), .A2(n4962), .B1(
        register_file_inst1_r0_16_), .B2(n5002), .ZN(n4555) );
  AOI22D1BWP12T U3648 ( .A1(register_file_inst1_r4_16_), .A2(n5003), .B1(
        register_file_inst1_r5_16_), .B2(n4990), .ZN(n4554) );
  AOI22D0BWP12T U3649 ( .A1(register_file_inst1_r6_16_), .A2(n5004), .B1(
        register_file_inst1_r7_16_), .B2(n4991), .ZN(n4553) );
  ND4D1BWP12T U3650 ( .A1(n4556), .A2(n4555), .A3(n4554), .A4(n4553), .ZN(
        n4561) );
  AOI22D1BWP12T U3651 ( .A1(register_file_inst1_lr_16_), .A2(n4437), .B1(
        register_file_inst1_r12_16_), .B2(n4510), .ZN(n4559) );
  AOI22D1BWP12T U3652 ( .A1(RF_next_sp[16]), .A2(n5010), .B1(
        register_file_inst1_r11_16_), .B2(n5009), .ZN(n4558) );
  AOI22D1BWP12T U3653 ( .A1(register_file_inst1_r9_16_), .A2(n6005), .B1(
        register_file_inst1_r10_16_), .B2(n5011), .ZN(n4557) );
  ND4D1BWP12T U3654 ( .A1(n6242), .A2(n4559), .A3(n4558), .A4(n4557), .ZN(
        n4560) );
  AO21D1BWP12T U3655 ( .A1(n3502), .A2(n4561), .B(n4560), .Z(
        RF_MEMCTRL_data_reg[16]) );
  AOI22D1BWP12T U3656 ( .A1(register_file_inst1_r1_3_), .A2(n5001), .B1(
        register_file_inst1_r3_3_), .B2(n4989), .ZN(n4565) );
  AOI22D0BWP12T U3657 ( .A1(register_file_inst1_r2_3_), .A2(n4962), .B1(
        register_file_inst1_r0_3_), .B2(n5002), .ZN(n4564) );
  AOI22D1BWP12T U3658 ( .A1(register_file_inst1_r4_3_), .A2(n5003), .B1(
        register_file_inst1_r5_3_), .B2(n4990), .ZN(n4563) );
  AOI22D1BWP12T U3659 ( .A1(register_file_inst1_r6_3_), .A2(n5004), .B1(
        register_file_inst1_r7_3_), .B2(n4991), .ZN(n4562) );
  ND4D1BWP12T U3660 ( .A1(n4565), .A2(n4564), .A3(n4563), .A4(n4562), .ZN(
        n4570) );
  AOI22D1BWP12T U3661 ( .A1(register_file_inst1_lr_3_), .A2(n4437), .B1(
        register_file_inst1_r12_3_), .B2(n4510), .ZN(n4568) );
  AOI22D1BWP12T U3662 ( .A1(register_file_inst1_r11_3_), .A2(n5009), .B1(
        RF_next_sp[3]), .B2(n5010), .ZN(n4567) );
  AOI22D1BWP12T U3663 ( .A1(register_file_inst1_r9_3_), .A2(n6005), .B1(
        register_file_inst1_r10_3_), .B2(n5011), .ZN(n4566) );
  ND4D1BWP12T U3664 ( .A1(n6241), .A2(n4568), .A3(n4567), .A4(n4566), .ZN(
        n4569) );
  AO21D1BWP12T U3665 ( .A1(n3502), .A2(n4570), .B(n4569), .Z(
        RF_MEMCTRL_data_reg[3]) );
  AOI22D1BWP12T U3666 ( .A1(register_file_inst1_r1_19_), .A2(n5001), .B1(
        register_file_inst1_r3_19_), .B2(n4989), .ZN(n4574) );
  AOI22D0BWP12T U3667 ( .A1(register_file_inst1_r2_19_), .A2(n4962), .B1(
        register_file_inst1_r0_19_), .B2(n5002), .ZN(n4573) );
  AOI22D0BWP12T U3668 ( .A1(register_file_inst1_r4_19_), .A2(n5003), .B1(
        register_file_inst1_r5_19_), .B2(n4990), .ZN(n4572) );
  AOI22D0BWP12T U3669 ( .A1(register_file_inst1_r6_19_), .A2(n5004), .B1(
        register_file_inst1_r7_19_), .B2(n4991), .ZN(n4571) );
  ND4D1BWP12T U3670 ( .A1(n4574), .A2(n4573), .A3(n4572), .A4(n4571), .ZN(
        n4579) );
  AOI22D1BWP12T U3671 ( .A1(register_file_inst1_lr_19_), .A2(n4437), .B1(
        register_file_inst1_r12_19_), .B2(n4510), .ZN(n4577) );
  AOI22D1BWP12T U3672 ( .A1(RF_next_sp[19]), .A2(n5010), .B1(
        register_file_inst1_r11_19_), .B2(n5009), .ZN(n4576) );
  AOI22D1BWP12T U3673 ( .A1(register_file_inst1_r9_19_), .A2(n6005), .B1(
        register_file_inst1_r10_19_), .B2(n5011), .ZN(n4575) );
  ND4D1BWP12T U3674 ( .A1(n6240), .A2(n4577), .A3(n4576), .A4(n4575), .ZN(
        n4578) );
  AO21D1BWP12T U3675 ( .A1(n3502), .A2(n4579), .B(n4578), .Z(
        RF_MEMCTRL_data_reg[19]) );
  AOI22D1BWP12T U3676 ( .A1(register_file_inst1_r1_6_), .A2(n5001), .B1(
        register_file_inst1_r3_6_), .B2(n4989), .ZN(n4583) );
  AOI22D0BWP12T U3677 ( .A1(register_file_inst1_r2_6_), .A2(n4962), .B1(
        register_file_inst1_r0_6_), .B2(n5002), .ZN(n4582) );
  AOI22D1BWP12T U3678 ( .A1(register_file_inst1_r4_6_), .A2(n5003), .B1(
        register_file_inst1_r5_6_), .B2(n4990), .ZN(n4581) );
  AOI22D0BWP12T U3679 ( .A1(register_file_inst1_r6_6_), .A2(n5004), .B1(
        register_file_inst1_r7_6_), .B2(n4991), .ZN(n4580) );
  ND4D1BWP12T U3680 ( .A1(n4583), .A2(n4582), .A3(n4581), .A4(n4580), .ZN(
        n4588) );
  AOI22D1BWP12T U3681 ( .A1(register_file_inst1_lr_6_), .A2(n4437), .B1(
        register_file_inst1_r12_6_), .B2(n4510), .ZN(n4586) );
  AOI22D1BWP12T U3682 ( .A1(register_file_inst1_r11_6_), .A2(n5009), .B1(
        RF_next_sp[6]), .B2(n5010), .ZN(n4585) );
  AOI22D1BWP12T U3683 ( .A1(register_file_inst1_r9_6_), .A2(n6005), .B1(
        register_file_inst1_r10_6_), .B2(n5011), .ZN(n4584) );
  ND4D1BWP12T U3684 ( .A1(n6245), .A2(n4586), .A3(n4585), .A4(n4584), .ZN(
        n4587) );
  AO21D1BWP12T U3685 ( .A1(n3502), .A2(n4588), .B(n4587), .Z(
        RF_MEMCTRL_data_reg[6]) );
  AOI22D0BWP12T U3686 ( .A1(register_file_inst1_r1_22_), .A2(n5001), .B1(
        register_file_inst1_r3_22_), .B2(n4989), .ZN(n4592) );
  AOI22D0BWP12T U3687 ( .A1(register_file_inst1_r2_22_), .A2(n4962), .B1(
        register_file_inst1_r0_22_), .B2(n5002), .ZN(n4591) );
  AOI22D0BWP12T U3688 ( .A1(register_file_inst1_r4_22_), .A2(n5003), .B1(
        register_file_inst1_r5_22_), .B2(n4990), .ZN(n4590) );
  AOI22D0BWP12T U3689 ( .A1(register_file_inst1_r6_22_), .A2(n5004), .B1(
        register_file_inst1_r7_22_), .B2(n4991), .ZN(n4589) );
  ND4D1BWP12T U3690 ( .A1(n4592), .A2(n4591), .A3(n4590), .A4(n4589), .ZN(
        n4597) );
  AOI22D1BWP12T U3691 ( .A1(register_file_inst1_lr_22_), .A2(n4437), .B1(
        register_file_inst1_r12_22_), .B2(n4510), .ZN(n4595) );
  AOI22D1BWP12T U3692 ( .A1(RF_next_sp[22]), .A2(n5010), .B1(
        register_file_inst1_r11_22_), .B2(n5009), .ZN(n4594) );
  AOI22D0BWP12T U3693 ( .A1(register_file_inst1_r9_22_), .A2(n6005), .B1(
        register_file_inst1_r10_22_), .B2(n5011), .ZN(n4593) );
  ND4D1BWP12T U3694 ( .A1(n6244), .A2(n4595), .A3(n4594), .A4(n4593), .ZN(
        n4596) );
  AO21D1BWP12T U3695 ( .A1(n3502), .A2(n4597), .B(n4596), .Z(
        RF_MEMCTRL_data_reg[22]) );
  AOI22D0BWP12T U3696 ( .A1(register_file_inst1_r1_4_), .A2(n5001), .B1(
        register_file_inst1_r3_4_), .B2(n4989), .ZN(n4601) );
  AOI22D0BWP12T U3697 ( .A1(register_file_inst1_r2_4_), .A2(n4962), .B1(
        register_file_inst1_r0_4_), .B2(n5002), .ZN(n4600) );
  AOI22D0BWP12T U3698 ( .A1(register_file_inst1_r4_4_), .A2(n5003), .B1(
        register_file_inst1_r5_4_), .B2(n4990), .ZN(n4599) );
  AOI22D0BWP12T U3699 ( .A1(register_file_inst1_r6_4_), .A2(n5004), .B1(
        register_file_inst1_r7_4_), .B2(n4991), .ZN(n4598) );
  ND4D1BWP12T U3700 ( .A1(n4601), .A2(n4600), .A3(n4599), .A4(n4598), .ZN(
        n4606) );
  AOI22D1BWP12T U3701 ( .A1(register_file_inst1_lr_4_), .A2(n4437), .B1(
        register_file_inst1_r12_4_), .B2(n4510), .ZN(n4604) );
  AOI22D1BWP12T U3702 ( .A1(register_file_inst1_r11_4_), .A2(n5009), .B1(
        RF_next_sp[4]), .B2(n5010), .ZN(n4603) );
  AOI22D0BWP12T U3703 ( .A1(register_file_inst1_r9_4_), .A2(n6005), .B1(
        register_file_inst1_r10_4_), .B2(n5011), .ZN(n4602) );
  ND4D1BWP12T U3704 ( .A1(n6270), .A2(n4604), .A3(n4603), .A4(n4602), .ZN(
        n4605) );
  AO21D1BWP12T U3705 ( .A1(n3502), .A2(n4606), .B(n4605), .Z(
        RF_MEMCTRL_data_reg[4]) );
  AOI22D1BWP12T U3706 ( .A1(register_file_inst1_r1_20_), .A2(n5001), .B1(
        register_file_inst1_r3_20_), .B2(n4989), .ZN(n4610) );
  AOI22D0BWP12T U3707 ( .A1(register_file_inst1_r2_20_), .A2(n4962), .B1(
        register_file_inst1_r0_20_), .B2(n5002), .ZN(n4609) );
  AOI22D1BWP12T U3708 ( .A1(register_file_inst1_r4_20_), .A2(n5003), .B1(
        register_file_inst1_r5_20_), .B2(n4990), .ZN(n4608) );
  AOI22D0BWP12T U3709 ( .A1(register_file_inst1_r6_20_), .A2(n5004), .B1(
        register_file_inst1_r7_20_), .B2(n4991), .ZN(n4607) );
  ND4D1BWP12T U3710 ( .A1(n4610), .A2(n4609), .A3(n4608), .A4(n4607), .ZN(
        n4615) );
  AOI22D1BWP12T U3711 ( .A1(register_file_inst1_lr_20_), .A2(n4437), .B1(
        register_file_inst1_r12_20_), .B2(n4510), .ZN(n4613) );
  AOI22D1BWP12T U3712 ( .A1(RF_next_sp[20]), .A2(n5010), .B1(
        register_file_inst1_r11_20_), .B2(n5009), .ZN(n4612) );
  AOI22D1BWP12T U3713 ( .A1(register_file_inst1_r9_20_), .A2(n6005), .B1(
        register_file_inst1_r10_20_), .B2(n5011), .ZN(n4611) );
  ND4D1BWP12T U3714 ( .A1(n6269), .A2(n4613), .A3(n4612), .A4(n4611), .ZN(
        n4614) );
  AO21D1BWP12T U3715 ( .A1(n3502), .A2(n4615), .B(n4614), .Z(
        RF_MEMCTRL_data_reg[20]) );
  BUFFD1BWP12T U3716 ( .I(n6394), .Z(n6007) );
  ND2D1BWP12T U3717 ( .A1(n2515), .A2(n6044), .ZN(n4627) );
  NR2D2BWP12T U3718 ( .A1(n6047), .A2(n4627), .ZN(n5963) );
  AOI22D1BWP12T U3719 ( .A1(RF_next_sp[0]), .A2(n5964), .B1(
        register_file_inst1_r12_0_), .B2(n5963), .ZN(n4616) );
  ND2D1BWP12T U3720 ( .A1(n4616), .A2(n6037), .ZN(n4625) );
  NR2D2BWP12T U3721 ( .A1(n6051), .A2(n6038), .ZN(n5996) );
  INVD1BWP12T U3722 ( .I(n5996), .ZN(n4767) );
  INVD1BWP12T U3723 ( .I(register_file_inst1_tmp1_0_), .ZN(n5018) );
  OAI22D1BWP12T U3724 ( .A1(n6040), .A2(n4767), .B1(n5018), .B2(n5981), .ZN(
        n4624) );
  ND2D1BWP12T U3725 ( .A1(n6042), .A2(n6044), .ZN(n4677) );
  INVD1BWP12T U3726 ( .I(n4677), .ZN(n4619) );
  ND2D1BWP12T U3727 ( .A1(n4619), .A2(n6043), .ZN(n5912) );
  INVD0BWP12T U3728 ( .I(n6046), .ZN(n4617) );
  ND2D1BWP12T U3729 ( .A1(n4617), .A2(n6043), .ZN(n5857) );
  INVD1BWP12T U3730 ( .I(n5857), .ZN(n5822) );
  INVD1BWP12T U3731 ( .I(n6045), .ZN(n4620) );
  ND2D1BWP12T U3732 ( .A1(n4620), .A2(n4619), .ZN(n5959) );
  INVD1BWP12T U3733 ( .I(n5959), .ZN(n5825) );
  ND2D1BWP12T U3734 ( .A1(n2516), .A2(n6044), .ZN(n4626) );
  NR2D1BWP12T U3735 ( .A1(n6047), .A2(n4626), .ZN(n5961) );
  INVD1BWP12T U3736 ( .I(n5961), .ZN(n5805) );
  NR4D0BWP12T U3737 ( .A1(n4625), .A2(n4624), .A3(n4623), .A4(n4622), .ZN(
        n4633) );
  ND2D1BWP12T U3738 ( .A1(n2515), .A2(n6036), .ZN(n4678) );
  AOI22D1BWP12T U3739 ( .A1(register_file_inst1_r9_0_), .A2(n5968), .B1(
        register_file_inst1_r3_0_), .B2(n5967), .ZN(n4631) );
  AOI22D1BWP12T U3740 ( .A1(register_file_inst1_r7_0_), .A2(n6001), .B1(
        register_file_inst1_r11_0_), .B2(n5969), .ZN(n4630) );
  NR2D2BWP12T U3741 ( .A1(n6048), .A2(n6047), .ZN(n6002) );
  AOI22D1BWP12T U3742 ( .A1(register_file_inst1_r5_0_), .A2(n6002), .B1(
        register_file_inst1_r10_0_), .B2(n5995), .ZN(n4629) );
  INVD1BWP12T U3743 ( .I(n6051), .ZN(n6050) );
  INVD1BWP12T U3744 ( .I(n5910), .ZN(n5823) );
  NR2D1BWP12T U3745 ( .A1(n6051), .A2(n4627), .ZN(n5970) );
  INVD1BWP12T U3746 ( .I(n5970), .ZN(n5653) );
  AOI22D1BWP12T U3747 ( .A1(register_file_inst1_r6_0_), .A2(n5823), .B1(
        register_file_inst1_lr_0_), .B2(n5970), .ZN(n4628) );
  AN4XD1BWP12T U3748 ( .A1(n4631), .A2(n4630), .A3(n4629), .A4(n4628), .Z(
        n4632) );
  CKND2D1BWP12T U3749 ( .A1(n4633), .A2(n4632), .ZN(RF_ALU_operand_b[0]) );
  AOI21D1BWP12T U3750 ( .A1(n6297), .A2(n6296), .B(n6008), .ZN(n6386) );
  CKND0BWP12T U3751 ( .I(n6386), .ZN(n6298) );
  TPNR2D0BWP12T U3752 ( .A1(n6364), .A2(n5233), .ZN(n6078) );
  ND2D1BWP12T U3753 ( .A1(n2470), .A2(n6402), .ZN(n4676) );
  ND2D1BWP12T U3754 ( .A1(n6147), .A2(n6150), .ZN(n4640) );
  AOI22D1BWP12T U3755 ( .A1(register_file_inst1_r0_10_), .A2(n6004), .B1(
        register_file_inst1_r6_10_), .B2(n6003), .ZN(n4636) );
  AOI22D1BWP12T U3756 ( .A1(register_file_inst1_r11_10_), .A2(n6229), .B1(
        register_file_inst1_r3_10_), .B2(n5946), .ZN(n4635) );
  INVD1BWP12T U3757 ( .I(n6155), .ZN(n4637) );
  NR2D1BWP12T U3758 ( .A1(n4637), .A2(n6157), .ZN(n5948) );
  AOI22D1BWP12T U3759 ( .A1(register_file_inst1_r5_10_), .A2(n5948), .B1(
        register_file_inst1_r8_10_), .B2(n5947), .ZN(n4634) );
  AN4XD1BWP12T U3760 ( .A1(n4636), .A2(n6180), .A3(n4635), .A4(n4634), .Z(
        n4646) );
  BUFFD2BWP12T U3761 ( .I(n6224), .Z(n5979) );
  INVD1BWP12T U3762 ( .I(n6223), .ZN(n5844) );
  AOI22D1BWP12T U3763 ( .A1(register_file_inst1_tmp1_10_), .A2(n5979), .B1(
        register_file_inst1_r10_10_), .B2(n6223), .ZN(n4639) );
  NR2D1BWP12T U3764 ( .A1(n4676), .A2(n4637), .ZN(n5900) );
  AOI22D1BWP12T U3765 ( .A1(register_file_inst1_r4_10_), .A2(n5900), .B1(
        register_file_inst1_r9_10_), .B2(n6225), .ZN(n4638) );
  AN3XD1BWP12T U3766 ( .A1(n4639), .A2(n4638), .A3(n6181), .Z(n4645) );
  INVD1BWP12T U3767 ( .I(n6154), .ZN(n6159) );
  INVD1BWP12T U3768 ( .I(n6157), .ZN(n4641) );
  ND2D1BWP12T U3769 ( .A1(n6159), .A2(n4641), .ZN(n5938) );
  INVD1BWP12T U3770 ( .I(n5938), .ZN(n5848) );
  INVD1BWP12T U3771 ( .I(n6222), .ZN(n5835) );
  AOI22D1BWP12T U3772 ( .A1(register_file_inst1_r7_10_), .A2(n5848), .B1(
        RF_next_sp[10]), .B2(n5835), .ZN(n4644) );
  INVD1BWP12T U3773 ( .I(n4640), .ZN(n4642) );
  ND2D1BWP12T U3774 ( .A1(n4642), .A2(n4641), .ZN(n5942) );
  INVD1BWP12T U3775 ( .I(n5942), .ZN(n5837) );
  INVD1BWP12T U3776 ( .I(n5940), .ZN(n5836) );
  AOI22D1BWP12T U3777 ( .A1(register_file_inst1_r1_10_), .A2(n5837), .B1(
        register_file_inst1_lr_10_), .B2(n5836), .ZN(n4643) );
  ND4D1BWP12T U3778 ( .A1(n4646), .A2(n4645), .A3(n4644), .A4(n4643), .ZN(
        RF_ALU_operand_a[10]) );
  CKND0BWP12T U3779 ( .I(n5143), .ZN(n5990) );
  OAI22D1BWP12T U3780 ( .A1(n4647), .A2(n5910), .B1(n5514), .B2(n5857), .ZN(
        n4658) );
  INVD1BWP12T U3781 ( .I(n5912), .ZN(n5824) );
  OAI22D1BWP12T U3782 ( .A1(n4649), .A2(n5959), .B1(n4648), .B2(n5912), .ZN(
        n4657) );
  AOI22D1BWP12T U3783 ( .A1(register_file_inst1_tmp1_17_), .A2(n5962), .B1(
        register_file_inst1_r4_17_), .B2(n5961), .ZN(n4651) );
  AOI22D1BWP12T U3784 ( .A1(RF_next_sp[17]), .A2(n5964), .B1(
        register_file_inst1_r12_17_), .B2(n5963), .ZN(n4650) );
  ND3D1BWP12T U3785 ( .A1(n4651), .A2(n4650), .A3(n6116), .ZN(n4656) );
  AOI22D1BWP12T U3786 ( .A1(register_file_inst1_r9_17_), .A2(n5968), .B1(
        register_file_inst1_r3_17_), .B2(n5967), .ZN(n4654) );
  AOI22D1BWP12T U3787 ( .A1(register_file_inst1_r7_17_), .A2(n6001), .B1(
        register_file_inst1_r11_17_), .B2(n5969), .ZN(n4653) );
  AOI22D1BWP12T U3788 ( .A1(register_file_inst1_r5_17_), .A2(n6002), .B1(
        register_file_inst1_lr_17_), .B2(n5970), .ZN(n4652) );
  ND4D1BWP12T U3789 ( .A1(n4654), .A2(n4653), .A3(n6117), .A4(n4652), .ZN(
        n4655) );
  OR4D4BWP12T U3790 ( .A1(n4658), .A2(n4657), .A3(n4656), .A4(n4655), .Z(
        RF_ALU_operand_b[17]) );
  AOI22D1BWP12T U3791 ( .A1(register_file_inst1_r0_2_), .A2(n6004), .B1(
        register_file_inst1_r6_2_), .B2(n6003), .ZN(n4661) );
  AOI22D1BWP12T U3792 ( .A1(register_file_inst1_r11_2_), .A2(n6229), .B1(
        register_file_inst1_r3_2_), .B2(n5946), .ZN(n4660) );
  AOI22D1BWP12T U3793 ( .A1(register_file_inst1_r5_2_), .A2(n5948), .B1(
        register_file_inst1_r8_2_), .B2(n5947), .ZN(n4659) );
  AN4XD1BWP12T U3794 ( .A1(n4661), .A2(n6164), .A3(n4660), .A4(n4659), .Z(
        n4667) );
  AOI22D1BWP12T U3795 ( .A1(register_file_inst1_tmp1_2_), .A2(n5979), .B1(
        register_file_inst1_r10_2_), .B2(n6223), .ZN(n4663) );
  AOI22D1BWP12T U3796 ( .A1(register_file_inst1_r4_2_), .A2(n5900), .B1(
        register_file_inst1_r9_2_), .B2(n6225), .ZN(n4662) );
  AN3XD2BWP12T U3797 ( .A1(n4663), .A2(n4662), .A3(n6165), .Z(n4666) );
  AOI22D1BWP12T U3798 ( .A1(register_file_inst1_r7_2_), .A2(n5848), .B1(
        RF_next_sp[2]), .B2(n5835), .ZN(n4665) );
  AOI22D1BWP12T U3799 ( .A1(register_file_inst1_r1_2_), .A2(n5837), .B1(
        register_file_inst1_lr_2_), .B2(n5836), .ZN(n4664) );
  CKND0BWP12T U3800 ( .I(n5074), .ZN(n5987) );
  CKND0BWP12T U3801 ( .I(n5145), .ZN(n5988) );
  CKND0BWP12T U3802 ( .I(n5140), .ZN(n5986) );
  CKND0BWP12T U3803 ( .I(n5238), .ZN(n5989) );
  INVD1BWP12T U3804 ( .I(register_file_inst1_r12_30_), .ZN(n5207) );
  INVD1BWP12T U3805 ( .I(register_file_inst1_r11_30_), .ZN(n5211) );
  OAI22D0BWP12T U3806 ( .A1(n4673), .A2(n5207), .B1(n5211), .B2(n4672), .ZN(
        n6257) );
  CKND0BWP12T U3807 ( .I(register_file_inst1_r12_24_), .ZN(n5139) );
  OAI22D0BWP12T U3808 ( .A1(n4673), .A2(n5139), .B1(n4668), .B2(n4672), .ZN(
        n6275) );
  INVD0BWP12T U3809 ( .I(register_file_inst1_r12_28_), .ZN(n5187) );
  INVD0BWP12T U3810 ( .I(register_file_inst1_r11_28_), .ZN(n4756) );
  OAI22D0BWP12T U3811 ( .A1(n4673), .A2(n5187), .B1(n4756), .B2(n4672), .ZN(
        n6253) );
  TPND2D0BWP12T U3812 ( .A1(n5985), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[7]), .ZN(n2265) );
  TPND2D0BWP12T U3813 ( .A1(n5985), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[6]), .ZN(n2266) );
  TPND2D0BWP12T U3814 ( .A1(n5985), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[8]), .ZN(n2261) );
  NR3D0BWP12T U3815 ( .A1(n5985), .A2(n6399), .A3(n6400), .ZN(n6237) );
  TPND2D0BWP12T U3816 ( .A1(n5985), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[9]), .ZN(n2259) );
  TPND2D0BWP12T U3817 ( .A1(n5985), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[10]), .ZN(n2257) );
  TPND2D0BWP12T U3818 ( .A1(n5985), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[11]), .ZN(n2255) );
  TPND2D0BWP12T U3819 ( .A1(n5985), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[12]), .ZN(n2253) );
  TPND2D0BWP12T U3820 ( .A1(n5985), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[13]), .ZN(n2251) );
  TPND2D0BWP12T U3821 ( .A1(n5985), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[14]), .ZN(n2249) );
  TPND2D0BWP12T U3822 ( .A1(n5985), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[15]), .ZN(n2247) );
  CKND1BWP12T U3823 ( .I(n2342), .ZN(n6406) );
  AOI31D0BWP12T U3824 ( .A1(n6282), .A2(n2348), .A3(n6406), .B(n6111), .ZN(
        n6112) );
  ND2XD0BWP12T U3825 ( .A1(memory_interface_inst1_fsm_state_0_), .A2(
        memory_interface_inst1_fsm_state_3_), .ZN(n4669) );
  NR2D0BWP12T U3826 ( .A1(n4090), .A2(n4669), .ZN(n4838) );
  AOI21D0BWP12T U3827 ( .A1(n6282), .A2(n2343), .B(n4838), .ZN(n6107) );
  INVD1BWP12T U3828 ( .I(memory_interface_inst1_fsm_state_3_), .ZN(n6401) );
  INVD1BWP12T U3829 ( .I(n4090), .ZN(n5181) );
  NR2D1BWP12T U3830 ( .A1(n4670), .A2(n4669), .ZN(n5180) );
  AOI31D0BWP12T U3831 ( .A1(n5181), .A2(memory_interface_inst1_fsm_state_0_), 
        .A3(n6401), .B(n5180), .ZN(n6108) );
  CKND0BWP12T U3832 ( .I(n4670), .ZN(n4671) );
  NR2D0BWP12T U3833 ( .A1(n4671), .A2(memory_interface_inst1_fsm_state_0_), 
        .ZN(n2244) );
  TPND2D0BWP12T U3834 ( .A1(n5985), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[0]), .ZN(n2269) );
  TPND2D0BWP12T U3835 ( .A1(n5985), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[4]), .ZN(n2268) );
  TPND2D0BWP12T U3836 ( .A1(n5985), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[5]), .ZN(n2267) );
  INVD1BWP12T U3837 ( .I(register_file_inst1_r12_31_), .ZN(n5241) );
  INVD1BWP12T U3838 ( .I(register_file_inst1_r11_31_), .ZN(n5218) );
  OAI22D0BWP12T U3839 ( .A1(n4673), .A2(n5241), .B1(n5218), .B2(n4672), .ZN(
        n6266) );
  CKND1BWP12T U3840 ( .I(register_file_inst1_r8_30_), .ZN(n5209) );
  TPNR2D0BWP12T U3841 ( .A1(n5209), .A2(n4674), .ZN(n6256) );
  CKND0BWP12T U3842 ( .I(register_file_inst1_r8_28_), .ZN(n5186) );
  TPNR2D0BWP12T U3843 ( .A1(n5186), .A2(n4674), .ZN(n6252) );
  INVD1BWP12T U3844 ( .I(n5234), .ZN(n5978) );
  INVD1BWP12T U3845 ( .I(register_file_inst1_r8_31_), .ZN(n5245) );
  TPNR2D0BWP12T U3846 ( .A1(n5245), .A2(n4674), .ZN(n6265) );
  NR2D1BWP12T U3847 ( .A1(n2911), .A2(n2919), .ZN(n6000) );
  BUFFD1BWP12T U3848 ( .I(n6226), .Z(n5997) );
  CKND0BWP12T U3849 ( .I(register_file_inst1_r8_24_), .ZN(n5144) );
  TPNR2D0BWP12T U3850 ( .A1(n5144), .A2(n4674), .ZN(n6274) );
  CKND0BWP12T U3851 ( .I(memory_interface_inst1_fsm_state_0_), .ZN(n4675) );
  AOI21D0BWP12T U3852 ( .A1(memory_interface_inst1_fsm_state_2_), .A2(
        memory_interface_inst1_fsm_state_1_), .B(n4675), .ZN(n2243) );
  CKND1BWP12T U3853 ( .I(n2471), .ZN(n6149) );
  INVD1BWP12T U3854 ( .I(n2874), .ZN(n6013) );
  CKND0BWP12T U3855 ( .I(n6286), .ZN(n6015) );
  CKND0BWP12T U3856 ( .I(n2469), .ZN(n6161) );
  CKND1BWP12T U3857 ( .I(n2516), .ZN(n6041) );
  OAI21D0BWP12T U3858 ( .A1(n6383), .A2(n6382), .B(n6381), .ZN(
        register_file_inst1_n2171) );
  INVD1BWP12T U3859 ( .I(n4754), .ZN(n4689) );
  CKND0BWP12T U3860 ( .I(register_file_inst1_r12_18_), .ZN(n4679) );
  OAI222D0BWP12T U3861 ( .A1(n4690), .A2(n5140), .B1(n5243), .B2(n4689), .C1(
        n5242), .C2(n4679), .ZN(register_file_inst1_n2251) );
  INVD1BWP12T U3862 ( .I(register_file_inst1_r1_18_), .ZN(n5501) );
  OAI222D0BWP12T U3863 ( .A1(n4690), .A2(n5074), .B1(n5240), .B2(n4689), .C1(
        n5239), .C2(n5501), .ZN(register_file_inst1_n2603) );
  CKND0BWP12T U3864 ( .I(register_file_inst1_r9_18_), .ZN(n4680) );
  OAI222D0BWP12T U3865 ( .A1(n4690), .A2(n5238), .B1(n5237), .B2(n4689), .C1(
        n5235), .C2(n4680), .ZN(register_file_inst1_n2347) );
  CKND0BWP12T U3866 ( .I(register_file_inst1_r8_18_), .ZN(n4681) );
  OAI222D0BWP12T U3867 ( .A1(n4690), .A2(n5145), .B1(n5246), .B2(n4689), .C1(
        n5244), .C2(n4681), .ZN(register_file_inst1_n2379) );
  CKND0BWP12T U3868 ( .I(register_file_inst1_r5_18_), .ZN(n4682) );
  OAI222D0BWP12T U3869 ( .A1(n4690), .A2(n5143), .B1(n5249), .B2(n4689), .C1(
        n5247), .C2(n4682), .ZN(register_file_inst1_n2475) );
  INVD1BWP12T U3870 ( .I(RF_next_sp[18]), .ZN(n5498) );
  OAI222D0BWP12T U3871 ( .A1(n4690), .A2(n5234), .B1(n5233), .B2(n4689), .C1(
        n5232), .C2(n5498), .ZN(register_file_inst1_spin[18]) );
  CKND0BWP12T U3872 ( .I(register_file_inst1_tmp1_18_), .ZN(n4684) );
  OAI222D0BWP12T U3873 ( .A1(n4690), .A2(n6144), .B1(n5212), .B2(n4689), .C1(
        n4683), .C2(n4684), .ZN(register_file_inst1_n2155) );
  INVD1BWP12T U3874 ( .I(register_file_inst1_lr_18_), .ZN(n5500) );
  OAI222D0BWP12T U3875 ( .A1(n4690), .A2(n5223), .B1(n5160), .B2(n4689), .C1(
        n5222), .C2(n5500), .ZN(register_file_inst1_n2219) );
  CKND0BWP12T U3876 ( .I(register_file_inst1_r4_18_), .ZN(n4685) );
  OAI222D0BWP12T U3877 ( .A1(n4690), .A2(n5226), .B1(n5205), .B2(n4689), .C1(
        n5225), .C2(n4685), .ZN(register_file_inst1_n2507) );
  INVD1BWP12T U3878 ( .I(register_file_inst1_r7_18_), .ZN(n5499) );
  OAI222D0BWP12T U3879 ( .A1(n4690), .A2(n5227), .B1(n5158), .B2(n4689), .C1(
        n5094), .C2(n5499), .ZN(register_file_inst1_n2411) );
  INVD1BWP12T U3880 ( .I(register_file_inst1_r2_18_), .ZN(n5488) );
  OAI222D0BWP12T U3881 ( .A1(n4690), .A2(n5257), .B1(n5256), .B2(n4689), .C1(
        n5254), .C2(n5488), .ZN(register_file_inst1_n2571) );
  INVD1BWP12T U3882 ( .I(register_file_inst1_r10_18_), .ZN(n4686) );
  OAI222D0BWP12T U3883 ( .A1(n4690), .A2(n5253), .B1(n5252), .B2(n4689), .C1(
        n5250), .C2(n4686), .ZN(register_file_inst1_n2315) );
  INVD1BWP12T U3884 ( .I(register_file_inst1_r0_18_), .ZN(n5487) );
  OAI222D0BWP12T U3885 ( .A1(n4690), .A2(n5231), .B1(n5230), .B2(n4689), .C1(
        n5096), .C2(n5487), .ZN(register_file_inst1_n2635) );
  INVD1BWP12T U3886 ( .I(register_file_inst1_r6_18_), .ZN(n5486) );
  OAI222D0BWP12T U3887 ( .A1(n4690), .A2(n5229), .B1(n5228), .B2(n4689), .C1(
        n5095), .C2(n5486), .ZN(register_file_inst1_n2443) );
  CKND0BWP12T U3888 ( .I(register_file_inst1_r11_18_), .ZN(n4687) );
  OAI222D0BWP12T U3889 ( .A1(n4690), .A2(n5220), .B1(n5219), .B2(n4689), .C1(
        n5217), .C2(n4687), .ZN(register_file_inst1_n2283) );
  CKND0BWP12T U3890 ( .I(register_file_inst1_r3_18_), .ZN(n4688) );
  OAI222D0BWP12T U3891 ( .A1(n4690), .A2(n5200), .B1(n5203), .B2(n4689), .C1(
        n4758), .C2(n4688), .ZN(register_file_inst1_n2539) );
  OAI21D0BWP12T U3892 ( .A1(n6375), .A2(n6374), .B(n6373), .ZN(
        register_file_inst1_n2173) );
  INVD1BWP12T U3893 ( .I(n6395), .ZN(n5270) );
  OAI222D0BWP12T U3894 ( .A1(n4691), .A2(n5269), .B1(n6369), .B2(n5270), .C1(
        n6364), .C2(n5267), .ZN(n6365) );
  OAI21D0BWP12T U3895 ( .A1(n6371), .A2(n5046), .B(n6370), .ZN(
        register_file_inst1_n2174) );
  OAI22D1BWP12T U3896 ( .A1(n4692), .A2(n5910), .B1(n5476), .B2(n5857), .ZN(
        n4703) );
  OAI22D1BWP12T U3897 ( .A1(n4694), .A2(n5959), .B1(n4693), .B2(n5912), .ZN(
        n4702) );
  AOI22D1BWP12T U3898 ( .A1(register_file_inst1_tmp1_19_), .A2(n5962), .B1(
        register_file_inst1_r4_19_), .B2(n5961), .ZN(n4696) );
  AOI22D1BWP12T U3899 ( .A1(RF_next_sp[19]), .A2(n5964), .B1(
        register_file_inst1_r12_19_), .B2(n5963), .ZN(n4695) );
  ND3D1BWP12T U3900 ( .A1(n4696), .A2(n4695), .A3(n6120), .ZN(n4701) );
  AOI22D1BWP12T U3901 ( .A1(register_file_inst1_r9_19_), .A2(n5968), .B1(
        register_file_inst1_r3_19_), .B2(n5967), .ZN(n4699) );
  AOI22D1BWP12T U3902 ( .A1(register_file_inst1_r7_19_), .A2(n6001), .B1(
        register_file_inst1_r11_19_), .B2(n5969), .ZN(n4698) );
  AOI22D1BWP12T U3903 ( .A1(register_file_inst1_r5_19_), .A2(n6002), .B1(
        register_file_inst1_lr_19_), .B2(n5970), .ZN(n4697) );
  ND4D1BWP12T U3904 ( .A1(n4699), .A2(n4698), .A3(n6121), .A4(n4697), .ZN(
        n4700) );
  OR4D4BWP12T U3905 ( .A1(n4703), .A2(n4702), .A3(n4701), .A4(n4700), .Z(
        RF_ALU_operand_b[19]) );
  OAI22D1BWP12T U3906 ( .A1(n4704), .A2(n5910), .B1(n5590), .B2(n5857), .ZN(
        n4715) );
  OAI22D1BWP12T U3907 ( .A1(n4706), .A2(n5959), .B1(n4705), .B2(n5912), .ZN(
        n4714) );
  AOI22D1BWP12T U3908 ( .A1(register_file_inst1_tmp1_13_), .A2(n5962), .B1(
        register_file_inst1_r4_13_), .B2(n5961), .ZN(n4708) );
  AOI22D1BWP12T U3909 ( .A1(RF_next_sp[13]), .A2(n5964), .B1(
        register_file_inst1_r12_13_), .B2(n5963), .ZN(n4707) );
  ND3D1BWP12T U3910 ( .A1(n4708), .A2(n4707), .A3(n6101), .ZN(n4713) );
  AOI22D1BWP12T U3911 ( .A1(register_file_inst1_r9_13_), .A2(n5968), .B1(
        register_file_inst1_r3_13_), .B2(n5967), .ZN(n4711) );
  AOI22D1BWP12T U3912 ( .A1(register_file_inst1_r7_13_), .A2(n6001), .B1(
        register_file_inst1_r11_13_), .B2(n5969), .ZN(n4710) );
  ND4D1BWP12T U3913 ( .A1(n4711), .A2(n4710), .A3(n6102), .A4(n4709), .ZN(
        n4712) );
  OR4D4BWP12T U3914 ( .A1(n4715), .A2(n4714), .A3(n4713), .A4(n4712), .Z(
        RF_ALU_operand_b[13]) );
  OAI21D0BWP12T U3915 ( .A1(n6363), .A2(n6362), .B(n6361), .ZN(
        register_file_inst1_n2177) );
  OAI21D0BWP12T U3916 ( .A1(n5984), .A2(n4716), .B(n6366), .ZN(n6360) );
  OAI21D0BWP12T U3917 ( .A1(n6359), .A2(n5117), .B(n6358), .ZN(
        register_file_inst1_n2178) );
  OAI222D0BWP12T U3918 ( .A1(n4717), .A2(n5269), .B1(n6357), .B2(n5270), .C1(
        n6352), .C2(n5267), .ZN(n6353) );
  OAI222D0BWP12T U3919 ( .A1(n5119), .A2(n5269), .B1(n5267), .B2(n5120), .C1(
        n5270), .C2(n6331), .ZN(n6328) );
  CKND0BWP12T U3920 ( .I(n5122), .ZN(n6354) );
  OAI222D0BWP12T U3921 ( .A1(n5084), .A2(n5269), .B1(n6351), .B2(n5270), .C1(
        n6346), .C2(n5267), .ZN(n6347) );
  OAI222D0BWP12T U3922 ( .A1(n5088), .A2(n5269), .B1(n6345), .B2(n5270), .C1(
        n6340), .C2(n5267), .ZN(n6341) );
  OAI222D0BWP12T U3923 ( .A1(n5098), .A2(n5269), .B1(n5267), .B2(n5099), .C1(
        n5270), .C2(n6339), .ZN(n6336) );
  OAI222D0BWP12T U3924 ( .A1(n5114), .A2(n5269), .B1(n5267), .B2(n5115), .C1(
        n5270), .C2(n6335), .ZN(n6332) );
  OAI222D0BWP12T U3925 ( .A1(n5136), .A2(n5269), .B1(n6327), .B2(n5270), .C1(
        n5135), .C2(n5267), .ZN(n6324) );
  CKND0BWP12T U3926 ( .I(n5137), .ZN(n6348) );
  CKND0BWP12T U3927 ( .I(n5215), .ZN(n6325) );
  CKND0BWP12T U3928 ( .I(n4752), .ZN(n6342) );
  CKND0BWP12T U3929 ( .I(n4755), .ZN(n6337) );
  CKND0BWP12T U3930 ( .I(n4760), .ZN(n6333) );
  INVD1BWP12T U3931 ( .I(n5267), .ZN(n6379) );
  AO222D0BWP12T U3932 ( .A1(n4749), .A2(n6379), .B1(n6376), .B2(
        ALU_MISC_OUT_result[22]), .C1(n6395), .C2(n4730), .Z(n6326) );
  OAI222D0BWP12T U3933 ( .A1(n5177), .A2(n5269), .B1(n5267), .B2(n5178), .C1(
        n5270), .C2(n6319), .ZN(n6316) );
  OAI22D1BWP12T U3934 ( .A1(n4718), .A2(n5910), .B1(n5577), .B2(n5857), .ZN(
        n4729) );
  OAI22D1BWP12T U3935 ( .A1(n4720), .A2(n5959), .B1(n4719), .B2(n5912), .ZN(
        n4728) );
  AOI22D1BWP12T U3936 ( .A1(register_file_inst1_tmp1_14_), .A2(n5962), .B1(
        register_file_inst1_r4_14_), .B2(n5961), .ZN(n4722) );
  AOI22D1BWP12T U3937 ( .A1(RF_next_sp[14]), .A2(n5964), .B1(
        register_file_inst1_r12_14_), .B2(n5963), .ZN(n4721) );
  ND3D1BWP12T U3938 ( .A1(n4722), .A2(n4721), .A3(n6103), .ZN(n4727) );
  AOI22D1BWP12T U3939 ( .A1(register_file_inst1_r9_14_), .A2(n5968), .B1(
        register_file_inst1_r3_14_), .B2(n5967), .ZN(n4725) );
  AOI22D1BWP12T U3940 ( .A1(register_file_inst1_r7_14_), .A2(n6001), .B1(
        register_file_inst1_r11_14_), .B2(n5969), .ZN(n4724) );
  AOI22D1BWP12T U3941 ( .A1(register_file_inst1_r5_14_), .A2(n6002), .B1(
        register_file_inst1_lr_14_), .B2(n5970), .ZN(n4723) );
  ND4D1BWP12T U3942 ( .A1(n4725), .A2(n4724), .A3(n6104), .A4(n4723), .ZN(
        n4726) );
  CKND0BWP12T U3943 ( .I(n4730), .ZN(n6329) );
  OAI22D1BWP12T U3944 ( .A1(n4731), .A2(n5910), .B1(n5874), .B2(n5857), .ZN(
        n4742) );
  OAI22D1BWP12T U3945 ( .A1(n4733), .A2(n5959), .B1(n4732), .B2(n5912), .ZN(
        n4741) );
  AOI22D1BWP12T U3946 ( .A1(register_file_inst1_tmp1_21_), .A2(n5962), .B1(
        register_file_inst1_r4_21_), .B2(n5961), .ZN(n4735) );
  AOI22D1BWP12T U3947 ( .A1(RF_next_sp[21]), .A2(n5964), .B1(
        register_file_inst1_r12_21_), .B2(n5963), .ZN(n4734) );
  ND3D1BWP12T U3948 ( .A1(n4735), .A2(n4734), .A3(n6124), .ZN(n4740) );
  AOI22D1BWP12T U3949 ( .A1(register_file_inst1_r9_21_), .A2(n5968), .B1(
        register_file_inst1_r3_21_), .B2(n5967), .ZN(n4738) );
  AOI22D1BWP12T U3950 ( .A1(register_file_inst1_r7_21_), .A2(n6001), .B1(
        register_file_inst1_r11_21_), .B2(n5969), .ZN(n4737) );
  AOI22D1BWP12T U3951 ( .A1(register_file_inst1_r5_21_), .A2(n6002), .B1(
        register_file_inst1_lr_21_), .B2(n5970), .ZN(n4736) );
  ND4D1BWP12T U3952 ( .A1(n4738), .A2(n4737), .A3(n6125), .A4(n4736), .ZN(
        n4739) );
  OR4XD1BWP12T U3953 ( .A1(n4742), .A2(n4741), .A3(n4740), .A4(n4739), .Z(
        RF_ALU_operand_b[21]) );
  OAI222D1BWP12T U3954 ( .A1(n3718), .A2(n5205), .B1(n5020), .B2(n5226), .C1(
        n5225), .C2(n4743), .ZN(register_file_inst1_n2489) );
  INVD1BWP12T U3955 ( .I(register_file_inst1_r3_6_), .ZN(n4744) );
  OAI222D1BWP12T U3956 ( .A1(n5034), .A2(n5200), .B1(n5203), .B2(n6367), .C1(
        n4758), .C2(n4744), .ZN(register_file_inst1_n2527) );
  INVD1BWP12T U3957 ( .I(register_file_inst1_r3_12_), .ZN(n4745) );
  OAI222D1BWP12T U3958 ( .A1(n5082), .A2(n5200), .B1(n5203), .B2(n6349), .C1(
        n4758), .C2(n4745), .ZN(register_file_inst1_n2533) );
  INVD1BWP12T U3959 ( .I(register_file_inst1_r11_16_), .ZN(n4746) );
  INVD1BWP12T U3960 ( .I(n4753), .ZN(n5103) );
  OAI222D1BWP12T U3961 ( .A1(n4746), .A2(n5217), .B1(n5219), .B2(n5103), .C1(
        n5102), .C2(n5220), .ZN(register_file_inst1_n2281) );
  INVD1BWP12T U3962 ( .I(register_file_inst1_r3_16_), .ZN(n4747) );
  OAI222D1BWP12T U3963 ( .A1(n4747), .A2(n4758), .B1(n5203), .B2(n5103), .C1(
        n5102), .C2(n5200), .ZN(register_file_inst1_n2537) );
  INVD1BWP12T U3964 ( .I(register_file_inst1_r3_20_), .ZN(n4748) );
  INVD1BWP12T U3965 ( .I(n4761), .ZN(n5112) );
  OAI222D1BWP12T U3966 ( .A1(n4748), .A2(n4758), .B1(n5203), .B2(n5112), .C1(
        n5111), .C2(n5200), .ZN(register_file_inst1_n2541) );
  CKND0BWP12T U3967 ( .I(register_file_inst1_r3_22_), .ZN(n4750) );
  INVD1BWP12T U3968 ( .I(n4749), .ZN(n5132) );
  INVD1BWP12T U3969 ( .I(register_file_inst1_r7_25_), .ZN(n5925) );
  OAI222D1BWP12T U3970 ( .A1(n5925), .A2(n5094), .B1(n5158), .B2(n5261), .C1(
        n5262), .C2(n5227), .ZN(register_file_inst1_n2418) );
  INVD1BWP12T U3971 ( .I(register_file_inst1_lr_25_), .ZN(n5926) );
  OAI222D1BWP12T U3972 ( .A1(n5926), .A2(n5222), .B1(n5160), .B2(n5261), .C1(
        n5262), .C2(n5223), .ZN(register_file_inst1_n2226) );
  CKND0BWP12T U3973 ( .I(register_file_inst1_r3_26_), .ZN(n4751) );
  OAI222D1BWP12T U3974 ( .A1(n4751), .A2(n4758), .B1(n5203), .B2(n5263), .C1(
        n5167), .C2(n5200), .ZN(register_file_inst1_n2547) );
  INVD1BWP12T U3975 ( .I(register_file_inst1_lr_27_), .ZN(n5387) );
  OAI222D1BWP12T U3976 ( .A1(n5387), .A2(n5222), .B1(n5160), .B2(n5178), .C1(
        n5177), .C2(n5223), .ZN(register_file_inst1_n2228) );
  INVD1BWP12T U3977 ( .I(register_file_inst1_r7_27_), .ZN(n5386) );
  OAI222D1BWP12T U3978 ( .A1(n5386), .A2(n5094), .B1(n5158), .B2(n5178), .C1(
        n5177), .C2(n5227), .ZN(register_file_inst1_n2420) );
  INVD1BWP12T U3979 ( .I(register_file_inst1_r0_27_), .ZN(n5374) );
  OAI222D1BWP12T U3980 ( .A1(n5374), .A2(n5096), .B1(n5230), .B2(n5178), .C1(
        n5177), .C2(n5231), .ZN(register_file_inst1_n2644) );
  INVD1BWP12T U3981 ( .I(register_file_inst1_r6_27_), .ZN(n5373) );
  OAI222D1BWP12T U3982 ( .A1(n5373), .A2(n5095), .B1(n5228), .B2(n5178), .C1(
        n5177), .C2(n5229), .ZN(register_file_inst1_n2452) );
  AO222D0BWP12T U3983 ( .A1(n4753), .A2(n6379), .B1(n6376), .B2(
        ALU_MISC_OUT_result[16]), .C1(n6395), .C2(n4752), .Z(n6338) );
  AO222D0BWP12T U3984 ( .A1(n6395), .A2(n4755), .B1(n6376), .B2(
        ALU_MISC_OUT_result[18]), .C1(n4754), .C2(n6379), .Z(n6334) );
  INVD3BWP12T U3985 ( .I(ALU_MISC_OUT_result[28]), .ZN(n5189) );
  OAI222D1BWP12T U3986 ( .A1(n4756), .A2(n5217), .B1(n5219), .B2(n5190), .C1(
        n5189), .C2(n5220), .ZN(register_file_inst1_n2293) );
  CKND0BWP12T U3987 ( .I(register_file_inst1_r3_28_), .ZN(n4757) );
  OAI222D1BWP12T U3988 ( .A1(n4757), .A2(n4758), .B1(n5203), .B2(n5190), .C1(
        n5189), .C2(n5200), .ZN(register_file_inst1_n2549) );
  INVD1BWP12T U3989 ( .I(register_file_inst1_r7_30_), .ZN(n5311) );
  INVD2BWP12T U3990 ( .I(ALU_MISC_OUT_result[30]), .ZN(n5268) );
  OAI222D1BWP12T U3991 ( .A1(n5311), .A2(n5094), .B1(n5158), .B2(n5266), .C1(
        n5268), .C2(n5227), .ZN(register_file_inst1_n2423) );
  INVD1BWP12T U3992 ( .I(register_file_inst1_r6_30_), .ZN(n5298) );
  OAI222D1BWP12T U3993 ( .A1(n5298), .A2(n5095), .B1(n5228), .B2(n5266), .C1(
        n5268), .C2(n5229), .ZN(register_file_inst1_n2455) );
  INVD1BWP12T U3994 ( .I(register_file_inst1_lr_30_), .ZN(n5312) );
  OAI222D1BWP12T U3995 ( .A1(n5312), .A2(n5222), .B1(n5160), .B2(n5266), .C1(
        n5268), .C2(n5223), .ZN(register_file_inst1_n2231) );
  INVD0BWP12T U3996 ( .I(register_file_inst1_r3_30_), .ZN(n4759) );
  OAI222D1BWP12T U3997 ( .A1(n4759), .A2(n4758), .B1(n5203), .B2(n5266), .C1(
        n5268), .C2(n5200), .ZN(register_file_inst1_n2551) );
  AO222D0BWP12T U3998 ( .A1(n4761), .A2(n6379), .B1(n6376), .B2(
        ALU_MISC_OUT_result[20]), .C1(n6395), .C2(n4760), .Z(n6330) );
  INVD0BWP12T U3999 ( .I(register_file_inst1_r3_31_), .ZN(n4762) );
  OAI222D1BWP12T U4000 ( .A1(n5258), .A2(n5200), .B1(n5203), .B2(n5255), .C1(
        n4758), .C2(n4762), .ZN(register_file_inst1_n2552) );
  INVD1BWP12T U4001 ( .I(n4763), .ZN(n6317) );
  OAI222D1BWP12T U4002 ( .A1(n5189), .A2(n5269), .B1(n5267), .B2(n5190), .C1(
        n5270), .C2(n6317), .ZN(n6314) );
  CKND2BWP12T U4003 ( .I(ALU_MISC_OUT_result[29]), .ZN(n5201) );
  INVD1BWP12T U4004 ( .I(n4764), .ZN(n5202) );
  OAI222D1BWP12T U4005 ( .A1(n5201), .A2(n5269), .B1(n5267), .B2(n5202), .C1(
        n5270), .C2(n6315), .ZN(n6312) );
  INR2D1BWP12T U4006 ( .A1(n2878), .B1(n6405), .ZN(n2871) );
  INVD1BWP12T U4007 ( .I(MEM_MEMCTRL_from_mem_data[8]), .ZN(n4096) );
  INVD1BWP12T U4008 ( .I(MEM_MEMCTRL_from_mem_data[12]), .ZN(n4095) );
  INVD1BWP12T U4009 ( .I(MEM_MEMCTRL_from_mem_data[13]), .ZN(n4094) );
  INVD1BWP12T U4010 ( .I(MEM_MEMCTRL_from_mem_data[14]), .ZN(n4093) );
  INVD1BWP12T U4011 ( .I(MEM_MEMCTRL_from_mem_data[0]), .ZN(n4104) );
  INVD1BWP12T U4012 ( .I(MEM_MEMCTRL_from_mem_data[1]), .ZN(n4103) );
  INVD1BWP12T U4013 ( .I(MEM_MEMCTRL_from_mem_data[2]), .ZN(n4102) );
  INVD1BWP12T U4014 ( .I(MEM_MEMCTRL_from_mem_data[3]), .ZN(n4101) );
  INVD1BWP12T U4015 ( .I(MEM_MEMCTRL_from_mem_data[4]), .ZN(n4100) );
  INVD1BWP12T U4016 ( .I(MEM_MEMCTRL_from_mem_data[6]), .ZN(n4098) );
  INVD1BWP12T U4017 ( .I(MEM_MEMCTRL_from_mem_data[7]), .ZN(n4097) );
  CKND0BWP12T U4018 ( .I(n5180), .ZN(n4822) );
  NR2D0BWP12T U4019 ( .A1(memory_interface_inst1_fsm_state_0_), .A2(
        memory_interface_inst1_fsm_state_1_), .ZN(n4766) );
  OAI21D1BWP12T U4020 ( .A1(n4766), .A2(n4765), .B(n6401), .ZN(n4841) );
  ND2D1BWP12T U4021 ( .A1(n4822), .A2(n4841), .ZN(n6232) );
  NR2D1BWP12T U4022 ( .A1(n3059), .A2(n3054), .ZN(n5992) );
  NR2D1BWP12T U4023 ( .A1(n6149), .A2(n6151), .ZN(n5999) );
  CKBD1BWP12T U4024 ( .I(n5999), .Z(n6006) );
  NR2D1BWP12T U4025 ( .A1(n3060), .A2(n3056), .ZN(n5991) );
  INVD1BWP12T U4026 ( .I(n5232), .ZN(n6097) );
  ND2D1BWP12T U4027 ( .A1(n3046), .A2(n3047), .ZN(n4773) );
  NR2D1BWP12T U4028 ( .A1(n3054), .A2(n4773), .ZN(n5058) );
  ND2D1BWP12T U4029 ( .A1(n3048), .A2(n3049), .ZN(n4768) );
  NR2D1BWP12T U4030 ( .A1(n3059), .A2(n4768), .ZN(n5057) );
  AOI22D1BWP12T U4031 ( .A1(n5058), .A2(register_file_inst1_r3_3_), .B1(
        register_file_inst1_r12_3_), .B2(n5057), .ZN(n4772) );
  NR2D1BWP12T U4032 ( .A1(n3060), .A2(n4768), .ZN(n5060) );
  NR2D1BWP12T U4033 ( .A1(n3055), .A2(n4768), .ZN(n5059) );
  AOI22D1BWP12T U4034 ( .A1(n5060), .A2(register_file_inst1_r4_3_), .B1(
        register_file_inst1_r8_3_), .B2(n5059), .ZN(n4771) );
  NR2D1BWP12T U4035 ( .A1(n4773), .A2(n4768), .ZN(n5062) );
  NR2D1BWP12T U4036 ( .A1(n3056), .A2(n4773), .ZN(n5061) );
  AOI22D0BWP12T U4037 ( .A1(n5062), .A2(register_file_inst1_r0_3_), .B1(
        register_file_inst1_r1_3_), .B2(n5061), .ZN(n4770) );
  NR2D1BWP12T U4038 ( .A1(n3061), .A2(n3055), .ZN(n5064) );
  NR2D1BWP12T U4039 ( .A1(n3055), .A2(n3054), .ZN(n5063) );
  AOI22D1BWP12T U4040 ( .A1(n5064), .A2(register_file_inst1_r10_3_), .B1(
        register_file_inst1_r11_3_), .B2(n5063), .ZN(n4769) );
  ND4D1BWP12T U4041 ( .A1(n4772), .A2(n4771), .A3(n4770), .A4(n4769), .ZN(
        n4778) );
  NR2D1BWP12T U4042 ( .A1(n3061), .A2(n3059), .ZN(n5049) );
  NR2D1BWP12T U4043 ( .A1(n3056), .A2(n3055), .ZN(n5048) );
  AOI22D1BWP12T U4044 ( .A1(n5049), .A2(register_file_inst1_lr_3_), .B1(
        register_file_inst1_r9_3_), .B2(n5048), .ZN(n4776) );
  NR2D1BWP12T U4045 ( .A1(n3059), .A2(n3056), .ZN(n5051) );
  NR2D1BWP12T U4046 ( .A1(n3060), .A2(n3054), .ZN(n5050) );
  AOI22D1BWP12T U4047 ( .A1(n5051), .A2(RF_next_sp[3]), .B1(
        register_file_inst1_r7_3_), .B2(n5050), .ZN(n4775) );
  NR2D1BWP12T U4048 ( .A1(n3060), .A2(n3061), .ZN(n5053) );
  NR2D1BWP12T U4049 ( .A1(n3061), .A2(n4773), .ZN(n5052) );
  AOI22D1BWP12T U4050 ( .A1(n5053), .A2(register_file_inst1_r6_3_), .B1(
        register_file_inst1_r2_3_), .B2(n5052), .ZN(n4774) );
  ND4D1BWP12T U4051 ( .A1(n6261), .A2(n4776), .A3(n4775), .A4(n4774), .ZN(
        n4777) );
  OAI21D1BWP12T U4052 ( .A1(n4778), .A2(n4777), .B(n6397), .ZN(n4779) );
  ND2D1BWP12T U4053 ( .A1(n3202), .A2(n4779), .ZN(MEMCTRL_IN_address[2]) );
  AOI22D1BWP12T U4054 ( .A1(memory_interface_inst1_delay_addr_single[2]), .A2(
        n6294), .B1(MEMCTRL_IN_address[2]), .B2(n6295), .ZN(n4781) );
  INVD1BWP12T U4055 ( .I(memory_interface_inst1_delay_addr_for_adder_0_), .ZN(
        n4821) );
  INR2D1BWP12T U4056 ( .A1(memory_interface_inst1_delay_addr_for_adder_1_), 
        .B1(n4821), .ZN(n4820) );
  NR2D1BWP12T U4057 ( .A1(n6295), .A2(n6294), .ZN(n4928) );
  ND2D1BWP12T U4058 ( .A1(n4820), .A2(
        memory_interface_inst1_delay_addr_for_adder_2_), .ZN(n4875) );
  OAI211D1BWP12T U4059 ( .A1(n4820), .A2(
        memory_interface_inst1_delay_addr_for_adder_2_), .B(n4928), .C(n4875), 
        .ZN(n4780) );
  ND2D1BWP12T U4060 ( .A1(n4781), .A2(n4780), .ZN(
        MEMCTRL_MEM_to_mem_address[2]) );
  AOI22D0BWP12T U4061 ( .A1(n5058), .A2(register_file_inst1_r3_8_), .B1(
        register_file_inst1_r12_8_), .B2(n5057), .ZN(n4785) );
  AOI22D0BWP12T U4062 ( .A1(n5060), .A2(register_file_inst1_r4_8_), .B1(
        register_file_inst1_r8_8_), .B2(n5059), .ZN(n4784) );
  AOI22D0BWP12T U4063 ( .A1(n5062), .A2(register_file_inst1_r0_8_), .B1(
        register_file_inst1_r1_8_), .B2(n5061), .ZN(n4783) );
  AOI22D0BWP12T U4064 ( .A1(n5064), .A2(register_file_inst1_r10_8_), .B1(
        register_file_inst1_r11_8_), .B2(n5063), .ZN(n4782) );
  ND4D1BWP12T U4065 ( .A1(n4785), .A2(n4784), .A3(n4783), .A4(n4782), .ZN(
        n4790) );
  AOI22D0BWP12T U4066 ( .A1(n5049), .A2(register_file_inst1_lr_8_), .B1(
        register_file_inst1_r9_8_), .B2(n5048), .ZN(n4788) );
  AOI22D0BWP12T U4067 ( .A1(n5051), .A2(RF_next_sp[8]), .B1(
        register_file_inst1_r7_8_), .B2(n5050), .ZN(n4787) );
  AOI22D0BWP12T U4068 ( .A1(n5053), .A2(register_file_inst1_r6_8_), .B1(
        register_file_inst1_r2_8_), .B2(n5052), .ZN(n4786) );
  ND4D1BWP12T U4069 ( .A1(n6260), .A2(n4788), .A3(n4787), .A4(n4786), .ZN(
        n4789) );
  OAI21D1BWP12T U4070 ( .A1(n4790), .A2(n4789), .B(n6397), .ZN(n4791) );
  ND2D1BWP12T U4071 ( .A1(n3217), .A2(n4791), .ZN(MEMCTRL_IN_address[7]) );
  AOI22D1BWP12T U4072 ( .A1(memory_interface_inst1_delay_addr_single[7]), .A2(
        n6294), .B1(MEMCTRL_IN_address[7]), .B2(n6295), .ZN(n4794) );
  INVD1BWP12T U4073 ( .I(memory_interface_inst1_delay_addr_for_adder_3_), .ZN(
        n4874) );
  NR2D1BWP12T U4074 ( .A1(n4875), .A2(n4874), .ZN(n4873) );
  ND2D1BWP12T U4075 ( .A1(n4873), .A2(
        memory_interface_inst1_delay_addr_for_adder_4_), .ZN(n4858) );
  INVD1BWP12T U4076 ( .I(memory_interface_inst1_delay_addr_for_adder_5_), .ZN(
        n4835) );
  NR2D1BWP12T U4077 ( .A1(n4858), .A2(n4835), .ZN(n4834) );
  ND2D1BWP12T U4078 ( .A1(n4834), .A2(
        memory_interface_inst1_delay_addr_for_adder_6_), .ZN(n4805) );
  INVD1BWP12T U4079 ( .I(memory_interface_inst1_delay_addr_for_adder_7_), .ZN(
        n4792) );
  NR2D1BWP12T U4080 ( .A1(n4805), .A2(n4792), .ZN(n4912) );
  INVD1BWP12T U4081 ( .I(n4928), .ZN(n4888) );
  AO211D1BWP12T U4082 ( .A1(n4805), .A2(n4792), .B(n4912), .C(n4888), .Z(n4793) );
  ND2D1BWP12T U4083 ( .A1(n4794), .A2(n4793), .ZN(
        MEMCTRL_MEM_to_mem_address[7]) );
  AOI22D1BWP12T U4084 ( .A1(n5058), .A2(register_file_inst1_r3_7_), .B1(
        register_file_inst1_r12_7_), .B2(n5057), .ZN(n4798) );
  AOI22D1BWP12T U4085 ( .A1(n5060), .A2(register_file_inst1_r4_7_), .B1(
        register_file_inst1_r8_7_), .B2(n5059), .ZN(n4797) );
  AOI22D0BWP12T U4086 ( .A1(n5062), .A2(register_file_inst1_r0_7_), .B1(
        register_file_inst1_r1_7_), .B2(n5061), .ZN(n4796) );
  AOI22D0BWP12T U4087 ( .A1(n5064), .A2(register_file_inst1_r10_7_), .B1(
        register_file_inst1_r11_7_), .B2(n5063), .ZN(n4795) );
  ND4D1BWP12T U4088 ( .A1(n4798), .A2(n4797), .A3(n4796), .A4(n4795), .ZN(
        n4803) );
  AOI22D1BWP12T U4089 ( .A1(n5049), .A2(register_file_inst1_lr_7_), .B1(
        register_file_inst1_r9_7_), .B2(n5048), .ZN(n4801) );
  AOI22D0BWP12T U4090 ( .A1(n5051), .A2(RF_next_sp[7]), .B1(
        register_file_inst1_r7_7_), .B2(n5050), .ZN(n4800) );
  AOI22D0BWP12T U4091 ( .A1(n5053), .A2(register_file_inst1_r6_7_), .B1(
        register_file_inst1_r2_7_), .B2(n5052), .ZN(n4799) );
  ND4D1BWP12T U4092 ( .A1(n6246), .A2(n4801), .A3(n4800), .A4(n4799), .ZN(
        n4802) );
  OAI21D1BWP12T U4093 ( .A1(n4803), .A2(n4802), .B(n6397), .ZN(n4804) );
  ND2D1BWP12T U4094 ( .A1(n3335), .A2(n4804), .ZN(MEMCTRL_IN_address[6]) );
  AOI22D1BWP12T U4095 ( .A1(memory_interface_inst1_delay_addr_single[6]), .A2(
        n6294), .B1(MEMCTRL_IN_address[6]), .B2(n6295), .ZN(n4807) );
  OAI211D1BWP12T U4096 ( .A1(n4834), .A2(
        memory_interface_inst1_delay_addr_for_adder_6_), .B(n4928), .C(n4805), 
        .ZN(n4806) );
  ND2D1BWP12T U4097 ( .A1(n4807), .A2(n4806), .ZN(
        MEMCTRL_MEM_to_mem_address[6]) );
  NR2D1BWP12T U4098 ( .A1(memory_interface_inst1_delay_addr_for_adder_0_), 
        .A2(memory_interface_inst1_delay_addr_for_adder_1_), .ZN(n4819) );
  AOI22D0BWP12T U4099 ( .A1(n5058), .A2(register_file_inst1_r3_2_), .B1(
        register_file_inst1_r12_2_), .B2(n5057), .ZN(n4811) );
  AOI22D0BWP12T U4100 ( .A1(n5060), .A2(register_file_inst1_r4_2_), .B1(
        register_file_inst1_r8_2_), .B2(n5059), .ZN(n4810) );
  AOI22D0BWP12T U4101 ( .A1(n5062), .A2(register_file_inst1_r0_2_), .B1(
        register_file_inst1_r1_2_), .B2(n5061), .ZN(n4809) );
  AOI22D0BWP12T U4102 ( .A1(n5064), .A2(register_file_inst1_r10_2_), .B1(
        register_file_inst1_r11_2_), .B2(n5063), .ZN(n4808) );
  ND4D1BWP12T U4103 ( .A1(n4811), .A2(n4810), .A3(n4809), .A4(n4808), .ZN(
        n4816) );
  AOI22D0BWP12T U4104 ( .A1(n5049), .A2(register_file_inst1_lr_2_), .B1(
        register_file_inst1_r9_2_), .B2(n5048), .ZN(n4814) );
  AOI22D0BWP12T U4105 ( .A1(n5051), .A2(RF_next_sp[2]), .B1(
        register_file_inst1_r7_2_), .B2(n5050), .ZN(n4813) );
  AOI22D0BWP12T U4106 ( .A1(n5053), .A2(register_file_inst1_r6_2_), .B1(
        register_file_inst1_r2_2_), .B2(n5052), .ZN(n4812) );
  ND4D1BWP12T U4107 ( .A1(n6273), .A2(n4814), .A3(n4813), .A4(n4812), .ZN(
        n4815) );
  OAI21D1BWP12T U4108 ( .A1(n4816), .A2(n4815), .B(n6397), .ZN(n4817) );
  ND2D1BWP12T U4109 ( .A1(n3095), .A2(n4817), .ZN(MEMCTRL_IN_address[1]) );
  AOI22D1BWP12T U4110 ( .A1(memory_interface_inst1_delay_addr_single[1]), .A2(
        n6294), .B1(MEMCTRL_IN_address[1]), .B2(n6295), .ZN(n4818) );
  OAI31D1BWP12T U4111 ( .A1(n4820), .A2(n4819), .A3(n4888), .B(n4818), .ZN(
        MEMCTRL_MEM_to_mem_address[1]) );
  AO222D1BWP12T U4112 ( .A1(n6295), .A2(MEMCTRL_IN_address[0]), .B1(n6294), 
        .B2(memory_interface_inst1_delay_addr_single[0]), .C1(n4821), .C2(
        n4928), .Z(MEMCTRL_MEM_to_mem_address[0]) );
  INVD1BWP12T U4113 ( .I(n5017), .ZN(n4823) );
  OAI21D1BWP12T U4114 ( .A1(n3018), .A2(n3017), .B(n4823), .ZN(
        MEMCTRL_MEM_to_mem_write_enable) );
  AOI22D1BWP12T U4115 ( .A1(n5058), .A2(register_file_inst1_r3_6_), .B1(
        register_file_inst1_r12_6_), .B2(n5057), .ZN(n4827) );
  AOI22D1BWP12T U4116 ( .A1(n5060), .A2(register_file_inst1_r4_6_), .B1(
        register_file_inst1_r8_6_), .B2(n5059), .ZN(n4826) );
  AOI22D0BWP12T U4117 ( .A1(n5062), .A2(register_file_inst1_r0_6_), .B1(
        register_file_inst1_r1_6_), .B2(n5061), .ZN(n4825) );
  AOI22D1BWP12T U4118 ( .A1(n5064), .A2(register_file_inst1_r10_6_), .B1(
        register_file_inst1_r11_6_), .B2(n5063), .ZN(n4824) );
  ND4D1BWP12T U4119 ( .A1(n4827), .A2(n4826), .A3(n4825), .A4(n4824), .ZN(
        n4832) );
  AOI22D1BWP12T U4120 ( .A1(n5049), .A2(register_file_inst1_lr_6_), .B1(
        register_file_inst1_r9_6_), .B2(n5048), .ZN(n4830) );
  AOI22D1BWP12T U4121 ( .A1(n5051), .A2(RF_next_sp[6]), .B1(
        register_file_inst1_r7_6_), .B2(n5050), .ZN(n4829) );
  AOI22D0BWP12T U4122 ( .A1(n5053), .A2(register_file_inst1_r6_6_), .B1(
        register_file_inst1_r2_6_), .B2(n5052), .ZN(n4828) );
  ND4D1BWP12T U4123 ( .A1(n6264), .A2(n4830), .A3(n4829), .A4(n4828), .ZN(
        n4831) );
  OAI21D1BWP12T U4124 ( .A1(n4832), .A2(n4831), .B(n6397), .ZN(n4833) );
  ND2D1BWP12T U4125 ( .A1(n3165), .A2(n4833), .ZN(MEMCTRL_IN_address[5]) );
  AOI22D1BWP12T U4126 ( .A1(memory_interface_inst1_delay_addr_single[5]), .A2(
        n6294), .B1(MEMCTRL_IN_address[5]), .B2(n6295), .ZN(n4837) );
  AO211D1BWP12T U4127 ( .A1(n4858), .A2(n4835), .B(n4834), .C(n4888), .Z(n4836) );
  ND2D1BWP12T U4128 ( .A1(n4837), .A2(n4836), .ZN(
        MEMCTRL_MEM_to_mem_address[5]) );
  INVD1BWP12T U4129 ( .I(n6398), .ZN(n4840) );
  IND3D1BWP12T U4130 ( .A1(n4838), .B1(n4841), .B2(n6235), .ZN(n4839) );
  ND2D1BWP12T U4131 ( .A1(n4840), .A2(n4839), .ZN(n4892) );
  INVD1BWP12T U4132 ( .I(n4892), .ZN(n4934) );
  AOI22D0BWP12T U4133 ( .A1(n5180), .A2(
        memory_interface_inst1_delay_data_in32[23]), .B1(n4934), .B2(
        memory_interface_inst1_delay_data_in32[7]), .ZN(n4843) );
  AN2D1BWP12T U4134 ( .A1(n6398), .A2(n4841), .Z(n4935) );
  AOI22D0BWP12T U4135 ( .A1(n6282), .A2(RF_MEMCTRL_data_reg[7]), .B1(n4935), 
        .B2(RF_MEMCTRL_data_reg[23]), .ZN(n4842) );
  ND2D1BWP12T U4136 ( .A1(n4843), .A2(n4842), .ZN(MEMCTRL_MEM_to_mem_data[15])
         );
  AOI22D0BWP12T U4137 ( .A1(n5180), .A2(
        memory_interface_inst1_delay_data_in32[22]), .B1(n4934), .B2(
        memory_interface_inst1_delay_data_in32[6]), .ZN(n4845) );
  AOI22D0BWP12T U4138 ( .A1(n6282), .A2(RF_MEMCTRL_data_reg[6]), .B1(n4935), 
        .B2(RF_MEMCTRL_data_reg[22]), .ZN(n4844) );
  ND2D1BWP12T U4139 ( .A1(n4845), .A2(n4844), .ZN(MEMCTRL_MEM_to_mem_data[14])
         );
  AOI22D0BWP12T U4140 ( .A1(n5180), .A2(
        memory_interface_inst1_delay_data_in32[21]), .B1(n4934), .B2(
        memory_interface_inst1_delay_data_in32[5]), .ZN(n4847) );
  AOI22D0BWP12T U4141 ( .A1(n6282), .A2(RF_MEMCTRL_data_reg[5]), .B1(n4935), 
        .B2(RF_MEMCTRL_data_reg[21]), .ZN(n4846) );
  ND2D1BWP12T U4142 ( .A1(n4847), .A2(n4846), .ZN(MEMCTRL_MEM_to_mem_data[13])
         );
  AOI22D1BWP12T U4143 ( .A1(n5058), .A2(register_file_inst1_r3_5_), .B1(
        register_file_inst1_r12_5_), .B2(n5057), .ZN(n4851) );
  AOI22D0BWP12T U4144 ( .A1(n5060), .A2(register_file_inst1_r4_5_), .B1(
        register_file_inst1_r8_5_), .B2(n5059), .ZN(n4850) );
  AOI22D0BWP12T U4145 ( .A1(n5062), .A2(register_file_inst1_r0_5_), .B1(
        register_file_inst1_r1_5_), .B2(n5061), .ZN(n4849) );
  AOI22D1BWP12T U4146 ( .A1(n5064), .A2(register_file_inst1_r10_5_), .B1(
        register_file_inst1_r11_5_), .B2(n5063), .ZN(n4848) );
  ND4D1BWP12T U4147 ( .A1(n4851), .A2(n4850), .A3(n4849), .A4(n4848), .ZN(
        n4856) );
  AOI22D0BWP12T U4148 ( .A1(n5049), .A2(register_file_inst1_lr_5_), .B1(
        register_file_inst1_r9_5_), .B2(n5048), .ZN(n4854) );
  AOI22D0BWP12T U4149 ( .A1(n5051), .A2(RF_next_sp[5]), .B1(
        register_file_inst1_r7_5_), .B2(n5050), .ZN(n4853) );
  AOI22D0BWP12T U4150 ( .A1(n5053), .A2(register_file_inst1_r6_5_), .B1(
        register_file_inst1_r2_5_), .B2(n5052), .ZN(n4852) );
  ND4D1BWP12T U4151 ( .A1(n6251), .A2(n4854), .A3(n4853), .A4(n4852), .ZN(
        n4855) );
  OAI21D1BWP12T U4152 ( .A1(n4856), .A2(n4855), .B(n6397), .ZN(n4857) );
  ND2D1BWP12T U4153 ( .A1(n3286), .A2(n4857), .ZN(MEMCTRL_IN_address[4]) );
  AOI22D1BWP12T U4154 ( .A1(memory_interface_inst1_delay_addr_single[4]), .A2(
        n6294), .B1(MEMCTRL_IN_address[4]), .B2(n6295), .ZN(n4860) );
  OAI211D1BWP12T U4155 ( .A1(n4873), .A2(
        memory_interface_inst1_delay_addr_for_adder_4_), .B(n4928), .C(n4858), 
        .ZN(n4859) );
  ND2D1BWP12T U4156 ( .A1(n4860), .A2(n4859), .ZN(
        MEMCTRL_MEM_to_mem_address[4]) );
  AOI22D0BWP12T U4157 ( .A1(n5180), .A2(
        memory_interface_inst1_delay_data_in32[20]), .B1(n4934), .B2(
        memory_interface_inst1_delay_data_in32[4]), .ZN(n4862) );
  AOI22D0BWP12T U4158 ( .A1(n6282), .A2(RF_MEMCTRL_data_reg[4]), .B1(n4935), 
        .B2(RF_MEMCTRL_data_reg[20]), .ZN(n4861) );
  ND2D1BWP12T U4159 ( .A1(n4862), .A2(n4861), .ZN(MEMCTRL_MEM_to_mem_data[12])
         );
  AOI22D0BWP12T U4160 ( .A1(n5058), .A2(register_file_inst1_r3_4_), .B1(
        register_file_inst1_r12_4_), .B2(n5057), .ZN(n4866) );
  AOI22D0BWP12T U4161 ( .A1(n5060), .A2(register_file_inst1_r4_4_), .B1(
        register_file_inst1_r8_4_), .B2(n5059), .ZN(n4865) );
  AOI22D0BWP12T U4162 ( .A1(n5062), .A2(register_file_inst1_r0_4_), .B1(
        register_file_inst1_r1_4_), .B2(n5061), .ZN(n4864) );
  AOI22D0BWP12T U4163 ( .A1(n5064), .A2(register_file_inst1_r10_4_), .B1(
        register_file_inst1_r11_4_), .B2(n5063), .ZN(n4863) );
  ND4D1BWP12T U4164 ( .A1(n4866), .A2(n4865), .A3(n4864), .A4(n4863), .ZN(
        n4871) );
  AOI22D0BWP12T U4165 ( .A1(n5049), .A2(register_file_inst1_lr_4_), .B1(
        register_file_inst1_r9_4_), .B2(n5048), .ZN(n4869) );
  AOI22D0BWP12T U4166 ( .A1(n5051), .A2(RF_next_sp[4]), .B1(
        register_file_inst1_r7_4_), .B2(n5050), .ZN(n4868) );
  AOI22D0BWP12T U4167 ( .A1(n5053), .A2(register_file_inst1_r6_4_), .B1(
        register_file_inst1_r2_4_), .B2(n5052), .ZN(n4867) );
  ND4D1BWP12T U4168 ( .A1(n6236), .A2(n4869), .A3(n4868), .A4(n4867), .ZN(
        n4870) );
  OAI21D1BWP12T U4169 ( .A1(n4871), .A2(n4870), .B(n6397), .ZN(n4872) );
  ND2D1BWP12T U4170 ( .A1(n3467), .A2(n4872), .ZN(MEMCTRL_IN_address[3]) );
  AOI22D1BWP12T U4171 ( .A1(memory_interface_inst1_delay_addr_single[3]), .A2(
        n6294), .B1(MEMCTRL_IN_address[3]), .B2(n6295), .ZN(n4877) );
  AO211D1BWP12T U4172 ( .A1(n4875), .A2(n4874), .B(n4873), .C(n4888), .Z(n4876) );
  ND2D1BWP12T U4173 ( .A1(n4877), .A2(n4876), .ZN(
        MEMCTRL_MEM_to_mem_address[3]) );
  AOI22D0BWP12T U4174 ( .A1(n5058), .A2(register_file_inst1_r3_10_), .B1(
        register_file_inst1_r12_10_), .B2(n5057), .ZN(n4881) );
  AOI22D0BWP12T U4175 ( .A1(n5060), .A2(register_file_inst1_r4_10_), .B1(
        register_file_inst1_r8_10_), .B2(n5059), .ZN(n4880) );
  AOI22D0BWP12T U4176 ( .A1(n5062), .A2(register_file_inst1_r0_10_), .B1(
        register_file_inst1_r1_10_), .B2(n5061), .ZN(n4879) );
  AOI22D0BWP12T U4177 ( .A1(n5064), .A2(register_file_inst1_r10_10_), .B1(
        register_file_inst1_r11_10_), .B2(n5063), .ZN(n4878) );
  ND4D1BWP12T U4178 ( .A1(n4881), .A2(n4880), .A3(n4879), .A4(n4878), .ZN(
        n4886) );
  AOI22D0BWP12T U4179 ( .A1(n5049), .A2(register_file_inst1_lr_10_), .B1(
        register_file_inst1_r9_10_), .B2(n5048), .ZN(n4884) );
  AOI22D0BWP12T U4180 ( .A1(n5051), .A2(RF_next_sp[10]), .B1(
        register_file_inst1_r7_10_), .B2(n5050), .ZN(n4883) );
  AOI22D0BWP12T U4181 ( .A1(n5053), .A2(register_file_inst1_r6_10_), .B1(
        register_file_inst1_r2_10_), .B2(n5052), .ZN(n4882) );
  ND4D1BWP12T U4182 ( .A1(n6239), .A2(n4884), .A3(n4883), .A4(n4882), .ZN(
        n4885) );
  OAI21D1BWP12T U4183 ( .A1(n4886), .A2(n4885), .B(n6397), .ZN(n4887) );
  ND2D1BWP12T U4184 ( .A1(n3420), .A2(n4887), .ZN(MEMCTRL_IN_address[9]) );
  AOI22D1BWP12T U4185 ( .A1(MEMCTRL_IN_address[9]), .A2(n6295), .B1(n6294), 
        .B2(memory_interface_inst1_delay_addr_single[9]), .ZN(n4891) );
  ND2D1BWP12T U4186 ( .A1(n4912), .A2(
        memory_interface_inst1_delay_addr_for_adder_8_), .ZN(n4911) );
  INVD1BWP12T U4187 ( .I(memory_interface_inst1_delay_addr_for_adder_9_), .ZN(
        n4889) );
  NR2D1BWP12T U4188 ( .A1(n4911), .A2(n4889), .ZN(n4927) );
  AO211D1BWP12T U4189 ( .A1(n4911), .A2(n4889), .B(n4927), .C(n4888), .Z(n4890) );
  ND2D1BWP12T U4190 ( .A1(n4891), .A2(n4890), .ZN(
        MEMCTRL_MEM_to_mem_address[9]) );
  AOI22D0BWP12T U4191 ( .A1(n5180), .A2(
        memory_interface_inst1_delay_data_in32[28]), .B1(
        MEM_MEMCTRL_from_mem_data[4]), .B2(n6294), .ZN(n4894) );
  NR2D1BWP12T U4192 ( .A1(n4892), .A2(n6294), .ZN(n4931) );
  AOI22D0BWP12T U4193 ( .A1(n6282), .A2(RF_MEMCTRL_data_reg[12]), .B1(n4931), 
        .B2(memory_interface_inst1_delay_data_in32[12]), .ZN(n4893) );
  ND2D1BWP12T U4194 ( .A1(n4894), .A2(n4893), .ZN(MEMCTRL_MEM_to_mem_data[4])
         );
  AOI22D0BWP12T U4195 ( .A1(n5180), .A2(
        memory_interface_inst1_delay_data_in32[27]), .B1(
        MEM_MEMCTRL_from_mem_data[3]), .B2(n6294), .ZN(n4896) );
  AOI22D0BWP12T U4196 ( .A1(n6282), .A2(RF_MEMCTRL_data_reg[11]), .B1(n4931), 
        .B2(memory_interface_inst1_delay_data_in32[11]), .ZN(n4895) );
  ND2D1BWP12T U4197 ( .A1(n4896), .A2(n4895), .ZN(MEMCTRL_MEM_to_mem_data[3])
         );
  AOI22D0BWP12T U4198 ( .A1(n5180), .A2(
        memory_interface_inst1_delay_data_in32[24]), .B1(
        MEM_MEMCTRL_from_mem_data[0]), .B2(n6294), .ZN(n4898) );
  AOI22D0BWP12T U4199 ( .A1(n6282), .A2(RF_MEMCTRL_data_reg[8]), .B1(n4931), 
        .B2(memory_interface_inst1_delay_data_in32[8]), .ZN(n4897) );
  ND2D1BWP12T U4200 ( .A1(n4898), .A2(n4897), .ZN(MEMCTRL_MEM_to_mem_data[0])
         );
  AOI22D0BWP12T U4201 ( .A1(n5180), .A2(
        memory_interface_inst1_delay_data_in32[25]), .B1(
        MEM_MEMCTRL_from_mem_data[1]), .B2(n6294), .ZN(n4900) );
  AOI22D0BWP12T U4202 ( .A1(n6282), .A2(RF_MEMCTRL_data_reg[9]), .B1(n4931), 
        .B2(memory_interface_inst1_delay_data_in32[9]), .ZN(n4899) );
  ND2D1BWP12T U4203 ( .A1(n4900), .A2(n4899), .ZN(MEMCTRL_MEM_to_mem_data[1])
         );
  AOI22D1BWP12T U4204 ( .A1(n5058), .A2(register_file_inst1_r3_9_), .B1(
        register_file_inst1_r12_9_), .B2(n5057), .ZN(n4904) );
  AOI22D0BWP12T U4205 ( .A1(n5060), .A2(register_file_inst1_r4_9_), .B1(
        register_file_inst1_r8_9_), .B2(n5059), .ZN(n4903) );
  AOI22D1BWP12T U4206 ( .A1(n5062), .A2(register_file_inst1_r0_9_), .B1(
        register_file_inst1_r1_9_), .B2(n5061), .ZN(n4902) );
  AOI22D1BWP12T U4207 ( .A1(n5064), .A2(register_file_inst1_r10_9_), .B1(
        register_file_inst1_r11_9_), .B2(n5063), .ZN(n4901) );
  ND4D1BWP12T U4208 ( .A1(n4904), .A2(n4903), .A3(n4902), .A4(n4901), .ZN(
        n4909) );
  AOI22D1BWP12T U4209 ( .A1(n5049), .A2(register_file_inst1_lr_9_), .B1(
        register_file_inst1_r9_9_), .B2(n5048), .ZN(n4907) );
  AOI22D0BWP12T U4210 ( .A1(n5051), .A2(RF_next_sp[9]), .B1(
        register_file_inst1_r2_9_), .B2(n5052), .ZN(n4906) );
  AOI22D0BWP12T U4211 ( .A1(n5050), .A2(register_file_inst1_r7_9_), .B1(
        register_file_inst1_r6_9_), .B2(n5053), .ZN(n4905) );
  ND4D1BWP12T U4212 ( .A1(n6278), .A2(n4907), .A3(n4906), .A4(n4905), .ZN(
        n4908) );
  OAI21D1BWP12T U4213 ( .A1(n4909), .A2(n4908), .B(n6397), .ZN(n4910) );
  ND2D1BWP12T U4214 ( .A1(n3068), .A2(n4910), .ZN(MEMCTRL_IN_address[8]) );
  AOI22D1BWP12T U4215 ( .A1(memory_interface_inst1_delay_addr_single[8]), .A2(
        n6294), .B1(MEMCTRL_IN_address[8]), .B2(n6295), .ZN(n4914) );
  OAI211D1BWP12T U4216 ( .A1(n4912), .A2(
        memory_interface_inst1_delay_addr_for_adder_8_), .B(n4928), .C(n4911), 
        .ZN(n4913) );
  ND2D1BWP12T U4217 ( .A1(n4914), .A2(n4913), .ZN(
        MEMCTRL_MEM_to_mem_address[8]) );
  AOI22D0BWP12T U4218 ( .A1(n5180), .A2(
        memory_interface_inst1_delay_data_in32[29]), .B1(
        MEM_MEMCTRL_from_mem_data[5]), .B2(n6294), .ZN(n4916) );
  AOI22D0BWP12T U4219 ( .A1(n6282), .A2(RF_MEMCTRL_data_reg[13]), .B1(n4931), 
        .B2(memory_interface_inst1_delay_data_in32[13]), .ZN(n4915) );
  ND2D1BWP12T U4220 ( .A1(n4916), .A2(n4915), .ZN(MEMCTRL_MEM_to_mem_data[5])
         );
  AOI22D0BWP12T U4221 ( .A1(n5180), .A2(
        memory_interface_inst1_delay_data_in32[16]), .B1(n4934), .B2(
        memory_interface_inst1_delay_data_in32[0]), .ZN(n4918) );
  AOI22D0BWP12T U4222 ( .A1(n6282), .A2(RF_MEMCTRL_data_reg[0]), .B1(n4935), 
        .B2(RF_MEMCTRL_data_reg[16]), .ZN(n4917) );
  ND2D1BWP12T U4223 ( .A1(n4918), .A2(n4917), .ZN(MEMCTRL_MEM_to_mem_data[8])
         );
  AOI22D0BWP12T U4224 ( .A1(n5180), .A2(
        memory_interface_inst1_delay_data_in32[19]), .B1(n4934), .B2(
        memory_interface_inst1_delay_data_in32[3]), .ZN(n4920) );
  AOI22D0BWP12T U4225 ( .A1(n6282), .A2(RF_MEMCTRL_data_reg[3]), .B1(n4935), 
        .B2(RF_MEMCTRL_data_reg[19]), .ZN(n4919) );
  ND2D1BWP12T U4226 ( .A1(n4920), .A2(n4919), .ZN(MEMCTRL_MEM_to_mem_data[11])
         );
  AOI22D0BWP12T U4227 ( .A1(n5180), .A2(
        memory_interface_inst1_delay_data_in32[30]), .B1(
        MEM_MEMCTRL_from_mem_data[6]), .B2(n6294), .ZN(n4922) );
  AOI22D0BWP12T U4228 ( .A1(n6282), .A2(RF_MEMCTRL_data_reg[14]), .B1(n4931), 
        .B2(memory_interface_inst1_delay_data_in32[14]), .ZN(n4921) );
  ND2D1BWP12T U4229 ( .A1(n4922), .A2(n4921), .ZN(MEMCTRL_MEM_to_mem_data[6])
         );
  AOI22D0BWP12T U4230 ( .A1(n5180), .A2(
        memory_interface_inst1_delay_data_in32[26]), .B1(
        MEM_MEMCTRL_from_mem_data[2]), .B2(n6294), .ZN(n4924) );
  AOI22D0BWP12T U4231 ( .A1(n6282), .A2(RF_MEMCTRL_data_reg[10]), .B1(n4931), 
        .B2(memory_interface_inst1_delay_data_in32[10]), .ZN(n4923) );
  ND2D1BWP12T U4232 ( .A1(n4924), .A2(n4923), .ZN(MEMCTRL_MEM_to_mem_data[2])
         );
  ND2D1BWP12T U4233 ( .A1(ALU_MISC_OUT_result[12]), .A2(n6396), .ZN(n4925) );
  ND2D1BWP12T U4234 ( .A1(n4925), .A2(n6293), .ZN(MEMCTRL_IN_address[11]) );
  ND2D1BWP12T U4235 ( .A1(ALU_MISC_OUT_result[11]), .A2(n6396), .ZN(n4926) );
  ND2D1BWP12T U4236 ( .A1(n4926), .A2(n6290), .ZN(MEMCTRL_IN_address[10]) );
  AOI22D0BWP12T U4237 ( .A1(n5180), .A2(
        memory_interface_inst1_delay_data_in32[17]), .B1(n4934), .B2(
        memory_interface_inst1_delay_data_in32[1]), .ZN(n4930) );
  AOI22D0BWP12T U4238 ( .A1(n6282), .A2(RF_MEMCTRL_data_reg[1]), .B1(n4935), 
        .B2(RF_MEMCTRL_data_reg[17]), .ZN(n4929) );
  ND2D1BWP12T U4239 ( .A1(n4930), .A2(n4929), .ZN(MEMCTRL_MEM_to_mem_data[9])
         );
  AOI22D0BWP12T U4240 ( .A1(n5180), .A2(
        memory_interface_inst1_delay_data_in32[31]), .B1(
        MEM_MEMCTRL_from_mem_data[7]), .B2(n6294), .ZN(n4933) );
  AOI22D0BWP12T U4241 ( .A1(n6282), .A2(RF_MEMCTRL_data_reg[15]), .B1(n4931), 
        .B2(memory_interface_inst1_delay_data_in32[15]), .ZN(n4932) );
  ND2D1BWP12T U4242 ( .A1(n4933), .A2(n4932), .ZN(MEMCTRL_MEM_to_mem_data[7])
         );
  AOI22D0BWP12T U4243 ( .A1(n5180), .A2(
        memory_interface_inst1_delay_data_in32[18]), .B1(n4934), .B2(
        memory_interface_inst1_delay_data_in32[2]), .ZN(n4937) );
  AOI22D0BWP12T U4244 ( .A1(n6282), .A2(RF_MEMCTRL_data_reg[2]), .B1(n4935), 
        .B2(RF_MEMCTRL_data_reg[18]), .ZN(n4936) );
  ND2D1BWP12T U4245 ( .A1(n4937), .A2(n4936), .ZN(MEMCTRL_MEM_to_mem_data[10])
         );
  AOI22D0BWP12T U4246 ( .A1(register_file_inst1_r1_24_), .A2(n5001), .B1(
        register_file_inst1_r3_24_), .B2(n4989), .ZN(n4941) );
  AOI22D0BWP12T U4247 ( .A1(register_file_inst1_r2_24_), .A2(n4962), .B1(
        register_file_inst1_r0_24_), .B2(n5002), .ZN(n4940) );
  AOI22D0BWP12T U4248 ( .A1(register_file_inst1_r4_24_), .A2(n5003), .B1(
        register_file_inst1_r5_24_), .B2(n4990), .ZN(n4939) );
  AOI22D0BWP12T U4249 ( .A1(register_file_inst1_r6_24_), .A2(n5004), .B1(
        register_file_inst1_r7_24_), .B2(n4991), .ZN(n4938) );
  ND4D1BWP12T U4250 ( .A1(n4941), .A2(n4940), .A3(n4939), .A4(n4938), .ZN(
        n4942) );
  ND2D1BWP12T U4251 ( .A1(n4942), .A2(n3502), .ZN(n4945) );
  AOI22D0BWP12T U4252 ( .A1(register_file_inst1_lr_24_), .A2(n4437), .B1(
        RF_next_sp[24]), .B2(n5010), .ZN(n4944) );
  AOI22D0BWP12T U4253 ( .A1(register_file_inst1_r9_24_), .A2(n6005), .B1(
        register_file_inst1_r10_24_), .B2(n5011), .ZN(n4943) );
  ND4D1BWP12T U4254 ( .A1(n4945), .A2(n6276), .A3(n4944), .A4(n4943), .ZN(
        RF_MEMCTRL_data_reg[24]) );
  AOI22D0BWP12T U4255 ( .A1(register_file_inst1_r1_28_), .A2(n5001), .B1(
        register_file_inst1_r3_28_), .B2(n4989), .ZN(n4949) );
  AOI22D0BWP12T U4256 ( .A1(register_file_inst1_r2_28_), .A2(n4962), .B1(
        register_file_inst1_r0_28_), .B2(n5002), .ZN(n4948) );
  AOI22D0BWP12T U4257 ( .A1(register_file_inst1_r4_28_), .A2(n5003), .B1(
        register_file_inst1_r5_28_), .B2(n4990), .ZN(n4947) );
  AOI22D0BWP12T U4258 ( .A1(register_file_inst1_r6_28_), .A2(n5004), .B1(
        register_file_inst1_r7_28_), .B2(n4991), .ZN(n4946) );
  ND4D1BWP12T U4259 ( .A1(n4949), .A2(n4948), .A3(n4947), .A4(n4946), .ZN(
        n4950) );
  ND2D1BWP12T U4260 ( .A1(n4950), .A2(n3502), .ZN(n4953) );
  AOI22D0BWP12T U4261 ( .A1(register_file_inst1_lr_28_), .A2(n4437), .B1(
        RF_next_sp[28]), .B2(n5010), .ZN(n4952) );
  AOI22D0BWP12T U4262 ( .A1(register_file_inst1_r9_28_), .A2(n6005), .B1(
        register_file_inst1_r10_28_), .B2(n5011), .ZN(n4951) );
  ND4D1BWP12T U4263 ( .A1(n4953), .A2(n6254), .A3(n4952), .A4(n4951), .ZN(
        RF_MEMCTRL_data_reg[28]) );
  AOI22D0BWP12T U4264 ( .A1(register_file_inst1_r1_30_), .A2(n5001), .B1(
        register_file_inst1_r3_30_), .B2(n4989), .ZN(n4957) );
  AOI22D0BWP12T U4265 ( .A1(register_file_inst1_r2_30_), .A2(n4962), .B1(
        register_file_inst1_r0_30_), .B2(n5002), .ZN(n4956) );
  AOI22D0BWP12T U4266 ( .A1(register_file_inst1_r4_30_), .A2(n5003), .B1(
        register_file_inst1_r5_30_), .B2(n4990), .ZN(n4955) );
  AOI22D0BWP12T U4267 ( .A1(register_file_inst1_r6_30_), .A2(n5004), .B1(
        register_file_inst1_r7_30_), .B2(n4991), .ZN(n4954) );
  ND4D1BWP12T U4268 ( .A1(n4957), .A2(n4956), .A3(n4955), .A4(n4954), .ZN(
        n4958) );
  ND2D1BWP12T U4269 ( .A1(n4958), .A2(n3502), .ZN(n4961) );
  AOI22D0BWP12T U4270 ( .A1(register_file_inst1_lr_30_), .A2(n4437), .B1(
        RF_next_sp[30]), .B2(n5010), .ZN(n4960) );
  AOI22D0BWP12T U4271 ( .A1(register_file_inst1_r9_30_), .A2(n6005), .B1(
        register_file_inst1_r10_30_), .B2(n5011), .ZN(n4959) );
  ND4D1BWP12T U4272 ( .A1(n4961), .A2(n6258), .A3(n4960), .A4(n4959), .ZN(
        RF_MEMCTRL_data_reg[30]) );
  AOI22D0BWP12T U4273 ( .A1(register_file_inst1_r1_31_), .A2(n5001), .B1(
        register_file_inst1_r3_31_), .B2(n4989), .ZN(n4966) );
  AOI22D0BWP12T U4274 ( .A1(register_file_inst1_r2_31_), .A2(n4962), .B1(
        register_file_inst1_r0_31_), .B2(n5002), .ZN(n4965) );
  AOI22D0BWP12T U4275 ( .A1(register_file_inst1_r4_31_), .A2(n5003), .B1(
        register_file_inst1_r5_31_), .B2(n4990), .ZN(n4964) );
  AOI22D0BWP12T U4276 ( .A1(register_file_inst1_r6_31_), .A2(n5004), .B1(
        register_file_inst1_r7_31_), .B2(n4991), .ZN(n4963) );
  ND4D1BWP12T U4277 ( .A1(n4966), .A2(n4965), .A3(n4964), .A4(n4963), .ZN(
        n4967) );
  ND2D1BWP12T U4278 ( .A1(n4967), .A2(n3502), .ZN(n4970) );
  AOI22D0BWP12T U4279 ( .A1(register_file_inst1_lr_31_), .A2(n4437), .B1(
        RF_next_sp[31]), .B2(n5010), .ZN(n4969) );
  AOI22D0BWP12T U4280 ( .A1(register_file_inst1_r9_31_), .A2(n6005), .B1(
        register_file_inst1_r10_31_), .B2(n5011), .ZN(n4968) );
  ND4D1BWP12T U4281 ( .A1(n4970), .A2(n6267), .A3(n4969), .A4(n4968), .ZN(
        RF_MEMCTRL_data_reg[31]) );
  AOI22D0BWP12T U4282 ( .A1(register_file_inst1_r1_26_), .A2(n5001), .B1(
        register_file_inst1_r3_26_), .B2(n4989), .ZN(n4974) );
  AOI22D0BWP12T U4283 ( .A1(register_file_inst1_r2_26_), .A2(n4962), .B1(
        register_file_inst1_r0_26_), .B2(n5002), .ZN(n4973) );
  AOI22D0BWP12T U4284 ( .A1(register_file_inst1_r4_26_), .A2(n5003), .B1(
        register_file_inst1_r5_26_), .B2(n4990), .ZN(n4972) );
  AOI22D0BWP12T U4285 ( .A1(register_file_inst1_r6_26_), .A2(n5004), .B1(
        register_file_inst1_r7_26_), .B2(n4991), .ZN(n4971) );
  ND4D1BWP12T U4286 ( .A1(n4974), .A2(n4973), .A3(n4972), .A4(n4971), .ZN(
        n4979) );
  AOI22D1BWP12T U4287 ( .A1(register_file_inst1_lr_26_), .A2(n4437), .B1(
        register_file_inst1_r12_26_), .B2(n4510), .ZN(n4977) );
  AOI22D1BWP12T U4288 ( .A1(RF_next_sp[26]), .A2(n5010), .B1(
        register_file_inst1_r11_26_), .B2(n5009), .ZN(n4976) );
  AOI22D0BWP12T U4289 ( .A1(register_file_inst1_r9_26_), .A2(n6005), .B1(
        register_file_inst1_r10_26_), .B2(n5011), .ZN(n4975) );
  ND4D1BWP12T U4290 ( .A1(n6249), .A2(n4977), .A3(n4976), .A4(n4975), .ZN(
        n4978) );
  AO21D1BWP12T U4291 ( .A1(n3502), .A2(n4979), .B(n4978), .Z(
        RF_MEMCTRL_data_reg[26]) );
  AOI22D0BWP12T U4292 ( .A1(register_file_inst1_r1_29_), .A2(n5001), .B1(
        register_file_inst1_r3_29_), .B2(n4989), .ZN(n4983) );
  AOI22D0BWP12T U4293 ( .A1(register_file_inst1_r2_29_), .A2(n4962), .B1(
        register_file_inst1_r0_29_), .B2(n5002), .ZN(n4982) );
  AOI22D0BWP12T U4294 ( .A1(register_file_inst1_r4_29_), .A2(n5003), .B1(
        register_file_inst1_r5_29_), .B2(n4990), .ZN(n4981) );
  AOI22D0BWP12T U4295 ( .A1(register_file_inst1_r6_29_), .A2(n5004), .B1(
        register_file_inst1_r7_29_), .B2(n4991), .ZN(n4980) );
  ND4D1BWP12T U4296 ( .A1(n4983), .A2(n4982), .A3(n4981), .A4(n4980), .ZN(
        n4988) );
  AOI22D1BWP12T U4297 ( .A1(register_file_inst1_lr_29_), .A2(n4437), .B1(
        register_file_inst1_r12_29_), .B2(n4510), .ZN(n4986) );
  AOI22D1BWP12T U4298 ( .A1(RF_next_sp[29]), .A2(n5010), .B1(
        register_file_inst1_r11_29_), .B2(n5009), .ZN(n4985) );
  AOI22D0BWP12T U4299 ( .A1(register_file_inst1_r9_29_), .A2(n6005), .B1(
        register_file_inst1_r10_29_), .B2(n5011), .ZN(n4984) );
  ND4D1BWP12T U4300 ( .A1(n6285), .A2(n4986), .A3(n4985), .A4(n4984), .ZN(
        n4987) );
  AO21D1BWP12T U4301 ( .A1(n3502), .A2(n4988), .B(n4987), .Z(
        RF_MEMCTRL_data_reg[29]) );
  AOI22D0BWP12T U4302 ( .A1(register_file_inst1_r1_27_), .A2(n5001), .B1(
        register_file_inst1_r3_27_), .B2(n4989), .ZN(n4995) );
  AOI22D0BWP12T U4303 ( .A1(register_file_inst1_r2_27_), .A2(n4962), .B1(
        register_file_inst1_r0_27_), .B2(n5002), .ZN(n4994) );
  AOI22D0BWP12T U4304 ( .A1(register_file_inst1_r4_27_), .A2(n5003), .B1(
        register_file_inst1_r5_27_), .B2(n4990), .ZN(n4993) );
  AOI22D0BWP12T U4305 ( .A1(register_file_inst1_r6_27_), .A2(n5004), .B1(
        register_file_inst1_r7_27_), .B2(n4991), .ZN(n4992) );
  ND4D1BWP12T U4306 ( .A1(n4995), .A2(n4994), .A3(n4993), .A4(n4992), .ZN(
        n5000) );
  AOI22D1BWP12T U4307 ( .A1(register_file_inst1_lr_27_), .A2(n4437), .B1(
        register_file_inst1_r12_27_), .B2(n4510), .ZN(n4998) );
  AOI22D1BWP12T U4308 ( .A1(RF_next_sp[27]), .A2(n5010), .B1(
        register_file_inst1_r11_27_), .B2(n5009), .ZN(n4997) );
  AOI22D0BWP12T U4309 ( .A1(register_file_inst1_r9_27_), .A2(n6005), .B1(
        register_file_inst1_r10_27_), .B2(n5011), .ZN(n4996) );
  ND4D1BWP12T U4310 ( .A1(n6284), .A2(n4998), .A3(n4997), .A4(n4996), .ZN(
        n4999) );
  AO21D1BWP12T U4311 ( .A1(n3502), .A2(n5000), .B(n4999), .Z(
        RF_MEMCTRL_data_reg[27]) );
  AOI22D0BWP12T U4312 ( .A1(register_file_inst1_r1_25_), .A2(n5001), .B1(
        register_file_inst1_r3_25_), .B2(n4989), .ZN(n5008) );
  AOI22D0BWP12T U4313 ( .A1(register_file_inst1_r2_25_), .A2(n4962), .B1(
        register_file_inst1_r0_25_), .B2(n5002), .ZN(n5007) );
  AOI22D0BWP12T U4314 ( .A1(register_file_inst1_r4_25_), .A2(n5003), .B1(
        register_file_inst1_r5_25_), .B2(n4990), .ZN(n5006) );
  AOI22D0BWP12T U4315 ( .A1(register_file_inst1_r6_25_), .A2(n5004), .B1(
        register_file_inst1_r7_25_), .B2(n4991), .ZN(n5005) );
  ND4D1BWP12T U4316 ( .A1(n5008), .A2(n5007), .A3(n5006), .A4(n5005), .ZN(
        n5016) );
  AOI22D1BWP12T U4317 ( .A1(register_file_inst1_lr_25_), .A2(n4437), .B1(
        register_file_inst1_r12_25_), .B2(n4510), .ZN(n5014) );
  AOI22D1BWP12T U4318 ( .A1(RF_next_sp[25]), .A2(n5010), .B1(
        register_file_inst1_r11_25_), .B2(n5009), .ZN(n5013) );
  AOI22D0BWP12T U4319 ( .A1(register_file_inst1_r9_25_), .A2(n6005), .B1(
        register_file_inst1_r10_25_), .B2(n5011), .ZN(n5012) );
  ND4D1BWP12T U4320 ( .A1(n6283), .A2(n5014), .A3(n5013), .A4(n5012), .ZN(
        n5015) );
  AO21D1BWP12T U4321 ( .A1(n3502), .A2(n5016), .B(n5015), .Z(
        RF_MEMCTRL_data_reg[25]) );
  OA21D1BWP12T U4322 ( .A1(n6111), .A2(n5017), .B(n6391), .Z(
        memory_interface_inst1_fsm_N35) );
  NR2D1BWP12T U4323 ( .A1(n6304), .A2(n5233), .ZN(n6070) );
  NR2D1BWP12T U4324 ( .A1(n6303), .A2(n5233), .ZN(n6066) );
  NR2D1BWP12T U4325 ( .A1(n6367), .A2(n5233), .ZN(n6074) );
  NR2D1BWP12T U4326 ( .A1(n6063), .A2(n5233), .ZN(n6061) );
  NR2D1BWP12T U4327 ( .A1(n6302), .A2(n5233), .ZN(n6057) );
  NR2D1BWP12T U4328 ( .A1(n6054), .A2(n5233), .ZN(n6052) );
  OAI222D1BWP12T U4329 ( .A1(n3718), .A2(n5212), .B1(n5020), .B2(n6144), .C1(
        n4683), .C2(n5018), .ZN(register_file_inst1_n2136) );
  INVD1BWP12T U4330 ( .I(n5021), .ZN(n5019) );
  OAI211D1BWP12T U4331 ( .A1(n6386), .A2(n5019), .B(n6385), .C(n6384), .ZN(
        register_file_inst1_n2170) );
  NR2D1BWP12T U4332 ( .A1(n6349), .A2(n5233), .ZN(n6096) );
  AOI22D1BWP12T U4333 ( .A1(n5984), .A2(n3718), .B1(n5020), .B2(n6008), .ZN(
        n2396) );
  NR2D1BWP12T U4334 ( .A1(n6307), .A2(n5233), .ZN(n6082) );
  NR2D1BWP12T U4335 ( .A1(n6352), .A2(n5233), .ZN(n6092) );
  OAI21D1BWP12T U4336 ( .A1(n5984), .A2(n5022), .B(n5021), .ZN(n6380) );
  OAI21D1BWP12T U4337 ( .A1(n5984), .A2(n5023), .B(n6378), .ZN(n6372) );
  OAI21D1BWP12T U4338 ( .A1(n5034), .A2(n5234), .B(n6075), .ZN(
        register_file_inst1_spin[6]) );
  INVD1BWP12T U4339 ( .I(register_file_inst1_r11_6_), .ZN(n5024) );
  OAI222D1BWP12T U4340 ( .A1(n5034), .A2(n5220), .B1(n5219), .B2(n6367), .C1(
        n5217), .C2(n5024), .ZN(register_file_inst1_n2271) );
  CKND0BWP12T U4341 ( .I(register_file_inst1_tmp1_6_), .ZN(n5025) );
  OAI222D1BWP12T U4342 ( .A1(n5034), .A2(n6144), .B1(n5212), .B2(n6367), .C1(
        n4683), .C2(n5025), .ZN(register_file_inst1_n2143) );
  INVD1BWP12T U4343 ( .I(register_file_inst1_lr_6_), .ZN(n5026) );
  OAI222D1BWP12T U4344 ( .A1(n5034), .A2(n5223), .B1(n5160), .B2(n6367), .C1(
        n5222), .C2(n5026), .ZN(register_file_inst1_n2207) );
  INVD1BWP12T U4345 ( .I(register_file_inst1_r6_6_), .ZN(n5718) );
  OAI222D1BWP12T U4346 ( .A1(n5034), .A2(n5229), .B1(n5228), .B2(n6367), .C1(
        n5095), .C2(n5718), .ZN(register_file_inst1_n2431) );
  INVD1BWP12T U4347 ( .I(register_file_inst1_r4_6_), .ZN(n5027) );
  OAI222D1BWP12T U4348 ( .A1(n5034), .A2(n5226), .B1(n5205), .B2(n6367), .C1(
        n5225), .C2(n5027), .ZN(register_file_inst1_n2495) );
  INVD1BWP12T U4349 ( .I(register_file_inst1_r0_6_), .ZN(n5719) );
  OAI222D1BWP12T U4350 ( .A1(n5034), .A2(n5231), .B1(n5230), .B2(n6367), .C1(
        n5096), .C2(n5719), .ZN(register_file_inst1_n2623) );
  CKND0BWP12T U4351 ( .I(register_file_inst1_r7_6_), .ZN(n5028) );
  OAI222D1BWP12T U4352 ( .A1(n5034), .A2(n5227), .B1(n5158), .B2(n6367), .C1(
        n5094), .C2(n5028), .ZN(register_file_inst1_n2399) );
  CKND0BWP12T U4353 ( .I(register_file_inst1_r5_6_), .ZN(n5029) );
  OAI222D1BWP12T U4354 ( .A1(n5034), .A2(n5143), .B1(n5249), .B2(n6367), .C1(
        n5247), .C2(n5029), .ZN(register_file_inst1_n2463) );
  INVD1BWP12T U4355 ( .I(register_file_inst1_r1_6_), .ZN(n5717) );
  OAI222D1BWP12T U4356 ( .A1(n5034), .A2(n5074), .B1(n5240), .B2(n6367), .C1(
        n5239), .C2(n5717), .ZN(register_file_inst1_n2591) );
  OAI222D1BWP12T U4357 ( .A1(n5034), .A2(n5140), .B1(n5243), .B2(n6367), .C1(
        n5242), .C2(n5030), .ZN(register_file_inst1_n2239) );
  CKND0BWP12T U4358 ( .I(register_file_inst1_r8_6_), .ZN(n5031) );
  OAI222D1BWP12T U4359 ( .A1(n5034), .A2(n5145), .B1(n5246), .B2(n6367), .C1(
        n5244), .C2(n5031), .ZN(register_file_inst1_n2367) );
  CKND0BWP12T U4360 ( .I(register_file_inst1_r9_6_), .ZN(n5032) );
  OAI222D1BWP12T U4361 ( .A1(n5034), .A2(n5238), .B1(n5237), .B2(n6367), .C1(
        n5235), .C2(n5032), .ZN(register_file_inst1_n2335) );
  INVD1BWP12T U4362 ( .I(register_file_inst1_r10_6_), .ZN(n5033) );
  OAI222D1BWP12T U4363 ( .A1(n5034), .A2(n5253), .B1(n5252), .B2(n6367), .C1(
        n5250), .C2(n5033), .ZN(register_file_inst1_n2303) );
  INVD1BWP12T U4364 ( .I(register_file_inst1_r2_6_), .ZN(n5720) );
  OAI222D1BWP12T U4365 ( .A1(n5034), .A2(n5257), .B1(n5256), .B2(n6367), .C1(
        n5254), .C2(n5720), .ZN(register_file_inst1_n2559) );
  ND2D1BWP12T U4366 ( .A1(ALU_MISC_OUT_result[9]), .A2(n5978), .ZN(n5035) );
  OAI211D1BWP12T U4367 ( .A1(n5233), .A2(n6308), .B(n5035), .C(n6086), .ZN(
        register_file_inst1_spin[9]) );
  ND2D1BWP12T U4368 ( .A1(ALU_MISC_OUT_result[10]), .A2(n5978), .ZN(n5036) );
  OAI211D1BWP12T U4369 ( .A1(n5233), .A2(n6355), .B(n5036), .C(n6089), .ZN(
        register_file_inst1_spin[10]) );
  AOI22D1BWP12T U4370 ( .A1(register_file_inst1_lr_12_), .A2(n5049), .B1(
        register_file_inst1_r9_12_), .B2(n5048), .ZN(n5039) );
  AOI22D0BWP12T U4371 ( .A1(RF_next_sp[12]), .A2(n5051), .B1(
        register_file_inst1_r7_12_), .B2(n5050), .ZN(n5038) );
  AOI22D0BWP12T U4372 ( .A1(register_file_inst1_r6_12_), .A2(n5053), .B1(
        register_file_inst1_r2_12_), .B2(n5052), .ZN(n5037) );
  AN4XD1BWP12T U4373 ( .A1(n6291), .A2(n5039), .A3(n5038), .A4(n5037), .Z(
        n5045) );
  AOI22D1BWP12T U4374 ( .A1(register_file_inst1_r3_12_), .A2(n5058), .B1(
        register_file_inst1_r12_12_), .B2(n5057), .ZN(n5043) );
  AOI22D1BWP12T U4375 ( .A1(register_file_inst1_r4_12_), .A2(n5060), .B1(
        register_file_inst1_r8_12_), .B2(n5059), .ZN(n5042) );
  AOI22D0BWP12T U4376 ( .A1(register_file_inst1_r0_12_), .A2(n5062), .B1(
        register_file_inst1_r1_12_), .B2(n5061), .ZN(n5041) );
  AOI22D1BWP12T U4377 ( .A1(register_file_inst1_r10_12_), .A2(n5064), .B1(
        register_file_inst1_r11_12_), .B2(n5063), .ZN(n5040) );
  AN4XD1BWP12T U4378 ( .A1(n5043), .A2(n5042), .A3(n5041), .A4(n5040), .Z(
        n5044) );
  ND2D1BWP12T U4379 ( .A1(n5045), .A2(n5044), .ZN(n6292) );
  AOI21D0BWP12T U4380 ( .A1(n6008), .A2(ALU_MISC_OUT_result[6]), .B(n5046), 
        .ZN(n5047) );
  OAI22D1BWP12T U4381 ( .A1(n5047), .A2(n5270), .B1(n5267), .B2(n6367), .ZN(
        n6368) );
  AOI22D1BWP12T U4382 ( .A1(n5049), .A2(register_file_inst1_lr_11_), .B1(
        register_file_inst1_r9_11_), .B2(n5048), .ZN(n5056) );
  AOI22D0BWP12T U4383 ( .A1(n5051), .A2(RF_next_sp[11]), .B1(
        register_file_inst1_r7_11_), .B2(n5050), .ZN(n5055) );
  AOI22D0BWP12T U4384 ( .A1(n5053), .A2(register_file_inst1_r6_11_), .B1(
        register_file_inst1_r2_11_), .B2(n5052), .ZN(n5054) );
  AN4XD1BWP12T U4385 ( .A1(n6288), .A2(n5056), .A3(n5055), .A4(n5054), .Z(
        n5070) );
  AOI22D1BWP12T U4386 ( .A1(n5058), .A2(register_file_inst1_r3_11_), .B1(
        register_file_inst1_r12_11_), .B2(n5057), .ZN(n5068) );
  AOI22D1BWP12T U4387 ( .A1(n5060), .A2(register_file_inst1_r4_11_), .B1(
        register_file_inst1_r8_11_), .B2(n5059), .ZN(n5067) );
  AOI22D0BWP12T U4388 ( .A1(n5062), .A2(register_file_inst1_r0_11_), .B1(
        register_file_inst1_r1_11_), .B2(n5061), .ZN(n5066) );
  AOI22D1BWP12T U4389 ( .A1(n5064), .A2(register_file_inst1_r10_11_), .B1(
        register_file_inst1_r11_11_), .B2(n5063), .ZN(n5065) );
  AN4XD1BWP12T U4390 ( .A1(n5068), .A2(n5067), .A3(n5066), .A4(n5065), .Z(
        n5069) );
  ND2D1BWP12T U4391 ( .A1(n5070), .A2(n5069), .ZN(n6289) );
  OAI21D1BWP12T U4392 ( .A1(n5082), .A2(n5234), .B(n6098), .ZN(
        register_file_inst1_spin[12]) );
  CKND0BWP12T U4393 ( .I(register_file_inst1_r8_12_), .ZN(n5071) );
  OAI222D1BWP12T U4394 ( .A1(n5082), .A2(n5145), .B1(n5246), .B2(n6349), .C1(
        n5244), .C2(n5071), .ZN(register_file_inst1_n2373) );
  INVD1BWP12T U4395 ( .I(register_file_inst1_r11_12_), .ZN(n5072) );
  OAI222D1BWP12T U4396 ( .A1(n5082), .A2(n5220), .B1(n5219), .B2(n6349), .C1(
        n5217), .C2(n5072), .ZN(register_file_inst1_n2277) );
  CKND0BWP12T U4397 ( .I(register_file_inst1_r9_12_), .ZN(n5073) );
  OAI222D1BWP12T U4398 ( .A1(n5082), .A2(n5238), .B1(n5237), .B2(n6349), .C1(
        n5235), .C2(n5073), .ZN(register_file_inst1_n2341) );
  INVD1BWP12T U4399 ( .I(register_file_inst1_r1_12_), .ZN(n5609) );
  OAI222D1BWP12T U4400 ( .A1(n5082), .A2(n5074), .B1(n5240), .B2(n6349), .C1(
        n5239), .C2(n5609), .ZN(register_file_inst1_n2597) );
  INVD1BWP12T U4401 ( .I(register_file_inst1_r5_12_), .ZN(n5075) );
  OAI222D1BWP12T U4402 ( .A1(n5082), .A2(n5143), .B1(n5249), .B2(n6349), .C1(
        n5247), .C2(n5075), .ZN(register_file_inst1_n2469) );
  INVD1BWP12T U4403 ( .I(register_file_inst1_r12_12_), .ZN(n5076) );
  OAI222D1BWP12T U4404 ( .A1(n5082), .A2(n5140), .B1(n5243), .B2(n6349), .C1(
        n5242), .C2(n5076), .ZN(register_file_inst1_n2245) );
  CKND0BWP12T U4405 ( .I(register_file_inst1_r7_12_), .ZN(n5077) );
  OAI222D1BWP12T U4406 ( .A1(n5082), .A2(n5227), .B1(n5158), .B2(n6349), .C1(
        n5094), .C2(n5077), .ZN(register_file_inst1_n2405) );
  INVD1BWP12T U4407 ( .I(register_file_inst1_r0_12_), .ZN(n5611) );
  OAI222D1BWP12T U4408 ( .A1(n5082), .A2(n5231), .B1(n5230), .B2(n6349), .C1(
        n5096), .C2(n5611), .ZN(register_file_inst1_n2629) );
  INVD1BWP12T U4409 ( .I(register_file_inst1_r6_12_), .ZN(n5610) );
  OAI222D1BWP12T U4410 ( .A1(n5082), .A2(n5229), .B1(n5228), .B2(n6349), .C1(
        n5095), .C2(n5610), .ZN(register_file_inst1_n2437) );
  INVD1BWP12T U4411 ( .I(register_file_inst1_r4_12_), .ZN(n5078) );
  OAI222D1BWP12T U4412 ( .A1(n5082), .A2(n5226), .B1(n5205), .B2(n6349), .C1(
        n5225), .C2(n5078), .ZN(register_file_inst1_n2501) );
  CKND0BWP12T U4413 ( .I(register_file_inst1_tmp1_12_), .ZN(n5079) );
  OAI222D1BWP12T U4414 ( .A1(n5082), .A2(n6144), .B1(n5212), .B2(n6349), .C1(
        n4683), .C2(n5079), .ZN(register_file_inst1_n2149) );
  INVD1BWP12T U4415 ( .I(register_file_inst1_lr_12_), .ZN(n5080) );
  OAI222D1BWP12T U4416 ( .A1(n5082), .A2(n5223), .B1(n5160), .B2(n6349), .C1(
        n5222), .C2(n5080), .ZN(register_file_inst1_n2213) );
  INVD1BWP12T U4417 ( .I(register_file_inst1_r2_12_), .ZN(n5612) );
  OAI222D1BWP12T U4418 ( .A1(n5082), .A2(n5257), .B1(n5256), .B2(n6349), .C1(
        n5254), .C2(n5612), .ZN(register_file_inst1_n2565) );
  INVD1BWP12T U4419 ( .I(register_file_inst1_r10_12_), .ZN(n5081) );
  OAI222D1BWP12T U4420 ( .A1(n5082), .A2(n5253), .B1(n5252), .B2(n6349), .C1(
        n5250), .C2(n5081), .ZN(register_file_inst1_n2309) );
  CKND0BWP12T U4421 ( .I(register_file_inst1_tmp1_13_), .ZN(n5083) );
  OAI222D1BWP12T U4422 ( .A1(n5084), .A2(n6144), .B1(n5212), .B2(n6346), .C1(
        n4683), .C2(n5083), .ZN(register_file_inst1_n2150) );
  CKND0BWP12T U4423 ( .I(register_file_inst1_tmp1_14_), .ZN(n5085) );
  OAI222D1BWP12T U4424 ( .A1(n5086), .A2(n6144), .B1(n5212), .B2(n6343), .C1(
        n4683), .C2(n5085), .ZN(register_file_inst1_n2151) );
  CKND0BWP12T U4425 ( .I(register_file_inst1_tmp1_15_), .ZN(n5087) );
  OAI222D1BWP12T U4426 ( .A1(n5088), .A2(n6144), .B1(n5212), .B2(n6340), .C1(
        n4683), .C2(n5087), .ZN(register_file_inst1_n2152) );
  CKND0BWP12T U4427 ( .I(register_file_inst1_tmp1_16_), .ZN(n5089) );
  OAI222D1BWP12T U4428 ( .A1(n5089), .A2(n4683), .B1(n5212), .B2(n5103), .C1(
        n5102), .C2(n6144), .ZN(register_file_inst1_n2153) );
  INVD1BWP12T U4429 ( .I(register_file_inst1_r5_16_), .ZN(n5090) );
  OAI222D1BWP12T U4430 ( .A1(n5090), .A2(n5247), .B1(n5249), .B2(n5103), .C1(
        n5102), .C2(n5143), .ZN(register_file_inst1_n2473) );
  INVD1BWP12T U4431 ( .I(register_file_inst1_r8_16_), .ZN(n5091) );
  OAI222D1BWP12T U4432 ( .A1(n5091), .A2(n5244), .B1(n5246), .B2(n5103), .C1(
        n5102), .C2(n5145), .ZN(register_file_inst1_n2377) );
  INVD1BWP12T U4433 ( .I(register_file_inst1_r9_16_), .ZN(n5092) );
  OAI222D1BWP12T U4434 ( .A1(n5092), .A2(n5235), .B1(n5237), .B2(n5103), .C1(
        n5102), .C2(n5238), .ZN(register_file_inst1_n2345) );
  INVD1BWP12T U4435 ( .I(register_file_inst1_r12_16_), .ZN(n5093) );
  OAI222D1BWP12T U4436 ( .A1(n5093), .A2(n5242), .B1(n5243), .B2(n5103), .C1(
        n5102), .C2(n5140), .ZN(register_file_inst1_n2249) );
  INVD1BWP12T U4437 ( .I(register_file_inst1_r1_16_), .ZN(n5539) );
  OAI222D1BWP12T U4438 ( .A1(n5539), .A2(n5239), .B1(n5240), .B2(n5103), .C1(
        n5102), .C2(n5074), .ZN(register_file_inst1_n2601) );
  INVD1BWP12T U4439 ( .I(register_file_inst1_r7_16_), .ZN(n5537) );
  OAI222D1BWP12T U4440 ( .A1(n5537), .A2(n5094), .B1(n5158), .B2(n5103), .C1(
        n5102), .C2(n5227), .ZN(register_file_inst1_n2409) );
  INVD1BWP12T U4441 ( .I(register_file_inst1_r6_16_), .ZN(n5524) );
  OAI222D1BWP12T U4442 ( .A1(n5524), .A2(n5095), .B1(n5228), .B2(n5103), .C1(
        n5102), .C2(n5229), .ZN(register_file_inst1_n2441) );
  INVD1BWP12T U4443 ( .I(register_file_inst1_r0_16_), .ZN(n5525) );
  OAI222D1BWP12T U4444 ( .A1(n5525), .A2(n5096), .B1(n5230), .B2(n5103), .C1(
        n5102), .C2(n5231), .ZN(register_file_inst1_n2633) );
  INVD1BWP12T U4445 ( .I(register_file_inst1_lr_16_), .ZN(n5538) );
  OAI222D1BWP12T U4446 ( .A1(n5538), .A2(n5222), .B1(n5160), .B2(n5103), .C1(
        n5102), .C2(n5223), .ZN(register_file_inst1_n2217) );
  INVD1BWP12T U4447 ( .I(register_file_inst1_r4_16_), .ZN(n5097) );
  OAI222D1BWP12T U4448 ( .A1(n5097), .A2(n5225), .B1(n5205), .B2(n5103), .C1(
        n5102), .C2(n5226), .ZN(register_file_inst1_n2505) );
  INVD1BWP12T U4449 ( .I(RF_next_sp[16]), .ZN(n5536) );
  OAI222D1BWP12T U4450 ( .A1(n5536), .A2(n5232), .B1(n5233), .B2(n5103), .C1(
        n5102), .C2(n5234), .ZN(register_file_inst1_spin[16]) );
  CKND0BWP12T U4451 ( .I(register_file_inst1_tmp1_17_), .ZN(n5100) );
  OAI222D1BWP12T U4452 ( .A1(n5100), .A2(n4683), .B1(n5212), .B2(n5099), .C1(
        n5098), .C2(n6144), .ZN(register_file_inst1_n2154) );
  INVD1BWP12T U4453 ( .I(register_file_inst1_r10_16_), .ZN(n5101) );
  OAI222D1BWP12T U4454 ( .A1(n5101), .A2(n5250), .B1(n5252), .B2(n5103), .C1(
        n5102), .C2(n5253), .ZN(register_file_inst1_n2313) );
  INVD1BWP12T U4455 ( .I(register_file_inst1_r2_16_), .ZN(n5526) );
  OAI222D1BWP12T U4456 ( .A1(n5526), .A2(n5254), .B1(n5256), .B2(n5103), .C1(
        n5102), .C2(n5257), .ZN(register_file_inst1_n2569) );
  INVD1BWP12T U4457 ( .I(register_file_inst1_r7_20_), .ZN(n5897) );
  OAI222D1BWP12T U4458 ( .A1(n5897), .A2(n5094), .B1(n5158), .B2(n5112), .C1(
        n5111), .C2(n5227), .ZN(register_file_inst1_n2413) );
  INVD1BWP12T U4459 ( .I(register_file_inst1_r6_20_), .ZN(n5884) );
  OAI222D1BWP12T U4460 ( .A1(n5884), .A2(n5095), .B1(n5228), .B2(n5112), .C1(
        n5111), .C2(n5229), .ZN(register_file_inst1_n2445) );
  INVD1BWP12T U4461 ( .I(register_file_inst1_r0_20_), .ZN(n5885) );
  OAI222D1BWP12T U4462 ( .A1(n5885), .A2(n5096), .B1(n5230), .B2(n5112), .C1(
        n5111), .C2(n5231), .ZN(register_file_inst1_n2637) );
  INVD1BWP12T U4463 ( .I(register_file_inst1_lr_20_), .ZN(n5898) );
  OAI222D1BWP12T U4464 ( .A1(n5898), .A2(n5222), .B1(n5160), .B2(n5112), .C1(
        n5111), .C2(n5223), .ZN(register_file_inst1_n2221) );
  INVD1BWP12T U4465 ( .I(register_file_inst1_r4_20_), .ZN(n5104) );
  OAI222D1BWP12T U4466 ( .A1(n5104), .A2(n5225), .B1(n5205), .B2(n5112), .C1(
        n5111), .C2(n5226), .ZN(register_file_inst1_n2509) );
  INVD1BWP12T U4467 ( .I(register_file_inst1_r12_20_), .ZN(n5105) );
  OAI222D1BWP12T U4468 ( .A1(n5105), .A2(n5242), .B1(n5243), .B2(n5112), .C1(
        n5111), .C2(n5140), .ZN(register_file_inst1_n2253) );
  CKND0BWP12T U4469 ( .I(register_file_inst1_r9_20_), .ZN(n5106) );
  OAI222D1BWP12T U4470 ( .A1(n5106), .A2(n5235), .B1(n5237), .B2(n5112), .C1(
        n5111), .C2(n5238), .ZN(register_file_inst1_n2349) );
  INVD1BWP12T U4471 ( .I(register_file_inst1_r8_20_), .ZN(n5107) );
  OAI222D1BWP12T U4472 ( .A1(n5107), .A2(n5244), .B1(n5246), .B2(n5112), .C1(
        n5111), .C2(n5145), .ZN(register_file_inst1_n2381) );
  INVD1BWP12T U4473 ( .I(register_file_inst1_r5_20_), .ZN(n5108) );
  OAI222D1BWP12T U4474 ( .A1(n5108), .A2(n5247), .B1(n5249), .B2(n5112), .C1(
        n5111), .C2(n5143), .ZN(register_file_inst1_n2477) );
  INVD1BWP12T U4475 ( .I(register_file_inst1_r1_20_), .ZN(n5899) );
  OAI222D1BWP12T U4476 ( .A1(n5899), .A2(n5239), .B1(n5240), .B2(n5112), .C1(
        n5111), .C2(n5074), .ZN(register_file_inst1_n2605) );
  INVD1BWP12T U4477 ( .I(RF_next_sp[20]), .ZN(n5896) );
  OAI222D1BWP12T U4478 ( .A1(n5896), .A2(n5232), .B1(n5233), .B2(n5112), .C1(
        n5111), .C2(n5234), .ZN(register_file_inst1_spin[20]) );
  INVD1BWP12T U4479 ( .I(register_file_inst1_r11_20_), .ZN(n5109) );
  OAI222D1BWP12T U4480 ( .A1(n5109), .A2(n5217), .B1(n5219), .B2(n5112), .C1(
        n5111), .C2(n5220), .ZN(register_file_inst1_n2285) );
  CKND0BWP12T U4481 ( .I(register_file_inst1_tmp1_20_), .ZN(n5110) );
  OAI222D1BWP12T U4482 ( .A1(n5110), .A2(n4683), .B1(n5212), .B2(n5112), .C1(
        n5111), .C2(n6144), .ZN(register_file_inst1_n2157) );
  INVD1BWP12T U4483 ( .I(register_file_inst1_r2_20_), .ZN(n5886) );
  OAI222D1BWP12T U4484 ( .A1(n5886), .A2(n5254), .B1(n5256), .B2(n5112), .C1(
        n5111), .C2(n5257), .ZN(register_file_inst1_n2573) );
  INVD1BWP12T U4485 ( .I(register_file_inst1_r10_20_), .ZN(n5113) );
  OAI222D1BWP12T U4486 ( .A1(n5113), .A2(n5250), .B1(n5252), .B2(n5112), .C1(
        n5111), .C2(n5253), .ZN(register_file_inst1_n2317) );
  CKND0BWP12T U4487 ( .I(register_file_inst1_tmp1_19_), .ZN(n5116) );
  OAI222D1BWP12T U4488 ( .A1(n5116), .A2(n4683), .B1(n5212), .B2(n5115), .C1(
        n5114), .C2(n6144), .ZN(register_file_inst1_n2156) );
  AOI21D0BWP12T U4489 ( .A1(n6008), .A2(ALU_MISC_OUT_result[10]), .B(n5117), 
        .ZN(n5118) );
  OAI22D1BWP12T U4490 ( .A1(n5118), .A2(n5270), .B1(n5267), .B2(n6355), .ZN(
        n6356) );
  CKND0BWP12T U4491 ( .I(register_file_inst1_tmp1_21_), .ZN(n5121) );
  OAI222D1BWP12T U4492 ( .A1(n5121), .A2(n4683), .B1(n5212), .B2(n5120), .C1(
        n5119), .C2(n6144), .ZN(register_file_inst1_n2158) );
  AOI21D0BWP12T U4493 ( .A1(n6008), .A2(ALU_MISC_OUT_result[12]), .B(n5122), 
        .ZN(n5123) );
  OAI22D1BWP12T U4494 ( .A1(n5123), .A2(n5270), .B1(n5267), .B2(n6349), .ZN(
        n6350) );
  CKND0BWP12T U4495 ( .I(register_file_inst1_tmp1_22_), .ZN(n5124) );
  INVD1BWP12T U4496 ( .I(register_file_inst1_r6_22_), .ZN(n5448) );
  INVD1BWP12T U4497 ( .I(register_file_inst1_r0_22_), .ZN(n5449) );
  CKND0BWP12T U4498 ( .I(register_file_inst1_r8_22_), .ZN(n5125) );
  CKND0BWP12T U4499 ( .I(register_file_inst1_r5_22_), .ZN(n5126) );
  CKND0BWP12T U4500 ( .I(register_file_inst1_r9_22_), .ZN(n5127) );
  INVD1BWP12T U4501 ( .I(register_file_inst1_r7_22_), .ZN(n5461) );
  INVD1BWP12T U4502 ( .I(register_file_inst1_r1_22_), .ZN(n5463) );
  INVD1BWP12T U4503 ( .I(register_file_inst1_lr_22_), .ZN(n5462) );
  CKND0BWP12T U4504 ( .I(register_file_inst1_r12_22_), .ZN(n5128) );
  CKND0BWP12T U4505 ( .I(register_file_inst1_r4_22_), .ZN(n5129) );
  INVD1BWP12T U4506 ( .I(RF_next_sp[22]), .ZN(n5460) );
  CKND0BWP12T U4507 ( .I(register_file_inst1_r11_22_), .ZN(n5130) );
  INVD1BWP12T U4508 ( .I(register_file_inst1_r2_22_), .ZN(n5450) );
  CKND0BWP12T U4509 ( .I(register_file_inst1_r10_22_), .ZN(n5133) );
  CKND0BWP12T U4510 ( .I(register_file_inst1_tmp1_23_), .ZN(n5134) );
  OAI222D1BWP12T U4511 ( .A1(n5136), .A2(n6144), .B1(n5212), .B2(n5135), .C1(
        n4683), .C2(n5134), .ZN(register_file_inst1_n2160) );
  AOI21D0BWP12T U4512 ( .A1(n6008), .A2(ALU_MISC_OUT_result[14]), .B(n5137), 
        .ZN(n5138) );
  OAI22D1BWP12T U4513 ( .A1(n5138), .A2(n5270), .B1(n5267), .B2(n6343), .ZN(
        n6344) );
  OAI222D1BWP12T U4514 ( .A1(n5140), .A2(n5260), .B1(n5243), .B2(n5259), .C1(
        n5242), .C2(n5139), .ZN(register_file_inst1_n2257) );
  CKND0BWP12T U4515 ( .I(register_file_inst1_r9_24_), .ZN(n5141) );
  OAI222D1BWP12T U4516 ( .A1(n5238), .A2(n5260), .B1(n5237), .B2(n5259), .C1(
        n5235), .C2(n5141), .ZN(register_file_inst1_n2353) );
  CKND0BWP12T U4517 ( .I(register_file_inst1_r5_24_), .ZN(n5142) );
  OAI222D1BWP12T U4518 ( .A1(n5143), .A2(n5260), .B1(n5249), .B2(n5259), .C1(
        n5247), .C2(n5142), .ZN(register_file_inst1_n2481) );
  OAI222D1BWP12T U4519 ( .A1(n5145), .A2(n5260), .B1(n5246), .B2(n5259), .C1(
        n5244), .C2(n5144), .ZN(register_file_inst1_n2385) );
  CKND0BWP12T U4520 ( .I(register_file_inst1_tmp1_24_), .ZN(n5146) );
  OAI222D1BWP12T U4521 ( .A1(n6144), .A2(n5260), .B1(n5212), .B2(n5259), .C1(
        n4683), .C2(n5146), .ZN(register_file_inst1_n2161) );
  CKND0BWP12T U4522 ( .I(register_file_inst1_r4_24_), .ZN(n5147) );
  OAI222D1BWP12T U4523 ( .A1(n5226), .A2(n5260), .B1(n5205), .B2(n5259), .C1(
        n5225), .C2(n5147), .ZN(register_file_inst1_n2513) );
  INVD1BWP12T U4524 ( .I(register_file_inst1_r6_25_), .ZN(n5911) );
  OAI222D1BWP12T U4525 ( .A1(n5911), .A2(n5095), .B1(n5228), .B2(n5261), .C1(
        n5262), .C2(n5229), .ZN(register_file_inst1_n2450) );
  INVD1BWP12T U4526 ( .I(register_file_inst1_r0_25_), .ZN(n5913) );
  OAI222D1BWP12T U4527 ( .A1(n5913), .A2(n5096), .B1(n5230), .B2(n5261), .C1(
        n5262), .C2(n5231), .ZN(register_file_inst1_n2642) );
  CKND0BWP12T U4528 ( .I(register_file_inst1_r4_25_), .ZN(n5148) );
  OAI222D1BWP12T U4529 ( .A1(n5148), .A2(n5225), .B1(n5205), .B2(n5261), .C1(
        n5262), .C2(n5226), .ZN(register_file_inst1_n2514) );
  CKND0BWP12T U4530 ( .I(register_file_inst1_r8_25_), .ZN(n5149) );
  OAI222D1BWP12T U4531 ( .A1(n5149), .A2(n5244), .B1(n5246), .B2(n5261), .C1(
        n5262), .C2(n5145), .ZN(register_file_inst1_n2386) );
  INVD1BWP12T U4532 ( .I(register_file_inst1_r1_25_), .ZN(n5927) );
  OAI222D1BWP12T U4533 ( .A1(n5927), .A2(n5239), .B1(n5240), .B2(n5261), .C1(
        n5262), .C2(n5074), .ZN(register_file_inst1_n2610) );
  CKND0BWP12T U4534 ( .I(register_file_inst1_r9_25_), .ZN(n5150) );
  OAI222D1BWP12T U4535 ( .A1(n5150), .A2(n5235), .B1(n5237), .B2(n5261), .C1(
        n5262), .C2(n5238), .ZN(register_file_inst1_n2354) );
  CKND0BWP12T U4536 ( .I(register_file_inst1_r12_25_), .ZN(n5151) );
  OAI222D1BWP12T U4537 ( .A1(n5151), .A2(n5242), .B1(n5243), .B2(n5261), .C1(
        n5262), .C2(n5140), .ZN(register_file_inst1_n2258) );
  CKND0BWP12T U4538 ( .I(register_file_inst1_r5_25_), .ZN(n5152) );
  OAI222D1BWP12T U4539 ( .A1(n5152), .A2(n5247), .B1(n5249), .B2(n5261), .C1(
        n5262), .C2(n5143), .ZN(register_file_inst1_n2482) );
  INVD1BWP12T U4540 ( .I(RF_next_sp[25]), .ZN(n5924) );
  OAI222D1BWP12T U4541 ( .A1(n5924), .A2(n5232), .B1(n5233), .B2(n5261), .C1(
        n5262), .C2(n5234), .ZN(register_file_inst1_spin[25]) );
  CKND0BWP12T U4542 ( .I(register_file_inst1_r11_25_), .ZN(n5153) );
  OAI222D1BWP12T U4543 ( .A1(n5153), .A2(n5217), .B1(n5219), .B2(n5261), .C1(
        n5262), .C2(n5220), .ZN(register_file_inst1_n2290) );
  CKND0BWP12T U4544 ( .I(register_file_inst1_tmp1_25_), .ZN(n5154) );
  OAI222D1BWP12T U4545 ( .A1(n5154), .A2(n4683), .B1(n5212), .B2(n5261), .C1(
        n5262), .C2(n6144), .ZN(register_file_inst1_n2162) );
  CKND0BWP12T U4546 ( .I(register_file_inst1_r10_25_), .ZN(n5155) );
  OAI222D1BWP12T U4547 ( .A1(n5155), .A2(n5250), .B1(n5252), .B2(n5261), .C1(
        n5262), .C2(n5253), .ZN(register_file_inst1_n2322) );
  INVD1BWP12T U4548 ( .I(register_file_inst1_r2_25_), .ZN(n5914) );
  OAI222D1BWP12T U4549 ( .A1(n5914), .A2(n5254), .B1(n5256), .B2(n5261), .C1(
        n5262), .C2(n5257), .ZN(register_file_inst1_n2578) );
  CKND0BWP12T U4550 ( .I(register_file_inst1_r3_25_), .ZN(n5156) );
  OAI222D1BWP12T U4551 ( .A1(n5156), .A2(n4758), .B1(n5203), .B2(n5261), .C1(
        n5262), .C2(n5200), .ZN(register_file_inst1_n2546) );
  INVD1BWP12T U4552 ( .I(register_file_inst1_r7_26_), .ZN(n5939) );
  OAI222D1BWP12T U4553 ( .A1(n5939), .A2(n5094), .B1(n5158), .B2(n5263), .C1(
        n5167), .C2(n5227), .ZN(register_file_inst1_n2419) );
  INVD1BWP12T U4554 ( .I(register_file_inst1_r6_26_), .ZN(n5957) );
  OAI222D1BWP12T U4555 ( .A1(n5957), .A2(n5095), .B1(n5228), .B2(n5263), .C1(
        n5167), .C2(n5229), .ZN(register_file_inst1_n2451) );
  INVD1BWP12T U4556 ( .I(register_file_inst1_r0_26_), .ZN(n5958) );
  OAI222D1BWP12T U4557 ( .A1(n5958), .A2(n5096), .B1(n5230), .B2(n5263), .C1(
        n5167), .C2(n5231), .ZN(register_file_inst1_n2643) );
  CKND0BWP12T U4558 ( .I(register_file_inst1_r4_26_), .ZN(n5159) );
  OAI222D1BWP12T U4559 ( .A1(n5159), .A2(n5225), .B1(n5205), .B2(n5263), .C1(
        n5167), .C2(n5226), .ZN(register_file_inst1_n2515) );
  INVD1BWP12T U4560 ( .I(register_file_inst1_lr_26_), .ZN(n5941) );
  OAI222D1BWP12T U4561 ( .A1(n5941), .A2(n5222), .B1(n5160), .B2(n5263), .C1(
        n5167), .C2(n5223), .ZN(register_file_inst1_n2227) );
  CKND0BWP12T U4562 ( .I(register_file_inst1_r8_26_), .ZN(n5161) );
  OAI222D1BWP12T U4563 ( .A1(n5161), .A2(n5244), .B1(n5246), .B2(n5263), .C1(
        n5167), .C2(n5145), .ZN(register_file_inst1_n2387) );
  CKND0BWP12T U4564 ( .I(register_file_inst1_r9_26_), .ZN(n5162) );
  OAI222D1BWP12T U4565 ( .A1(n5162), .A2(n5235), .B1(n5237), .B2(n5263), .C1(
        n5167), .C2(n5238), .ZN(register_file_inst1_n2355) );
  CKND0BWP12T U4566 ( .I(register_file_inst1_r12_26_), .ZN(n5163) );
  OAI222D1BWP12T U4567 ( .A1(n5163), .A2(n5242), .B1(n5243), .B2(n5263), .C1(
        n5167), .C2(n5140), .ZN(register_file_inst1_n2259) );
  CKND0BWP12T U4568 ( .I(register_file_inst1_r5_26_), .ZN(n5164) );
  OAI222D1BWP12T U4569 ( .A1(n5164), .A2(n5247), .B1(n5249), .B2(n5263), .C1(
        n5167), .C2(n5143), .ZN(register_file_inst1_n2483) );
  INVD1BWP12T U4570 ( .I(register_file_inst1_r1_26_), .ZN(n5956) );
  OAI222D1BWP12T U4571 ( .A1(n5956), .A2(n5239), .B1(n5240), .B2(n5263), .C1(
        n5167), .C2(n5074), .ZN(register_file_inst1_n2611) );
  INVD1BWP12T U4572 ( .I(RF_next_sp[26]), .ZN(n5937) );
  OAI222D1BWP12T U4573 ( .A1(n5937), .A2(n5232), .B1(n5233), .B2(n5263), .C1(
        n5167), .C2(n5234), .ZN(register_file_inst1_spin[26]) );
  CKND0BWP12T U4574 ( .I(register_file_inst1_r11_26_), .ZN(n5165) );
  OAI222D1BWP12T U4575 ( .A1(n5165), .A2(n5217), .B1(n5219), .B2(n5263), .C1(
        n5167), .C2(n5220), .ZN(register_file_inst1_n2291) );
  CKND0BWP12T U4576 ( .I(register_file_inst1_tmp1_26_), .ZN(n5166) );
  OAI222D1BWP12T U4577 ( .A1(n5166), .A2(n4683), .B1(n5212), .B2(n5263), .C1(
        n5167), .C2(n6144), .ZN(register_file_inst1_n2163) );
  INVD1BWP12T U4578 ( .I(register_file_inst1_r2_26_), .ZN(n5960) );
  OAI222D1BWP12T U4579 ( .A1(n5960), .A2(n5254), .B1(n5256), .B2(n5263), .C1(
        n5167), .C2(n5257), .ZN(register_file_inst1_n2579) );
  CKND0BWP12T U4580 ( .I(register_file_inst1_r10_26_), .ZN(n5168) );
  OAI222D1BWP12T U4581 ( .A1(n5168), .A2(n5250), .B1(n5252), .B2(n5263), .C1(
        n5167), .C2(n5253), .ZN(register_file_inst1_n2323) );
  CKND0BWP12T U4582 ( .I(register_file_inst1_r4_27_), .ZN(n5169) );
  OAI222D1BWP12T U4583 ( .A1(n5169), .A2(n5225), .B1(n5205), .B2(n5178), .C1(
        n5177), .C2(n5226), .ZN(register_file_inst1_n2516) );
  CKND0BWP12T U4584 ( .I(register_file_inst1_r8_27_), .ZN(n5170) );
  OAI222D1BWP12T U4585 ( .A1(n5170), .A2(n5244), .B1(n5246), .B2(n5178), .C1(
        n5177), .C2(n5145), .ZN(register_file_inst1_n2388) );
  CKND0BWP12T U4586 ( .I(register_file_inst1_r5_27_), .ZN(n5171) );
  OAI222D1BWP12T U4587 ( .A1(n5171), .A2(n5247), .B1(n5249), .B2(n5178), .C1(
        n5177), .C2(n5143), .ZN(register_file_inst1_n2484) );
  CKND0BWP12T U4588 ( .I(register_file_inst1_r9_27_), .ZN(n5172) );
  OAI222D1BWP12T U4589 ( .A1(n5172), .A2(n5235), .B1(n5237), .B2(n5178), .C1(
        n5177), .C2(n5238), .ZN(register_file_inst1_n2356) );
  INVD1BWP12T U4590 ( .I(register_file_inst1_r1_27_), .ZN(n5388) );
  OAI222D1BWP12T U4591 ( .A1(n5388), .A2(n5239), .B1(n5240), .B2(n5178), .C1(
        n5177), .C2(n5074), .ZN(register_file_inst1_n2612) );
  CKND0BWP12T U4592 ( .I(register_file_inst1_r12_27_), .ZN(n5173) );
  OAI222D1BWP12T U4593 ( .A1(n5173), .A2(n5242), .B1(n5243), .B2(n5178), .C1(
        n5177), .C2(n5140), .ZN(register_file_inst1_n2260) );
  INVD1BWP12T U4594 ( .I(RF_next_sp[27]), .ZN(n5385) );
  OAI222D1BWP12T U4595 ( .A1(n5385), .A2(n5232), .B1(n5233), .B2(n5178), .C1(
        n5177), .C2(n5234), .ZN(register_file_inst1_spin[27]) );
  CKND0BWP12T U4596 ( .I(register_file_inst1_r11_27_), .ZN(n5174) );
  OAI222D1BWP12T U4597 ( .A1(n5174), .A2(n5217), .B1(n5219), .B2(n5178), .C1(
        n5177), .C2(n5220), .ZN(register_file_inst1_n2292) );
  CKND0BWP12T U4598 ( .I(register_file_inst1_tmp1_27_), .ZN(n5175) );
  OAI222D1BWP12T U4599 ( .A1(n5175), .A2(n4683), .B1(n5212), .B2(n5178), .C1(
        n5177), .C2(n6144), .ZN(register_file_inst1_n2164) );
  CKND0BWP12T U4600 ( .I(register_file_inst1_r10_27_), .ZN(n5176) );
  OAI222D1BWP12T U4601 ( .A1(n5176), .A2(n5250), .B1(n5252), .B2(n5178), .C1(
        n5177), .C2(n5253), .ZN(register_file_inst1_n2324) );
  INVD1BWP12T U4602 ( .I(register_file_inst1_r2_27_), .ZN(n5375) );
  OAI222D1BWP12T U4603 ( .A1(n5375), .A2(n5254), .B1(n5256), .B2(n5178), .C1(
        n5177), .C2(n5257), .ZN(register_file_inst1_n2580) );
  CKND0BWP12T U4604 ( .I(register_file_inst1_r3_27_), .ZN(n5179) );
  OAI222D1BWP12T U4605 ( .A1(n5179), .A2(n4758), .B1(n5203), .B2(n5178), .C1(
        n5177), .C2(n5200), .ZN(register_file_inst1_n2548) );
  AOI21D1BWP12T U4606 ( .A1(n5181), .A2(memory_interface_inst1_fsm_state_0_), 
        .B(n5180), .ZN(n6113) );
  OAI21D1BWP12T U4607 ( .A1(n6234), .A2(n6400), .B(n5182), .ZN(n2264) );
  CKND0BWP12T U4608 ( .I(register_file_inst1_tmp1_28_), .ZN(n5183) );
  OAI222D1BWP12T U4609 ( .A1(n5183), .A2(n4683), .B1(n5212), .B2(n5190), .C1(
        n5189), .C2(n6144), .ZN(register_file_inst1_n2165) );
  INVD1BWP12T U4610 ( .I(register_file_inst1_r7_28_), .ZN(n5361) );
  OAI222D1BWP12T U4611 ( .A1(n5361), .A2(n5094), .B1(n5158), .B2(n5190), .C1(
        n5189), .C2(n5227), .ZN(register_file_inst1_n2421) );
  CKND0BWP12T U4612 ( .I(register_file_inst1_r9_28_), .ZN(n5184) );
  OAI222D1BWP12T U4613 ( .A1(n5184), .A2(n5235), .B1(n5237), .B2(n5190), .C1(
        n5189), .C2(n5238), .ZN(register_file_inst1_n2357) );
  CKND0BWP12T U4614 ( .I(register_file_inst1_r5_28_), .ZN(n5185) );
  OAI222D1BWP12T U4615 ( .A1(n5185), .A2(n5247), .B1(n5249), .B2(n5190), .C1(
        n5189), .C2(n5143), .ZN(register_file_inst1_n2485) );
  INVD1BWP12T U4616 ( .I(register_file_inst1_r6_28_), .ZN(n5348) );
  OAI222D1BWP12T U4617 ( .A1(n5348), .A2(n5095), .B1(n5228), .B2(n5190), .C1(
        n5189), .C2(n5229), .ZN(register_file_inst1_n2453) );
  INVD1BWP12T U4618 ( .I(register_file_inst1_r0_28_), .ZN(n5349) );
  OAI222D1BWP12T U4619 ( .A1(n5349), .A2(n5096), .B1(n5230), .B2(n5190), .C1(
        n5189), .C2(n5231), .ZN(register_file_inst1_n2645) );
  OAI222D1BWP12T U4620 ( .A1(n5186), .A2(n5244), .B1(n5246), .B2(n5190), .C1(
        n5189), .C2(n5145), .ZN(register_file_inst1_n2389) );
  INVD1BWP12T U4621 ( .I(register_file_inst1_r1_28_), .ZN(n5363) );
  OAI222D1BWP12T U4622 ( .A1(n5363), .A2(n5239), .B1(n5240), .B2(n5190), .C1(
        n5189), .C2(n5074), .ZN(register_file_inst1_n2613) );
  INVD1BWP12T U4623 ( .I(register_file_inst1_lr_28_), .ZN(n5362) );
  OAI222D1BWP12T U4624 ( .A1(n5362), .A2(n5222), .B1(n5160), .B2(n5190), .C1(
        n5189), .C2(n5223), .ZN(register_file_inst1_n2229) );
  OAI222D1BWP12T U4625 ( .A1(n5187), .A2(n5242), .B1(n5243), .B2(n5190), .C1(
        n5189), .C2(n5140), .ZN(register_file_inst1_n2261) );
  CKND0BWP12T U4626 ( .I(register_file_inst1_r4_28_), .ZN(n5188) );
  OAI222D1BWP12T U4627 ( .A1(n5188), .A2(n5225), .B1(n5205), .B2(n5190), .C1(
        n5189), .C2(n5226), .ZN(register_file_inst1_n2517) );
  INVD1BWP12T U4628 ( .I(RF_next_sp[28]), .ZN(n5360) );
  OAI222D1BWP12T U4629 ( .A1(n5360), .A2(n5232), .B1(n5233), .B2(n5190), .C1(
        n5189), .C2(n5234), .ZN(register_file_inst1_spin[28]) );
  INVD1BWP12T U4630 ( .I(register_file_inst1_r2_28_), .ZN(n5350) );
  OAI222D1BWP12T U4631 ( .A1(n5350), .A2(n5254), .B1(n5256), .B2(n5190), .C1(
        n5189), .C2(n5257), .ZN(register_file_inst1_n2581) );
  CKND0BWP12T U4632 ( .I(register_file_inst1_r10_28_), .ZN(n5191) );
  OAI222D1BWP12T U4633 ( .A1(n5191), .A2(n5250), .B1(n5252), .B2(n5190), .C1(
        n5189), .C2(n5253), .ZN(register_file_inst1_n2325) );
  INVD1BWP12T U4634 ( .I(register_file_inst1_r6_29_), .ZN(n5323) );
  OAI222D1BWP12T U4635 ( .A1(n5323), .A2(n5095), .B1(n5228), .B2(n5202), .C1(
        n5201), .C2(n5229), .ZN(register_file_inst1_n2454) );
  INVD1BWP12T U4636 ( .I(register_file_inst1_r0_29_), .ZN(n5324) );
  OAI222D1BWP12T U4637 ( .A1(n5324), .A2(n5096), .B1(n5230), .B2(n5202), .C1(
        n5201), .C2(n5231), .ZN(register_file_inst1_n2646) );
  INVD1BWP12T U4638 ( .I(register_file_inst1_r7_29_), .ZN(n5336) );
  OAI222D1BWP12T U4639 ( .A1(n5336), .A2(n5094), .B1(n5158), .B2(n5202), .C1(
        n5201), .C2(n5227), .ZN(register_file_inst1_n2422) );
  INVD1BWP12T U4640 ( .I(register_file_inst1_lr_29_), .ZN(n5337) );
  OAI222D1BWP12T U4641 ( .A1(n5337), .A2(n5222), .B1(n5160), .B2(n5202), .C1(
        n5201), .C2(n5223), .ZN(register_file_inst1_n2230) );
  CKND0BWP12T U4642 ( .I(register_file_inst1_r4_29_), .ZN(n5192) );
  OAI222D1BWP12T U4643 ( .A1(n5192), .A2(n5225), .B1(n5205), .B2(n5202), .C1(
        n5201), .C2(n5226), .ZN(register_file_inst1_n2518) );
  CKND0BWP12T U4644 ( .I(register_file_inst1_tmp1_29_), .ZN(n5193) );
  OAI222D1BWP12T U4645 ( .A1(n5193), .A2(n4683), .B1(n5212), .B2(n5202), .C1(
        n5201), .C2(n6144), .ZN(register_file_inst1_n2166) );
  CKND0BWP12T U4646 ( .I(register_file_inst1_r8_29_), .ZN(n5194) );
  OAI222D1BWP12T U4647 ( .A1(n5194), .A2(n5244), .B1(n5246), .B2(n5202), .C1(
        n5201), .C2(n5145), .ZN(register_file_inst1_n2390) );
  CKND0BWP12T U4648 ( .I(register_file_inst1_r12_29_), .ZN(n5195) );
  OAI222D1BWP12T U4649 ( .A1(n5195), .A2(n5242), .B1(n5243), .B2(n5202), .C1(
        n5201), .C2(n5140), .ZN(register_file_inst1_n2262) );
  INVD0BWP12T U4650 ( .I(register_file_inst1_r5_29_), .ZN(n5196) );
  OAI222D1BWP12T U4651 ( .A1(n5196), .A2(n5247), .B1(n5249), .B2(n5202), .C1(
        n5201), .C2(n5143), .ZN(register_file_inst1_n2486) );
  CKND0BWP12T U4652 ( .I(register_file_inst1_r9_29_), .ZN(n5197) );
  OAI222D1BWP12T U4653 ( .A1(n5197), .A2(n5235), .B1(n5237), .B2(n5202), .C1(
        n5201), .C2(n5238), .ZN(register_file_inst1_n2358) );
  INVD1BWP12T U4654 ( .I(register_file_inst1_r1_29_), .ZN(n5338) );
  OAI222D1BWP12T U4655 ( .A1(n5338), .A2(n5239), .B1(n5240), .B2(n5202), .C1(
        n5201), .C2(n5074), .ZN(register_file_inst1_n2614) );
  INVD1BWP12T U4656 ( .I(RF_next_sp[29]), .ZN(n5335) );
  OAI222D1BWP12T U4657 ( .A1(n5335), .A2(n5232), .B1(n5233), .B2(n5202), .C1(
        n5201), .C2(n5234), .ZN(register_file_inst1_spin[29]) );
  INVD0BWP12T U4658 ( .I(register_file_inst1_r11_29_), .ZN(n5198) );
  OAI222D1BWP12T U4659 ( .A1(n5198), .A2(n5217), .B1(n5219), .B2(n5202), .C1(
        n5201), .C2(n5220), .ZN(register_file_inst1_n2294) );
  INVD0BWP12T U4660 ( .I(register_file_inst1_r10_29_), .ZN(n5199) );
  OAI222D1BWP12T U4661 ( .A1(n5199), .A2(n5250), .B1(n5252), .B2(n5202), .C1(
        n5201), .C2(n5253), .ZN(register_file_inst1_n2326) );
  INVD1BWP12T U4662 ( .I(register_file_inst1_r2_29_), .ZN(n5325) );
  OAI222D1BWP12T U4663 ( .A1(n5325), .A2(n5254), .B1(n5256), .B2(n5202), .C1(
        n5201), .C2(n5257), .ZN(register_file_inst1_n2582) );
  INVD0BWP12T U4664 ( .I(register_file_inst1_r3_29_), .ZN(n5204) );
  OAI222D1BWP12T U4665 ( .A1(n5204), .A2(n4758), .B1(n5203), .B2(n5202), .C1(
        n5201), .C2(n5200), .ZN(register_file_inst1_n2550) );
  INVD1BWP12T U4666 ( .I(register_file_inst1_r0_30_), .ZN(n5299) );
  OAI222D1BWP12T U4667 ( .A1(n5299), .A2(n5096), .B1(n5230), .B2(n5266), .C1(
        n5268), .C2(n5231), .ZN(register_file_inst1_n2647) );
  INVD0BWP12T U4668 ( .I(register_file_inst1_r4_30_), .ZN(n5206) );
  OAI222D1BWP12T U4669 ( .A1(n5206), .A2(n5225), .B1(n5205), .B2(n5266), .C1(
        n5268), .C2(n5226), .ZN(register_file_inst1_n2519) );
  OAI222D1BWP12T U4670 ( .A1(n5207), .A2(n5242), .B1(n5243), .B2(n5266), .C1(
        n5268), .C2(n5140), .ZN(register_file_inst1_n2263) );
  INVD1BWP12T U4671 ( .I(register_file_inst1_r1_30_), .ZN(n5313) );
  OAI222D1BWP12T U4672 ( .A1(n5313), .A2(n5239), .B1(n5240), .B2(n5266), .C1(
        n5268), .C2(n5074), .ZN(register_file_inst1_n2615) );
  INVD0BWP12T U4673 ( .I(register_file_inst1_r9_30_), .ZN(n5208) );
  OAI222D1BWP12T U4674 ( .A1(n5208), .A2(n5235), .B1(n5237), .B2(n5266), .C1(
        n5268), .C2(n5238), .ZN(register_file_inst1_n2359) );
  OAI222D1BWP12T U4675 ( .A1(n5209), .A2(n5244), .B1(n5246), .B2(n5266), .C1(
        n5268), .C2(n5145), .ZN(register_file_inst1_n2391) );
  INVD0BWP12T U4676 ( .I(register_file_inst1_r5_30_), .ZN(n5210) );
  OAI222D1BWP12T U4677 ( .A1(n5210), .A2(n5247), .B1(n5249), .B2(n5266), .C1(
        n5268), .C2(n5143), .ZN(register_file_inst1_n2487) );
  INVD1BWP12T U4678 ( .I(RF_next_sp[30]), .ZN(n5310) );
  OAI222D1BWP12T U4679 ( .A1(n5310), .A2(n5232), .B1(n5233), .B2(n5266), .C1(
        n5268), .C2(n5234), .ZN(register_file_inst1_spin[30]) );
  OAI222D1BWP12T U4680 ( .A1(n5211), .A2(n5217), .B1(n5219), .B2(n5266), .C1(
        n5268), .C2(n5220), .ZN(register_file_inst1_n2295) );
  INVD0BWP12T U4681 ( .I(register_file_inst1_tmp1_30_), .ZN(n5213) );
  OAI222D1BWP12T U4682 ( .A1(n5213), .A2(n4683), .B1(n5212), .B2(n5266), .C1(
        n5268), .C2(n6144), .ZN(register_file_inst1_n2167) );
  INVD0BWP12T U4683 ( .I(register_file_inst1_r10_30_), .ZN(n5214) );
  OAI222D1BWP12T U4684 ( .A1(n5214), .A2(n5250), .B1(n5252), .B2(n5266), .C1(
        n5268), .C2(n5253), .ZN(register_file_inst1_n2327) );
  INVD1BWP12T U4685 ( .I(register_file_inst1_r2_30_), .ZN(n5300) );
  OAI222D1BWP12T U4686 ( .A1(n5300), .A2(n5254), .B1(n5256), .B2(n5266), .C1(
        n5268), .C2(n5257), .ZN(register_file_inst1_n2583) );
  NR2D1BWP12T U4687 ( .A1(n6323), .A2(n5216), .ZN(n5264) );
  INVD1BWP12T U4688 ( .I(n5264), .ZN(n6321) );
  OAI222D1BWP12T U4689 ( .A1(n5258), .A2(n5220), .B1(n5219), .B2(n5255), .C1(
        n5218), .C2(n5217), .ZN(register_file_inst1_n2296) );
  INVD0BWP12T U4690 ( .I(register_file_inst1_tmp1_31_), .ZN(n5221) );
  OAI222D1BWP12T U4691 ( .A1(n5258), .A2(n6144), .B1(n5212), .B2(n5255), .C1(
        n4683), .C2(n5221), .ZN(register_file_inst1_n2168) );
  INVD1BWP12T U4692 ( .I(register_file_inst1_lr_31_), .ZN(n5275) );
  OAI222D1BWP12T U4693 ( .A1(n5258), .A2(n5223), .B1(n5160), .B2(n5255), .C1(
        n5222), .C2(n5275), .ZN(register_file_inst1_n2232) );
  INVD0BWP12T U4694 ( .I(register_file_inst1_r4_31_), .ZN(n5224) );
  OAI222D1BWP12T U4695 ( .A1(n5258), .A2(n5226), .B1(n5205), .B2(n5255), .C1(
        n5225), .C2(n5224), .ZN(register_file_inst1_n2520) );
  INVD1BWP12T U4696 ( .I(register_file_inst1_r7_31_), .ZN(n5274) );
  OAI222D1BWP12T U4697 ( .A1(n5258), .A2(n5227), .B1(n5158), .B2(n5255), .C1(
        n5274), .C2(n5094), .ZN(register_file_inst1_n2424) );
  INVD1BWP12T U4698 ( .I(register_file_inst1_r6_31_), .ZN(n5286) );
  OAI222D1BWP12T U4699 ( .A1(n5258), .A2(n5229), .B1(n5228), .B2(n5255), .C1(
        n5286), .C2(n5095), .ZN(register_file_inst1_n2456) );
  INVD1BWP12T U4700 ( .I(register_file_inst1_r0_31_), .ZN(n5287) );
  OAI222D1BWP12T U4701 ( .A1(n5258), .A2(n5231), .B1(n5230), .B2(n5255), .C1(
        n5287), .C2(n5096), .ZN(register_file_inst1_n2648) );
  INVD1BWP12T U4702 ( .I(RF_next_sp[31]), .ZN(n5273) );
  OAI222D1BWP12T U4703 ( .A1(n5258), .A2(n5234), .B1(n5233), .B2(n5255), .C1(
        n5273), .C2(n5232), .ZN(register_file_inst1_spin[31]) );
  INVD0BWP12T U4704 ( .I(register_file_inst1_r9_31_), .ZN(n5236) );
  OAI222D1BWP12T U4705 ( .A1(n5258), .A2(n5238), .B1(n5237), .B2(n5255), .C1(
        n5236), .C2(n5235), .ZN(register_file_inst1_n2360) );
  INVD1BWP12T U4706 ( .I(register_file_inst1_r1_31_), .ZN(n5285) );
  OAI222D1BWP12T U4707 ( .A1(n5258), .A2(n5074), .B1(n5240), .B2(n5255), .C1(
        n5285), .C2(n5239), .ZN(register_file_inst1_n2616) );
  OAI222D1BWP12T U4708 ( .A1(n5258), .A2(n5140), .B1(n5243), .B2(n5255), .C1(
        n5242), .C2(n5241), .ZN(register_file_inst1_n2264) );
  OAI222D1BWP12T U4709 ( .A1(n5258), .A2(n5145), .B1(n5246), .B2(n5255), .C1(
        n5245), .C2(n5244), .ZN(register_file_inst1_n2392) );
  INVD0BWP12T U4710 ( .I(register_file_inst1_r5_31_), .ZN(n5248) );
  OAI222D1BWP12T U4711 ( .A1(n5258), .A2(n5143), .B1(n5249), .B2(n5255), .C1(
        n5248), .C2(n5247), .ZN(register_file_inst1_n2488) );
  INVD1BWP12T U4712 ( .I(n2871), .ZN(n6016) );
  INVD0BWP12T U4713 ( .I(register_file_inst1_r10_31_), .ZN(n5251) );
  OAI222D1BWP12T U4714 ( .A1(n5258), .A2(n5253), .B1(n5252), .B2(n5255), .C1(
        n5251), .C2(n5250), .ZN(register_file_inst1_n2328) );
  INVD1BWP12T U4715 ( .I(register_file_inst1_r2_31_), .ZN(n5288) );
  OAI222D1BWP12T U4716 ( .A1(n5258), .A2(n5257), .B1(n5256), .B2(n5255), .C1(
        n5288), .C2(n5254), .ZN(register_file_inst1_n2584) );
  INVD1BWP12T U4717 ( .I(ALU_OUT_z), .ZN(n6390) );
  OAI222D1BWP12T U4718 ( .A1(n5260), .A2(n5269), .B1(n5267), .B2(n5259), .C1(
        n5270), .C2(n6325), .ZN(n6322) );
  OAI222D1BWP12T U4719 ( .A1(n5262), .A2(n5269), .B1(n5267), .B2(n5261), .C1(
        n5270), .C2(n6323), .ZN(n6320) );
  CKND0BWP12T U4720 ( .I(n5263), .ZN(n5265) );
  AO222D1BWP12T U4721 ( .A1(n5265), .A2(n6379), .B1(n6376), .B2(
        ALU_MISC_OUT_result[26]), .C1(n6395), .C2(n5264), .Z(n6318) );
  OAI21D1BWP12T U4722 ( .A1(n5272), .A2(n5271), .B(n6311), .ZN(
        register_file_inst1_n2199) );
  OAI22D1BWP12T U4723 ( .A1(n5274), .A2(n5938), .B1(n5273), .B2(n6222), .ZN(
        n5284) );
  OAI22D1BWP12T U4724 ( .A1(n5285), .A2(n5942), .B1(n5275), .B2(n5940), .ZN(
        n5283) );
  AOI22D1BWP12T U4725 ( .A1(register_file_inst1_tmp1_31_), .A2(n5979), .B1(
        register_file_inst1_r10_31_), .B2(n6223), .ZN(n5277) );
  AOI22D1BWP12T U4726 ( .A1(register_file_inst1_r4_31_), .A2(n5900), .B1(
        register_file_inst1_r9_31_), .B2(n6225), .ZN(n5276) );
  ND3D1BWP12T U4727 ( .A1(n5277), .A2(n5276), .A3(n6227), .ZN(n5282) );
  AOI22D1BWP12T U4728 ( .A1(register_file_inst1_r0_31_), .A2(n6004), .B1(
        register_file_inst1_r6_31_), .B2(n6003), .ZN(n5280) );
  AOI22D1BWP12T U4729 ( .A1(register_file_inst1_r11_31_), .A2(n6229), .B1(
        register_file_inst1_r3_31_), .B2(n5946), .ZN(n5279) );
  AOI22D1BWP12T U4730 ( .A1(register_file_inst1_r5_31_), .A2(n5948), .B1(
        register_file_inst1_r8_31_), .B2(n5947), .ZN(n5278) );
  ND4D1BWP12T U4731 ( .A1(n5280), .A2(n6231), .A3(n5279), .A4(n5278), .ZN(
        n5281) );
  OR4XD1BWP12T U4732 ( .A1(n5284), .A2(n5283), .A3(n5282), .A4(n5281), .Z(
        RF_ALU_operand_a[31]) );
  OAI22D1BWP12T U4733 ( .A1(n5286), .A2(n5910), .B1(n5285), .B2(n5857), .ZN(
        n5297) );
  OAI22D1BWP12T U4734 ( .A1(n5288), .A2(n5959), .B1(n5287), .B2(n5912), .ZN(
        n5296) );
  AOI22D1BWP12T U4735 ( .A1(register_file_inst1_tmp1_31_), .A2(n5962), .B1(
        register_file_inst1_r4_31_), .B2(n5961), .ZN(n5290) );
  AOI22D1BWP12T U4736 ( .A1(RF_next_sp[31]), .A2(n5964), .B1(
        register_file_inst1_r12_31_), .B2(n5963), .ZN(n5289) );
  ND3D1BWP12T U4737 ( .A1(n5290), .A2(n5289), .A3(n6145), .ZN(n5295) );
  AOI22D1BWP12T U4738 ( .A1(register_file_inst1_r9_31_), .A2(n5968), .B1(
        register_file_inst1_r3_31_), .B2(n5967), .ZN(n5293) );
  AOI22D1BWP12T U4739 ( .A1(register_file_inst1_r7_31_), .A2(n6001), .B1(
        register_file_inst1_r11_31_), .B2(n5969), .ZN(n5292) );
  AOI22D1BWP12T U4740 ( .A1(register_file_inst1_r5_31_), .A2(n6002), .B1(
        register_file_inst1_lr_31_), .B2(n5970), .ZN(n5291) );
  ND4D1BWP12T U4741 ( .A1(n5293), .A2(n5292), .A3(n6146), .A4(n5291), .ZN(
        n5294) );
  OR4XD1BWP12T U4742 ( .A1(n5297), .A2(n5296), .A3(n5295), .A4(n5294), .Z(
        RF_ALU_operand_b[31]) );
  OAI22D1BWP12T U4743 ( .A1(n5298), .A2(n5910), .B1(n5313), .B2(n5857), .ZN(
        n5309) );
  OAI22D1BWP12T U4744 ( .A1(n5300), .A2(n5959), .B1(n5299), .B2(n5912), .ZN(
        n5308) );
  AOI22D1BWP12T U4745 ( .A1(register_file_inst1_tmp1_30_), .A2(n5962), .B1(
        register_file_inst1_r4_30_), .B2(n5961), .ZN(n5302) );
  AOI22D1BWP12T U4746 ( .A1(RF_next_sp[30]), .A2(n5964), .B1(
        register_file_inst1_r12_30_), .B2(n5963), .ZN(n5301) );
  ND3D1BWP12T U4747 ( .A1(n5302), .A2(n5301), .A3(n6142), .ZN(n5307) );
  AOI22D1BWP12T U4748 ( .A1(register_file_inst1_r9_30_), .A2(n5968), .B1(
        register_file_inst1_r3_30_), .B2(n5967), .ZN(n5305) );
  AOI22D1BWP12T U4749 ( .A1(register_file_inst1_r7_30_), .A2(n6001), .B1(
        register_file_inst1_r11_30_), .B2(n5969), .ZN(n5304) );
  AOI22D1BWP12T U4750 ( .A1(register_file_inst1_r5_30_), .A2(n6002), .B1(
        register_file_inst1_lr_30_), .B2(n5970), .ZN(n5303) );
  ND4D1BWP12T U4751 ( .A1(n5305), .A2(n5304), .A3(n6143), .A4(n5303), .ZN(
        n5306) );
  OR4XD1BWP12T U4752 ( .A1(n5309), .A2(n5308), .A3(n5307), .A4(n5306), .Z(
        RF_ALU_operand_b[30]) );
  OAI22D1BWP12T U4753 ( .A1(n5311), .A2(n5938), .B1(n5310), .B2(n6222), .ZN(
        n5322) );
  OAI22D1BWP12T U4754 ( .A1(n5313), .A2(n5942), .B1(n5312), .B2(n5940), .ZN(
        n5321) );
  AOI22D1BWP12T U4755 ( .A1(register_file_inst1_tmp1_30_), .A2(n5979), .B1(
        register_file_inst1_r10_30_), .B2(n6223), .ZN(n5315) );
  BUFFD1BWP12T U4756 ( .I(n6225), .Z(n5943) );
  AOI22D1BWP12T U4757 ( .A1(register_file_inst1_r4_30_), .A2(n5900), .B1(
        register_file_inst1_r9_30_), .B2(n5943), .ZN(n5314) );
  ND3D1BWP12T U4758 ( .A1(n5315), .A2(n5314), .A3(n6220), .ZN(n5320) );
  AOI22D1BWP12T U4759 ( .A1(register_file_inst1_r0_30_), .A2(n6004), .B1(
        register_file_inst1_r6_30_), .B2(n6003), .ZN(n5318) );
  AOI22D1BWP12T U4760 ( .A1(register_file_inst1_r11_30_), .A2(n6229), .B1(
        register_file_inst1_r3_30_), .B2(n5946), .ZN(n5317) );
  AOI22D1BWP12T U4761 ( .A1(register_file_inst1_r5_30_), .A2(n5948), .B1(
        register_file_inst1_r8_30_), .B2(n5947), .ZN(n5316) );
  ND4D1BWP12T U4762 ( .A1(n5318), .A2(n6221), .A3(n5317), .A4(n5316), .ZN(
        n5319) );
  OR4XD1BWP12T U4763 ( .A1(n5322), .A2(n5321), .A3(n5320), .A4(n5319), .Z(
        RF_ALU_operand_a[30]) );
  OAI22D1BWP12T U4764 ( .A1(n5323), .A2(n5910), .B1(n5338), .B2(n5857), .ZN(
        n5334) );
  OAI22D1BWP12T U4765 ( .A1(n5325), .A2(n5959), .B1(n5324), .B2(n5912), .ZN(
        n5333) );
  AOI22D1BWP12T U4766 ( .A1(register_file_inst1_tmp1_29_), .A2(n5962), .B1(
        register_file_inst1_r4_29_), .B2(n5961), .ZN(n5327) );
  AOI22D1BWP12T U4767 ( .A1(RF_next_sp[29]), .A2(n5964), .B1(
        register_file_inst1_r12_29_), .B2(n5963), .ZN(n5326) );
  ND3D1BWP12T U4768 ( .A1(n5327), .A2(n5326), .A3(n6140), .ZN(n5332) );
  AOI22D1BWP12T U4769 ( .A1(register_file_inst1_r9_29_), .A2(n5968), .B1(
        register_file_inst1_r3_29_), .B2(n5967), .ZN(n5330) );
  AOI22D1BWP12T U4770 ( .A1(register_file_inst1_r7_29_), .A2(n6001), .B1(
        register_file_inst1_r11_29_), .B2(n5969), .ZN(n5329) );
  AOI22D1BWP12T U4771 ( .A1(register_file_inst1_r5_29_), .A2(n6002), .B1(
        register_file_inst1_lr_29_), .B2(n5970), .ZN(n5328) );
  ND4D1BWP12T U4772 ( .A1(n5330), .A2(n5329), .A3(n6141), .A4(n5328), .ZN(
        n5331) );
  OR4XD1BWP12T U4773 ( .A1(n5334), .A2(n5333), .A3(n5332), .A4(n5331), .Z(
        RF_ALU_operand_b[29]) );
  OAI22D1BWP12T U4774 ( .A1(n5336), .A2(n5938), .B1(n5335), .B2(n6222), .ZN(
        n5347) );
  OAI22D1BWP12T U4775 ( .A1(n5338), .A2(n5942), .B1(n5337), .B2(n5940), .ZN(
        n5346) );
  AOI22D1BWP12T U4776 ( .A1(register_file_inst1_tmp1_29_), .A2(n5979), .B1(
        register_file_inst1_r10_29_), .B2(n6223), .ZN(n5340) );
  AOI22D1BWP12T U4777 ( .A1(register_file_inst1_r4_29_), .A2(n5900), .B1(
        register_file_inst1_r9_29_), .B2(n5943), .ZN(n5339) );
  ND3D1BWP12T U4778 ( .A1(n5340), .A2(n5339), .A3(n6218), .ZN(n5345) );
  AOI22D1BWP12T U4779 ( .A1(register_file_inst1_r0_29_), .A2(n6004), .B1(
        register_file_inst1_r6_29_), .B2(n6003), .ZN(n5343) );
  AOI22D1BWP12T U4780 ( .A1(register_file_inst1_r11_29_), .A2(n6229), .B1(
        register_file_inst1_r3_29_), .B2(n5946), .ZN(n5342) );
  AOI22D1BWP12T U4781 ( .A1(register_file_inst1_r5_29_), .A2(n5948), .B1(
        register_file_inst1_r8_29_), .B2(n5947), .ZN(n5341) );
  ND4D1BWP12T U4782 ( .A1(n5343), .A2(n6219), .A3(n5342), .A4(n5341), .ZN(
        n5344) );
  OR4XD1BWP12T U4783 ( .A1(n5347), .A2(n5346), .A3(n5345), .A4(n5344), .Z(
        RF_ALU_operand_a[29]) );
  OAI22D1BWP12T U4784 ( .A1(n5348), .A2(n5910), .B1(n5363), .B2(n5857), .ZN(
        n5359) );
  OAI22D1BWP12T U4785 ( .A1(n5350), .A2(n5959), .B1(n5349), .B2(n5912), .ZN(
        n5358) );
  AOI22D1BWP12T U4786 ( .A1(register_file_inst1_tmp1_28_), .A2(n5962), .B1(
        register_file_inst1_r4_28_), .B2(n5961), .ZN(n5352) );
  AOI22D1BWP12T U4787 ( .A1(RF_next_sp[28]), .A2(n5964), .B1(
        register_file_inst1_r12_28_), .B2(n5963), .ZN(n5351) );
  ND3D1BWP12T U4788 ( .A1(n5352), .A2(n5351), .A3(n6138), .ZN(n5357) );
  AOI22D1BWP12T U4789 ( .A1(register_file_inst1_r9_28_), .A2(n5968), .B1(
        register_file_inst1_r3_28_), .B2(n5967), .ZN(n5355) );
  AOI22D1BWP12T U4790 ( .A1(register_file_inst1_r7_28_), .A2(n6001), .B1(
        register_file_inst1_r11_28_), .B2(n5969), .ZN(n5354) );
  AOI22D1BWP12T U4791 ( .A1(register_file_inst1_r5_28_), .A2(n6002), .B1(
        register_file_inst1_lr_28_), .B2(n5970), .ZN(n5353) );
  ND4D1BWP12T U4792 ( .A1(n5355), .A2(n5354), .A3(n6139), .A4(n5353), .ZN(
        n5356) );
  OR4XD1BWP12T U4793 ( .A1(n5359), .A2(n5358), .A3(n5357), .A4(n5356), .Z(
        RF_ALU_operand_b[28]) );
  OAI22D1BWP12T U4794 ( .A1(n5361), .A2(n5938), .B1(n5360), .B2(n6222), .ZN(
        n5372) );
  OAI22D1BWP12T U4795 ( .A1(n5363), .A2(n5942), .B1(n5362), .B2(n5940), .ZN(
        n5371) );
  AOI22D1BWP12T U4796 ( .A1(register_file_inst1_tmp1_28_), .A2(n5979), .B1(
        register_file_inst1_r10_28_), .B2(n6223), .ZN(n5365) );
  AOI22D1BWP12T U4797 ( .A1(register_file_inst1_r4_28_), .A2(n5900), .B1(
        register_file_inst1_r9_28_), .B2(n5943), .ZN(n5364) );
  ND3D1BWP12T U4798 ( .A1(n5365), .A2(n5364), .A3(n6216), .ZN(n5370) );
  AOI22D1BWP12T U4799 ( .A1(register_file_inst1_r0_28_), .A2(n6004), .B1(
        register_file_inst1_r6_28_), .B2(n6003), .ZN(n5368) );
  AOI22D1BWP12T U4800 ( .A1(register_file_inst1_r11_28_), .A2(n6229), .B1(
        register_file_inst1_r3_28_), .B2(n5946), .ZN(n5367) );
  AOI22D1BWP12T U4801 ( .A1(register_file_inst1_r5_28_), .A2(n5948), .B1(
        register_file_inst1_r8_28_), .B2(n5947), .ZN(n5366) );
  ND4D1BWP12T U4802 ( .A1(n5368), .A2(n6217), .A3(n5367), .A4(n5366), .ZN(
        n5369) );
  OR4XD1BWP12T U4803 ( .A1(n5372), .A2(n5371), .A3(n5370), .A4(n5369), .Z(
        RF_ALU_operand_a[28]) );
  OAI22D1BWP12T U4804 ( .A1(n5373), .A2(n5910), .B1(n5388), .B2(n5857), .ZN(
        n5384) );
  OAI22D1BWP12T U4805 ( .A1(n5375), .A2(n5959), .B1(n5374), .B2(n5912), .ZN(
        n5383) );
  AOI22D1BWP12T U4806 ( .A1(register_file_inst1_tmp1_27_), .A2(n5962), .B1(
        register_file_inst1_r4_27_), .B2(n5961), .ZN(n5377) );
  AOI22D1BWP12T U4807 ( .A1(RF_next_sp[27]), .A2(n5964), .B1(
        register_file_inst1_r12_27_), .B2(n5963), .ZN(n5376) );
  ND3D1BWP12T U4808 ( .A1(n5377), .A2(n5376), .A3(n6136), .ZN(n5382) );
  AOI22D1BWP12T U4809 ( .A1(register_file_inst1_r9_27_), .A2(n5968), .B1(
        register_file_inst1_r3_27_), .B2(n5967), .ZN(n5380) );
  AOI22D1BWP12T U4810 ( .A1(register_file_inst1_r7_27_), .A2(n6001), .B1(
        register_file_inst1_r11_27_), .B2(n5969), .ZN(n5379) );
  AOI22D1BWP12T U4811 ( .A1(register_file_inst1_r5_27_), .A2(n6002), .B1(
        register_file_inst1_lr_27_), .B2(n5970), .ZN(n5378) );
  ND4D1BWP12T U4812 ( .A1(n5380), .A2(n5379), .A3(n6137), .A4(n5378), .ZN(
        n5381) );
  OR4XD1BWP12T U4813 ( .A1(n5384), .A2(n5383), .A3(n5382), .A4(n5381), .Z(
        RF_ALU_operand_b[27]) );
  OAI22D1BWP12T U4814 ( .A1(n5386), .A2(n5938), .B1(n5385), .B2(n6222), .ZN(
        n5397) );
  OAI22D1BWP12T U4815 ( .A1(n5388), .A2(n5942), .B1(n5387), .B2(n5940), .ZN(
        n5396) );
  AOI22D1BWP12T U4816 ( .A1(register_file_inst1_tmp1_27_), .A2(n6224), .B1(
        register_file_inst1_r10_27_), .B2(n6223), .ZN(n5390) );
  AOI22D1BWP12T U4817 ( .A1(register_file_inst1_r4_27_), .A2(n5900), .B1(
        register_file_inst1_r9_27_), .B2(n5943), .ZN(n5389) );
  ND3D1BWP12T U4818 ( .A1(n5390), .A2(n5389), .A3(n6214), .ZN(n5395) );
  AOI22D1BWP12T U4819 ( .A1(register_file_inst1_r0_27_), .A2(n6004), .B1(
        register_file_inst1_r6_27_), .B2(n6003), .ZN(n5393) );
  AOI22D1BWP12T U4820 ( .A1(register_file_inst1_r11_27_), .A2(n6229), .B1(
        register_file_inst1_r3_27_), .B2(n5946), .ZN(n5392) );
  AOI22D1BWP12T U4821 ( .A1(register_file_inst1_r5_27_), .A2(n5948), .B1(
        register_file_inst1_r8_27_), .B2(n5947), .ZN(n5391) );
  ND4D1BWP12T U4822 ( .A1(n5393), .A2(n6215), .A3(n5392), .A4(n5391), .ZN(
        n5394) );
  OR4XD1BWP12T U4823 ( .A1(n5397), .A2(n5396), .A3(n5395), .A4(n5394), .Z(
        RF_ALU_operand_a[27]) );
  OAI22D1BWP12T U4824 ( .A1(n5399), .A2(n5938), .B1(n5398), .B2(n6222), .ZN(
        n5409) );
  OAI22D1BWP12T U4825 ( .A1(n5410), .A2(n5942), .B1(n5400), .B2(n5940), .ZN(
        n5408) );
  AOI22D1BWP12T U4826 ( .A1(register_file_inst1_tmp1_24_), .A2(n5979), .B1(
        register_file_inst1_r10_24_), .B2(n6223), .ZN(n5402) );
  AOI22D1BWP12T U4827 ( .A1(register_file_inst1_r4_24_), .A2(n5900), .B1(
        register_file_inst1_r9_24_), .B2(n5943), .ZN(n5401) );
  ND3D1BWP12T U4828 ( .A1(n5402), .A2(n5401), .A3(n6208), .ZN(n5407) );
  AOI22D1BWP12T U4829 ( .A1(register_file_inst1_r0_24_), .A2(n6004), .B1(
        register_file_inst1_r6_24_), .B2(n6003), .ZN(n5405) );
  AOI22D1BWP12T U4830 ( .A1(register_file_inst1_r11_24_), .A2(n6229), .B1(
        register_file_inst1_r3_24_), .B2(n5946), .ZN(n5404) );
  AOI22D1BWP12T U4831 ( .A1(register_file_inst1_r5_24_), .A2(n5948), .B1(
        register_file_inst1_r8_24_), .B2(n5947), .ZN(n5403) );
  ND4D1BWP12T U4832 ( .A1(n5405), .A2(n6209), .A3(n5404), .A4(n5403), .ZN(
        n5406) );
  OR4XD1BWP12T U4833 ( .A1(n5409), .A2(n5408), .A3(n5407), .A4(n5406), .Z(
        RF_ALU_operand_a[24]) );
  OAI22D1BWP12T U4834 ( .A1(n5411), .A2(n5910), .B1(n5410), .B2(n5857), .ZN(
        n5422) );
  OAI22D1BWP12T U4835 ( .A1(n5413), .A2(n5959), .B1(n5412), .B2(n5912), .ZN(
        n5421) );
  AOI22D1BWP12T U4836 ( .A1(register_file_inst1_tmp1_24_), .A2(n5962), .B1(
        register_file_inst1_r4_24_), .B2(n5961), .ZN(n5415) );
  AOI22D1BWP12T U4837 ( .A1(RF_next_sp[24]), .A2(n5964), .B1(
        register_file_inst1_r12_24_), .B2(n5963), .ZN(n5414) );
  ND3D1BWP12T U4838 ( .A1(n5415), .A2(n5414), .A3(n6130), .ZN(n5420) );
  AOI22D1BWP12T U4839 ( .A1(register_file_inst1_r9_24_), .A2(n5968), .B1(
        register_file_inst1_r3_24_), .B2(n5967), .ZN(n5418) );
  AOI22D1BWP12T U4840 ( .A1(register_file_inst1_r7_24_), .A2(n6001), .B1(
        register_file_inst1_r11_24_), .B2(n5969), .ZN(n5417) );
  AOI22D1BWP12T U4841 ( .A1(register_file_inst1_r5_24_), .A2(n6002), .B1(
        register_file_inst1_lr_24_), .B2(n5970), .ZN(n5416) );
  ND4D1BWP12T U4842 ( .A1(n5418), .A2(n5417), .A3(n6131), .A4(n5416), .ZN(
        n5419) );
  OR4XD1BWP12T U4843 ( .A1(n5422), .A2(n5421), .A3(n5420), .A4(n5419), .Z(
        RF_ALU_operand_b[24]) );
  OAI22D1BWP12T U4844 ( .A1(n5423), .A2(n5910), .B1(n5438), .B2(n5857), .ZN(
        n5434) );
  OAI22D1BWP12T U4845 ( .A1(n5425), .A2(n5959), .B1(n5424), .B2(n5912), .ZN(
        n5433) );
  AOI22D1BWP12T U4846 ( .A1(register_file_inst1_tmp1_23_), .A2(n5962), .B1(
        register_file_inst1_r4_23_), .B2(n5961), .ZN(n5427) );
  AOI22D1BWP12T U4847 ( .A1(RF_next_sp[23]), .A2(n5964), .B1(
        register_file_inst1_r12_23_), .B2(n5963), .ZN(n5426) );
  ND3D1BWP12T U4848 ( .A1(n5427), .A2(n5426), .A3(n6128), .ZN(n5432) );
  AOI22D1BWP12T U4849 ( .A1(register_file_inst1_r9_23_), .A2(n5968), .B1(
        register_file_inst1_r3_23_), .B2(n5967), .ZN(n5430) );
  AOI22D1BWP12T U4850 ( .A1(register_file_inst1_r7_23_), .A2(n6001), .B1(
        register_file_inst1_r11_23_), .B2(n5969), .ZN(n5429) );
  AOI22D1BWP12T U4851 ( .A1(register_file_inst1_r5_23_), .A2(n6002), .B1(
        register_file_inst1_lr_23_), .B2(n5970), .ZN(n5428) );
  ND4D1BWP12T U4852 ( .A1(n5430), .A2(n5429), .A3(n6129), .A4(n5428), .ZN(
        n5431) );
  OR4XD1BWP12T U4853 ( .A1(n5434), .A2(n5433), .A3(n5432), .A4(n5431), .Z(
        RF_ALU_operand_b[23]) );
  OAI22D1BWP12T U4854 ( .A1(n5436), .A2(n5938), .B1(n5435), .B2(n6222), .ZN(
        n5447) );
  OAI22D1BWP12T U4855 ( .A1(n5438), .A2(n5942), .B1(n5437), .B2(n5940), .ZN(
        n5446) );
  AOI22D1BWP12T U4856 ( .A1(register_file_inst1_tmp1_23_), .A2(n5979), .B1(
        register_file_inst1_r10_23_), .B2(n6223), .ZN(n5440) );
  AOI22D1BWP12T U4857 ( .A1(register_file_inst1_r4_23_), .A2(n5900), .B1(
        register_file_inst1_r9_23_), .B2(n6225), .ZN(n5439) );
  ND3D1BWP12T U4858 ( .A1(n5440), .A2(n5439), .A3(n6206), .ZN(n5445) );
  AOI22D1BWP12T U4859 ( .A1(register_file_inst1_r0_23_), .A2(n6004), .B1(
        register_file_inst1_r6_23_), .B2(n6003), .ZN(n5443) );
  AOI22D1BWP12T U4860 ( .A1(register_file_inst1_r11_23_), .A2(n6229), .B1(
        register_file_inst1_r3_23_), .B2(n5946), .ZN(n5442) );
  AOI22D1BWP12T U4861 ( .A1(register_file_inst1_r5_23_), .A2(n5948), .B1(
        register_file_inst1_r8_23_), .B2(n5947), .ZN(n5441) );
  ND4D1BWP12T U4862 ( .A1(n5443), .A2(n6207), .A3(n5442), .A4(n5441), .ZN(
        n5444) );
  OR4XD1BWP12T U4863 ( .A1(n5447), .A2(n5446), .A3(n5445), .A4(n5444), .Z(
        RF_ALU_operand_a[23]) );
  OAI22D1BWP12T U4864 ( .A1(n5448), .A2(n5910), .B1(n5463), .B2(n5857), .ZN(
        n5459) );
  OAI22D1BWP12T U4865 ( .A1(n5450), .A2(n5959), .B1(n5449), .B2(n5912), .ZN(
        n5458) );
  AOI22D1BWP12T U4866 ( .A1(register_file_inst1_tmp1_22_), .A2(n5962), .B1(
        register_file_inst1_r4_22_), .B2(n5961), .ZN(n5452) );
  AOI22D1BWP12T U4867 ( .A1(RF_next_sp[22]), .A2(n5964), .B1(
        register_file_inst1_r12_22_), .B2(n5963), .ZN(n5451) );
  ND3D1BWP12T U4868 ( .A1(n5452), .A2(n5451), .A3(n6126), .ZN(n5457) );
  AOI22D1BWP12T U4869 ( .A1(register_file_inst1_r9_22_), .A2(n5968), .B1(
        register_file_inst1_r3_22_), .B2(n5967), .ZN(n5455) );
  AOI22D1BWP12T U4870 ( .A1(register_file_inst1_r7_22_), .A2(n6001), .B1(
        register_file_inst1_r11_22_), .B2(n5969), .ZN(n5454) );
  AOI22D1BWP12T U4871 ( .A1(register_file_inst1_r5_22_), .A2(n6002), .B1(
        register_file_inst1_lr_22_), .B2(n5970), .ZN(n5453) );
  ND4D1BWP12T U4872 ( .A1(n5455), .A2(n5454), .A3(n6127), .A4(n5453), .ZN(
        n5456) );
  OR4XD1BWP12T U4873 ( .A1(n5459), .A2(n5458), .A3(n5457), .A4(n5456), .Z(
        RF_ALU_operand_b[22]) );
  OAI22D1BWP12T U4874 ( .A1(n5461), .A2(n5938), .B1(n5460), .B2(n6222), .ZN(
        n5472) );
  OAI22D1BWP12T U4875 ( .A1(n5463), .A2(n5942), .B1(n5462), .B2(n5940), .ZN(
        n5471) );
  AOI22D1BWP12T U4876 ( .A1(register_file_inst1_tmp1_22_), .A2(n5979), .B1(
        register_file_inst1_r10_22_), .B2(n6223), .ZN(n5465) );
  AOI22D1BWP12T U4877 ( .A1(register_file_inst1_r4_22_), .A2(n5900), .B1(
        register_file_inst1_r9_22_), .B2(n5943), .ZN(n5464) );
  ND3D1BWP12T U4878 ( .A1(n5465), .A2(n5464), .A3(n6204), .ZN(n5470) );
  AOI22D1BWP12T U4879 ( .A1(register_file_inst1_r0_22_), .A2(n6004), .B1(
        register_file_inst1_r6_22_), .B2(n6003), .ZN(n5468) );
  AOI22D1BWP12T U4880 ( .A1(register_file_inst1_r11_22_), .A2(n6229), .B1(
        register_file_inst1_r3_22_), .B2(n5946), .ZN(n5467) );
  AOI22D1BWP12T U4881 ( .A1(register_file_inst1_r5_22_), .A2(n5948), .B1(
        register_file_inst1_r8_22_), .B2(n6230), .ZN(n5466) );
  ND4D1BWP12T U4882 ( .A1(n5468), .A2(n6205), .A3(n5467), .A4(n5466), .ZN(
        n5469) );
  OR4XD1BWP12T U4883 ( .A1(n5472), .A2(n5471), .A3(n5470), .A4(n5469), .Z(
        RF_ALU_operand_a[22]) );
  OAI22D1BWP12T U4884 ( .A1(n5474), .A2(n5938), .B1(n5473), .B2(n6222), .ZN(
        n5485) );
  OAI22D1BWP12T U4885 ( .A1(n5476), .A2(n5942), .B1(n5475), .B2(n5940), .ZN(
        n5484) );
  AOI22D1BWP12T U4886 ( .A1(register_file_inst1_tmp1_19_), .A2(n5979), .B1(
        register_file_inst1_r10_19_), .B2(n6223), .ZN(n5478) );
  AOI22D1BWP12T U4887 ( .A1(register_file_inst1_r4_19_), .A2(n5900), .B1(
        register_file_inst1_r9_19_), .B2(n6225), .ZN(n5477) );
  ND3D1BWP12T U4888 ( .A1(n5478), .A2(n5477), .A3(n6198), .ZN(n5483) );
  AOI22D1BWP12T U4889 ( .A1(register_file_inst1_r0_19_), .A2(n6004), .B1(
        register_file_inst1_r6_19_), .B2(n6003), .ZN(n5481) );
  AOI22D1BWP12T U4890 ( .A1(register_file_inst1_r11_19_), .A2(n6229), .B1(
        register_file_inst1_r3_19_), .B2(n5946), .ZN(n5480) );
  AOI22D1BWP12T U4891 ( .A1(register_file_inst1_r5_19_), .A2(n5948), .B1(
        register_file_inst1_r8_19_), .B2(n5947), .ZN(n5479) );
  ND4D1BWP12T U4892 ( .A1(n5481), .A2(n6199), .A3(n5480), .A4(n5479), .ZN(
        n5482) );
  OR4XD1BWP12T U4893 ( .A1(n5485), .A2(n5484), .A3(n5483), .A4(n5482), .Z(
        RF_ALU_operand_a[19]) );
  OAI22D1BWP12T U4894 ( .A1(n5486), .A2(n5910), .B1(n5501), .B2(n5857), .ZN(
        n5497) );
  OAI22D1BWP12T U4895 ( .A1(n5488), .A2(n5959), .B1(n5487), .B2(n5912), .ZN(
        n5496) );
  AOI22D1BWP12T U4896 ( .A1(register_file_inst1_tmp1_18_), .A2(n5962), .B1(
        register_file_inst1_r4_18_), .B2(n5961), .ZN(n5490) );
  AOI22D1BWP12T U4897 ( .A1(RF_next_sp[18]), .A2(n5964), .B1(
        register_file_inst1_r12_18_), .B2(n5963), .ZN(n5489) );
  ND3D1BWP12T U4898 ( .A1(n5490), .A2(n5489), .A3(n6118), .ZN(n5495) );
  AOI22D1BWP12T U4899 ( .A1(register_file_inst1_r9_18_), .A2(n5968), .B1(
        register_file_inst1_r3_18_), .B2(n5967), .ZN(n5493) );
  AOI22D1BWP12T U4900 ( .A1(register_file_inst1_r7_18_), .A2(n6001), .B1(
        register_file_inst1_r11_18_), .B2(n5969), .ZN(n5492) );
  AOI22D1BWP12T U4901 ( .A1(register_file_inst1_r5_18_), .A2(n6002), .B1(
        register_file_inst1_lr_18_), .B2(n5970), .ZN(n5491) );
  ND4D1BWP12T U4902 ( .A1(n5493), .A2(n5492), .A3(n6119), .A4(n5491), .ZN(
        n5494) );
  OR4XD1BWP12T U4903 ( .A1(n5497), .A2(n5496), .A3(n5495), .A4(n5494), .Z(
        RF_ALU_operand_b[18]) );
  OAI22D1BWP12T U4904 ( .A1(n5499), .A2(n5938), .B1(n5498), .B2(n6222), .ZN(
        n5510) );
  OAI22D1BWP12T U4905 ( .A1(n5501), .A2(n5942), .B1(n5500), .B2(n5940), .ZN(
        n5509) );
  AOI22D1BWP12T U4906 ( .A1(register_file_inst1_tmp1_18_), .A2(n5979), .B1(
        register_file_inst1_r10_18_), .B2(n6223), .ZN(n5503) );
  AOI22D1BWP12T U4907 ( .A1(register_file_inst1_r4_18_), .A2(n5900), .B1(
        register_file_inst1_r9_18_), .B2(n5943), .ZN(n5502) );
  ND3D1BWP12T U4908 ( .A1(n5503), .A2(n5502), .A3(n6196), .ZN(n5508) );
  AOI22D1BWP12T U4909 ( .A1(register_file_inst1_r0_18_), .A2(n6004), .B1(
        register_file_inst1_r6_18_), .B2(n6003), .ZN(n5506) );
  AOI22D1BWP12T U4910 ( .A1(register_file_inst1_r11_18_), .A2(n6229), .B1(
        register_file_inst1_r3_18_), .B2(n5946), .ZN(n5505) );
  AOI22D1BWP12T U4911 ( .A1(register_file_inst1_r5_18_), .A2(n5948), .B1(
        register_file_inst1_r8_18_), .B2(n6230), .ZN(n5504) );
  ND4D1BWP12T U4912 ( .A1(n5506), .A2(n6197), .A3(n5505), .A4(n5504), .ZN(
        n5507) );
  OR4XD1BWP12T U4913 ( .A1(n5510), .A2(n5509), .A3(n5508), .A4(n5507), .Z(
        RF_ALU_operand_a[18]) );
  OAI22D1BWP12T U4914 ( .A1(n5512), .A2(n5938), .B1(n5511), .B2(n6222), .ZN(
        n5523) );
  OAI22D1BWP12T U4915 ( .A1(n5514), .A2(n5942), .B1(n5513), .B2(n5940), .ZN(
        n5522) );
  AOI22D1BWP12T U4916 ( .A1(register_file_inst1_tmp1_17_), .A2(n5979), .B1(
        register_file_inst1_r10_17_), .B2(n6223), .ZN(n5516) );
  AOI22D1BWP12T U4917 ( .A1(register_file_inst1_r4_17_), .A2(n5900), .B1(
        register_file_inst1_r9_17_), .B2(n6225), .ZN(n5515) );
  ND3D1BWP12T U4918 ( .A1(n5516), .A2(n5515), .A3(n6194), .ZN(n5521) );
  AOI22D1BWP12T U4919 ( .A1(register_file_inst1_r0_17_), .A2(n6004), .B1(
        register_file_inst1_r6_17_), .B2(n6003), .ZN(n5519) );
  AOI22D1BWP12T U4920 ( .A1(register_file_inst1_r11_17_), .A2(n6229), .B1(
        register_file_inst1_r3_17_), .B2(n5946), .ZN(n5518) );
  AOI22D1BWP12T U4921 ( .A1(register_file_inst1_r5_17_), .A2(n5948), .B1(
        register_file_inst1_r8_17_), .B2(n5947), .ZN(n5517) );
  ND4D1BWP12T U4922 ( .A1(n5519), .A2(n6195), .A3(n5518), .A4(n5517), .ZN(
        n5520) );
  OR4XD1BWP12T U4923 ( .A1(n5523), .A2(n5522), .A3(n5521), .A4(n5520), .Z(
        RF_ALU_operand_a[17]) );
  OAI22D1BWP12T U4924 ( .A1(n5524), .A2(n5910), .B1(n5539), .B2(n5857), .ZN(
        n5535) );
  OAI22D1BWP12T U4925 ( .A1(n5526), .A2(n5959), .B1(n5525), .B2(n5912), .ZN(
        n5534) );
  AOI22D1BWP12T U4926 ( .A1(register_file_inst1_tmp1_16_), .A2(n5962), .B1(
        register_file_inst1_r4_16_), .B2(n5961), .ZN(n5528) );
  AOI22D1BWP12T U4927 ( .A1(RF_next_sp[16]), .A2(n5964), .B1(
        register_file_inst1_r12_16_), .B2(n5963), .ZN(n5527) );
  ND3D1BWP12T U4928 ( .A1(n5528), .A2(n5527), .A3(n6114), .ZN(n5533) );
  AOI22D1BWP12T U4929 ( .A1(register_file_inst1_r9_16_), .A2(n5968), .B1(
        register_file_inst1_r3_16_), .B2(n5967), .ZN(n5531) );
  AOI22D1BWP12T U4930 ( .A1(register_file_inst1_r7_16_), .A2(n6001), .B1(
        register_file_inst1_r11_16_), .B2(n5969), .ZN(n5530) );
  AOI22D1BWP12T U4931 ( .A1(register_file_inst1_r5_16_), .A2(n6002), .B1(
        register_file_inst1_lr_16_), .B2(n5970), .ZN(n5529) );
  ND4D1BWP12T U4932 ( .A1(n5531), .A2(n5530), .A3(n6115), .A4(n5529), .ZN(
        n5532) );
  OR4XD1BWP12T U4933 ( .A1(n5535), .A2(n5534), .A3(n5533), .A4(n5532), .Z(
        RF_ALU_operand_b[16]) );
  OAI22D1BWP12T U4934 ( .A1(n5537), .A2(n5938), .B1(n5536), .B2(n6222), .ZN(
        n5548) );
  OAI22D1BWP12T U4935 ( .A1(n5539), .A2(n5942), .B1(n5538), .B2(n5940), .ZN(
        n5547) );
  AOI22D1BWP12T U4936 ( .A1(register_file_inst1_tmp1_16_), .A2(n5979), .B1(
        register_file_inst1_r10_16_), .B2(n6223), .ZN(n5541) );
  AOI22D1BWP12T U4937 ( .A1(register_file_inst1_r4_16_), .A2(n5900), .B1(
        register_file_inst1_r9_16_), .B2(n5943), .ZN(n5540) );
  ND3D1BWP12T U4938 ( .A1(n5541), .A2(n5540), .A3(n6192), .ZN(n5546) );
  AOI22D1BWP12T U4939 ( .A1(register_file_inst1_r0_16_), .A2(n6004), .B1(
        register_file_inst1_r6_16_), .B2(n6003), .ZN(n5544) );
  AOI22D1BWP12T U4940 ( .A1(register_file_inst1_r11_16_), .A2(n6229), .B1(
        register_file_inst1_r3_16_), .B2(n5946), .ZN(n5543) );
  AOI22D1BWP12T U4941 ( .A1(register_file_inst1_r5_16_), .A2(n5948), .B1(
        register_file_inst1_r8_16_), .B2(n6230), .ZN(n5542) );
  ND4D1BWP12T U4942 ( .A1(n5544), .A2(n6193), .A3(n5543), .A4(n5542), .ZN(
        n5545) );
  OAI22D1BWP12T U4943 ( .A1(n5549), .A2(n5910), .B1(n5564), .B2(n5857), .ZN(
        n5560) );
  OAI22D1BWP12T U4944 ( .A1(n5551), .A2(n5959), .B1(n5550), .B2(n5912), .ZN(
        n5559) );
  AOI22D1BWP12T U4945 ( .A1(register_file_inst1_tmp1_15_), .A2(n5962), .B1(
        register_file_inst1_r4_15_), .B2(n5961), .ZN(n5553) );
  AOI22D1BWP12T U4946 ( .A1(RF_next_sp[15]), .A2(n5964), .B1(
        register_file_inst1_r12_15_), .B2(n5963), .ZN(n5552) );
  AOI22D1BWP12T U4947 ( .A1(register_file_inst1_r9_15_), .A2(n5968), .B1(
        register_file_inst1_r3_15_), .B2(n5967), .ZN(n5556) );
  AOI22D1BWP12T U4948 ( .A1(register_file_inst1_r7_15_), .A2(n6001), .B1(
        register_file_inst1_r11_15_), .B2(n5969), .ZN(n5555) );
  AOI22D1BWP12T U4949 ( .A1(register_file_inst1_r5_15_), .A2(n6002), .B1(
        register_file_inst1_lr_15_), .B2(n5970), .ZN(n5554) );
  ND4D1BWP12T U4950 ( .A1(n5556), .A2(n5555), .A3(n6106), .A4(n5554), .ZN(
        n5557) );
  OR4XD1BWP12T U4951 ( .A1(n5560), .A2(n5559), .A3(n5558), .A4(n5557), .Z(
        RF_ALU_operand_b[15]) );
  OAI22D1BWP12T U4952 ( .A1(n5562), .A2(n5938), .B1(n5561), .B2(n6222), .ZN(
        n5573) );
  OAI22D1BWP12T U4953 ( .A1(n5564), .A2(n5942), .B1(n5563), .B2(n5940), .ZN(
        n5572) );
  AOI22D1BWP12T U4954 ( .A1(register_file_inst1_tmp1_15_), .A2(n5979), .B1(
        register_file_inst1_r10_15_), .B2(n6223), .ZN(n5566) );
  AOI22D1BWP12T U4955 ( .A1(register_file_inst1_r4_15_), .A2(n5900), .B1(
        register_file_inst1_r9_15_), .B2(n6225), .ZN(n5565) );
  AOI22D1BWP12T U4956 ( .A1(register_file_inst1_r0_15_), .A2(n6004), .B1(
        register_file_inst1_r6_15_), .B2(n6003), .ZN(n5569) );
  AOI22D1BWP12T U4957 ( .A1(register_file_inst1_r11_15_), .A2(n6229), .B1(
        register_file_inst1_r3_15_), .B2(n5946), .ZN(n5568) );
  AOI22D1BWP12T U4958 ( .A1(register_file_inst1_r5_15_), .A2(n5948), .B1(
        register_file_inst1_r8_15_), .B2(n5947), .ZN(n5567) );
  ND4D1BWP12T U4959 ( .A1(n5569), .A2(n6191), .A3(n5568), .A4(n5567), .ZN(
        n5570) );
  OR4XD1BWP12T U4960 ( .A1(n5573), .A2(n5572), .A3(n5571), .A4(n5570), .Z(
        RF_ALU_operand_a[15]) );
  OAI22D1BWP12T U4961 ( .A1(n5575), .A2(n5938), .B1(n5574), .B2(n6222), .ZN(
        n5586) );
  OAI22D1BWP12T U4962 ( .A1(n5577), .A2(n5942), .B1(n5576), .B2(n5940), .ZN(
        n5585) );
  AOI22D1BWP12T U4963 ( .A1(register_file_inst1_tmp1_14_), .A2(n5979), .B1(
        register_file_inst1_r10_14_), .B2(n6223), .ZN(n5579) );
  AOI22D1BWP12T U4964 ( .A1(register_file_inst1_r4_14_), .A2(n5900), .B1(
        register_file_inst1_r9_14_), .B2(n6225), .ZN(n5578) );
  ND3D1BWP12T U4965 ( .A1(n5579), .A2(n5578), .A3(n6188), .ZN(n5584) );
  AOI22D1BWP12T U4966 ( .A1(register_file_inst1_r0_14_), .A2(n6004), .B1(
        register_file_inst1_r6_14_), .B2(n6003), .ZN(n5582) );
  AOI22D1BWP12T U4967 ( .A1(register_file_inst1_r11_14_), .A2(n6229), .B1(
        register_file_inst1_r3_14_), .B2(n5946), .ZN(n5581) );
  AOI22D1BWP12T U4968 ( .A1(register_file_inst1_r5_14_), .A2(n5948), .B1(
        register_file_inst1_r8_14_), .B2(n6230), .ZN(n5580) );
  ND4D1BWP12T U4969 ( .A1(n5582), .A2(n6189), .A3(n5581), .A4(n5580), .ZN(
        n5583) );
  OR4XD1BWP12T U4970 ( .A1(n5586), .A2(n5585), .A3(n5584), .A4(n5583), .Z(
        RF_ALU_operand_a[14]) );
  OAI22D1BWP12T U4971 ( .A1(n5588), .A2(n5938), .B1(n5587), .B2(n6222), .ZN(
        n5599) );
  OAI22D1BWP12T U4972 ( .A1(n5590), .A2(n5942), .B1(n5589), .B2(n5940), .ZN(
        n5598) );
  AOI22D1BWP12T U4973 ( .A1(register_file_inst1_tmp1_13_), .A2(n5979), .B1(
        register_file_inst1_r10_13_), .B2(n6223), .ZN(n5592) );
  AOI22D1BWP12T U4974 ( .A1(register_file_inst1_r4_13_), .A2(n5900), .B1(
        register_file_inst1_r9_13_), .B2(n5943), .ZN(n5591) );
  ND3D1BWP12T U4975 ( .A1(n5592), .A2(n5591), .A3(n6186), .ZN(n5597) );
  AOI22D1BWP12T U4976 ( .A1(register_file_inst1_r0_13_), .A2(n6004), .B1(
        register_file_inst1_r6_13_), .B2(n6003), .ZN(n5595) );
  AOI22D1BWP12T U4977 ( .A1(register_file_inst1_r11_13_), .A2(n6229), .B1(
        register_file_inst1_r3_13_), .B2(n5946), .ZN(n5594) );
  ND4D1BWP12T U4978 ( .A1(n5595), .A2(n6187), .A3(n5594), .A4(n5593), .ZN(
        n5596) );
  OR4XD1BWP12T U4979 ( .A1(n5599), .A2(n5598), .A3(n5597), .A4(n5596), .Z(
        RF_ALU_operand_a[13]) );
  AOI22D1BWP12T U4980 ( .A1(register_file_inst1_r6_12_), .A2(n6003), .B1(
        register_file_inst1_r0_12_), .B2(n6004), .ZN(n5602) );
  AOI22D1BWP12T U4981 ( .A1(register_file_inst1_r3_12_), .A2(n5946), .B1(
        register_file_inst1_r11_12_), .B2(n6229), .ZN(n5601) );
  AOI22D1BWP12T U4982 ( .A1(register_file_inst1_r5_12_), .A2(n5948), .B1(
        register_file_inst1_r8_12_), .B2(n5947), .ZN(n5600) );
  AN4XD1BWP12T U4983 ( .A1(n5602), .A2(n6184), .A3(n5601), .A4(n5600), .Z(
        n5608) );
  AOI22D1BWP12T U4984 ( .A1(register_file_inst1_tmp1_12_), .A2(n5979), .B1(
        register_file_inst1_r10_12_), .B2(n6223), .ZN(n5604) );
  AOI22D1BWP12T U4985 ( .A1(register_file_inst1_r9_12_), .A2(n5943), .B1(
        register_file_inst1_r4_12_), .B2(n5900), .ZN(n5603) );
  AN3XD1BWP12T U4986 ( .A1(n5604), .A2(n5603), .A3(n6185), .Z(n5607) );
  AOI22D1BWP12T U4987 ( .A1(RF_next_sp[12]), .A2(n5835), .B1(
        register_file_inst1_r7_12_), .B2(n5848), .ZN(n5606) );
  AOI22D1BWP12T U4988 ( .A1(register_file_inst1_lr_12_), .A2(n5836), .B1(
        register_file_inst1_r1_12_), .B2(n5837), .ZN(n5605) );
  ND4D1BWP12T U4989 ( .A1(n5608), .A2(n5607), .A3(n5606), .A4(n5605), .ZN(
        RF_ALU_operand_a[12]) );
  OAI22D1BWP12T U4990 ( .A1(n5610), .A2(n5910), .B1(n5609), .B2(n5857), .ZN(
        n5621) );
  OAI22D1BWP12T U4991 ( .A1(n5612), .A2(n5959), .B1(n5611), .B2(n5912), .ZN(
        n5620) );
  AOI22D1BWP12T U4992 ( .A1(register_file_inst1_tmp1_12_), .A2(n5962), .B1(
        register_file_inst1_r4_12_), .B2(n5961), .ZN(n5614) );
  AOI22D1BWP12T U4993 ( .A1(RF_next_sp[12]), .A2(n5964), .B1(
        register_file_inst1_r12_12_), .B2(n5963), .ZN(n5613) );
  TPND3D0BWP12T U4994 ( .A1(n5614), .A2(n5613), .A3(n6099), .ZN(n5619) );
  AOI22D1BWP12T U4995 ( .A1(register_file_inst1_r9_12_), .A2(n5968), .B1(
        register_file_inst1_r3_12_), .B2(n5967), .ZN(n5617) );
  AOI22D1BWP12T U4996 ( .A1(register_file_inst1_r7_12_), .A2(n6001), .B1(
        register_file_inst1_r11_12_), .B2(n5969), .ZN(n5616) );
  AOI22D1BWP12T U4997 ( .A1(register_file_inst1_r5_12_), .A2(n6002), .B1(
        register_file_inst1_lr_12_), .B2(n5970), .ZN(n5615) );
  ND4D1BWP12T U4998 ( .A1(n5617), .A2(n5616), .A3(n6100), .A4(n5615), .ZN(
        n5618) );
  OR4XD1BWP12T U4999 ( .A1(n5621), .A2(n5620), .A3(n5619), .A4(n5618), .Z(
        RF_ALU_operand_b[12]) );
  AOI22D1BWP12T U5000 ( .A1(register_file_inst1_r6_11_), .A2(n6003), .B1(
        register_file_inst1_r0_11_), .B2(n6004), .ZN(n5624) );
  AOI22D1BWP12T U5001 ( .A1(register_file_inst1_r3_11_), .A2(n5946), .B1(
        register_file_inst1_r11_11_), .B2(n6229), .ZN(n5623) );
  AOI22D1BWP12T U5002 ( .A1(register_file_inst1_r5_11_), .A2(n5948), .B1(
        register_file_inst1_r8_11_), .B2(n5947), .ZN(n5622) );
  AN4XD1BWP12T U5003 ( .A1(n5624), .A2(n6182), .A3(n5623), .A4(n5622), .Z(
        n5630) );
  AOI22D1BWP12T U5004 ( .A1(register_file_inst1_tmp1_11_), .A2(n5979), .B1(
        register_file_inst1_r10_11_), .B2(n6223), .ZN(n5626) );
  AOI22D1BWP12T U5005 ( .A1(register_file_inst1_r9_11_), .A2(n5943), .B1(
        register_file_inst1_r4_11_), .B2(n5900), .ZN(n5625) );
  AN3XD1BWP12T U5006 ( .A1(n5626), .A2(n5625), .A3(n6183), .Z(n5629) );
  AOI22D1BWP12T U5007 ( .A1(RF_next_sp[11]), .A2(n5835), .B1(
        register_file_inst1_r7_11_), .B2(n5848), .ZN(n5628) );
  AOI22D1BWP12T U5008 ( .A1(register_file_inst1_lr_11_), .A2(n5836), .B1(
        register_file_inst1_r1_11_), .B2(n5837), .ZN(n5627) );
  ND4D1BWP12T U5009 ( .A1(n5630), .A2(n5629), .A3(n5628), .A4(n5627), .ZN(
        RF_ALU_operand_a[11]) );
  OAI22D1BWP12T U5010 ( .A1(n5632), .A2(n5910), .B1(n5631), .B2(n5857), .ZN(
        n5643) );
  OAI22D1BWP12T U5011 ( .A1(n5634), .A2(n5959), .B1(n5633), .B2(n5912), .ZN(
        n5642) );
  AOI22D1BWP12T U5012 ( .A1(register_file_inst1_tmp1_11_), .A2(n5962), .B1(
        register_file_inst1_r4_11_), .B2(n5961), .ZN(n5636) );
  AOI22D1BWP12T U5013 ( .A1(RF_next_sp[11]), .A2(n5964), .B1(
        register_file_inst1_r12_11_), .B2(n5963), .ZN(n5635) );
  ND3D1BWP12T U5014 ( .A1(n5636), .A2(n5635), .A3(n6094), .ZN(n5641) );
  AOI22D1BWP12T U5015 ( .A1(register_file_inst1_r9_11_), .A2(n5968), .B1(
        register_file_inst1_r3_11_), .B2(n5967), .ZN(n5639) );
  AOI22D1BWP12T U5016 ( .A1(register_file_inst1_r7_11_), .A2(n6001), .B1(
        register_file_inst1_r11_11_), .B2(n5969), .ZN(n5638) );
  AOI22D1BWP12T U5017 ( .A1(register_file_inst1_r5_11_), .A2(n6002), .B1(
        register_file_inst1_lr_11_), .B2(n5970), .ZN(n5637) );
  ND4D1BWP12T U5018 ( .A1(n5639), .A2(n5638), .A3(n6095), .A4(n5637), .ZN(
        n5640) );
  OR4XD1BWP12T U5019 ( .A1(n5643), .A2(n5642), .A3(n5641), .A4(n5640), .Z(
        RF_ALU_operand_b[11]) );
  AOI22D1BWP12T U5020 ( .A1(register_file_inst1_r4_9_), .A2(n5900), .B1(
        register_file_inst1_r9_9_), .B2(n5943), .ZN(n5646) );
  AOI22D1BWP12T U5021 ( .A1(register_file_inst1_r12_9_), .A2(n6228), .B1(
        register_file_inst1_r3_9_), .B2(n5946), .ZN(n5645) );
  AOI22D1BWP12T U5022 ( .A1(register_file_inst1_r5_9_), .A2(n5948), .B1(
        register_file_inst1_r11_9_), .B2(n6229), .ZN(n5644) );
  AN4XD1BWP12T U5023 ( .A1(n5646), .A2(n6178), .A3(n5645), .A4(n5644), .Z(
        n5652) );
  AOI22D1BWP12T U5024 ( .A1(register_file_inst1_tmp1_9_), .A2(n5979), .B1(
        register_file_inst1_r10_9_), .B2(n6223), .ZN(n5648) );
  AOI22D1BWP12T U5025 ( .A1(register_file_inst1_r2_9_), .A2(n5998), .B1(
        register_file_inst1_r7_9_), .B2(n5848), .ZN(n5647) );
  AN3XD1BWP12T U5026 ( .A1(n5648), .A2(n6179), .A3(n5647), .Z(n5651) );
  AOI22D1BWP12T U5027 ( .A1(register_file_inst1_r8_9_), .A2(n5947), .B1(
        RF_next_sp[9]), .B2(n5835), .ZN(n5650) );
  AOI22D1BWP12T U5028 ( .A1(register_file_inst1_r1_9_), .A2(n5837), .B1(
        register_file_inst1_lr_9_), .B2(n5836), .ZN(n5649) );
  ND4D1BWP12T U5029 ( .A1(n5652), .A2(n5651), .A3(n5650), .A4(n5649), .ZN(
        RF_ALU_operand_a[9]) );
  OAI22D1BWP12T U5030 ( .A1(n5655), .A2(n5857), .B1(n5654), .B2(n5653), .ZN(
        n5666) );
  OAI22D1BWP12T U5031 ( .A1(n5657), .A2(n5959), .B1(n5656), .B2(n5912), .ZN(
        n5665) );
  AOI22D1BWP12T U5032 ( .A1(register_file_inst1_tmp1_9_), .A2(n5962), .B1(
        register_file_inst1_r4_9_), .B2(n5961), .ZN(n5659) );
  AOI22D1BWP12T U5033 ( .A1(register_file_inst1_r8_9_), .A2(n5994), .B1(
        register_file_inst1_r6_9_), .B2(n5823), .ZN(n5658) );
  ND3D1BWP12T U5034 ( .A1(n5659), .A2(n6087), .A3(n5658), .ZN(n5664) );
  AOI22D1BWP12T U5035 ( .A1(register_file_inst1_r12_9_), .A2(n5963), .B1(
        RF_next_sp[9]), .B2(n5964), .ZN(n5662) );
  AOI22D1BWP12T U5036 ( .A1(register_file_inst1_r9_9_), .A2(n5968), .B1(
        register_file_inst1_r3_9_), .B2(n5967), .ZN(n5661) );
  AOI22D1BWP12T U5037 ( .A1(register_file_inst1_r10_9_), .A2(n5995), .B1(
        register_file_inst1_r11_9_), .B2(n5969), .ZN(n5660) );
  ND4D1BWP12T U5038 ( .A1(n5662), .A2(n5661), .A3(n5660), .A4(n6088), .ZN(
        n5663) );
  OAI22D1BWP12T U5039 ( .A1(n5667), .A2(n5910), .B1(n5682), .B2(n5857), .ZN(
        n5678) );
  OAI22D1BWP12T U5040 ( .A1(n5669), .A2(n5959), .B1(n5668), .B2(n5912), .ZN(
        n5677) );
  AOI22D1BWP12T U5041 ( .A1(register_file_inst1_tmp1_8_), .A2(n5962), .B1(
        register_file_inst1_r4_8_), .B2(n5961), .ZN(n5671) );
  AOI22D1BWP12T U5042 ( .A1(register_file_inst1_r12_8_), .A2(n5963), .B1(
        RF_next_sp[8]), .B2(n5964), .ZN(n5670) );
  ND3D1BWP12T U5043 ( .A1(n5671), .A2(n5670), .A3(n6084), .ZN(n5676) );
  AOI22D1BWP12T U5044 ( .A1(register_file_inst1_r9_8_), .A2(n5968), .B1(
        register_file_inst1_r3_8_), .B2(n5967), .ZN(n5674) );
  AOI22D1BWP12T U5045 ( .A1(register_file_inst1_r7_8_), .A2(n6001), .B1(
        register_file_inst1_r11_8_), .B2(n5969), .ZN(n5673) );
  AOI22D1BWP12T U5046 ( .A1(register_file_inst1_r5_8_), .A2(n6002), .B1(
        register_file_inst1_lr_8_), .B2(n5970), .ZN(n5672) );
  ND4D1BWP12T U5047 ( .A1(n5674), .A2(n5673), .A3(n6085), .A4(n5672), .ZN(
        n5675) );
  OR4XD1BWP12T U5048 ( .A1(n5678), .A2(n5677), .A3(n5676), .A4(n5675), .Z(
        RF_ALU_operand_b[8]) );
  INVD1BWP12T U5049 ( .I(RF_next_sp[8]), .ZN(n5679) );
  OAI22D1BWP12T U5050 ( .A1(n5680), .A2(n5938), .B1(n5679), .B2(n6222), .ZN(
        n5691) );
  OAI22D1BWP12T U5051 ( .A1(n5682), .A2(n5942), .B1(n5681), .B2(n5940), .ZN(
        n5690) );
  AOI22D1BWP12T U5052 ( .A1(register_file_inst1_tmp1_8_), .A2(n5979), .B1(
        register_file_inst1_r10_8_), .B2(n6223), .ZN(n5684) );
  AOI22D1BWP12T U5053 ( .A1(register_file_inst1_r4_8_), .A2(n5900), .B1(
        register_file_inst1_r9_8_), .B2(n6225), .ZN(n5683) );
  ND3D1BWP12T U5054 ( .A1(n5684), .A2(n5683), .A3(n6176), .ZN(n5689) );
  AOI22D1BWP12T U5055 ( .A1(register_file_inst1_r0_8_), .A2(n6004), .B1(
        register_file_inst1_r6_8_), .B2(n6003), .ZN(n5687) );
  AOI22D1BWP12T U5056 ( .A1(register_file_inst1_r11_8_), .A2(n6229), .B1(
        register_file_inst1_r3_8_), .B2(n5946), .ZN(n5686) );
  AOI22D1BWP12T U5057 ( .A1(register_file_inst1_r5_8_), .A2(n5948), .B1(
        register_file_inst1_r8_8_), .B2(n5947), .ZN(n5685) );
  ND4D1BWP12T U5058 ( .A1(n5687), .A2(n6177), .A3(n5686), .A4(n5685), .ZN(
        n5688) );
  OR4XD1BWP12T U5059 ( .A1(n5691), .A2(n5690), .A3(n5689), .A4(n5688), .Z(
        RF_ALU_operand_a[8]) );
  INVD1BWP12T U5060 ( .I(RF_next_sp[7]), .ZN(n5692) );
  OAI22D1BWP12T U5061 ( .A1(n5693), .A2(n5938), .B1(n5692), .B2(n6222), .ZN(
        n5703) );
  OAI22D1BWP12T U5062 ( .A1(n5704), .A2(n5942), .B1(n5694), .B2(n5940), .ZN(
        n5702) );
  AOI22D1BWP12T U5063 ( .A1(register_file_inst1_tmp1_7_), .A2(n5979), .B1(
        register_file_inst1_r10_7_), .B2(n6223), .ZN(n5696) );
  AOI22D1BWP12T U5064 ( .A1(register_file_inst1_r4_7_), .A2(n5900), .B1(
        register_file_inst1_r9_7_), .B2(n6225), .ZN(n5695) );
  ND3D1BWP12T U5065 ( .A1(n5696), .A2(n5695), .A3(n6174), .ZN(n5701) );
  AOI22D1BWP12T U5066 ( .A1(register_file_inst1_r0_7_), .A2(n6004), .B1(
        register_file_inst1_r6_7_), .B2(n6003), .ZN(n5699) );
  AOI22D1BWP12T U5067 ( .A1(register_file_inst1_r11_7_), .A2(n6229), .B1(
        register_file_inst1_r3_7_), .B2(n5946), .ZN(n5698) );
  AOI22D1BWP12T U5068 ( .A1(register_file_inst1_r5_7_), .A2(n5948), .B1(
        register_file_inst1_r8_7_), .B2(n5947), .ZN(n5697) );
  ND4D1BWP12T U5069 ( .A1(n5699), .A2(n6175), .A3(n5698), .A4(n5697), .ZN(
        n5700) );
  OR4XD1BWP12T U5070 ( .A1(n5703), .A2(n5702), .A3(n5701), .A4(n5700), .Z(
        RF_ALU_operand_a[7]) );
  OAI22D1BWP12T U5071 ( .A1(n5705), .A2(n5910), .B1(n5704), .B2(n5857), .ZN(
        n5716) );
  OAI22D1BWP12T U5072 ( .A1(n5707), .A2(n5959), .B1(n5706), .B2(n5912), .ZN(
        n5715) );
  AOI22D1BWP12T U5073 ( .A1(register_file_inst1_tmp1_7_), .A2(n5962), .B1(
        register_file_inst1_r4_7_), .B2(n5961), .ZN(n5709) );
  AOI22D1BWP12T U5074 ( .A1(register_file_inst1_r12_7_), .A2(n5963), .B1(
        RF_next_sp[7]), .B2(n5964), .ZN(n5708) );
  ND3D1BWP12T U5075 ( .A1(n5709), .A2(n5708), .A3(n6080), .ZN(n5714) );
  AOI22D1BWP12T U5076 ( .A1(register_file_inst1_r9_7_), .A2(n5968), .B1(
        register_file_inst1_r3_7_), .B2(n5967), .ZN(n5712) );
  AOI22D1BWP12T U5077 ( .A1(register_file_inst1_r7_7_), .A2(n6001), .B1(
        register_file_inst1_r11_7_), .B2(n5969), .ZN(n5711) );
  AOI22D1BWP12T U5078 ( .A1(register_file_inst1_r5_7_), .A2(n6002), .B1(
        register_file_inst1_lr_7_), .B2(n5970), .ZN(n5710) );
  ND4D1BWP12T U5079 ( .A1(n5712), .A2(n5711), .A3(n6081), .A4(n5710), .ZN(
        n5713) );
  OR4XD1BWP12T U5080 ( .A1(n5716), .A2(n5715), .A3(n5714), .A4(n5713), .Z(
        RF_ALU_operand_b[7]) );
  OAI22D1BWP12T U5081 ( .A1(n5718), .A2(n5910), .B1(n5717), .B2(n5857), .ZN(
        n5729) );
  OAI22D1BWP12T U5082 ( .A1(n5720), .A2(n5959), .B1(n5719), .B2(n5912), .ZN(
        n5728) );
  AOI22D1BWP12T U5083 ( .A1(register_file_inst1_tmp1_6_), .A2(n5962), .B1(
        register_file_inst1_r4_6_), .B2(n5961), .ZN(n5722) );
  AOI22D1BWP12T U5084 ( .A1(register_file_inst1_r12_6_), .A2(n5963), .B1(
        RF_next_sp[6]), .B2(n5964), .ZN(n5721) );
  ND3D1BWP12T U5085 ( .A1(n5722), .A2(n5721), .A3(n6076), .ZN(n5727) );
  AOI22D1BWP12T U5086 ( .A1(register_file_inst1_r9_6_), .A2(n5968), .B1(
        register_file_inst1_r3_6_), .B2(n5967), .ZN(n5725) );
  AOI22D1BWP12T U5087 ( .A1(register_file_inst1_r7_6_), .A2(n6001), .B1(
        register_file_inst1_r11_6_), .B2(n5969), .ZN(n5724) );
  AOI22D1BWP12T U5088 ( .A1(register_file_inst1_r5_6_), .A2(n6002), .B1(
        register_file_inst1_lr_6_), .B2(n5970), .ZN(n5723) );
  ND4D1BWP12T U5089 ( .A1(n5725), .A2(n5724), .A3(n6077), .A4(n5723), .ZN(
        n5726) );
  OR4XD1BWP12T U5090 ( .A1(n5729), .A2(n5728), .A3(n5727), .A4(n5726), .Z(
        RF_ALU_operand_b[6]) );
  AOI22D1BWP12T U5091 ( .A1(register_file_inst1_r0_6_), .A2(n6004), .B1(
        register_file_inst1_r6_6_), .B2(n6003), .ZN(n5732) );
  AOI22D1BWP12T U5092 ( .A1(register_file_inst1_r11_6_), .A2(n6229), .B1(
        register_file_inst1_r3_6_), .B2(n5946), .ZN(n5731) );
  AOI22D1BWP12T U5093 ( .A1(register_file_inst1_r5_6_), .A2(n5948), .B1(
        register_file_inst1_r8_6_), .B2(n5947), .ZN(n5730) );
  AOI22D1BWP12T U5094 ( .A1(register_file_inst1_tmp1_6_), .A2(n5979), .B1(
        register_file_inst1_r10_6_), .B2(n6223), .ZN(n5734) );
  AOI22D1BWP12T U5095 ( .A1(register_file_inst1_r4_6_), .A2(n5900), .B1(
        register_file_inst1_r9_6_), .B2(n5943), .ZN(n5733) );
  OAI22D1BWP12T U5096 ( .A1(n5736), .A2(n5910), .B1(n5735), .B2(n5857), .ZN(
        n5747) );
  OAI22D1BWP12T U5097 ( .A1(n5738), .A2(n5959), .B1(n5737), .B2(n5912), .ZN(
        n5746) );
  AOI22D1BWP12T U5098 ( .A1(register_file_inst1_tmp1_5_), .A2(n5962), .B1(
        register_file_inst1_r4_5_), .B2(n5961), .ZN(n5740) );
  AOI22D1BWP12T U5099 ( .A1(register_file_inst1_r12_5_), .A2(n5963), .B1(
        RF_next_sp[5]), .B2(n5964), .ZN(n5739) );
  ND3D1BWP12T U5100 ( .A1(n5740), .A2(n5739), .A3(n6072), .ZN(n5745) );
  AOI22D1BWP12T U5101 ( .A1(register_file_inst1_r9_5_), .A2(n5968), .B1(
        register_file_inst1_r3_5_), .B2(n5967), .ZN(n5743) );
  AOI22D1BWP12T U5102 ( .A1(register_file_inst1_r7_5_), .A2(n6001), .B1(
        register_file_inst1_r11_5_), .B2(n5969), .ZN(n5742) );
  AOI22D1BWP12T U5103 ( .A1(register_file_inst1_r5_5_), .A2(n6002), .B1(
        register_file_inst1_lr_5_), .B2(n5970), .ZN(n5741) );
  ND4D1BWP12T U5104 ( .A1(n5743), .A2(n5742), .A3(n6073), .A4(n5741), .ZN(
        n5744) );
  OR4XD1BWP12T U5105 ( .A1(n5747), .A2(n5746), .A3(n5745), .A4(n5744), .Z(
        RF_ALU_operand_b[5]) );
  AOI22D1BWP12T U5106 ( .A1(register_file_inst1_r0_5_), .A2(n6004), .B1(
        register_file_inst1_r6_5_), .B2(n6003), .ZN(n5750) );
  AOI22D1BWP12T U5107 ( .A1(register_file_inst1_r11_5_), .A2(n6229), .B1(
        register_file_inst1_r3_5_), .B2(n5946), .ZN(n5749) );
  AOI22D1BWP12T U5108 ( .A1(register_file_inst1_r5_5_), .A2(n5948), .B1(
        register_file_inst1_r8_5_), .B2(n5947), .ZN(n5748) );
  AN4XD1BWP12T U5109 ( .A1(n5750), .A2(n6170), .A3(n5749), .A4(n5748), .Z(
        n5756) );
  AOI22D1BWP12T U5110 ( .A1(register_file_inst1_tmp1_5_), .A2(n5979), .B1(
        register_file_inst1_r10_5_), .B2(n6223), .ZN(n5752) );
  AOI22D1BWP12T U5111 ( .A1(register_file_inst1_r4_5_), .A2(n5900), .B1(
        register_file_inst1_r9_5_), .B2(n6225), .ZN(n5751) );
  AN3XD1BWP12T U5112 ( .A1(n5752), .A2(n5751), .A3(n6171), .Z(n5755) );
  AOI22D1BWP12T U5113 ( .A1(register_file_inst1_r7_5_), .A2(n5848), .B1(
        RF_next_sp[5]), .B2(n5835), .ZN(n5754) );
  AOI22D1BWP12T U5114 ( .A1(register_file_inst1_r1_5_), .A2(n5837), .B1(
        register_file_inst1_lr_5_), .B2(n5836), .ZN(n5753) );
  ND4D1BWP12T U5115 ( .A1(n5756), .A2(n5755), .A3(n5754), .A4(n5753), .ZN(
        RF_ALU_operand_a[5]) );
  AOI22D1BWP12T U5116 ( .A1(register_file_inst1_r12_4_), .A2(n5963), .B1(
        RF_next_sp[4]), .B2(n5964), .ZN(n5757) );
  CKND2D1BWP12T U5117 ( .A1(n5757), .A2(n6068), .ZN(n5767) );
  OAI22D1BWP12T U5118 ( .A1(n5759), .A2(n5910), .B1(n5758), .B2(n5857), .ZN(
        n5766) );
  OAI22D1BWP12T U5119 ( .A1(n5761), .A2(n5959), .B1(n5760), .B2(n5912), .ZN(
        n5765) );
  OAI22D1BWP12T U5120 ( .A1(n5763), .A2(n5981), .B1(n5762), .B2(n5805), .ZN(
        n5764) );
  NR4D0BWP12T U5121 ( .A1(n5767), .A2(n5766), .A3(n5765), .A4(n5764), .ZN(
        n5772) );
  AOI22D1BWP12T U5122 ( .A1(register_file_inst1_r9_4_), .A2(n5968), .B1(
        register_file_inst1_r3_4_), .B2(n5967), .ZN(n5770) );
  AOI22D1BWP12T U5123 ( .A1(register_file_inst1_r7_4_), .A2(n6001), .B1(
        register_file_inst1_r11_4_), .B2(n5969), .ZN(n5769) );
  AOI22D1BWP12T U5124 ( .A1(register_file_inst1_r5_4_), .A2(n6002), .B1(
        register_file_inst1_lr_4_), .B2(n5970), .ZN(n5768) );
  AN4XD1BWP12T U5125 ( .A1(n5770), .A2(n5769), .A3(n6069), .A4(n5768), .Z(
        n5771) );
  ND2D1BWP12T U5126 ( .A1(n5772), .A2(n5771), .ZN(RF_ALU_operand_b[4]) );
  AOI22D1BWP12T U5127 ( .A1(register_file_inst1_r0_4_), .A2(n6004), .B1(
        register_file_inst1_r6_4_), .B2(n6003), .ZN(n5775) );
  AOI22D1BWP12T U5128 ( .A1(register_file_inst1_r11_4_), .A2(n6229), .B1(
        register_file_inst1_r3_4_), .B2(n5946), .ZN(n5774) );
  AOI22D1BWP12T U5129 ( .A1(register_file_inst1_r5_4_), .A2(n5948), .B1(
        register_file_inst1_r8_4_), .B2(n5947), .ZN(n5773) );
  AN4XD1BWP12T U5130 ( .A1(n5775), .A2(n6168), .A3(n5774), .A4(n5773), .Z(
        n5781) );
  AOI22D1BWP12T U5131 ( .A1(register_file_inst1_tmp1_4_), .A2(n5979), .B1(
        register_file_inst1_r10_4_), .B2(n6223), .ZN(n5777) );
  AOI22D1BWP12T U5132 ( .A1(register_file_inst1_r4_4_), .A2(n5900), .B1(
        register_file_inst1_r9_4_), .B2(n6225), .ZN(n5776) );
  AN3XD1BWP12T U5133 ( .A1(n5777), .A2(n5776), .A3(n6169), .Z(n5780) );
  AOI22D1BWP12T U5134 ( .A1(register_file_inst1_r7_4_), .A2(n5848), .B1(
        RF_next_sp[4]), .B2(n5835), .ZN(n5779) );
  AOI22D1BWP12T U5135 ( .A1(register_file_inst1_r1_4_), .A2(n5837), .B1(
        register_file_inst1_lr_4_), .B2(n5836), .ZN(n5778) );
  ND4D1BWP12T U5136 ( .A1(n5781), .A2(n5780), .A3(n5779), .A4(n5778), .ZN(
        RF_ALU_operand_a[4]) );
  AOI22D1BWP12T U5137 ( .A1(register_file_inst1_r0_3_), .A2(n6004), .B1(
        register_file_inst1_r6_3_), .B2(n6003), .ZN(n5784) );
  AOI22D1BWP12T U5138 ( .A1(register_file_inst1_r11_3_), .A2(n6229), .B1(
        register_file_inst1_r3_3_), .B2(n5946), .ZN(n5783) );
  AN4XD1BWP12T U5139 ( .A1(n5784), .A2(n6166), .A3(n5783), .A4(n5782), .Z(
        n5790) );
  AOI22D1BWP12T U5140 ( .A1(register_file_inst1_tmp1_3_), .A2(n5979), .B1(
        register_file_inst1_r10_3_), .B2(n6223), .ZN(n5786) );
  AN3XD1BWP12T U5141 ( .A1(n5786), .A2(n5785), .A3(n6167), .Z(n5789) );
  AOI22D1BWP12T U5142 ( .A1(register_file_inst1_r7_3_), .A2(n5848), .B1(
        RF_next_sp[3]), .B2(n5835), .ZN(n5788) );
  AOI22D1BWP12T U5143 ( .A1(register_file_inst1_r1_3_), .A2(n5837), .B1(
        register_file_inst1_lr_3_), .B2(n5836), .ZN(n5787) );
  AOI22D1BWP12T U5144 ( .A1(register_file_inst1_r9_3_), .A2(n5968), .B1(
        register_file_inst1_r3_3_), .B2(n5967), .ZN(n5793) );
  AOI22D1BWP12T U5145 ( .A1(register_file_inst1_r7_3_), .A2(n6001), .B1(
        register_file_inst1_r11_3_), .B2(n5969), .ZN(n5792) );
  AOI22D1BWP12T U5146 ( .A1(register_file_inst1_r5_3_), .A2(n6002), .B1(
        register_file_inst1_lr_3_), .B2(n5970), .ZN(n5791) );
  AN4XD1BWP12T U5147 ( .A1(n5793), .A2(n5792), .A3(n6064), .A4(n5791), .Z(
        n5799) );
  AOI22D1BWP12T U5148 ( .A1(register_file_inst1_tmp1_3_), .A2(n5962), .B1(
        register_file_inst1_r4_3_), .B2(n5961), .ZN(n5795) );
  AOI22D1BWP12T U5149 ( .A1(register_file_inst1_r12_3_), .A2(n5963), .B1(
        RF_next_sp[3]), .B2(n5964), .ZN(n5794) );
  AN3XD1BWP12T U5150 ( .A1(n5795), .A2(n5794), .A3(n6065), .Z(n5798) );
  AOI22D1BWP12T U5151 ( .A1(register_file_inst1_r6_3_), .A2(n5823), .B1(
        register_file_inst1_r1_3_), .B2(n5822), .ZN(n5797) );
  AOI22D1BWP12T U5152 ( .A1(register_file_inst1_r2_3_), .A2(n5825), .B1(
        register_file_inst1_r0_3_), .B2(n5824), .ZN(n5796) );
  ND4D1BWP12T U5153 ( .A1(n5799), .A2(n5798), .A3(n5797), .A4(n5796), .ZN(
        RF_ALU_operand_b[3]) );
  AOI22D1BWP12T U5154 ( .A1(register_file_inst1_r12_2_), .A2(n5963), .B1(
        RF_next_sp[2]), .B2(n5964), .ZN(n5800) );
  CKND2D1BWP12T U5155 ( .A1(n5800), .A2(n6059), .ZN(n5811) );
  OAI22D1BWP12T U5156 ( .A1(n5802), .A2(n5910), .B1(n5801), .B2(n5857), .ZN(
        n5810) );
  OAI22D1BWP12T U5157 ( .A1(n5807), .A2(n5981), .B1(n5806), .B2(n5805), .ZN(
        n5808) );
  NR4D0BWP12T U5158 ( .A1(n5811), .A2(n5810), .A3(n5809), .A4(n5808), .ZN(
        n5816) );
  AOI22D1BWP12T U5159 ( .A1(register_file_inst1_r9_2_), .A2(n5968), .B1(
        register_file_inst1_r3_2_), .B2(n5967), .ZN(n5814) );
  AOI22D1BWP12T U5160 ( .A1(register_file_inst1_r7_2_), .A2(n6001), .B1(
        register_file_inst1_r11_2_), .B2(n5969), .ZN(n5813) );
  AOI22D1BWP12T U5161 ( .A1(register_file_inst1_r5_2_), .A2(n6002), .B1(
        register_file_inst1_lr_2_), .B2(n5970), .ZN(n5812) );
  AN4XD1BWP12T U5162 ( .A1(n5814), .A2(n5813), .A3(n6060), .A4(n5812), .Z(
        n5815) );
  ND2D1BWP12T U5163 ( .A1(n5816), .A2(n5815), .ZN(RF_ALU_operand_b[2]) );
  AOI22D1BWP12T U5164 ( .A1(register_file_inst1_r9_1_), .A2(n5968), .B1(
        register_file_inst1_r3_1_), .B2(n5967), .ZN(n5819) );
  AOI22D1BWP12T U5165 ( .A1(register_file_inst1_r7_1_), .A2(n6001), .B1(
        register_file_inst1_r11_1_), .B2(n5969), .ZN(n5818) );
  AOI22D1BWP12T U5166 ( .A1(register_file_inst1_r5_1_), .A2(n6002), .B1(
        register_file_inst1_lr_1_), .B2(n5970), .ZN(n5817) );
  AN4XD1BWP12T U5167 ( .A1(n5819), .A2(n5818), .A3(n6055), .A4(n5817), .Z(
        n5829) );
  AOI22D1BWP12T U5168 ( .A1(register_file_inst1_tmp1_1_), .A2(n5962), .B1(
        register_file_inst1_r4_1_), .B2(n5961), .ZN(n5821) );
  AOI22D1BWP12T U5169 ( .A1(register_file_inst1_r12_1_), .A2(n5963), .B1(
        RF_next_sp[1]), .B2(n5964), .ZN(n5820) );
  AN3XD1BWP12T U5170 ( .A1(n5821), .A2(n5820), .A3(n6056), .Z(n5828) );
  AOI22D1BWP12T U5171 ( .A1(register_file_inst1_r6_1_), .A2(n5823), .B1(
        register_file_inst1_r1_1_), .B2(n5822), .ZN(n5827) );
  AOI22D1BWP12T U5172 ( .A1(register_file_inst1_r2_1_), .A2(n5825), .B1(
        register_file_inst1_r0_1_), .B2(n5824), .ZN(n5826) );
  AOI22D1BWP12T U5173 ( .A1(register_file_inst1_r0_1_), .A2(n6004), .B1(
        register_file_inst1_r6_1_), .B2(n6003), .ZN(n5832) );
  AOI22D1BWP12T U5174 ( .A1(register_file_inst1_r11_1_), .A2(n6229), .B1(
        register_file_inst1_r3_1_), .B2(n5946), .ZN(n5831) );
  AOI22D1BWP12T U5175 ( .A1(register_file_inst1_r5_1_), .A2(n5948), .B1(
        register_file_inst1_r8_1_), .B2(n5947), .ZN(n5830) );
  AN4XD1BWP12T U5176 ( .A1(n5832), .A2(n6162), .A3(n5831), .A4(n5830), .Z(
        n5841) );
  AOI22D1BWP12T U5177 ( .A1(register_file_inst1_tmp1_1_), .A2(n5979), .B1(
        register_file_inst1_r10_1_), .B2(n6223), .ZN(n5834) );
  AOI22D1BWP12T U5178 ( .A1(register_file_inst1_r4_1_), .A2(n5900), .B1(
        register_file_inst1_r9_1_), .B2(n6225), .ZN(n5833) );
  AN3XD1BWP12T U5179 ( .A1(n5834), .A2(n5833), .A3(n6163), .Z(n5840) );
  AOI22D1BWP12T U5180 ( .A1(register_file_inst1_r7_1_), .A2(n5848), .B1(
        RF_next_sp[1]), .B2(n5835), .ZN(n5839) );
  AOI22D1BWP12T U5181 ( .A1(register_file_inst1_r1_1_), .A2(n5837), .B1(
        register_file_inst1_lr_1_), .B2(n5836), .ZN(n5838) );
  OAI22D1BWP12T U5182 ( .A1(n5843), .A2(n5942), .B1(n5842), .B2(n6222), .ZN(
        n5856) );
  OAI22D1BWP12T U5183 ( .A1(n5846), .A2(n5940), .B1(n5845), .B2(n5844), .ZN(
        n5855) );
  AOI22D1BWP12T U5184 ( .A1(register_file_inst1_r4_0_), .A2(n5900), .B1(
        register_file_inst1_r9_0_), .B2(n6225), .ZN(n5847) );
  ND3D1BWP12T U5185 ( .A1(n6153), .A2(n5847), .A3(n6152), .ZN(n5854) );
  AOI22D1BWP12T U5186 ( .A1(register_file_inst1_r0_0_), .A2(n6004), .B1(
        register_file_inst1_r6_0_), .B2(n6003), .ZN(n5852) );
  AOI22D1BWP12T U5187 ( .A1(register_file_inst1_r12_0_), .A2(n6228), .B1(
        register_file_inst1_r3_0_), .B2(n5946), .ZN(n5851) );
  AOI22D1BWP12T U5188 ( .A1(register_file_inst1_r5_0_), .A2(n5948), .B1(
        register_file_inst1_r11_0_), .B2(n6229), .ZN(n5850) );
  AOI22D1BWP12T U5189 ( .A1(register_file_inst1_r7_0_), .A2(n5848), .B1(
        register_file_inst1_r8_0_), .B2(n6230), .ZN(n5849) );
  ND4D1BWP12T U5190 ( .A1(n5852), .A2(n5851), .A3(n5850), .A4(n5849), .ZN(
        n5853) );
  OAI22D1BWP12T U5191 ( .A1(n5859), .A2(n5910), .B1(n5858), .B2(n5857), .ZN(
        n5870) );
  OAI22D1BWP12T U5192 ( .A1(n5861), .A2(n5959), .B1(n5860), .B2(n5912), .ZN(
        n5869) );
  AOI22D1BWP12T U5193 ( .A1(register_file_inst1_tmp1_10_), .A2(n5962), .B1(
        register_file_inst1_r4_10_), .B2(n5961), .ZN(n5863) );
  AOI22D1BWP12T U5194 ( .A1(register_file_inst1_r12_10_), .A2(n5963), .B1(
        RF_next_sp[10]), .B2(n5964), .ZN(n5862) );
  ND3D1BWP12T U5195 ( .A1(n5863), .A2(n5862), .A3(n6090), .ZN(n5868) );
  AOI22D1BWP12T U5196 ( .A1(register_file_inst1_r9_10_), .A2(n5968), .B1(
        register_file_inst1_r3_10_), .B2(n5967), .ZN(n5866) );
  AOI22D1BWP12T U5197 ( .A1(register_file_inst1_r7_10_), .A2(n6001), .B1(
        register_file_inst1_r11_10_), .B2(n5969), .ZN(n5865) );
  AOI22D1BWP12T U5198 ( .A1(register_file_inst1_r5_10_), .A2(n6002), .B1(
        register_file_inst1_lr_10_), .B2(n5970), .ZN(n5864) );
  ND4D1BWP12T U5199 ( .A1(n5866), .A2(n5865), .A3(n6091), .A4(n5864), .ZN(
        n5867) );
  OR4XD1BWP12T U5200 ( .A1(n5870), .A2(n5869), .A3(n5868), .A4(n5867), .Z(
        RF_ALU_operand_b[10]) );
  OAI22D1BWP12T U5201 ( .A1(n5872), .A2(n5938), .B1(n5871), .B2(n6222), .ZN(
        n5883) );
  OAI22D1BWP12T U5202 ( .A1(n5874), .A2(n5942), .B1(n5873), .B2(n5940), .ZN(
        n5882) );
  AOI22D1BWP12T U5203 ( .A1(register_file_inst1_tmp1_21_), .A2(n5979), .B1(
        register_file_inst1_r10_21_), .B2(n6223), .ZN(n5876) );
  AOI22D1BWP12T U5204 ( .A1(register_file_inst1_r4_21_), .A2(n5900), .B1(
        register_file_inst1_r9_21_), .B2(n6225), .ZN(n5875) );
  ND3D1BWP12T U5205 ( .A1(n5876), .A2(n5875), .A3(n6202), .ZN(n5881) );
  AOI22D1BWP12T U5206 ( .A1(register_file_inst1_r0_21_), .A2(n6004), .B1(
        register_file_inst1_r6_21_), .B2(n6003), .ZN(n5879) );
  AOI22D1BWP12T U5207 ( .A1(register_file_inst1_r11_21_), .A2(n6229), .B1(
        register_file_inst1_r3_21_), .B2(n5946), .ZN(n5878) );
  AOI22D1BWP12T U5208 ( .A1(register_file_inst1_r5_21_), .A2(n5948), .B1(
        register_file_inst1_r8_21_), .B2(n5947), .ZN(n5877) );
  ND4D1BWP12T U5209 ( .A1(n5879), .A2(n6203), .A3(n5878), .A4(n5877), .ZN(
        n5880) );
  OR4XD1BWP12T U5210 ( .A1(n5883), .A2(n5882), .A3(n5881), .A4(n5880), .Z(
        RF_ALU_operand_a[21]) );
  OAI22D1BWP12T U5211 ( .A1(n5884), .A2(n5910), .B1(n5899), .B2(n5857), .ZN(
        n5895) );
  OAI22D1BWP12T U5212 ( .A1(n5886), .A2(n5959), .B1(n5885), .B2(n5912), .ZN(
        n5894) );
  AOI22D1BWP12T U5213 ( .A1(register_file_inst1_tmp1_20_), .A2(n5962), .B1(
        register_file_inst1_r4_20_), .B2(n5961), .ZN(n5888) );
  AOI22D1BWP12T U5214 ( .A1(RF_next_sp[20]), .A2(n5964), .B1(
        register_file_inst1_r12_20_), .B2(n5963), .ZN(n5887) );
  ND3D1BWP12T U5215 ( .A1(n5888), .A2(n5887), .A3(n6122), .ZN(n5893) );
  AOI22D1BWP12T U5216 ( .A1(register_file_inst1_r9_20_), .A2(n5968), .B1(
        register_file_inst1_r3_20_), .B2(n5967), .ZN(n5891) );
  AOI22D1BWP12T U5217 ( .A1(register_file_inst1_r7_20_), .A2(n6001), .B1(
        register_file_inst1_r11_20_), .B2(n5969), .ZN(n5890) );
  AOI22D1BWP12T U5218 ( .A1(register_file_inst1_r5_20_), .A2(n6002), .B1(
        register_file_inst1_lr_20_), .B2(n5970), .ZN(n5889) );
  ND4D1BWP12T U5219 ( .A1(n5891), .A2(n5890), .A3(n6123), .A4(n5889), .ZN(
        n5892) );
  OR4XD1BWP12T U5220 ( .A1(n5895), .A2(n5894), .A3(n5893), .A4(n5892), .Z(
        RF_ALU_operand_b[20]) );
  OAI22D1BWP12T U5221 ( .A1(n5897), .A2(n5938), .B1(n5896), .B2(n6222), .ZN(
        n5909) );
  OAI22D1BWP12T U5222 ( .A1(n5899), .A2(n5942), .B1(n5898), .B2(n5940), .ZN(
        n5908) );
  AOI22D1BWP12T U5223 ( .A1(register_file_inst1_tmp1_20_), .A2(n5979), .B1(
        register_file_inst1_r10_20_), .B2(n6223), .ZN(n5902) );
  AOI22D1BWP12T U5224 ( .A1(register_file_inst1_r4_20_), .A2(n5900), .B1(
        register_file_inst1_r9_20_), .B2(n5943), .ZN(n5901) );
  ND3D1BWP12T U5225 ( .A1(n5902), .A2(n5901), .A3(n6200), .ZN(n5907) );
  AOI22D1BWP12T U5226 ( .A1(register_file_inst1_r0_20_), .A2(n6004), .B1(
        register_file_inst1_r6_20_), .B2(n6003), .ZN(n5905) );
  AOI22D1BWP12T U5227 ( .A1(register_file_inst1_r11_20_), .A2(n6229), .B1(
        register_file_inst1_r3_20_), .B2(n5946), .ZN(n5904) );
  AOI22D1BWP12T U5228 ( .A1(register_file_inst1_r5_20_), .A2(n5948), .B1(
        register_file_inst1_r8_20_), .B2(n6230), .ZN(n5903) );
  ND4D1BWP12T U5229 ( .A1(n5905), .A2(n6201), .A3(n5904), .A4(n5903), .ZN(
        n5906) );
  OR4XD1BWP12T U5230 ( .A1(n5909), .A2(n5908), .A3(n5907), .A4(n5906), .Z(
        RF_ALU_operand_a[20]) );
  OAI22D1BWP12T U5231 ( .A1(n5911), .A2(n5910), .B1(n5927), .B2(n5857), .ZN(
        n5923) );
  OAI22D1BWP12T U5232 ( .A1(n5914), .A2(n5959), .B1(n5913), .B2(n5912), .ZN(
        n5922) );
  AOI22D1BWP12T U5233 ( .A1(register_file_inst1_tmp1_25_), .A2(n5962), .B1(
        register_file_inst1_r4_25_), .B2(n5961), .ZN(n5916) );
  AOI22D1BWP12T U5234 ( .A1(RF_next_sp[25]), .A2(n5964), .B1(
        register_file_inst1_r12_25_), .B2(n5963), .ZN(n5915) );
  ND3D1BWP12T U5235 ( .A1(n5916), .A2(n5915), .A3(n6132), .ZN(n5921) );
  AOI22D1BWP12T U5236 ( .A1(register_file_inst1_r9_25_), .A2(n5968), .B1(
        register_file_inst1_r3_25_), .B2(n5967), .ZN(n5919) );
  AOI22D1BWP12T U5237 ( .A1(register_file_inst1_r7_25_), .A2(n6001), .B1(
        register_file_inst1_r11_25_), .B2(n5969), .ZN(n5918) );
  AOI22D1BWP12T U5238 ( .A1(register_file_inst1_r5_25_), .A2(n6002), .B1(
        register_file_inst1_lr_25_), .B2(n5970), .ZN(n5917) );
  ND4D1BWP12T U5239 ( .A1(n5919), .A2(n5918), .A3(n6133), .A4(n5917), .ZN(
        n5920) );
  OR4XD1BWP12T U5240 ( .A1(n5923), .A2(n5922), .A3(n5921), .A4(n5920), .Z(
        RF_ALU_operand_b[25]) );
  OAI22D1BWP12T U5241 ( .A1(n5925), .A2(n5938), .B1(n5924), .B2(n6222), .ZN(
        n5936) );
  OAI22D1BWP12T U5242 ( .A1(n5927), .A2(n5942), .B1(n5926), .B2(n5940), .ZN(
        n5935) );
  AOI22D1BWP12T U5243 ( .A1(register_file_inst1_tmp1_25_), .A2(n5979), .B1(
        register_file_inst1_r10_25_), .B2(n6223), .ZN(n5929) );
  AOI22D1BWP12T U5244 ( .A1(register_file_inst1_r4_25_), .A2(n5900), .B1(
        register_file_inst1_r9_25_), .B2(n5943), .ZN(n5928) );
  ND3D1BWP12T U5245 ( .A1(n5929), .A2(n5928), .A3(n6210), .ZN(n5934) );
  AOI22D1BWP12T U5246 ( .A1(register_file_inst1_r0_25_), .A2(n6004), .B1(
        register_file_inst1_r6_25_), .B2(n6003), .ZN(n5932) );
  AOI22D1BWP12T U5247 ( .A1(register_file_inst1_r11_25_), .A2(n6229), .B1(
        register_file_inst1_r3_25_), .B2(n5946), .ZN(n5931) );
  AOI22D1BWP12T U5248 ( .A1(register_file_inst1_r5_25_), .A2(n5948), .B1(
        register_file_inst1_r8_25_), .B2(n5947), .ZN(n5930) );
  ND4D1BWP12T U5249 ( .A1(n5932), .A2(n6211), .A3(n5931), .A4(n5930), .ZN(
        n5933) );
  OR4XD1BWP12T U5250 ( .A1(n5936), .A2(n5935), .A3(n5934), .A4(n5933), .Z(
        RF_ALU_operand_a[25]) );
  OAI22D1BWP12T U5251 ( .A1(n5939), .A2(n5938), .B1(n5937), .B2(n6222), .ZN(
        n5955) );
  OAI22D1BWP12T U5252 ( .A1(n5956), .A2(n5942), .B1(n5941), .B2(n5940), .ZN(
        n5954) );
  AOI22D1BWP12T U5253 ( .A1(register_file_inst1_tmp1_26_), .A2(n6224), .B1(
        register_file_inst1_r10_26_), .B2(n6223), .ZN(n5945) );
  AOI22D1BWP12T U5254 ( .A1(register_file_inst1_r4_26_), .A2(n5900), .B1(
        register_file_inst1_r9_26_), .B2(n5943), .ZN(n5944) );
  ND3D1BWP12T U5255 ( .A1(n5945), .A2(n5944), .A3(n6212), .ZN(n5953) );
  AOI22D1BWP12T U5256 ( .A1(register_file_inst1_r0_26_), .A2(n6004), .B1(
        register_file_inst1_r6_26_), .B2(n6003), .ZN(n5951) );
  AOI22D1BWP12T U5257 ( .A1(register_file_inst1_r11_26_), .A2(n6229), .B1(
        register_file_inst1_r3_26_), .B2(n5946), .ZN(n5950) );
  AOI22D1BWP12T U5258 ( .A1(register_file_inst1_r5_26_), .A2(n5948), .B1(
        register_file_inst1_r8_26_), .B2(n5947), .ZN(n5949) );
  ND4D1BWP12T U5259 ( .A1(n5951), .A2(n6213), .A3(n5950), .A4(n5949), .ZN(
        n5952) );
  OR4XD1BWP12T U5260 ( .A1(n5955), .A2(n5954), .A3(n5953), .A4(n5952), .Z(
        RF_ALU_operand_a[26]) );
  INVD1BWP12T U5261 ( .I(n6158), .ZN(n6160) );
  OAI22D1BWP12T U5262 ( .A1(n5957), .A2(n5910), .B1(n5956), .B2(n5857), .ZN(
        n5977) );
  OAI22D1BWP12T U5263 ( .A1(n5960), .A2(n5959), .B1(n5958), .B2(n5912), .ZN(
        n5976) );
  AOI22D1BWP12T U5264 ( .A1(register_file_inst1_tmp1_26_), .A2(n5962), .B1(
        register_file_inst1_r4_26_), .B2(n5961), .ZN(n5966) );
  AOI22D1BWP12T U5265 ( .A1(RF_next_sp[26]), .A2(n5964), .B1(
        register_file_inst1_r12_26_), .B2(n5963), .ZN(n5965) );
  ND3D1BWP12T U5266 ( .A1(n5966), .A2(n5965), .A3(n6134), .ZN(n5975) );
  AOI22D1BWP12T U5267 ( .A1(register_file_inst1_r9_26_), .A2(n5968), .B1(
        register_file_inst1_r3_26_), .B2(n5967), .ZN(n5973) );
  AOI22D1BWP12T U5268 ( .A1(register_file_inst1_r7_26_), .A2(n6001), .B1(
        register_file_inst1_r11_26_), .B2(n5969), .ZN(n5972) );
  AOI22D1BWP12T U5269 ( .A1(register_file_inst1_r5_26_), .A2(n6002), .B1(
        register_file_inst1_lr_26_), .B2(n5970), .ZN(n5971) );
  ND4D1BWP12T U5270 ( .A1(n5973), .A2(n5972), .A3(n6135), .A4(n5971), .ZN(
        n5974) );
  OR4XD1BWP12T U5271 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .Z(
        RF_ALU_operand_b[26]) );
  AO222D1BWP12T U5272 ( .A1(n6317), .A2(n6316), .B1(RF_pc_out[27]), .B2(n6007), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[27]), .Z(
        register_file_inst1_n2196) );
  AO222D1BWP12T U5273 ( .A1(n6321), .A2(n6320), .B1(RF_pc_out[25]), .B2(n6394), 
        .C1(IF_RF_incremented_pc_out[25]), .C2(n6393), .Z(
        register_file_inst1_n2194) );
  IND2XD1BWP12T U5274 ( .A1(ALU_OUT_n), .B1(DEC_CPSR_update_flag_n), .ZN(n6387) );
  IND2XD1BWP12T U5275 ( .A1(ALU_OUT_c), .B1(DEC_CPSR_update_flag_c), .ZN(n6388) );
  IND2XD1BWP12T U5276 ( .A1(ALU_OUT_v), .B1(DEC_CPSR_update_flag_v), .ZN(n6392) );
  AOI22D1BWP12T U5277 ( .A1(n6360), .A2(n6395), .B1(n6379), .B2(
        MEMCTRL_RF_IF_data_in[8]), .ZN(n6363) );
  AOI22D1BWP12T U5278 ( .A1(n6372), .A2(n6395), .B1(n6379), .B2(
        MEMCTRL_RF_IF_data_in[4]), .ZN(n6375) );
  AOI22D1BWP12T U5279 ( .A1(n6380), .A2(n6395), .B1(n6379), .B2(
        MEMCTRL_RF_IF_data_in[2]), .ZN(n6383) );
  RCAOI211D0BWP12T U5280 ( .A1(n6097), .A2(RF_next_sp[8]), .B(n6082), .C(reset), .ZN(n6083) );
  RCAOI211D0BWP12T U5281 ( .A1(n6097), .A2(RF_next_sp[11]), .B(n6092), .C(
        reset), .ZN(n6093) );
  RCAOI211D0BWP12T U5282 ( .A1(n6097), .A2(RF_next_sp[12]), .B(n6096), .C(
        reset), .ZN(n6098) );
  CKND2D1BWP12T U5283 ( .A1(n6393), .A2(IF_RF_incremented_pc_out[1]), .ZN(
        n6384) );
  TPAOI21D0BWP12T U5284 ( .A1(RF_next_sp[10]), .A2(n6097), .B(reset), .ZN(
        n6089) );
  RCAOI211D0BWP12T U5285 ( .A1(n6097), .A2(RF_next_sp[7]), .B(n6078), .C(reset), .ZN(n6079) );
  RCAOI211D0BWP12T U5286 ( .A1(n6097), .A2(RF_next_sp[6]), .B(n6074), .C(reset), .ZN(n6075) );
  RCAOI211D0BWP12T U5287 ( .A1(n6097), .A2(RF_next_sp[5]), .B(n6070), .C(reset), .ZN(n6071) );
  RCAOI211D0BWP12T U5288 ( .A1(n6097), .A2(RF_next_sp[4]), .B(n6066), .C(reset), .ZN(n6067) );
  RCAOI211D0BWP12T U5289 ( .A1(n6097), .A2(RF_next_sp[3]), .B(n6061), .C(reset), .ZN(n6062) );
  TPAOI21D0BWP12T U5290 ( .A1(RF_next_sp[9]), .A2(n6097), .B(reset), .ZN(n6086) );
  RCAOI211D0BWP12T U5291 ( .A1(n6097), .A2(RF_next_sp[1]), .B(n6052), .C(reset), .ZN(n6053) );
  RCAOI211D0BWP12T U5292 ( .A1(n6097), .A2(RF_next_sp[2]), .B(n6057), .C(reset), .ZN(n6058) );
  TPNR2D0BWP12T U5293 ( .A1(n6234), .A2(MEMCTRL_read_finished), .ZN(n6398) );
  NR2XD0BWP12T U5294 ( .A1(n6112), .A2(reset), .ZN(
        memory_interface_inst1_fsm_N32) );
  NR2XD0BWP12T U5295 ( .A1(n6107), .A2(reset), .ZN(
        memory_interface_inst1_fsm_N33) );
  TPAOI21D0BWP12T U5296 ( .A1(n6109), .A2(n6108), .B(reset), .ZN(
        memory_interface_inst1_fsm_N34) );
  AN2XD1BWP12T U5297 ( .A1(MEMCTRL_RF_IF_data_in[1]), .A2(n5984), .Z(n5982) );
  AOI22D1BWP12T U5298 ( .A1(RF_pc_out[2]), .A2(n5996), .B1(
        register_file_inst1_r10_2_), .B2(n5995), .ZN(n6060) );
  AOI22D1BWP12T U5299 ( .A1(RF_pc_out[9]), .A2(n5999), .B1(
        register_file_inst1_r0_9_), .B2(n6004), .ZN(n6178) );
  ND4D0BWP12T U5300 ( .A1(n6282), .A2(n2342), .A3(
        DEC_MEMCTRL_memory_store_request), .A4(n2348), .ZN(n6109) );
  AN4D0BWP12T U5301 ( .A1(n6282), .A2(n2342), .A3(
        DEC_MEMCTRL_memory_store_request), .A4(n6110), .Z(n6111) );
  AOI22D1BWP12T U5302 ( .A1(RF_pc_out[18]), .A2(n5999), .B1(
        register_file_inst1_r12_18_), .B2(n6228), .ZN(n6197) );
  AN2XD1BWP12T U5303 ( .A1(DEC_RF_alu_write_to_reg[3]), .A2(n2871), .Z(n6287)
         );
  NR2XD0BWP12T U5304 ( .A1(reset), .A2(n6015), .ZN(n6027) );
  ND3D1BWP12T U5305 ( .A1(DEC_RF_memory_write_to_reg[1]), .A2(n6391), .A3(
        n6021), .ZN(n6025) );
  AN2XD1BWP12T U5306 ( .A1(DEC_RF_alu_write_to_reg[2]), .A2(n2874), .Z(n6034)
         );
  CKND2D1BWP12T U5307 ( .A1(DEC_RF_alu_write_to_reg[3]), .A2(n6405), .ZN(n6019) );
  NR2XD0BWP12T U5308 ( .A1(DEC_RF_operand_a[2]), .A2(n6148), .ZN(n6158) );
  AN2XD1BWP12T U5309 ( .A1(DEC_RF_alu_write_to_reg[2]), .A2(
        DEC_RF_alu_write_to_reg[1]), .Z(n6286) );
  AN2XD1BWP12T U5310 ( .A1(DEC_RF_memory_write_to_reg[1]), .A2(
        DEC_RF_memory_write_to_reg[2]), .Z(n6296) );
  INVD0BWP12T U5311 ( .I(DEC_RF_operand_a[3]), .ZN(n6148) );
  CKND2D1BWP12T U5312 ( .A1(DEC_MEMCTRL_load_store_width[1]), .A2(
        DEC_MEMCTRL_load_store_width[0]), .ZN(n6110) );
  AOI22D1BWP12T U5313 ( .A1(RF_pc_out[14]), .A2(n5996), .B1(
        register_file_inst1_r10_14_), .B2(n5995), .ZN(n6104) );
  AOI22D0BWP12T U5314 ( .A1(RF_pc_out[18]), .A2(n5996), .B1(
        register_file_inst1_r10_18_), .B2(n5995), .ZN(n6119) );
  AOI22D1BWP12T U5315 ( .A1(RF_pc_out[24]), .A2(n5996), .B1(
        register_file_inst1_r10_24_), .B2(n5995), .ZN(n6131) );
  AOI22D1BWP12T U5316 ( .A1(RF_pc_out[22]), .A2(n5996), .B1(
        register_file_inst1_r10_22_), .B2(n5995), .ZN(n6127) );
  AOI22D1BWP12T U5317 ( .A1(RF_pc_out[7]), .A2(n5996), .B1(
        register_file_inst1_r10_7_), .B2(n5995), .ZN(n6081) );
  AOI22D1BWP12T U5318 ( .A1(RF_pc_out[8]), .A2(n5996), .B1(
        register_file_inst1_r10_8_), .B2(n5995), .ZN(n6085) );
  AOI22D1BWP12T U5319 ( .A1(RF_pc_out[10]), .A2(n5996), .B1(
        register_file_inst1_r10_10_), .B2(n5995), .ZN(n6091) );
  AOI22D1BWP12T U5320 ( .A1(RF_pc_out[11]), .A2(n5996), .B1(
        register_file_inst1_r10_11_), .B2(n5995), .ZN(n6095) );
  AOI22D1BWP12T U5321 ( .A1(RF_pc_out[12]), .A2(n5996), .B1(
        register_file_inst1_r10_12_), .B2(n5995), .ZN(n6100) );
  AO222D0BWP12T U5322 ( .A1(n6313), .A2(n6312), .B1(RF_pc_out[29]), .B2(n6394), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[29]), .Z(
        register_file_inst1_n2198) );
  AOI222D0BWP12T U5323 ( .A1(ALU_MISC_OUT_result[5]), .A2(n6376), .B1(n6395), 
        .B2(n6374), .C1(n6379), .C2(MEMCTRL_RF_IF_data_in[5]), .ZN(n6371) );
  OR2XD1BWP12T U5324 ( .A1(DEC_RF_operand_b[0]), .A2(n6039), .Z(n5981) );
  IND4D1BWP12T U5325 ( .A1(n6019), .B1(n6027), .B2(
        DEC_RF_alu_write_to_reg_enable), .B3(DEC_RF_alu_write_to_reg[4]), .ZN(
        n6144) );
  NR2D1BWP12T U5326 ( .A1(DEC_RF_alu_write_to_reg[2]), .A2(n6013), .ZN(n6030)
         );
  INVD1BWP12T U5327 ( .I(DEC_RF_memory_write_to_reg[1]), .ZN(n6014) );
  INVD1BWP12T U5328 ( .I(DEC_RF_memory_write_to_reg[3]), .ZN(n6403) );
  NR2D1BWP12T U5329 ( .A1(DEC_RF_alu_write_to_reg[3]), .A2(n6016), .ZN(n6026)
         );
  INVD1BWP12T U5330 ( .I(DEC_RF_memory_write_to_reg[0]), .ZN(n6404) );
  INVD1BWP12T U5331 ( .I(DEC_RF_memory_write_to_reg[2]), .ZN(n6021) );
  INVD1BWP12T U5332 ( .I(DEC_RF_alu_write_to_reg[0]), .ZN(n6405) );
  INVD1BWP12T U5333 ( .I(DEC_RF_alu_write_to_reg_enable), .ZN(n3519) );
  AOI22D1BWP12T U5334 ( .A1(n6292), .A2(n6397), .B1(IF_memory_load_req), .B2(
        IF_instruction_memory_address[11]), .ZN(n6293) );
  AOI22D1BWP12T U5335 ( .A1(n6289), .A2(n6397), .B1(IF_memory_load_req), .B2(
        IF_instruction_memory_address[10]), .ZN(n6290) );
  NR2D1BWP12T U5336 ( .A1(IF_memory_load_req), .A2(
        DEC_MISC_OUT_memory_address_source_is_reg), .ZN(n6396) );
  AN4XD1BWP12T U5337 ( .A1(n6296), .A2(DEC_RF_memory_write_to_reg[4]), .A3(
        n3521), .A4(DEC_RF_memory_write_to_reg_enable), .Z(n6020) );
  ND2D1BWP12T U5338 ( .A1(DEC_RF_memory_write_to_reg[2]), .A2(n6014), .ZN(
        n6033) );
  IND3D1BWP12T U5339 ( .A1(n2880), .B1(DEC_RF_memory_write_to_reg[3]), .B2(
        n6404), .ZN(n6032) );
  IND3D1BWP12T U5340 ( .A1(DEC_RF_alu_write_to_reg[3]), .B1(n2878), .B2(n6405), 
        .ZN(n6012) );
  OAI21D1BWP12T U5341 ( .A1(n6011), .A2(DEC_ALU_alu_opcode[4]), .B(n6010), 
        .ZN(ALU_IN_c) );
  ND4D1BWP12T U5342 ( .A1(DEC_ALU_alu_opcode[2]), .A2(DEC_ALU_alu_opcode[1]), 
        .A3(DEC_ALU_alu_opcode[4]), .A4(n6009), .ZN(n6010) );
  NR2D1BWP12T U5343 ( .A1(DEC_ALU_alu_opcode[3]), .A2(DEC_ALU_alu_opcode[0]), 
        .ZN(n6009) );
  AOI22D1BWP12T U5344 ( .A1(register_file_inst1_r2_31_), .A2(n5998), .B1(n6226), .B2(DEC_RF_offset_a[31]), .ZN(n6227) );
  AOI22D1BWP12T U5345 ( .A1(register_file_inst1_r8_31_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[31]), .ZN(n6145) );
  AOI22D1BWP12T U5346 ( .A1(register_file_inst1_r8_30_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[30]), .ZN(n6142) );
  AOI22D1BWP12T U5347 ( .A1(register_file_inst1_r2_30_), .A2(n5998), .B1(n5997), .B2(DEC_RF_offset_a[30]), .ZN(n6220) );
  AOI22D1BWP12T U5348 ( .A1(register_file_inst1_r8_29_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[29]), .ZN(n6140) );
  AOI22D1BWP12T U5349 ( .A1(register_file_inst1_r2_29_), .A2(n5998), .B1(n6226), .B2(DEC_RF_offset_a[29]), .ZN(n6218) );
  AOI22D1BWP12T U5350 ( .A1(register_file_inst1_r8_28_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[28]), .ZN(n6138) );
  AOI22D1BWP12T U5351 ( .A1(register_file_inst1_r2_28_), .A2(n5998), .B1(n5997), .B2(DEC_RF_offset_a[28]), .ZN(n6216) );
  AOI22D1BWP12T U5352 ( .A1(register_file_inst1_r8_27_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[27]), .ZN(n6136) );
  AOI22D1BWP12T U5353 ( .A1(register_file_inst1_r2_27_), .A2(n5998), .B1(n6226), .B2(DEC_RF_offset_a[27]), .ZN(n6214) );
  AOI22D1BWP12T U5354 ( .A1(register_file_inst1_r2_24_), .A2(n5998), .B1(n5997), .B2(DEC_RF_offset_a[24]), .ZN(n6208) );
  AOI22D1BWP12T U5355 ( .A1(register_file_inst1_r8_24_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[24]), .ZN(n6130) );
  AOI22D1BWP12T U5356 ( .A1(register_file_inst1_r8_23_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[23]), .ZN(n6128) );
  AOI22D1BWP12T U5357 ( .A1(register_file_inst1_r2_23_), .A2(n5998), .B1(n6226), .B2(DEC_RF_offset_a[23]), .ZN(n6206) );
  AOI22D1BWP12T U5358 ( .A1(register_file_inst1_r8_22_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[22]), .ZN(n6126) );
  AOI22D1BWP12T U5359 ( .A1(register_file_inst1_r2_22_), .A2(n5998), .B1(n5997), .B2(DEC_RF_offset_a[22]), .ZN(n6204) );
  AOI22D1BWP12T U5360 ( .A1(register_file_inst1_r8_19_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[19]), .ZN(n6120) );
  AOI22D1BWP12T U5361 ( .A1(register_file_inst1_r2_19_), .A2(n5998), .B1(n5997), .B2(DEC_RF_offset_a[19]), .ZN(n6198) );
  AOI22D1BWP12T U5362 ( .A1(register_file_inst1_r8_18_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[18]), .ZN(n6118) );
  AOI22D1BWP12T U5363 ( .A1(register_file_inst1_r2_18_), .A2(n5998), .B1(n5997), .B2(DEC_RF_offset_a[18]), .ZN(n6196) );
  AOI22D1BWP12T U5364 ( .A1(register_file_inst1_r8_17_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[17]), .ZN(n6116) );
  AOI22D1BWP12T U5365 ( .A1(register_file_inst1_r2_17_), .A2(n5998), .B1(n6226), .B2(DEC_RF_offset_a[17]), .ZN(n6194) );
  AOI22D1BWP12T U5366 ( .A1(register_file_inst1_r8_16_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[16]), .ZN(n6114) );
  AOI22D1BWP12T U5367 ( .A1(register_file_inst1_r2_16_), .A2(n5998), .B1(n6226), .B2(DEC_RF_offset_a[16]), .ZN(n6192) );
  AOI22D1BWP12T U5368 ( .A1(register_file_inst1_r8_15_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[15]), .ZN(n6105) );
  AOI22D1BWP12T U5369 ( .A1(register_file_inst1_r2_15_), .A2(n5998), .B1(n6226), .B2(DEC_RF_offset_a[15]), .ZN(n6190) );
  AOI22D1BWP12T U5370 ( .A1(register_file_inst1_r8_14_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[14]), .ZN(n6103) );
  AOI22D1BWP12T U5371 ( .A1(register_file_inst1_r2_14_), .A2(n5998), .B1(n6226), .B2(DEC_RF_offset_a[14]), .ZN(n6188) );
  AOI22D1BWP12T U5372 ( .A1(register_file_inst1_r8_13_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[13]), .ZN(n6101) );
  AOI22D1BWP12T U5373 ( .A1(register_file_inst1_r2_13_), .A2(n5998), .B1(n5997), .B2(DEC_RF_offset_a[13]), .ZN(n6186) );
  AOI22D1BWP12T U5374 ( .A1(register_file_inst1_r2_12_), .A2(n5998), .B1(n5997), .B2(DEC_RF_offset_a[12]), .ZN(n6185) );
  AOI22D1BWP12T U5375 ( .A1(register_file_inst1_r8_12_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[12]), .ZN(n6099) );
  AOI22D1BWP12T U5376 ( .A1(register_file_inst1_r2_11_), .A2(n5998), .B1(n6226), .B2(DEC_RF_offset_a[11]), .ZN(n6183) );
  AOI22D1BWP12T U5377 ( .A1(register_file_inst1_r8_11_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[11]), .ZN(n6094) );
  AOI22D1BWP12T U5378 ( .A1(register_file_inst1_r6_9_), .A2(n6003), .B1(n6226), 
        .B2(DEC_RF_offset_a[9]), .ZN(n6179) );
  AOI22D1BWP12T U5379 ( .A1(register_file_inst1_r7_9_), .A2(n6001), .B1(n5993), 
        .B2(DEC_RF_offset_b[9]), .ZN(n6087) );
  AOI22D1BWP12T U5380 ( .A1(register_file_inst1_r8_8_), .A2(n5994), .B1(n5993), 
        .B2(DEC_RF_offset_b[8]), .ZN(n6084) );
  AOI22D1BWP12T U5381 ( .A1(register_file_inst1_r2_8_), .A2(n5998), .B1(n5997), 
        .B2(DEC_RF_offset_a[8]), .ZN(n6176) );
  AOI22D1BWP12T U5382 ( .A1(register_file_inst1_r2_7_), .A2(n5998), .B1(n6226), 
        .B2(DEC_RF_offset_a[7]), .ZN(n6174) );
  AOI22D1BWP12T U5383 ( .A1(register_file_inst1_r8_7_), .A2(n5994), .B1(n5993), 
        .B2(DEC_RF_offset_b[7]), .ZN(n6080) );
  AOI22D1BWP12T U5384 ( .A1(register_file_inst1_r8_6_), .A2(n5994), .B1(n5993), 
        .B2(DEC_RF_offset_b[6]), .ZN(n6076) );
  AOI22D1BWP12T U5385 ( .A1(register_file_inst1_r2_6_), .A2(n5998), .B1(n5997), 
        .B2(DEC_RF_offset_a[6]), .ZN(n6173) );
  AOI22D1BWP12T U5386 ( .A1(register_file_inst1_r8_5_), .A2(n5994), .B1(n5993), 
        .B2(DEC_RF_offset_b[5]), .ZN(n6072) );
  AOI22D1BWP12T U5387 ( .A1(register_file_inst1_r2_5_), .A2(n5998), .B1(n6226), 
        .B2(DEC_RF_offset_a[5]), .ZN(n6171) );
  AOI22D1BWP12T U5388 ( .A1(register_file_inst1_r8_4_), .A2(n5994), .B1(n5993), 
        .B2(DEC_RF_offset_b[4]), .ZN(n6068) );
  AOI22D1BWP12T U5389 ( .A1(register_file_inst1_r2_4_), .A2(n5998), .B1(n5997), 
        .B2(DEC_RF_offset_a[4]), .ZN(n6169) );
  AOI22D1BWP12T U5390 ( .A1(register_file_inst1_r2_3_), .A2(n5998), .B1(n6226), 
        .B2(DEC_RF_offset_a[3]), .ZN(n6167) );
  AOI22D1BWP12T U5391 ( .A1(register_file_inst1_r8_3_), .A2(n5994), .B1(n5993), 
        .B2(DEC_RF_offset_b[3]), .ZN(n6065) );
  AOI22D1BWP12T U5392 ( .A1(register_file_inst1_r8_2_), .A2(n5994), .B1(n5993), 
        .B2(DEC_RF_offset_b[2]), .ZN(n6059) );
  AOI22D1BWP12T U5393 ( .A1(register_file_inst1_r2_2_), .A2(n5998), .B1(n5997), 
        .B2(DEC_RF_offset_a[2]), .ZN(n6165) );
  AOI22D1BWP12T U5394 ( .A1(register_file_inst1_r8_1_), .A2(n5994), .B1(n5993), 
        .B2(DEC_RF_offset_b[1]), .ZN(n6056) );
  AOI22D1BWP12T U5395 ( .A1(register_file_inst1_r2_1_), .A2(n5998), .B1(n6226), 
        .B2(DEC_RF_offset_a[1]), .ZN(n6163) );
  AOI22D1BWP12T U5396 ( .A1(register_file_inst1_r8_0_), .A2(n5994), .B1(n5993), 
        .B2(DEC_RF_offset_b[0]), .ZN(n6037) );
  AOI22D1BWP12T U5397 ( .A1(register_file_inst1_r2_0_), .A2(n5998), .B1(n5997), 
        .B2(DEC_RF_offset_a[0]), .ZN(n6152) );
  AOI22D1BWP12T U5398 ( .A1(register_file_inst1_r8_10_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[10]), .ZN(n6090) );
  AOI22D1BWP12T U5399 ( .A1(register_file_inst1_r2_10_), .A2(n5998), .B1(n5997), .B2(DEC_RF_offset_a[10]), .ZN(n6181) );
  AOI22D1BWP12T U5400 ( .A1(register_file_inst1_r2_21_), .A2(n5998), .B1(n6226), .B2(DEC_RF_offset_a[21]), .ZN(n6202) );
  AOI22D1BWP12T U5401 ( .A1(register_file_inst1_r8_21_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[21]), .ZN(n6124) );
  AOI22D1BWP12T U5402 ( .A1(register_file_inst1_r8_20_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[20]), .ZN(n6122) );
  AOI22D1BWP12T U5403 ( .A1(register_file_inst1_r2_20_), .A2(n5998), .B1(n5997), .B2(DEC_RF_offset_a[20]), .ZN(n6200) );
  AOI22D1BWP12T U5404 ( .A1(register_file_inst1_r8_25_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[25]), .ZN(n6132) );
  AOI22D1BWP12T U5405 ( .A1(register_file_inst1_r2_25_), .A2(n5998), .B1(n6226), .B2(DEC_RF_offset_a[25]), .ZN(n6210) );
  NR3D1BWP12T U5406 ( .A1(DEC_RF_operand_a[1]), .A2(n6161), .A3(n6160), .ZN(
        n6230) );
  AOI22D1BWP12T U5407 ( .A1(register_file_inst1_r2_26_), .A2(n5998), .B1(n5997), .B2(DEC_RF_offset_a[26]), .ZN(n6212) );
  ND2D1BWP12T U5408 ( .A1(DEC_RF_operand_a[1]), .A2(n6150), .ZN(n6156) );
  NR3D1BWP12T U5409 ( .A1(DEC_RF_operand_a[1]), .A2(n6149), .A3(n6160), .ZN(
        n6225) );
  AN3XD1BWP12T U5410 ( .A1(DEC_RF_operand_a[1]), .A2(n2469), .A3(n6158), .Z(
        n6223) );
  ND2D1BWP12T U5411 ( .A1(n6159), .A2(DEC_RF_operand_a[3]), .ZN(n6151) );
  INVD1BWP12T U5412 ( .I(DEC_RF_operand_a[1]), .ZN(n6147) );
  ND3D1BWP12T U5413 ( .A1(n2471), .A2(DEC_RF_operand_a[3]), .A3(n6155), .ZN(
        n6222) );
  NR2D1BWP12T U5414 ( .A1(DEC_RF_operand_a[1]), .A2(n6150), .ZN(n6155) );
  INVD1BWP12T U5415 ( .I(DEC_RF_operand_a[2]), .ZN(n6150) );
  INVD1BWP12T U5416 ( .I(DEC_RF_operand_a[0]), .ZN(n6402) );
  ND2D1BWP12T U5417 ( .A1(n2470), .A2(DEC_RF_operand_a[0]), .ZN(n6157) );
  ND2D1BWP12T U5418 ( .A1(DEC_RF_operand_a[1]), .A2(DEC_RF_operand_a[2]), .ZN(
        n6154) );
  ND2D1BWP12T U5419 ( .A1(n2515), .A2(DEC_RF_operand_b[1]), .ZN(n6049) );
  ND2D1BWP12T U5420 ( .A1(DEC_RF_operand_b[0]), .A2(n2516), .ZN(n6048) );
  AOI22D1BWP12T U5421 ( .A1(register_file_inst1_r8_26_), .A2(n5994), .B1(n5993), .B2(DEC_RF_offset_b[26]), .ZN(n6134) );
  ND2D1BWP12T U5422 ( .A1(n2515), .A2(DEC_RF_operand_b[0]), .ZN(n6038) );
  ND2D1BWP12T U5423 ( .A1(DEC_RF_operand_b[2]), .A2(n6036), .ZN(n6047) );
  INVD1BWP12T U5424 ( .I(DEC_RF_operand_b[1]), .ZN(n6036) );
  ND3D1BWP12T U5425 ( .A1(n6050), .A2(DEC_RF_operand_b[3]), .A3(
        DEC_RF_operand_b[4]), .ZN(n6039) );
  ND2D1BWP12T U5426 ( .A1(DEC_RF_operand_b[1]), .A2(n2516), .ZN(n6045) );
  NR2D1BWP12T U5427 ( .A1(DEC_RF_operand_b[1]), .A2(n6041), .ZN(n6043) );
  ND2D1BWP12T U5428 ( .A1(DEC_RF_operand_b[0]), .A2(n6042), .ZN(n6046) );
  INVD1BWP12T U5429 ( .I(DEC_RF_operand_b[2]), .ZN(n6042) );
  ND2D1BWP12T U5430 ( .A1(DEC_RF_operand_b[1]), .A2(DEC_RF_operand_b[2]), .ZN(
        n6051) );
  AN3XD1BWP12T U5431 ( .A1(DEC_RF_memory_write_to_reg[1]), .A2(n6297), .A3(
        n6021), .Z(n6023) );
  INVD1BWP12T U5432 ( .I(DEC_RF_operand_b[0]), .ZN(n6044) );
  INR3D0BWP12T U5433 ( .A1(DEC_MISC_OUT_memory_address_source_is_reg), .B1(
        IF_memory_load_req), .B2(DEC_RF_memory_store_address_reg[4]), .ZN(
        n6397) );
  INR3D0BWP12T U5434 ( .A1(DEC_RF_operand_a[4]), .B1(n6151), .B2(n6402), .ZN(
        n6226) );
  AOI22D1BWP12T U5435 ( .A1(RF_pc_out[3]), .A2(n5996), .B1(
        register_file_inst1_r10_3_), .B2(n5995), .ZN(n6064) );
  AOI22D0BWP12T U5436 ( .A1(RF_pc_out[0]), .A2(n6000), .B1(
        register_file_inst1_r9_0_), .B2(n6005), .ZN(n6243) );
  AOI22D0BWP12T U5437 ( .A1(RF_pc_out[8]), .A2(n5999), .B1(
        register_file_inst1_r12_8_), .B2(n6228), .ZN(n6177) );
  AOI22D0BWP12T U5438 ( .A1(RF_pc_out[14]), .A2(n5999), .B1(
        register_file_inst1_r12_14_), .B2(n6228), .ZN(n6189) );
  AOI22D0BWP12T U5439 ( .A1(RF_pc_out[16]), .A2(n5999), .B1(
        register_file_inst1_r12_16_), .B2(n6228), .ZN(n6193) );
  AOI22D0BWP12T U5440 ( .A1(RF_pc_out[20]), .A2(n5999), .B1(
        register_file_inst1_r12_20_), .B2(n6228), .ZN(n6201) );
  AOI22D0BWP12T U5441 ( .A1(RF_pc_out[21]), .A2(n5999), .B1(
        register_file_inst1_r12_21_), .B2(n6228), .ZN(n6203) );
  AOI22D0BWP12T U5442 ( .A1(RF_pc_out[22]), .A2(n5999), .B1(
        register_file_inst1_r12_22_), .B2(n6228), .ZN(n6205) );
  AOI22D1BWP12T U5443 ( .A1(RF_pc_out[23]), .A2(n5999), .B1(
        register_file_inst1_r12_23_), .B2(n6228), .ZN(n6207) );
  AOI22D1BWP12T U5444 ( .A1(RF_pc_out[24]), .A2(n5999), .B1(
        register_file_inst1_r12_24_), .B2(n6228), .ZN(n6209) );
  AOI22D1BWP12T U5445 ( .A1(RF_pc_out[25]), .A2(n5999), .B1(
        register_file_inst1_r12_25_), .B2(n6228), .ZN(n6211) );
  AOI22D0BWP12T U5446 ( .A1(RF_pc_out[27]), .A2(n5999), .B1(
        register_file_inst1_r12_27_), .B2(n6228), .ZN(n6215) );
  AOI22D0BWP12T U5447 ( .A1(RF_pc_out[19]), .A2(n6006), .B1(
        register_file_inst1_r12_19_), .B2(n6228), .ZN(n6199) );
  AOI22D0BWP12T U5448 ( .A1(RF_pc_out[26]), .A2(n6006), .B1(
        register_file_inst1_r12_26_), .B2(n6228), .ZN(n6213) );
  AOI22D0BWP12T U5449 ( .A1(RF_pc_out[28]), .A2(n6006), .B1(
        register_file_inst1_r12_28_), .B2(n6228), .ZN(n6217) );
  AOI22D0BWP12T U5450 ( .A1(RF_pc_out[29]), .A2(n6006), .B1(
        register_file_inst1_r12_29_), .B2(n6228), .ZN(n6219) );
  AOI22D0BWP12T U5451 ( .A1(RF_pc_out[30]), .A2(n6006), .B1(
        register_file_inst1_r12_30_), .B2(n6228), .ZN(n6221) );
  AOI22D0BWP12T U5452 ( .A1(RF_pc_out[31]), .A2(n6006), .B1(
        register_file_inst1_r12_31_), .B2(n6228), .ZN(n6231) );
  AOI22D0BWP12T U5453 ( .A1(n5991), .A2(register_file_inst1_r5_4_), .B1(
        RF_pc_out[4]), .B2(n5992), .ZN(n6236) );
  AOI22D0BWP12T U5454 ( .A1(n5991), .A2(register_file_inst1_r5_7_), .B1(
        RF_pc_out[7]), .B2(n5992), .ZN(n6246) );
  AOI22D0BWP12T U5455 ( .A1(n5991), .A2(register_file_inst1_r5_5_), .B1(
        RF_pc_out[5]), .B2(n5992), .ZN(n6251) );
  AOI22D0BWP12T U5456 ( .A1(n5991), .A2(register_file_inst1_r5_8_), .B1(
        RF_pc_out[8]), .B2(n5992), .ZN(n6260) );
  AOI22D0BWP12T U5457 ( .A1(n5991), .A2(register_file_inst1_r5_3_), .B1(
        RF_pc_out[3]), .B2(n5992), .ZN(n6261) );
  AOI22D0BWP12T U5458 ( .A1(n5991), .A2(register_file_inst1_r5_6_), .B1(
        RF_pc_out[6]), .B2(n5992), .ZN(n6264) );
  AOI22D0BWP12T U5459 ( .A1(n5991), .A2(register_file_inst1_r5_2_), .B1(
        RF_pc_out[2]), .B2(n5992), .ZN(n6273) );
  AOI22D0BWP12T U5460 ( .A1(n5991), .A2(register_file_inst1_r5_9_), .B1(
        RF_pc_out[9]), .B2(n5992), .ZN(n6278) );
  AOI22D0BWP12T U5461 ( .A1(RF_pc_out[4]), .A2(n5996), .B1(
        register_file_inst1_r10_4_), .B2(n5995), .ZN(n6069) );
  AOI22D0BWP12T U5462 ( .A1(RF_pc_out[10]), .A2(n5999), .B1(
        register_file_inst1_r12_10_), .B2(n6228), .ZN(n6180) );
  AOI22D0BWP12T U5463 ( .A1(RF_pc_out[12]), .A2(n5999), .B1(
        register_file_inst1_r12_12_), .B2(n6228), .ZN(n6184) );
  AOI22D0BWP12T U5464 ( .A1(RF_pc_out[0]), .A2(n6006), .B1(
        register_file_inst1_tmp1_0_), .B2(n5979), .ZN(n6153) );
  AOI22D0BWP12T U5465 ( .A1(RF_pc_out[9]), .A2(n6000), .B1(
        register_file_inst1_r8_9_), .B2(n5980), .ZN(n6233) );
  AOI22D0BWP12T U5466 ( .A1(RF_pc_out[13]), .A2(n6000), .B1(
        register_file_inst1_r8_13_), .B2(n5980), .ZN(n6238) );
  AOI22D0BWP12T U5467 ( .A1(RF_pc_out[19]), .A2(n6000), .B1(
        register_file_inst1_r8_19_), .B2(n5980), .ZN(n6240) );
  AOI22D0BWP12T U5468 ( .A1(RF_pc_out[16]), .A2(n6000), .B1(
        register_file_inst1_r8_16_), .B2(n5980), .ZN(n6242) );
  AOI22D0BWP12T U5469 ( .A1(RF_pc_out[22]), .A2(n6000), .B1(
        register_file_inst1_r8_22_), .B2(n5980), .ZN(n6244) );
  AOI22D0BWP12T U5470 ( .A1(RF_pc_out[6]), .A2(n6000), .B1(
        register_file_inst1_r8_6_), .B2(n5980), .ZN(n6245) );
  AOI22D0BWP12T U5471 ( .A1(RF_pc_out[17]), .A2(n6000), .B1(
        register_file_inst1_r8_17_), .B2(n5980), .ZN(n6247) );
  AOI22D0BWP12T U5472 ( .A1(RF_pc_out[26]), .A2(n6000), .B1(
        register_file_inst1_r8_26_), .B2(n5980), .ZN(n6249) );
  AOI22D0BWP12T U5473 ( .A1(RF_pc_out[10]), .A2(n6000), .B1(
        register_file_inst1_r8_10_), .B2(n5980), .ZN(n6250) );
  AOI22D0BWP12T U5474 ( .A1(RF_pc_out[14]), .A2(n6000), .B1(
        register_file_inst1_r8_14_), .B2(n5980), .ZN(n6259) );
  AOI22D0BWP12T U5475 ( .A1(RF_pc_out[10]), .A2(n5992), .B1(
        register_file_inst1_r5_10_), .B2(n5991), .ZN(n6239) );
  INVD1BWP12T U5476 ( .I(MEMCTRL_RF_IF_data_in[7]), .ZN(n6364) );
  AOI22D0BWP12T U5477 ( .A1(RF_pc_out[12]), .A2(n6000), .B1(
        register_file_inst1_r8_12_), .B2(n5980), .ZN(n6255) );
  AOI22D0BWP12T U5478 ( .A1(RF_pc_out[21]), .A2(n6000), .B1(
        register_file_inst1_r8_21_), .B2(n5980), .ZN(n6262) );
  AOI22D0BWP12T U5479 ( .A1(RF_pc_out[5]), .A2(n6000), .B1(
        register_file_inst1_r8_5_), .B2(n5980), .ZN(n6263) );
  AOI22D0BWP12T U5480 ( .A1(RF_pc_out[15]), .A2(n6000), .B1(
        register_file_inst1_r8_15_), .B2(n5980), .ZN(n6268) );
  AOI22D0BWP12T U5481 ( .A1(RF_pc_out[20]), .A2(n6000), .B1(
        register_file_inst1_r8_20_), .B2(n5980), .ZN(n6269) );
  AOI22D0BWP12T U5482 ( .A1(RF_pc_out[18]), .A2(n6000), .B1(
        register_file_inst1_r8_18_), .B2(n5980), .ZN(n6271) );
  AOI22D0BWP12T U5483 ( .A1(RF_pc_out[2]), .A2(n6000), .B1(
        register_file_inst1_r8_2_), .B2(n5980), .ZN(n6272) );
  AOI22D0BWP12T U5484 ( .A1(RF_pc_out[8]), .A2(n6000), .B1(
        register_file_inst1_r8_8_), .B2(n5980), .ZN(n6277) );
  AOI22D0BWP12T U5485 ( .A1(RF_pc_out[23]), .A2(n6000), .B1(
        register_file_inst1_r8_23_), .B2(n5980), .ZN(n6279) );
  AOI22D0BWP12T U5486 ( .A1(RF_pc_out[11]), .A2(n6000), .B1(
        register_file_inst1_r8_11_), .B2(n5980), .ZN(n6281) );
  AOI22D0BWP12T U5487 ( .A1(RF_pc_out[25]), .A2(n6000), .B1(
        register_file_inst1_r8_25_), .B2(n5980), .ZN(n6283) );
  AOI22D0BWP12T U5488 ( .A1(RF_pc_out[27]), .A2(n6000), .B1(
        register_file_inst1_r8_27_), .B2(n5980), .ZN(n6284) );
  AOI22D0BWP12T U5489 ( .A1(RF_pc_out[29]), .A2(n6000), .B1(
        register_file_inst1_r8_29_), .B2(n5980), .ZN(n6285) );
  NR2D1BWP12T U5490 ( .A1(MEMCTRL_RF_IF_data_in[12]), .A2(n6008), .ZN(n6309)
         );
  AOI211D1BWP12T U5491 ( .A1(n6000), .A2(RF_pc_out[28]), .B(n6253), .C(n6252), 
        .ZN(n6254) );
  AOI211D1BWP12T U5492 ( .A1(n6000), .A2(RF_pc_out[30]), .B(n6257), .C(n6256), 
        .ZN(n6258) );
  AOI211D1BWP12T U5493 ( .A1(n6000), .A2(RF_pc_out[31]), .B(n6266), .C(n6265), 
        .ZN(n6267) );
  AOI211D1BWP12T U5494 ( .A1(n6000), .A2(RF_pc_out[24]), .B(n6275), .C(n6274), 
        .ZN(n6276) );
  AOI22D0BWP12T U5495 ( .A1(RF_pc_out[3]), .A2(n6000), .B1(
        register_file_inst1_r8_3_), .B2(n5980), .ZN(n6241) );
  AOI22D0BWP12T U5496 ( .A1(RF_pc_out[1]), .A2(n6000), .B1(
        register_file_inst1_r8_1_), .B2(n5980), .ZN(n6248) );
  AOI22D0BWP12T U5497 ( .A1(RF_pc_out[4]), .A2(n6000), .B1(
        register_file_inst1_r8_4_), .B2(n5980), .ZN(n6270) );
  AOI22D0BWP12T U5498 ( .A1(RF_pc_out[7]), .A2(n6000), .B1(
        register_file_inst1_r8_7_), .B2(n5980), .ZN(n6280) );
  AOI22D1BWP12T U5499 ( .A1(RF_pc_out[2]), .A2(n6007), .B1(n6393), .B2(
        IF_RF_incremented_pc_out[2]), .ZN(n6381) );
  AOI22D0BWP12T U5500 ( .A1(RF_pc_out[11]), .A2(n5992), .B1(
        register_file_inst1_r5_11_), .B2(n5991), .ZN(n6288) );
  AOI22D0BWP12T U5501 ( .A1(RF_pc_out[12]), .A2(n5992), .B1(
        register_file_inst1_r5_12_), .B2(n5991), .ZN(n6291) );
  NR2D1BWP12T U5502 ( .A1(MEMCTRL_RF_IF_data_in[6]), .A2(n6008), .ZN(n6305) );
  AOI22D1BWP12T U5503 ( .A1(RF_pc_out[31]), .A2(n6394), .B1(n6393), .B2(
        IF_RF_incremented_pc_out[31]), .ZN(n6310) );
  AOI22D1BWP12T U5504 ( .A1(RF_pc_out[8]), .A2(n6394), .B1(n6393), .B2(
        IF_RF_incremented_pc_out[8]), .ZN(n6361) );
  AOI22D1BWP12T U5505 ( .A1(RF_pc_out[5]), .A2(n6007), .B1(n6393), .B2(
        IF_RF_incremented_pc_out[5]), .ZN(n6370) );
  AOI22D1BWP12T U5506 ( .A1(RF_pc_out[9]), .A2(n6007), .B1(n6393), .B2(
        IF_RF_incremented_pc_out[9]), .ZN(n6358) );
  AOI22D1BWP12T U5507 ( .A1(RF_pc_out[4]), .A2(n6394), .B1(n6393), .B2(
        IF_RF_incremented_pc_out[4]), .ZN(n6373) );
  AOI22D1BWP12T U5508 ( .A1(RF_pc_out[30]), .A2(n6394), .B1(n6393), .B2(
        IF_RF_incremented_pc_out[30]), .ZN(n6311) );
  NR2D1BWP12T U5509 ( .A1(MEMCTRL_RF_IF_data_in[3]), .A2(n6008), .ZN(n6301) );
  NR2D1BWP12T U5510 ( .A1(MEMCTRL_RF_IF_data_in[10]), .A2(n6008), .ZN(n6300)
         );
  NR2D1BWP12T U5511 ( .A1(MEMCTRL_RF_IF_data_in[7]), .A2(n6008), .ZN(n6306) );
  NR2D1BWP12T U5512 ( .A1(MEMCTRL_RF_IF_data_in[14]), .A2(n6008), .ZN(n6299)
         );
  AOI21D1BWP12T U5513 ( .A1(RF_pc_out[1]), .A2(n6007), .B(reset), .ZN(n6385)
         );
  IND2D1BWP12T U5514 ( .A1(MEMCTRL_write_finished), .B1(n6113), .ZN(n6234) );
  AO222D0BWP12T U5515 ( .A1(n6395), .A2(n6382), .B1(n6376), .B2(
        ALU_MISC_OUT_result[3]), .C1(MEMCTRL_RF_IF_data_in[3]), .C2(n6379), 
        .Z(n6377) );
  AO222D1BWP12T U5516 ( .A1(n6325), .A2(n6324), .B1(RF_pc_out[23]), .B2(n6394), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[23]), .Z(
        register_file_inst1_n2192) );
  AO222D1BWP12T U5517 ( .A1(n6329), .A2(n6328), .B1(RF_pc_out[21]), .B2(n6394), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[21]), .Z(
        register_file_inst1_n2190) );
  AO222D1BWP12T U5518 ( .A1(n6333), .A2(n6332), .B1(RF_pc_out[19]), .B2(n6007), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[19]), .Z(
        register_file_inst1_n2188) );
  AO222D0BWP12T U5519 ( .A1(n6335), .A2(n6334), .B1(RF_pc_out[18]), .B2(n6007), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[18]), .Z(
        register_file_inst1_n2187) );
  AO222D1BWP12T U5520 ( .A1(n6337), .A2(n6336), .B1(RF_pc_out[17]), .B2(n6394), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[17]), .Z(
        register_file_inst1_n2186) );
  AO222D1BWP12T U5521 ( .A1(n6342), .A2(n6341), .B1(RF_pc_out[15]), .B2(n6007), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[15]), .Z(
        register_file_inst1_n2184) );
  AO222D1BWP12T U5522 ( .A1(n6348), .A2(n6347), .B1(RF_pc_out[13]), .B2(n6394), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[13]), .Z(
        register_file_inst1_n2182) );
  AO222D1BWP12T U5523 ( .A1(n6354), .A2(n6353), .B1(RF_pc_out[11]), .B2(n6007), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[11]), .Z(
        register_file_inst1_n2180) );
  AO222D0BWP12T U5524 ( .A1(n6357), .A2(n6356), .B1(RF_pc_out[10]), .B2(n6007), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[10]), .Z(
        register_file_inst1_n2179) );
  AO222D0BWP12T U5525 ( .A1(n6369), .A2(n6368), .B1(RF_pc_out[6]), .B2(n6007), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[6]), .Z(
        register_file_inst1_n2175) );
  AOI211D1BWP12T U5526 ( .A1(n6390), .A2(DEC_CPSR_update_flag_z), .B(reset), 
        .C(n6389), .ZN(register_file_inst1_cpsrin[1]) );
  NR2D1BWP12T U5527 ( .A1(RF_OUT_z), .A2(DEC_CPSR_update_flag_z), .ZN(n6389)
         );
  AO222D0BWP12T U5528 ( .A1(n6323), .A2(n6322), .B1(RF_pc_out[24]), .B2(n6007), 
        .C1(IF_RF_incremented_pc_out[24]), .C2(n6393), .Z(
        register_file_inst1_n2193) );
  INVD1BWP12T U5529 ( .I(RF_OUT_c), .ZN(n6011) );
  NR2D1BWP12T U5530 ( .A1(MEMCTRL_write_finished), .A2(n6232), .ZN(n6294) );
  NR3D1BWP12T U5531 ( .A1(reset), .A2(IF_RF_incremented_pc_write_enable), .A3(
        n6298), .ZN(n6394) );
  IND2D1BWP12T U5532 ( .A1(MEMCTRL_write_finished), .B1(n6237), .ZN(n6295) );
  NR2D1BWP12T U5533 ( .A1(reset), .A2(n6386), .ZN(n6395) );
  NR2D1BWP12T U5534 ( .A1(reset), .A2(n5978), .ZN(n6028) );
  INVD1BWP12T U5535 ( .I(MEMCTRL_write_finished), .ZN(n6235) );
  NR2D1BWP12T U5536 ( .A1(reset), .A2(n5986), .ZN(n6035) );
  NR2D1BWP12T U5537 ( .A1(reset), .A2(n5987), .ZN(n6017) );
  NR2D1BWP12T U5538 ( .A1(reset), .A2(n5990), .ZN(n6018) );
  NR2D1BWP12T U5539 ( .A1(reset), .A2(n5988), .ZN(n6031) );
  NR2D1BWP12T U5540 ( .A1(reset), .A2(n5989), .ZN(n6029) );
  AOI21D1BWP12T U5541 ( .A1(n6287), .A2(n6022), .B(reset), .ZN(n6024) );
  INR3D0BWP12T U5542 ( .A1(DEC_RF_operand_a[4]), .B1(DEC_RF_operand_a[0]), 
        .B2(n6151), .ZN(n6224) );
  AO222D0BWP12T U5543 ( .A1(n6351), .A2(n6350), .B1(RF_pc_out[12]), .B2(n6007), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[12]), .Z(
        register_file_inst1_n2181) );
  AO222D0BWP12T U5544 ( .A1(n6378), .A2(n6377), .B1(RF_pc_out[3]), .B2(n6007), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[3]), .Z(
        register_file_inst1_n2172) );
  AO222D0BWP12T U5545 ( .A1(n6339), .A2(n6338), .B1(RF_pc_out[16]), .B2(n6394), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[16]), .Z(
        register_file_inst1_n2185) );
  AO222D0BWP12T U5546 ( .A1(n6331), .A2(n6330), .B1(RF_pc_out[20]), .B2(n6394), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[20]), .Z(
        register_file_inst1_n2189) );
  AO222D0BWP12T U5547 ( .A1(n6345), .A2(n6344), .B1(RF_pc_out[14]), .B2(n6007), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[14]), .Z(
        register_file_inst1_n2183) );
  AO222D0BWP12T U5548 ( .A1(n6366), .A2(n6365), .B1(RF_pc_out[7]), .B2(n6007), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[7]), .Z(
        register_file_inst1_n2176) );
  AO222D0BWP12T U5549 ( .A1(n6327), .A2(n6326), .B1(RF_pc_out[22]), .B2(n6007), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[22]), .Z(
        register_file_inst1_n2191) );
  AO222D0BWP12T U5550 ( .A1(n6319), .A2(n6318), .B1(RF_pc_out[26]), .B2(n6394), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[26]), .Z(
        register_file_inst1_n2195) );
  AO222D0BWP12T U5551 ( .A1(n6315), .A2(n6314), .B1(RF_pc_out[28]), .B2(n6007), 
        .C1(n6393), .C2(IF_RF_incremented_pc_out[28]), .Z(
        register_file_inst1_n2197) );
  OA211D1BWP12T U5552 ( .A1(DEC_CPSR_update_flag_n), .A2(RF_OUT_n), .B(n6387), 
        .C(n6391), .Z(register_file_inst1_cpsrin[3]) );
  OA211D1BWP12T U5553 ( .A1(DEC_CPSR_update_flag_c), .A2(RF_OUT_c), .B(n6388), 
        .C(n6391), .Z(register_file_inst1_cpsrin[2]) );
  OA211D1BWP12T U5554 ( .A1(DEC_CPSR_update_flag_v), .A2(RF_OUT_v), .B(n6392), 
        .C(n6391), .Z(register_file_inst1_cpsrin[0]) );
endmodule

