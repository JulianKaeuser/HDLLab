// AUTHORS: Group 06
// Tuesday 08/01/2017

module stack ();

localparam WIDE = 16;
localparam LARGE = 32;
localparam STACK_SIZE = 32; //words of 32 bit






endmodule
