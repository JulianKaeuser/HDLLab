
module register_file ( readA_sel, readB_sel, readC_sel, readD_sel, write1_sel, 
        write2_sel, write1_en, write2_en, write1_in, write2_in, immediate1_in, 
        immediate2_in, next_pc_in, next_cpsr_in, next_sp_in, next_pc_en, clk, 
        regA_out, regB_out, regC_out, regD_out, pc_out, cpsr_out, sp_out );
  input [4:0] readA_sel;
  input [4:0] readB_sel;
  input [4:0] readC_sel;
  input [4:0] readD_sel;
  input [4:0] write1_sel;
  input [4:0] write2_sel;
  input [31:0] write1_in;
  input [31:0] write2_in;
  input [31:0] immediate1_in;
  input [31:0] immediate2_in;
  input [31:0] next_pc_in;
  input [3:0] next_cpsr_in;
  input [31:0] next_sp_in;
  output [31:0] regA_out;
  output [31:0] regB_out;
  output [31:0] regC_out;
  output [31:0] regD_out;
  output [31:0] pc_out;
  output [3:0] cpsr_out;
  output [31:0] sp_out;
  input write1_en, write2_en, next_pc_en, clk;
  wire   n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888;
  wire   [31:0] r0;
  wire   [31:0] r1;
  wire   [31:0] r2;
  wire   [31:0] r3;
  wire   [31:0] r4;
  wire   [31:0] r5;
  wire   [31:0] r6;
  wire   [31:0] r7;
  wire   [31:0] r8;
  wire   [31:0] r9;
  wire   [31:0] r10;
  wire   [31:0] r11;
  wire   [31:0] r12;
  wire   [31:0] lr;
  wire   [31:0] tmp1;
  wire   [31:0] spin;

  DFQD1BWP12T r0_reg_31_ ( .D(n2680), .CP(clk), .Q(r0[31]) );
  DFQD1BWP12T r0_reg_30_ ( .D(n2679), .CP(clk), .Q(r0[30]) );
  DFQD1BWP12T r0_reg_29_ ( .D(n2678), .CP(clk), .Q(r0[29]) );
  DFQD1BWP12T r0_reg_28_ ( .D(n2677), .CP(clk), .Q(r0[28]) );
  DFQD1BWP12T r0_reg_27_ ( .D(n2676), .CP(clk), .Q(r0[27]) );
  DFQD1BWP12T r0_reg_26_ ( .D(n2675), .CP(clk), .Q(r0[26]) );
  DFQD1BWP12T r0_reg_25_ ( .D(n2674), .CP(clk), .Q(r0[25]) );
  DFQD1BWP12T r0_reg_24_ ( .D(n2673), .CP(clk), .Q(r0[24]) );
  DFQD1BWP12T r0_reg_23_ ( .D(n2672), .CP(clk), .Q(r0[23]) );
  DFQD1BWP12T r0_reg_22_ ( .D(n2671), .CP(clk), .Q(r0[22]) );
  DFQD1BWP12T r0_reg_21_ ( .D(n2670), .CP(clk), .Q(r0[21]) );
  DFQD1BWP12T r0_reg_20_ ( .D(n2669), .CP(clk), .Q(r0[20]) );
  DFQD1BWP12T r0_reg_19_ ( .D(n2668), .CP(clk), .Q(r0[19]) );
  DFQD1BWP12T r0_reg_18_ ( .D(n2667), .CP(clk), .Q(r0[18]) );
  DFQD1BWP12T r0_reg_17_ ( .D(n2666), .CP(clk), .Q(r0[17]) );
  DFQD1BWP12T r0_reg_16_ ( .D(n2665), .CP(clk), .Q(r0[16]) );
  DFQD1BWP12T r0_reg_15_ ( .D(n2664), .CP(clk), .Q(r0[15]) );
  DFQD1BWP12T r0_reg_14_ ( .D(n2663), .CP(clk), .Q(r0[14]) );
  DFQD1BWP12T r0_reg_13_ ( .D(n2662), .CP(clk), .Q(r0[13]) );
  DFQD1BWP12T r0_reg_12_ ( .D(n2661), .CP(clk), .Q(r0[12]) );
  DFQD1BWP12T r0_reg_11_ ( .D(n2660), .CP(clk), .Q(r0[11]) );
  DFQD1BWP12T r0_reg_10_ ( .D(n2659), .CP(clk), .Q(r0[10]) );
  DFQD1BWP12T r0_reg_9_ ( .D(n2658), .CP(clk), .Q(r0[9]) );
  DFQD1BWP12T r0_reg_8_ ( .D(n2657), .CP(clk), .Q(r0[8]) );
  DFQD1BWP12T r0_reg_7_ ( .D(n2656), .CP(clk), .Q(r0[7]) );
  DFQD1BWP12T r0_reg_6_ ( .D(n2655), .CP(clk), .Q(r0[6]) );
  DFQD1BWP12T r0_reg_5_ ( .D(n2654), .CP(clk), .Q(r0[5]) );
  DFQD1BWP12T r0_reg_4_ ( .D(n2653), .CP(clk), .Q(r0[4]) );
  DFQD1BWP12T r0_reg_3_ ( .D(n2652), .CP(clk), .Q(r0[3]) );
  DFQD1BWP12T r0_reg_2_ ( .D(n2651), .CP(clk), .Q(r0[2]) );
  DFQD1BWP12T r0_reg_1_ ( .D(n2650), .CP(clk), .Q(r0[1]) );
  DFQD1BWP12T r0_reg_0_ ( .D(n2649), .CP(clk), .Q(r0[0]) );
  DFQD1BWP12T r1_reg_31_ ( .D(n2648), .CP(clk), .Q(r1[31]) );
  DFQD1BWP12T r1_reg_30_ ( .D(n2647), .CP(clk), .Q(r1[30]) );
  DFQD1BWP12T r1_reg_29_ ( .D(n2646), .CP(clk), .Q(r1[29]) );
  DFQD1BWP12T r1_reg_28_ ( .D(n2645), .CP(clk), .Q(r1[28]) );
  DFQD1BWP12T r1_reg_27_ ( .D(n2644), .CP(clk), .Q(r1[27]) );
  DFQD1BWP12T r1_reg_26_ ( .D(n2643), .CP(clk), .Q(r1[26]) );
  DFQD1BWP12T r1_reg_25_ ( .D(n2642), .CP(clk), .Q(r1[25]) );
  DFQD1BWP12T r1_reg_24_ ( .D(n2641), .CP(clk), .Q(r1[24]) );
  DFQD1BWP12T r1_reg_23_ ( .D(n2640), .CP(clk), .Q(r1[23]) );
  DFQD1BWP12T r1_reg_22_ ( .D(n2639), .CP(clk), .Q(r1[22]) );
  DFQD1BWP12T r1_reg_21_ ( .D(n2638), .CP(clk), .Q(r1[21]) );
  DFQD1BWP12T r1_reg_20_ ( .D(n2637), .CP(clk), .Q(r1[20]) );
  DFQD1BWP12T r1_reg_19_ ( .D(n2636), .CP(clk), .Q(r1[19]) );
  DFQD1BWP12T r1_reg_18_ ( .D(n2635), .CP(clk), .Q(r1[18]) );
  DFQD1BWP12T r1_reg_17_ ( .D(n2634), .CP(clk), .Q(r1[17]) );
  DFQD1BWP12T r1_reg_16_ ( .D(n2633), .CP(clk), .Q(r1[16]) );
  DFQD1BWP12T r1_reg_15_ ( .D(n2632), .CP(clk), .Q(r1[15]) );
  DFQD1BWP12T r1_reg_14_ ( .D(n2631), .CP(clk), .Q(r1[14]) );
  DFQD1BWP12T r1_reg_13_ ( .D(n2630), .CP(clk), .Q(r1[13]) );
  DFQD1BWP12T r1_reg_12_ ( .D(n2629), .CP(clk), .Q(r1[12]) );
  DFQD1BWP12T r1_reg_11_ ( .D(n2628), .CP(clk), .Q(r1[11]) );
  DFQD1BWP12T r1_reg_10_ ( .D(n2627), .CP(clk), .Q(r1[10]) );
  DFQD1BWP12T r1_reg_9_ ( .D(n2626), .CP(clk), .Q(r1[9]) );
  DFQD1BWP12T r1_reg_8_ ( .D(n2625), .CP(clk), .Q(r1[8]) );
  DFQD1BWP12T r1_reg_7_ ( .D(n2624), .CP(clk), .Q(r1[7]) );
  DFQD1BWP12T r1_reg_6_ ( .D(n2623), .CP(clk), .Q(r1[6]) );
  DFQD1BWP12T r1_reg_5_ ( .D(n2622), .CP(clk), .Q(r1[5]) );
  DFQD1BWP12T r1_reg_4_ ( .D(n2621), .CP(clk), .Q(r1[4]) );
  DFQD1BWP12T r1_reg_3_ ( .D(n2620), .CP(clk), .Q(r1[3]) );
  DFQD1BWP12T r1_reg_2_ ( .D(n2619), .CP(clk), .Q(r1[2]) );
  DFQD1BWP12T r1_reg_1_ ( .D(n2618), .CP(clk), .Q(r1[1]) );
  DFQD1BWP12T r1_reg_0_ ( .D(n2617), .CP(clk), .Q(r1[0]) );
  DFQD1BWP12T r2_reg_31_ ( .D(n2616), .CP(clk), .Q(r2[31]) );
  DFQD1BWP12T r2_reg_30_ ( .D(n2615), .CP(clk), .Q(r2[30]) );
  DFQD1BWP12T r2_reg_29_ ( .D(n2614), .CP(clk), .Q(r2[29]) );
  DFQD1BWP12T r2_reg_28_ ( .D(n2613), .CP(clk), .Q(r2[28]) );
  DFQD1BWP12T r2_reg_27_ ( .D(n2612), .CP(clk), .Q(r2[27]) );
  DFQD1BWP12T r2_reg_26_ ( .D(n2611), .CP(clk), .Q(r2[26]) );
  DFQD1BWP12T r2_reg_25_ ( .D(n2610), .CP(clk), .Q(r2[25]) );
  DFQD1BWP12T r2_reg_24_ ( .D(n2609), .CP(clk), .Q(r2[24]) );
  DFQD1BWP12T r2_reg_23_ ( .D(n2608), .CP(clk), .Q(r2[23]) );
  DFQD1BWP12T r2_reg_22_ ( .D(n2607), .CP(clk), .Q(r2[22]) );
  DFQD1BWP12T r2_reg_21_ ( .D(n2606), .CP(clk), .Q(r2[21]) );
  DFQD1BWP12T r2_reg_20_ ( .D(n2605), .CP(clk), .Q(r2[20]) );
  DFQD1BWP12T r2_reg_19_ ( .D(n2604), .CP(clk), .Q(r2[19]) );
  DFQD1BWP12T r2_reg_18_ ( .D(n2603), .CP(clk), .Q(r2[18]) );
  DFQD1BWP12T r2_reg_17_ ( .D(n2602), .CP(clk), .Q(r2[17]) );
  DFQD1BWP12T r2_reg_16_ ( .D(n2601), .CP(clk), .Q(r2[16]) );
  DFQD1BWP12T r2_reg_15_ ( .D(n2600), .CP(clk), .Q(r2[15]) );
  DFQD1BWP12T r2_reg_14_ ( .D(n2599), .CP(clk), .Q(r2[14]) );
  DFQD1BWP12T r2_reg_13_ ( .D(n2598), .CP(clk), .Q(r2[13]) );
  DFQD1BWP12T r2_reg_12_ ( .D(n2597), .CP(clk), .Q(r2[12]) );
  DFQD1BWP12T r2_reg_11_ ( .D(n2596), .CP(clk), .Q(r2[11]) );
  DFQD1BWP12T r2_reg_10_ ( .D(n2595), .CP(clk), .Q(r2[10]) );
  DFQD1BWP12T r2_reg_9_ ( .D(n2594), .CP(clk), .Q(r2[9]) );
  DFQD1BWP12T r2_reg_8_ ( .D(n2593), .CP(clk), .Q(r2[8]) );
  DFQD1BWP12T r2_reg_7_ ( .D(n2592), .CP(clk), .Q(r2[7]) );
  DFQD1BWP12T r2_reg_6_ ( .D(n2591), .CP(clk), .Q(r2[6]) );
  DFQD1BWP12T r2_reg_5_ ( .D(n2590), .CP(clk), .Q(r2[5]) );
  DFQD1BWP12T r2_reg_4_ ( .D(n2589), .CP(clk), .Q(r2[4]) );
  DFQD1BWP12T r2_reg_3_ ( .D(n2588), .CP(clk), .Q(r2[3]) );
  DFQD1BWP12T r2_reg_2_ ( .D(n2587), .CP(clk), .Q(r2[2]) );
  DFQD1BWP12T r2_reg_1_ ( .D(n2586), .CP(clk), .Q(r2[1]) );
  DFQD1BWP12T r2_reg_0_ ( .D(n2585), .CP(clk), .Q(r2[0]) );
  DFQD1BWP12T r3_reg_31_ ( .D(n2584), .CP(clk), .Q(r3[31]) );
  DFQD1BWP12T r3_reg_30_ ( .D(n2583), .CP(clk), .Q(r3[30]) );
  DFQD1BWP12T r3_reg_29_ ( .D(n2582), .CP(clk), .Q(r3[29]) );
  DFQD1BWP12T r3_reg_28_ ( .D(n2581), .CP(clk), .Q(r3[28]) );
  DFQD1BWP12T r3_reg_27_ ( .D(n2580), .CP(clk), .Q(r3[27]) );
  DFQD1BWP12T r3_reg_26_ ( .D(n2579), .CP(clk), .Q(r3[26]) );
  DFQD1BWP12T r3_reg_25_ ( .D(n2578), .CP(clk), .Q(r3[25]) );
  DFQD1BWP12T r3_reg_24_ ( .D(n2577), .CP(clk), .Q(r3[24]) );
  DFQD1BWP12T r3_reg_23_ ( .D(n2576), .CP(clk), .Q(r3[23]) );
  DFQD1BWP12T r3_reg_22_ ( .D(n2575), .CP(clk), .Q(r3[22]) );
  DFQD1BWP12T r3_reg_21_ ( .D(n2574), .CP(clk), .Q(r3[21]) );
  DFQD1BWP12T r3_reg_20_ ( .D(n2573), .CP(clk), .Q(r3[20]) );
  DFQD1BWP12T r3_reg_19_ ( .D(n2572), .CP(clk), .Q(r3[19]) );
  DFQD1BWP12T r3_reg_18_ ( .D(n2571), .CP(clk), .Q(r3[18]) );
  DFQD1BWP12T r3_reg_17_ ( .D(n2570), .CP(clk), .Q(r3[17]) );
  DFQD1BWP12T r3_reg_16_ ( .D(n2569), .CP(clk), .Q(r3[16]) );
  DFQD1BWP12T r3_reg_15_ ( .D(n2568), .CP(clk), .Q(r3[15]) );
  DFQD1BWP12T r3_reg_14_ ( .D(n2567), .CP(clk), .Q(r3[14]) );
  DFQD1BWP12T r3_reg_13_ ( .D(n2566), .CP(clk), .Q(r3[13]) );
  DFQD1BWP12T r3_reg_12_ ( .D(n2565), .CP(clk), .Q(r3[12]) );
  DFQD1BWP12T r3_reg_11_ ( .D(n2564), .CP(clk), .Q(r3[11]) );
  DFQD1BWP12T r3_reg_10_ ( .D(n2563), .CP(clk), .Q(r3[10]) );
  DFQD1BWP12T r3_reg_9_ ( .D(n2562), .CP(clk), .Q(r3[9]) );
  DFQD1BWP12T r3_reg_8_ ( .D(n2561), .CP(clk), .Q(r3[8]) );
  DFQD1BWP12T r3_reg_7_ ( .D(n2560), .CP(clk), .Q(r3[7]) );
  DFQD1BWP12T r3_reg_6_ ( .D(n2559), .CP(clk), .Q(r3[6]) );
  DFQD1BWP12T r3_reg_5_ ( .D(n2558), .CP(clk), .Q(r3[5]) );
  DFQD1BWP12T r3_reg_4_ ( .D(n2557), .CP(clk), .Q(r3[4]) );
  DFQD1BWP12T r3_reg_3_ ( .D(n2556), .CP(clk), .Q(r3[3]) );
  DFQD1BWP12T r3_reg_2_ ( .D(n2555), .CP(clk), .Q(r3[2]) );
  DFQD1BWP12T r3_reg_1_ ( .D(n2554), .CP(clk), .Q(r3[1]) );
  DFQD1BWP12T r3_reg_0_ ( .D(n2553), .CP(clk), .Q(r3[0]) );
  DFQD1BWP12T r4_reg_31_ ( .D(n2552), .CP(clk), .Q(r4[31]) );
  DFQD1BWP12T r4_reg_30_ ( .D(n2551), .CP(clk), .Q(r4[30]) );
  DFQD1BWP12T r4_reg_29_ ( .D(n2550), .CP(clk), .Q(r4[29]) );
  DFQD1BWP12T r4_reg_28_ ( .D(n2549), .CP(clk), .Q(r4[28]) );
  DFQD1BWP12T r4_reg_27_ ( .D(n2548), .CP(clk), .Q(r4[27]) );
  DFQD1BWP12T r4_reg_26_ ( .D(n2547), .CP(clk), .Q(r4[26]) );
  DFQD1BWP12T r4_reg_25_ ( .D(n2546), .CP(clk), .Q(r4[25]) );
  DFQD1BWP12T r4_reg_24_ ( .D(n2545), .CP(clk), .Q(r4[24]) );
  DFQD1BWP12T r4_reg_23_ ( .D(n2544), .CP(clk), .Q(r4[23]) );
  DFQD1BWP12T r4_reg_22_ ( .D(n2543), .CP(clk), .Q(r4[22]) );
  DFQD1BWP12T r4_reg_21_ ( .D(n2542), .CP(clk), .Q(r4[21]) );
  DFQD1BWP12T r4_reg_20_ ( .D(n2541), .CP(clk), .Q(r4[20]) );
  DFQD1BWP12T r4_reg_19_ ( .D(n2540), .CP(clk), .Q(r4[19]) );
  DFQD1BWP12T r4_reg_18_ ( .D(n2539), .CP(clk), .Q(r4[18]) );
  DFQD1BWP12T r4_reg_17_ ( .D(n2538), .CP(clk), .Q(r4[17]) );
  DFQD1BWP12T r4_reg_16_ ( .D(n2537), .CP(clk), .Q(r4[16]) );
  DFQD1BWP12T r4_reg_15_ ( .D(n2536), .CP(clk), .Q(r4[15]) );
  DFQD1BWP12T r4_reg_14_ ( .D(n2535), .CP(clk), .Q(r4[14]) );
  DFQD1BWP12T r4_reg_13_ ( .D(n2534), .CP(clk), .Q(r4[13]) );
  DFQD1BWP12T r4_reg_12_ ( .D(n2533), .CP(clk), .Q(r4[12]) );
  DFQD1BWP12T r4_reg_11_ ( .D(n2532), .CP(clk), .Q(r4[11]) );
  DFQD1BWP12T r4_reg_10_ ( .D(n2531), .CP(clk), .Q(r4[10]) );
  DFQD1BWP12T r4_reg_9_ ( .D(n2530), .CP(clk), .Q(r4[9]) );
  DFQD1BWP12T r4_reg_8_ ( .D(n2529), .CP(clk), .Q(r4[8]) );
  DFQD1BWP12T r4_reg_7_ ( .D(n2528), .CP(clk), .Q(r4[7]) );
  DFQD1BWP12T r4_reg_6_ ( .D(n2527), .CP(clk), .Q(r4[6]) );
  DFQD1BWP12T r4_reg_5_ ( .D(n2526), .CP(clk), .Q(r4[5]) );
  DFQD1BWP12T r4_reg_4_ ( .D(n2525), .CP(clk), .Q(r4[4]) );
  DFQD1BWP12T r4_reg_3_ ( .D(n2524), .CP(clk), .Q(r4[3]) );
  DFQD1BWP12T r4_reg_2_ ( .D(n2523), .CP(clk), .Q(r4[2]) );
  DFQD1BWP12T r4_reg_1_ ( .D(n2522), .CP(clk), .Q(r4[1]) );
  DFQD1BWP12T r4_reg_0_ ( .D(n2521), .CP(clk), .Q(r4[0]) );
  DFQD1BWP12T r5_reg_31_ ( .D(n2520), .CP(clk), .Q(r5[31]) );
  DFQD1BWP12T r5_reg_30_ ( .D(n2519), .CP(clk), .Q(r5[30]) );
  DFQD1BWP12T r5_reg_29_ ( .D(n2518), .CP(clk), .Q(r5[29]) );
  DFQD1BWP12T r5_reg_28_ ( .D(n2517), .CP(clk), .Q(r5[28]) );
  DFQD1BWP12T r5_reg_27_ ( .D(n2516), .CP(clk), .Q(r5[27]) );
  DFQD1BWP12T r5_reg_26_ ( .D(n2515), .CP(clk), .Q(r5[26]) );
  DFQD1BWP12T r5_reg_25_ ( .D(n2514), .CP(clk), .Q(r5[25]) );
  DFQD1BWP12T r5_reg_24_ ( .D(n2513), .CP(clk), .Q(r5[24]) );
  DFQD1BWP12T r5_reg_23_ ( .D(n2512), .CP(clk), .Q(r5[23]) );
  DFQD1BWP12T r5_reg_22_ ( .D(n2511), .CP(clk), .Q(r5[22]) );
  DFQD1BWP12T r5_reg_21_ ( .D(n2510), .CP(clk), .Q(r5[21]) );
  DFQD1BWP12T r5_reg_20_ ( .D(n2509), .CP(clk), .Q(r5[20]) );
  DFQD1BWP12T r5_reg_19_ ( .D(n2508), .CP(clk), .Q(r5[19]) );
  DFQD1BWP12T r5_reg_18_ ( .D(n2507), .CP(clk), .Q(r5[18]) );
  DFQD1BWP12T r5_reg_17_ ( .D(n2506), .CP(clk), .Q(r5[17]) );
  DFQD1BWP12T r5_reg_16_ ( .D(n2505), .CP(clk), .Q(r5[16]) );
  DFQD1BWP12T r5_reg_15_ ( .D(n2504), .CP(clk), .Q(r5[15]) );
  DFQD1BWP12T r5_reg_14_ ( .D(n2503), .CP(clk), .Q(r5[14]) );
  DFQD1BWP12T r5_reg_13_ ( .D(n2502), .CP(clk), .Q(r5[13]) );
  DFQD1BWP12T r5_reg_12_ ( .D(n2501), .CP(clk), .Q(r5[12]) );
  DFQD1BWP12T r5_reg_11_ ( .D(n2500), .CP(clk), .Q(r5[11]) );
  DFQD1BWP12T r5_reg_10_ ( .D(n2499), .CP(clk), .Q(r5[10]) );
  DFQD1BWP12T r5_reg_9_ ( .D(n2498), .CP(clk), .Q(r5[9]) );
  DFQD1BWP12T r5_reg_8_ ( .D(n2497), .CP(clk), .Q(r5[8]) );
  DFQD1BWP12T r5_reg_7_ ( .D(n2496), .CP(clk), .Q(r5[7]) );
  DFQD1BWP12T r5_reg_6_ ( .D(n2495), .CP(clk), .Q(r5[6]) );
  DFQD1BWP12T r5_reg_5_ ( .D(n2494), .CP(clk), .Q(r5[5]) );
  DFQD1BWP12T r5_reg_4_ ( .D(n2493), .CP(clk), .Q(r5[4]) );
  DFQD1BWP12T r5_reg_3_ ( .D(n2492), .CP(clk), .Q(r5[3]) );
  DFQD1BWP12T r5_reg_2_ ( .D(n2491), .CP(clk), .Q(r5[2]) );
  DFQD1BWP12T r5_reg_1_ ( .D(n2490), .CP(clk), .Q(r5[1]) );
  DFQD1BWP12T r5_reg_0_ ( .D(n2489), .CP(clk), .Q(r5[0]) );
  DFQD1BWP12T r6_reg_31_ ( .D(n2488), .CP(clk), .Q(r6[31]) );
  DFQD1BWP12T r6_reg_30_ ( .D(n2487), .CP(clk), .Q(r6[30]) );
  DFQD1BWP12T r6_reg_29_ ( .D(n2486), .CP(clk), .Q(r6[29]) );
  DFQD1BWP12T r6_reg_28_ ( .D(n2485), .CP(clk), .Q(r6[28]) );
  DFQD1BWP12T r6_reg_27_ ( .D(n2484), .CP(clk), .Q(r6[27]) );
  DFQD1BWP12T r6_reg_26_ ( .D(n2483), .CP(clk), .Q(r6[26]) );
  DFQD1BWP12T r6_reg_25_ ( .D(n2482), .CP(clk), .Q(r6[25]) );
  DFQD1BWP12T r6_reg_24_ ( .D(n2481), .CP(clk), .Q(r6[24]) );
  DFQD1BWP12T r6_reg_23_ ( .D(n2480), .CP(clk), .Q(r6[23]) );
  DFQD1BWP12T r6_reg_22_ ( .D(n2479), .CP(clk), .Q(r6[22]) );
  DFQD1BWP12T r6_reg_21_ ( .D(n2478), .CP(clk), .Q(r6[21]) );
  DFQD1BWP12T r6_reg_20_ ( .D(n2477), .CP(clk), .Q(r6[20]) );
  DFQD1BWP12T r6_reg_19_ ( .D(n2476), .CP(clk), .Q(r6[19]) );
  DFQD1BWP12T r6_reg_18_ ( .D(n2475), .CP(clk), .Q(r6[18]) );
  DFQD1BWP12T r6_reg_17_ ( .D(n2474), .CP(clk), .Q(r6[17]) );
  DFQD1BWP12T r6_reg_16_ ( .D(n2473), .CP(clk), .Q(r6[16]) );
  DFQD1BWP12T r6_reg_15_ ( .D(n2472), .CP(clk), .Q(r6[15]) );
  DFQD1BWP12T r6_reg_14_ ( .D(n2471), .CP(clk), .Q(r6[14]) );
  DFQD1BWP12T r6_reg_13_ ( .D(n2470), .CP(clk), .Q(r6[13]) );
  DFQD1BWP12T r6_reg_12_ ( .D(n2469), .CP(clk), .Q(r6[12]) );
  DFQD1BWP12T r6_reg_11_ ( .D(n2468), .CP(clk), .Q(r6[11]) );
  DFQD1BWP12T r6_reg_10_ ( .D(n2467), .CP(clk), .Q(r6[10]) );
  DFQD1BWP12T r6_reg_9_ ( .D(n2466), .CP(clk), .Q(r6[9]) );
  DFQD1BWP12T r6_reg_8_ ( .D(n2465), .CP(clk), .Q(r6[8]) );
  DFQD1BWP12T r6_reg_7_ ( .D(n2464), .CP(clk), .Q(r6[7]) );
  DFQD1BWP12T r6_reg_6_ ( .D(n2463), .CP(clk), .Q(r6[6]) );
  DFQD1BWP12T r6_reg_5_ ( .D(n2462), .CP(clk), .Q(r6[5]) );
  DFQD1BWP12T r6_reg_4_ ( .D(n2461), .CP(clk), .Q(r6[4]) );
  DFQD1BWP12T r6_reg_3_ ( .D(n2460), .CP(clk), .Q(r6[3]) );
  DFQD1BWP12T r6_reg_2_ ( .D(n2459), .CP(clk), .Q(r6[2]) );
  DFQD1BWP12T r6_reg_1_ ( .D(n2458), .CP(clk), .Q(r6[1]) );
  DFQD1BWP12T r6_reg_0_ ( .D(n2457), .CP(clk), .Q(r6[0]) );
  DFQD1BWP12T r7_reg_31_ ( .D(n2456), .CP(clk), .Q(r7[31]) );
  DFQD1BWP12T r7_reg_30_ ( .D(n2455), .CP(clk), .Q(r7[30]) );
  DFQD1BWP12T r7_reg_29_ ( .D(n2454), .CP(clk), .Q(r7[29]) );
  DFQD1BWP12T r7_reg_28_ ( .D(n2453), .CP(clk), .Q(r7[28]) );
  DFQD1BWP12T r7_reg_27_ ( .D(n2452), .CP(clk), .Q(r7[27]) );
  DFQD1BWP12T r7_reg_26_ ( .D(n2451), .CP(clk), .Q(r7[26]) );
  DFQD1BWP12T r7_reg_25_ ( .D(n2450), .CP(clk), .Q(r7[25]) );
  DFQD1BWP12T r7_reg_24_ ( .D(n2449), .CP(clk), .Q(r7[24]) );
  DFQD1BWP12T r7_reg_23_ ( .D(n2448), .CP(clk), .Q(r7[23]) );
  DFQD1BWP12T r7_reg_22_ ( .D(n2447), .CP(clk), .Q(r7[22]) );
  DFQD1BWP12T r7_reg_21_ ( .D(n2446), .CP(clk), .Q(r7[21]) );
  DFQD1BWP12T r7_reg_20_ ( .D(n2445), .CP(clk), .Q(r7[20]) );
  DFQD1BWP12T r7_reg_19_ ( .D(n2444), .CP(clk), .Q(r7[19]) );
  DFQD1BWP12T r7_reg_18_ ( .D(n2443), .CP(clk), .Q(r7[18]) );
  DFQD1BWP12T r7_reg_17_ ( .D(n2442), .CP(clk), .Q(r7[17]) );
  DFQD1BWP12T r7_reg_16_ ( .D(n2441), .CP(clk), .Q(r7[16]) );
  DFQD1BWP12T r7_reg_15_ ( .D(n2440), .CP(clk), .Q(r7[15]) );
  DFQD1BWP12T r7_reg_14_ ( .D(n2439), .CP(clk), .Q(r7[14]) );
  DFQD1BWP12T r7_reg_13_ ( .D(n2438), .CP(clk), .Q(r7[13]) );
  DFQD1BWP12T r7_reg_12_ ( .D(n2437), .CP(clk), .Q(r7[12]) );
  DFQD1BWP12T r7_reg_11_ ( .D(n2436), .CP(clk), .Q(r7[11]) );
  DFQD1BWP12T r7_reg_10_ ( .D(n2435), .CP(clk), .Q(r7[10]) );
  DFQD1BWP12T r7_reg_9_ ( .D(n2434), .CP(clk), .Q(r7[9]) );
  DFQD1BWP12T r7_reg_8_ ( .D(n2433), .CP(clk), .Q(r7[8]) );
  DFQD1BWP12T r7_reg_7_ ( .D(n2432), .CP(clk), .Q(r7[7]) );
  DFQD1BWP12T r7_reg_6_ ( .D(n2431), .CP(clk), .Q(r7[6]) );
  DFQD1BWP12T r7_reg_5_ ( .D(n2430), .CP(clk), .Q(r7[5]) );
  DFQD1BWP12T r7_reg_4_ ( .D(n2429), .CP(clk), .Q(r7[4]) );
  DFQD1BWP12T r7_reg_3_ ( .D(n2428), .CP(clk), .Q(r7[3]) );
  DFQD1BWP12T r7_reg_2_ ( .D(n2427), .CP(clk), .Q(r7[2]) );
  DFQD1BWP12T r7_reg_1_ ( .D(n2426), .CP(clk), .Q(r7[1]) );
  DFQD1BWP12T r7_reg_0_ ( .D(n2425), .CP(clk), .Q(r7[0]) );
  DFQD1BWP12T r8_reg_31_ ( .D(n2424), .CP(clk), .Q(r8[31]) );
  DFQD1BWP12T r8_reg_30_ ( .D(n2423), .CP(clk), .Q(r8[30]) );
  DFQD1BWP12T r8_reg_29_ ( .D(n2422), .CP(clk), .Q(r8[29]) );
  DFQD1BWP12T r8_reg_28_ ( .D(n2421), .CP(clk), .Q(r8[28]) );
  DFQD1BWP12T r8_reg_27_ ( .D(n2420), .CP(clk), .Q(r8[27]) );
  DFQD1BWP12T r8_reg_26_ ( .D(n2419), .CP(clk), .Q(r8[26]) );
  DFQD1BWP12T r8_reg_25_ ( .D(n2418), .CP(clk), .Q(r8[25]) );
  DFQD1BWP12T r8_reg_24_ ( .D(n2417), .CP(clk), .Q(r8[24]) );
  DFQD1BWP12T r8_reg_23_ ( .D(n2416), .CP(clk), .Q(r8[23]) );
  DFQD1BWP12T r8_reg_22_ ( .D(n2415), .CP(clk), .Q(r8[22]) );
  DFQD1BWP12T r8_reg_21_ ( .D(n2414), .CP(clk), .Q(r8[21]) );
  DFQD1BWP12T r8_reg_20_ ( .D(n2413), .CP(clk), .Q(r8[20]) );
  DFQD1BWP12T r8_reg_19_ ( .D(n2412), .CP(clk), .Q(r8[19]) );
  DFQD1BWP12T r8_reg_18_ ( .D(n2411), .CP(clk), .Q(r8[18]) );
  DFQD1BWP12T r8_reg_17_ ( .D(n2410), .CP(clk), .Q(r8[17]) );
  DFQD1BWP12T r8_reg_16_ ( .D(n2409), .CP(clk), .Q(r8[16]) );
  DFQD1BWP12T r8_reg_15_ ( .D(n2408), .CP(clk), .Q(r8[15]) );
  DFQD1BWP12T r8_reg_14_ ( .D(n2407), .CP(clk), .Q(r8[14]) );
  DFQD1BWP12T r8_reg_13_ ( .D(n2406), .CP(clk), .Q(r8[13]) );
  DFQD1BWP12T r8_reg_12_ ( .D(n2405), .CP(clk), .Q(r8[12]) );
  DFQD1BWP12T r8_reg_11_ ( .D(n2404), .CP(clk), .Q(r8[11]) );
  DFQD1BWP12T r8_reg_10_ ( .D(n2403), .CP(clk), .Q(r8[10]) );
  DFQD1BWP12T r8_reg_9_ ( .D(n2402), .CP(clk), .Q(r8[9]) );
  DFQD1BWP12T r8_reg_8_ ( .D(n2401), .CP(clk), .Q(r8[8]) );
  DFQD1BWP12T r8_reg_7_ ( .D(n2400), .CP(clk), .Q(r8[7]) );
  DFQD1BWP12T r8_reg_6_ ( .D(n2399), .CP(clk), .Q(r8[6]) );
  DFQD1BWP12T r8_reg_5_ ( .D(n2398), .CP(clk), .Q(r8[5]) );
  DFQD1BWP12T r8_reg_4_ ( .D(n2397), .CP(clk), .Q(r8[4]) );
  DFQD1BWP12T r8_reg_3_ ( .D(n2396), .CP(clk), .Q(r8[3]) );
  DFQD1BWP12T r8_reg_2_ ( .D(n2395), .CP(clk), .Q(r8[2]) );
  DFQD1BWP12T r8_reg_1_ ( .D(n2394), .CP(clk), .Q(r8[1]) );
  DFQD1BWP12T r8_reg_0_ ( .D(n2393), .CP(clk), .Q(r8[0]) );
  DFQD1BWP12T r9_reg_31_ ( .D(n2392), .CP(clk), .Q(r9[31]) );
  DFQD1BWP12T r9_reg_30_ ( .D(n2391), .CP(clk), .Q(r9[30]) );
  DFQD1BWP12T r9_reg_29_ ( .D(n2390), .CP(clk), .Q(r9[29]) );
  DFQD1BWP12T r9_reg_28_ ( .D(n2389), .CP(clk), .Q(r9[28]) );
  DFQD1BWP12T r9_reg_27_ ( .D(n2388), .CP(clk), .Q(r9[27]) );
  DFQD1BWP12T r9_reg_26_ ( .D(n2387), .CP(clk), .Q(r9[26]) );
  DFQD1BWP12T r9_reg_25_ ( .D(n2386), .CP(clk), .Q(r9[25]) );
  DFQD1BWP12T r9_reg_24_ ( .D(n2385), .CP(clk), .Q(r9[24]) );
  DFQD1BWP12T r9_reg_23_ ( .D(n2384), .CP(clk), .Q(r9[23]) );
  DFQD1BWP12T r9_reg_22_ ( .D(n2383), .CP(clk), .Q(r9[22]) );
  DFQD1BWP12T r9_reg_21_ ( .D(n2382), .CP(clk), .Q(r9[21]) );
  DFQD1BWP12T r9_reg_20_ ( .D(n2381), .CP(clk), .Q(r9[20]) );
  DFQD1BWP12T r9_reg_19_ ( .D(n2380), .CP(clk), .Q(r9[19]) );
  DFQD1BWP12T r9_reg_18_ ( .D(n2379), .CP(clk), .Q(r9[18]) );
  DFQD1BWP12T r9_reg_17_ ( .D(n2378), .CP(clk), .Q(r9[17]) );
  DFQD1BWP12T r9_reg_16_ ( .D(n2377), .CP(clk), .Q(r9[16]) );
  DFQD1BWP12T r9_reg_15_ ( .D(n2376), .CP(clk), .Q(r9[15]) );
  DFQD1BWP12T r9_reg_14_ ( .D(n2375), .CP(clk), .Q(r9[14]) );
  DFQD1BWP12T r9_reg_13_ ( .D(n2374), .CP(clk), .Q(r9[13]) );
  DFQD1BWP12T r9_reg_12_ ( .D(n2373), .CP(clk), .Q(r9[12]) );
  DFQD1BWP12T r9_reg_11_ ( .D(n2372), .CP(clk), .Q(r9[11]) );
  DFQD1BWP12T r9_reg_10_ ( .D(n2371), .CP(clk), .Q(r9[10]) );
  DFQD1BWP12T r9_reg_9_ ( .D(n2370), .CP(clk), .Q(r9[9]) );
  DFQD1BWP12T r9_reg_8_ ( .D(n2369), .CP(clk), .Q(r9[8]) );
  DFQD1BWP12T r9_reg_7_ ( .D(n2368), .CP(clk), .Q(r9[7]) );
  DFQD1BWP12T r9_reg_6_ ( .D(n2367), .CP(clk), .Q(r9[6]) );
  DFQD1BWP12T r9_reg_5_ ( .D(n2366), .CP(clk), .Q(r9[5]) );
  DFQD1BWP12T r9_reg_4_ ( .D(n2365), .CP(clk), .Q(r9[4]) );
  DFQD1BWP12T r9_reg_3_ ( .D(n2364), .CP(clk), .Q(r9[3]) );
  DFQD1BWP12T r9_reg_2_ ( .D(n2363), .CP(clk), .Q(r9[2]) );
  DFQD1BWP12T r9_reg_1_ ( .D(n2362), .CP(clk), .Q(r9[1]) );
  DFQD1BWP12T r9_reg_0_ ( .D(n2361), .CP(clk), .Q(r9[0]) );
  DFQD1BWP12T r10_reg_31_ ( .D(n2360), .CP(clk), .Q(r10[31]) );
  DFQD1BWP12T r10_reg_30_ ( .D(n2359), .CP(clk), .Q(r10[30]) );
  DFQD1BWP12T r10_reg_29_ ( .D(n2358), .CP(clk), .Q(r10[29]) );
  DFQD1BWP12T r10_reg_28_ ( .D(n2357), .CP(clk), .Q(r10[28]) );
  DFQD1BWP12T r10_reg_27_ ( .D(n2356), .CP(clk), .Q(r10[27]) );
  DFQD1BWP12T r10_reg_26_ ( .D(n2355), .CP(clk), .Q(r10[26]) );
  DFQD1BWP12T r10_reg_25_ ( .D(n2354), .CP(clk), .Q(r10[25]) );
  DFQD1BWP12T r10_reg_24_ ( .D(n2353), .CP(clk), .Q(r10[24]) );
  DFQD1BWP12T r10_reg_23_ ( .D(n2352), .CP(clk), .Q(r10[23]) );
  DFQD1BWP12T r10_reg_22_ ( .D(n2351), .CP(clk), .Q(r10[22]) );
  DFQD1BWP12T r10_reg_21_ ( .D(n2350), .CP(clk), .Q(r10[21]) );
  DFQD1BWP12T r10_reg_20_ ( .D(n2349), .CP(clk), .Q(r10[20]) );
  DFQD1BWP12T r10_reg_19_ ( .D(n2348), .CP(clk), .Q(r10[19]) );
  DFQD1BWP12T r10_reg_18_ ( .D(n2347), .CP(clk), .Q(r10[18]) );
  DFQD1BWP12T r10_reg_17_ ( .D(n2346), .CP(clk), .Q(r10[17]) );
  DFQD1BWP12T r10_reg_16_ ( .D(n2345), .CP(clk), .Q(r10[16]) );
  DFQD1BWP12T r10_reg_15_ ( .D(n2344), .CP(clk), .Q(r10[15]) );
  DFQD1BWP12T r10_reg_14_ ( .D(n2343), .CP(clk), .Q(r10[14]) );
  DFQD1BWP12T r10_reg_13_ ( .D(n2342), .CP(clk), .Q(r10[13]) );
  DFQD1BWP12T r10_reg_12_ ( .D(n2341), .CP(clk), .Q(r10[12]) );
  DFQD1BWP12T r10_reg_11_ ( .D(n2340), .CP(clk), .Q(r10[11]) );
  DFQD1BWP12T r10_reg_10_ ( .D(n2339), .CP(clk), .Q(r10[10]) );
  DFQD1BWP12T r10_reg_9_ ( .D(n2338), .CP(clk), .Q(r10[9]) );
  DFQD1BWP12T r10_reg_8_ ( .D(n2337), .CP(clk), .Q(r10[8]) );
  DFQD1BWP12T r10_reg_7_ ( .D(n2336), .CP(clk), .Q(r10[7]) );
  DFQD1BWP12T r10_reg_6_ ( .D(n2335), .CP(clk), .Q(r10[6]) );
  DFQD1BWP12T r10_reg_5_ ( .D(n2334), .CP(clk), .Q(r10[5]) );
  DFQD1BWP12T r10_reg_4_ ( .D(n2333), .CP(clk), .Q(r10[4]) );
  DFQD1BWP12T r10_reg_3_ ( .D(n2332), .CP(clk), .Q(r10[3]) );
  DFQD1BWP12T r10_reg_2_ ( .D(n2331), .CP(clk), .Q(r10[2]) );
  DFQD1BWP12T r10_reg_1_ ( .D(n2330), .CP(clk), .Q(r10[1]) );
  DFQD1BWP12T r10_reg_0_ ( .D(n2329), .CP(clk), .Q(r10[0]) );
  DFQD1BWP12T r11_reg_31_ ( .D(n2328), .CP(clk), .Q(r11[31]) );
  DFQD1BWP12T r11_reg_30_ ( .D(n2327), .CP(clk), .Q(r11[30]) );
  DFQD1BWP12T r11_reg_29_ ( .D(n2326), .CP(clk), .Q(r11[29]) );
  DFQD1BWP12T r11_reg_28_ ( .D(n2325), .CP(clk), .Q(r11[28]) );
  DFQD1BWP12T r11_reg_27_ ( .D(n2324), .CP(clk), .Q(r11[27]) );
  DFQD1BWP12T r11_reg_26_ ( .D(n2323), .CP(clk), .Q(r11[26]) );
  DFQD1BWP12T r11_reg_25_ ( .D(n2322), .CP(clk), .Q(r11[25]) );
  DFQD1BWP12T r11_reg_24_ ( .D(n2321), .CP(clk), .Q(r11[24]) );
  DFQD1BWP12T r11_reg_23_ ( .D(n2320), .CP(clk), .Q(r11[23]) );
  DFQD1BWP12T r11_reg_22_ ( .D(n2319), .CP(clk), .Q(r11[22]) );
  DFQD1BWP12T r11_reg_21_ ( .D(n2318), .CP(clk), .Q(r11[21]) );
  DFQD1BWP12T r11_reg_20_ ( .D(n2317), .CP(clk), .Q(r11[20]) );
  DFQD1BWP12T r11_reg_19_ ( .D(n2316), .CP(clk), .Q(r11[19]) );
  DFQD1BWP12T r11_reg_18_ ( .D(n2315), .CP(clk), .Q(r11[18]) );
  DFQD1BWP12T r11_reg_17_ ( .D(n2314), .CP(clk), .Q(r11[17]) );
  DFQD1BWP12T r11_reg_16_ ( .D(n2313), .CP(clk), .Q(r11[16]) );
  DFQD1BWP12T r11_reg_15_ ( .D(n2312), .CP(clk), .Q(r11[15]) );
  DFQD1BWP12T r11_reg_14_ ( .D(n2311), .CP(clk), .Q(r11[14]) );
  DFQD1BWP12T r11_reg_13_ ( .D(n2310), .CP(clk), .Q(r11[13]) );
  DFQD1BWP12T r11_reg_12_ ( .D(n2309), .CP(clk), .Q(r11[12]) );
  DFQD1BWP12T r11_reg_11_ ( .D(n2308), .CP(clk), .Q(r11[11]) );
  DFQD1BWP12T r11_reg_10_ ( .D(n2307), .CP(clk), .Q(r11[10]) );
  DFQD1BWP12T r11_reg_9_ ( .D(n2306), .CP(clk), .Q(r11[9]) );
  DFQD1BWP12T r11_reg_8_ ( .D(n2305), .CP(clk), .Q(r11[8]) );
  DFQD1BWP12T r11_reg_7_ ( .D(n2304), .CP(clk), .Q(r11[7]) );
  DFQD1BWP12T r11_reg_6_ ( .D(n2303), .CP(clk), .Q(r11[6]) );
  DFQD1BWP12T r11_reg_5_ ( .D(n2302), .CP(clk), .Q(r11[5]) );
  DFQD1BWP12T r11_reg_4_ ( .D(n2301), .CP(clk), .Q(r11[4]) );
  DFQD1BWP12T r11_reg_3_ ( .D(n2300), .CP(clk), .Q(r11[3]) );
  DFQD1BWP12T r11_reg_2_ ( .D(n2299), .CP(clk), .Q(r11[2]) );
  DFQD1BWP12T r11_reg_1_ ( .D(n2298), .CP(clk), .Q(r11[1]) );
  DFQD1BWP12T r11_reg_0_ ( .D(n2297), .CP(clk), .Q(r11[0]) );
  DFQD1BWP12T r12_reg_31_ ( .D(n2296), .CP(clk), .Q(r12[31]) );
  DFQD1BWP12T r12_reg_30_ ( .D(n2295), .CP(clk), .Q(r12[30]) );
  DFQD1BWP12T r12_reg_29_ ( .D(n2294), .CP(clk), .Q(r12[29]) );
  DFQD1BWP12T r12_reg_28_ ( .D(n2293), .CP(clk), .Q(r12[28]) );
  DFQD1BWP12T r12_reg_27_ ( .D(n2292), .CP(clk), .Q(r12[27]) );
  DFQD1BWP12T r12_reg_26_ ( .D(n2291), .CP(clk), .Q(r12[26]) );
  DFQD1BWP12T r12_reg_25_ ( .D(n2290), .CP(clk), .Q(r12[25]) );
  DFQD1BWP12T r12_reg_24_ ( .D(n2289), .CP(clk), .Q(r12[24]) );
  DFQD1BWP12T r12_reg_23_ ( .D(n2288), .CP(clk), .Q(r12[23]) );
  DFQD1BWP12T r12_reg_22_ ( .D(n2287), .CP(clk), .Q(r12[22]) );
  DFQD1BWP12T r12_reg_21_ ( .D(n2286), .CP(clk), .Q(r12[21]) );
  DFQD1BWP12T r12_reg_20_ ( .D(n2285), .CP(clk), .Q(r12[20]) );
  DFQD1BWP12T r12_reg_19_ ( .D(n2284), .CP(clk), .Q(r12[19]) );
  DFQD1BWP12T r12_reg_18_ ( .D(n2283), .CP(clk), .Q(r12[18]) );
  DFQD1BWP12T r12_reg_17_ ( .D(n2282), .CP(clk), .Q(r12[17]) );
  DFQD1BWP12T r12_reg_16_ ( .D(n2281), .CP(clk), .Q(r12[16]) );
  DFQD1BWP12T r12_reg_15_ ( .D(n2280), .CP(clk), .Q(r12[15]) );
  DFQD1BWP12T r12_reg_14_ ( .D(n2279), .CP(clk), .Q(r12[14]) );
  DFQD1BWP12T r12_reg_13_ ( .D(n2278), .CP(clk), .Q(r12[13]) );
  DFQD1BWP12T r12_reg_12_ ( .D(n2277), .CP(clk), .Q(r12[12]) );
  DFQD1BWP12T r12_reg_11_ ( .D(n2276), .CP(clk), .Q(r12[11]) );
  DFQD1BWP12T r12_reg_10_ ( .D(n2275), .CP(clk), .Q(r12[10]) );
  DFQD1BWP12T r12_reg_9_ ( .D(n2274), .CP(clk), .Q(r12[9]) );
  DFQD1BWP12T r12_reg_8_ ( .D(n2273), .CP(clk), .Q(r12[8]) );
  DFQD1BWP12T r12_reg_7_ ( .D(n2272), .CP(clk), .Q(r12[7]) );
  DFQD1BWP12T r12_reg_6_ ( .D(n2271), .CP(clk), .Q(r12[6]) );
  DFQD1BWP12T r12_reg_5_ ( .D(n2270), .CP(clk), .Q(r12[5]) );
  DFQD1BWP12T r12_reg_4_ ( .D(n2269), .CP(clk), .Q(r12[4]) );
  DFQD1BWP12T r12_reg_3_ ( .D(n2268), .CP(clk), .Q(r12[3]) );
  DFQD1BWP12T r12_reg_2_ ( .D(n2267), .CP(clk), .Q(r12[2]) );
  DFQD1BWP12T r12_reg_1_ ( .D(n2266), .CP(clk), .Q(r12[1]) );
  DFQD1BWP12T r12_reg_0_ ( .D(n2265), .CP(clk), .Q(r12[0]) );
  DFQD1BWP12T lr_reg_31_ ( .D(n2264), .CP(clk), .Q(lr[31]) );
  DFQD1BWP12T lr_reg_30_ ( .D(n2263), .CP(clk), .Q(lr[30]) );
  DFQD1BWP12T lr_reg_29_ ( .D(n2262), .CP(clk), .Q(lr[29]) );
  DFQD1BWP12T lr_reg_28_ ( .D(n2261), .CP(clk), .Q(lr[28]) );
  DFQD1BWP12T lr_reg_27_ ( .D(n2260), .CP(clk), .Q(lr[27]) );
  DFQD1BWP12T lr_reg_26_ ( .D(n2259), .CP(clk), .Q(lr[26]) );
  DFQD1BWP12T lr_reg_25_ ( .D(n2258), .CP(clk), .Q(lr[25]) );
  DFQD1BWP12T lr_reg_24_ ( .D(n2257), .CP(clk), .Q(lr[24]) );
  DFQD1BWP12T lr_reg_23_ ( .D(n2256), .CP(clk), .Q(lr[23]) );
  DFQD1BWP12T lr_reg_22_ ( .D(n2255), .CP(clk), .Q(lr[22]) );
  DFQD1BWP12T lr_reg_21_ ( .D(n2254), .CP(clk), .Q(lr[21]) );
  DFQD1BWP12T lr_reg_20_ ( .D(n2253), .CP(clk), .Q(lr[20]) );
  DFQD1BWP12T lr_reg_19_ ( .D(n2252), .CP(clk), .Q(lr[19]) );
  DFQD1BWP12T lr_reg_18_ ( .D(n2251), .CP(clk), .Q(lr[18]) );
  DFQD1BWP12T lr_reg_17_ ( .D(n2250), .CP(clk), .Q(lr[17]) );
  DFQD1BWP12T lr_reg_16_ ( .D(n2249), .CP(clk), .Q(lr[16]) );
  DFQD1BWP12T lr_reg_15_ ( .D(n2248), .CP(clk), .Q(lr[15]) );
  DFQD1BWP12T lr_reg_14_ ( .D(n2247), .CP(clk), .Q(lr[14]) );
  DFQD1BWP12T lr_reg_13_ ( .D(n2246), .CP(clk), .Q(lr[13]) );
  DFQD1BWP12T lr_reg_12_ ( .D(n2245), .CP(clk), .Q(lr[12]) );
  DFQD1BWP12T lr_reg_11_ ( .D(n2244), .CP(clk), .Q(lr[11]) );
  DFQD1BWP12T lr_reg_10_ ( .D(n2243), .CP(clk), .Q(lr[10]) );
  DFQD1BWP12T lr_reg_9_ ( .D(n2242), .CP(clk), .Q(lr[9]) );
  DFQD1BWP12T lr_reg_8_ ( .D(n2241), .CP(clk), .Q(lr[8]) );
  DFQD1BWP12T lr_reg_7_ ( .D(n2240), .CP(clk), .Q(lr[7]) );
  DFQD1BWP12T lr_reg_6_ ( .D(n2239), .CP(clk), .Q(lr[6]) );
  DFQD1BWP12T lr_reg_5_ ( .D(n2238), .CP(clk), .Q(lr[5]) );
  DFQD1BWP12T lr_reg_4_ ( .D(n2237), .CP(clk), .Q(lr[4]) );
  DFQD1BWP12T lr_reg_3_ ( .D(n2236), .CP(clk), .Q(lr[3]) );
  DFQD1BWP12T lr_reg_2_ ( .D(n2235), .CP(clk), .Q(lr[2]) );
  DFQD1BWP12T lr_reg_1_ ( .D(n2234), .CP(clk), .Q(lr[1]) );
  DFQD1BWP12T lr_reg_0_ ( .D(n2233), .CP(clk), .Q(lr[0]) );
  DFQD1BWP12T sp_reg_31_ ( .D(spin[31]), .CP(clk), .Q(sp_out[31]) );
  DFQD1BWP12T sp_reg_30_ ( .D(spin[30]), .CP(clk), .Q(sp_out[30]) );
  DFQD1BWP12T sp_reg_29_ ( .D(spin[29]), .CP(clk), .Q(sp_out[29]) );
  DFQD1BWP12T sp_reg_28_ ( .D(spin[28]), .CP(clk), .Q(sp_out[28]) );
  DFQD1BWP12T sp_reg_27_ ( .D(spin[27]), .CP(clk), .Q(sp_out[27]) );
  DFQD1BWP12T sp_reg_26_ ( .D(spin[26]), .CP(clk), .Q(sp_out[26]) );
  DFQD1BWP12T sp_reg_25_ ( .D(spin[25]), .CP(clk), .Q(sp_out[25]) );
  DFQD1BWP12T sp_reg_24_ ( .D(spin[24]), .CP(clk), .Q(sp_out[24]) );
  DFQD1BWP12T sp_reg_23_ ( .D(spin[23]), .CP(clk), .Q(sp_out[23]) );
  DFQD1BWP12T sp_reg_22_ ( .D(spin[22]), .CP(clk), .Q(sp_out[22]) );
  DFQD1BWP12T sp_reg_21_ ( .D(spin[21]), .CP(clk), .Q(sp_out[21]) );
  DFQD1BWP12T sp_reg_20_ ( .D(spin[20]), .CP(clk), .Q(sp_out[20]) );
  DFQD1BWP12T sp_reg_19_ ( .D(spin[19]), .CP(clk), .Q(sp_out[19]) );
  DFQD1BWP12T sp_reg_18_ ( .D(spin[18]), .CP(clk), .Q(sp_out[18]) );
  DFQD1BWP12T sp_reg_17_ ( .D(spin[17]), .CP(clk), .Q(sp_out[17]) );
  DFQD1BWP12T sp_reg_16_ ( .D(spin[16]), .CP(clk), .Q(sp_out[16]) );
  DFQD1BWP12T sp_reg_15_ ( .D(spin[15]), .CP(clk), .Q(sp_out[15]) );
  DFQD1BWP12T sp_reg_14_ ( .D(spin[14]), .CP(clk), .Q(sp_out[14]) );
  DFQD1BWP12T sp_reg_13_ ( .D(spin[13]), .CP(clk), .Q(sp_out[13]) );
  DFQD1BWP12T sp_reg_12_ ( .D(spin[12]), .CP(clk), .Q(sp_out[12]) );
  DFQD1BWP12T sp_reg_11_ ( .D(spin[11]), .CP(clk), .Q(sp_out[11]) );
  DFQD1BWP12T sp_reg_10_ ( .D(spin[10]), .CP(clk), .Q(sp_out[10]) );
  DFQD1BWP12T sp_reg_9_ ( .D(spin[9]), .CP(clk), .Q(sp_out[9]) );
  DFQD1BWP12T sp_reg_8_ ( .D(spin[8]), .CP(clk), .Q(sp_out[8]) );
  DFQD1BWP12T sp_reg_7_ ( .D(spin[7]), .CP(clk), .Q(sp_out[7]) );
  DFQD1BWP12T sp_reg_6_ ( .D(spin[6]), .CP(clk), .Q(sp_out[6]) );
  DFQD1BWP12T sp_reg_5_ ( .D(spin[5]), .CP(clk), .Q(sp_out[5]) );
  DFQD1BWP12T sp_reg_4_ ( .D(spin[4]), .CP(clk), .Q(sp_out[4]) );
  DFQD1BWP12T sp_reg_3_ ( .D(spin[3]), .CP(clk), .Q(sp_out[3]) );
  DFQD1BWP12T sp_reg_2_ ( .D(spin[2]), .CP(clk), .Q(sp_out[2]) );
  DFQD1BWP12T sp_reg_1_ ( .D(spin[1]), .CP(clk), .Q(sp_out[1]) );
  DFQD1BWP12T sp_reg_0_ ( .D(spin[0]), .CP(clk), .Q(sp_out[0]) );
  DFQD1BWP12T pc_reg_31_ ( .D(n2232), .CP(clk), .Q(pc_out[31]) );
  DFQD1BWP12T pc_reg_30_ ( .D(n2231), .CP(clk), .Q(pc_out[30]) );
  DFQD1BWP12T pc_reg_29_ ( .D(n2230), .CP(clk), .Q(pc_out[29]) );
  DFQD1BWP12T pc_reg_28_ ( .D(n2229), .CP(clk), .Q(pc_out[28]) );
  DFQD1BWP12T pc_reg_27_ ( .D(n2228), .CP(clk), .Q(pc_out[27]) );
  DFQD1BWP12T pc_reg_26_ ( .D(n2227), .CP(clk), .Q(pc_out[26]) );
  DFQD1BWP12T pc_reg_25_ ( .D(n2226), .CP(clk), .Q(pc_out[25]) );
  DFQD1BWP12T pc_reg_24_ ( .D(n2225), .CP(clk), .Q(pc_out[24]) );
  DFQD1BWP12T pc_reg_23_ ( .D(n2224), .CP(clk), .Q(pc_out[23]) );
  DFQD1BWP12T pc_reg_22_ ( .D(n2223), .CP(clk), .Q(pc_out[22]) );
  DFQD1BWP12T pc_reg_21_ ( .D(n2222), .CP(clk), .Q(pc_out[21]) );
  DFQD1BWP12T pc_reg_20_ ( .D(n2221), .CP(clk), .Q(pc_out[20]) );
  DFQD1BWP12T pc_reg_19_ ( .D(n2220), .CP(clk), .Q(pc_out[19]) );
  DFQD1BWP12T pc_reg_18_ ( .D(n2219), .CP(clk), .Q(pc_out[18]) );
  DFQD1BWP12T pc_reg_17_ ( .D(n2218), .CP(clk), .Q(pc_out[17]) );
  DFQD1BWP12T pc_reg_16_ ( .D(n2217), .CP(clk), .Q(pc_out[16]) );
  DFQD1BWP12T pc_reg_14_ ( .D(n2215), .CP(clk), .Q(pc_out[14]) );
  DFQD1BWP12T pc_reg_13_ ( .D(n2214), .CP(clk), .Q(pc_out[13]) );
  DFQD1BWP12T pc_reg_12_ ( .D(n2213), .CP(clk), .Q(pc_out[12]) );
  DFQD1BWP12T pc_reg_11_ ( .D(n2212), .CP(clk), .Q(pc_out[11]) );
  DFQD1BWP12T pc_reg_10_ ( .D(n2211), .CP(clk), .Q(pc_out[10]) );
  DFQD1BWP12T pc_reg_9_ ( .D(n2210), .CP(clk), .Q(pc_out[9]) );
  DFQD1BWP12T pc_reg_8_ ( .D(n2209), .CP(clk), .Q(pc_out[8]) );
  DFQD1BWP12T pc_reg_7_ ( .D(n2208), .CP(clk), .Q(pc_out[7]) );
  DFQD1BWP12T pc_reg_6_ ( .D(n2207), .CP(clk), .Q(pc_out[6]) );
  DFQD1BWP12T pc_reg_5_ ( .D(n2206), .CP(clk), .Q(pc_out[5]) );
  DFQD1BWP12T pc_reg_4_ ( .D(n2205), .CP(clk), .Q(pc_out[4]) );
  DFQD1BWP12T pc_reg_3_ ( .D(n2204), .CP(clk), .Q(pc_out[3]) );
  DFQD1BWP12T pc_reg_2_ ( .D(n2203), .CP(clk), .Q(pc_out[2]) );
  DFQD1BWP12T pc_reg_1_ ( .D(n2202), .CP(clk), .Q(pc_out[1]) );
  DFQD1BWP12T pc_reg_0_ ( .D(n2201), .CP(clk), .Q(pc_out[0]) );
  DFQD1BWP12T cpsr_reg_3_ ( .D(next_cpsr_in[3]), .CP(clk), .Q(cpsr_out[3]) );
  DFQD1BWP12T cpsr_reg_2_ ( .D(next_cpsr_in[2]), .CP(clk), .Q(cpsr_out[2]) );
  DFQD1BWP12T cpsr_reg_1_ ( .D(next_cpsr_in[1]), .CP(clk), .Q(cpsr_out[1]) );
  DFQD1BWP12T cpsr_reg_0_ ( .D(next_cpsr_in[0]), .CP(clk), .Q(cpsr_out[0]) );
  DFQD1BWP12T tmp1_reg_31_ ( .D(n2200), .CP(clk), .Q(tmp1[31]) );
  DFQD1BWP12T tmp1_reg_30_ ( .D(n2199), .CP(clk), .Q(tmp1[30]) );
  DFQD1BWP12T tmp1_reg_29_ ( .D(n2198), .CP(clk), .Q(tmp1[29]) );
  DFQD1BWP12T tmp1_reg_28_ ( .D(n2197), .CP(clk), .Q(tmp1[28]) );
  DFQD1BWP12T tmp1_reg_27_ ( .D(n2196), .CP(clk), .Q(tmp1[27]) );
  DFQD1BWP12T tmp1_reg_26_ ( .D(n2195), .CP(clk), .Q(tmp1[26]) );
  DFQD1BWP12T tmp1_reg_25_ ( .D(n2194), .CP(clk), .Q(tmp1[25]) );
  DFQD1BWP12T tmp1_reg_24_ ( .D(n2193), .CP(clk), .Q(tmp1[24]) );
  DFQD1BWP12T tmp1_reg_23_ ( .D(n2192), .CP(clk), .Q(tmp1[23]) );
  DFQD1BWP12T tmp1_reg_22_ ( .D(n2191), .CP(clk), .Q(tmp1[22]) );
  DFQD1BWP12T tmp1_reg_21_ ( .D(n2190), .CP(clk), .Q(tmp1[21]) );
  DFQD1BWP12T tmp1_reg_20_ ( .D(n2189), .CP(clk), .Q(tmp1[20]) );
  DFQD1BWP12T tmp1_reg_19_ ( .D(n2188), .CP(clk), .Q(tmp1[19]) );
  DFQD1BWP12T tmp1_reg_18_ ( .D(n2187), .CP(clk), .Q(tmp1[18]) );
  DFQD1BWP12T tmp1_reg_17_ ( .D(n2186), .CP(clk), .Q(tmp1[17]) );
  DFQD1BWP12T tmp1_reg_16_ ( .D(n2185), .CP(clk), .Q(tmp1[16]) );
  DFQD1BWP12T tmp1_reg_15_ ( .D(n2184), .CP(clk), .Q(tmp1[15]) );
  DFQD1BWP12T tmp1_reg_14_ ( .D(n2183), .CP(clk), .Q(tmp1[14]) );
  DFQD1BWP12T tmp1_reg_13_ ( .D(n2182), .CP(clk), .Q(tmp1[13]) );
  DFQD1BWP12T tmp1_reg_12_ ( .D(n2181), .CP(clk), .Q(tmp1[12]) );
  DFQD1BWP12T tmp1_reg_11_ ( .D(n2180), .CP(clk), .Q(tmp1[11]) );
  DFQD1BWP12T tmp1_reg_10_ ( .D(n2179), .CP(clk), .Q(tmp1[10]) );
  DFQD1BWP12T tmp1_reg_9_ ( .D(n2178), .CP(clk), .Q(tmp1[9]) );
  DFQD1BWP12T tmp1_reg_8_ ( .D(n2177), .CP(clk), .Q(tmp1[8]) );
  DFQD1BWP12T tmp1_reg_7_ ( .D(n2176), .CP(clk), .Q(tmp1[7]) );
  DFQD1BWP12T tmp1_reg_6_ ( .D(n2175), .CP(clk), .Q(tmp1[6]) );
  DFQD1BWP12T tmp1_reg_5_ ( .D(n2174), .CP(clk), .Q(tmp1[5]) );
  DFQD1BWP12T tmp1_reg_4_ ( .D(n2173), .CP(clk), .Q(tmp1[4]) );
  DFQD1BWP12T tmp1_reg_3_ ( .D(n2172), .CP(clk), .Q(tmp1[3]) );
  DFQD1BWP12T tmp1_reg_2_ ( .D(n2171), .CP(clk), .Q(tmp1[2]) );
  DFQD1BWP12T tmp1_reg_1_ ( .D(n2170), .CP(clk), .Q(tmp1[1]) );
  DFQD1BWP12T tmp1_reg_0_ ( .D(n2169), .CP(clk), .Q(tmp1[0]) );
  DFKCNXD1BWP12T pc_reg_15_ ( .CN(n4887), .D(n4888), .CP(clk), .Q(n4886), .QN(
        pc_out[15]) );
  ND2D1BWP12T U2843 ( .A1(write2_sel[2]), .A2(write2_sel[3]), .ZN(n4679) );
  INVD1BWP12T U2844 ( .I(write2_sel[2]), .ZN(n3124) );
  INVD1BWP12T U2845 ( .I(write2_sel[0]), .ZN(n3133) );
  INR3D0BWP12T U2846 ( .A1(write2_en), .B1(write2_sel[1]), .B2(write2_sel[4]), 
        .ZN(n3134) );
  INVD1BWP12T U2847 ( .I(write2_sel[3]), .ZN(n3147) );
  IND2D1BWP12T U2848 ( .A1(write1_sel[4]), .B1(write1_en), .ZN(n3125) );
  ND2D1BWP12T U2849 ( .A1(n3134), .A2(n3133), .ZN(n4762) );
  ND2D1BWP12T U2850 ( .A1(n3124), .A2(n3147), .ZN(n4756) );
  INVD1BWP12T U2851 ( .I(write1_sel[0]), .ZN(n3142) );
  IND4D1BWP12T U2852 ( .A1(n4679), .B1(write2_sel[1]), .B2(write2_en), .B3(
        n3133), .ZN(n3146) );
  INVD1BWP12T U2853 ( .I(write2_sel[4]), .ZN(n3145) );
  NR2D1BWP12T U2854 ( .A1(write2_sel[4]), .A2(n3146), .ZN(n3132) );
  NR2D1BWP12T U2855 ( .A1(n4679), .A2(n4762), .ZN(n3138) );
  ND4D1BWP12T U2856 ( .A1(write2_sel[0]), .A2(write2_sel[1]), .A3(write2_en), 
        .A4(n3145), .ZN(n4752) );
  NR2D1BWP12T U2857 ( .A1(n3142), .A2(n3128), .ZN(n4678) );
  ND2D1BWP12T U2858 ( .A1(write2_sel[3]), .A2(n3124), .ZN(n3135) );
  NR2D1BWP12T U2859 ( .A1(n4762), .A2(n3135), .ZN(n3136) );
  NR2D1BWP12T U2860 ( .A1(n4752), .A2(n4761), .ZN(n4754) );
  ND4D1BWP12T U2861 ( .A1(write2_sel[1]), .A2(write2_en), .A3(n3133), .A4(
        n3145), .ZN(n3149) );
  ND2D1BWP12T U2862 ( .A1(write2_sel[0]), .A2(n3134), .ZN(n4757) );
  ND2D1BWP12T U2863 ( .A1(write2_sel[2]), .A2(n3147), .ZN(n4761) );
  INR2D1BWP12T U2864 ( .A1(write1_sel[2]), .B1(write1_sel[1]), .ZN(n4764) );
  NR2D1BWP12T U2865 ( .A1(n4762), .A2(n4761), .ZN(n4765) );
  NR2D1BWP12T U2866 ( .A1(n4756), .A2(n3149), .ZN(n3126) );
  NR3D1BWP12T U2867 ( .A1(write1_sel[3]), .A2(n3142), .A3(n3125), .ZN(n4758)
         );
  NR2D1BWP12T U2868 ( .A1(n4757), .A2(n4756), .ZN(n4760) );
  NR3D1BWP12T U2869 ( .A1(write1_sel[0]), .A2(write1_sel[3]), .A3(n3125), .ZN(
        n4763) );
  NR2D1BWP12T U2870 ( .A1(write1_sel[1]), .A2(write1_sel[2]), .ZN(n4759) );
  NR2D1BWP12T U2871 ( .A1(n4762), .A2(n4756), .ZN(n4755) );
  INVD1BWP12T U2872 ( .I(n4601), .ZN(n4653) );
  ND2D1BWP12T U2873 ( .A1(write1_en), .A2(n3143), .ZN(n4751) );
  OAI21D1BWP12T U2874 ( .A1(n3146), .A2(n3145), .B(n4751), .ZN(n4750) );
  ND2D1BWP12T U2875 ( .A1(n3144), .A2(n4751), .ZN(n4749) );
  NR2D1BWP12T U2876 ( .A1(n3145), .A2(n3146), .ZN(n3144) );
  NR2D1BWP12T U2877 ( .A1(n4742), .A2(n4682), .ZN(n4741) );
  INVD1BWP12T U2878 ( .I(n4681), .ZN(n4742) );
  NR2D1BWP12T U2879 ( .A1(next_pc_en), .A2(n4680), .ZN(n4744) );
  INR2D1BWP12T U2880 ( .A1(next_pc_en), .B1(n4680), .ZN(n4743) );
  INVD1BWP12T U2881 ( .I(lr[2]), .ZN(n3850) );
  INVD1BWP12T U2882 ( .I(lr[4]), .ZN(n4330) );
  INVD1BWP12T U2883 ( .I(lr[8]), .ZN(n4377) );
  INVD1BWP12T U2884 ( .I(lr[9]), .ZN(n4827) );
  INVD1BWP12T U2885 ( .I(lr[11]), .ZN(n4870) );
  INVD1BWP12T U2886 ( .I(lr[12]), .ZN(n4851) );
  INVD1BWP12T U2887 ( .I(lr[13]), .ZN(n4857) );
  INVD1BWP12T U2888 ( .I(lr[14]), .ZN(n4243) );
  INVD1BWP12T U2889 ( .I(lr[18]), .ZN(n4504) );
  INVD1BWP12T U2890 ( .I(lr[19]), .ZN(n4516) );
  INVD1BWP12T U2891 ( .I(lr[26]), .ZN(n4602) );
  ND2D1BWP12T U2892 ( .A1(n4753), .A2(n3137), .ZN(n4873) );
  ND2D1BWP12T U2893 ( .A1(n3132), .A2(n4873), .ZN(n4869) );
  INVD1BWP12T U2894 ( .I(r12[0]), .ZN(n4860) );
  INVD1BWP12T U2895 ( .I(r12[2]), .ZN(n4864) );
  INVD1BWP12T U2896 ( .I(r12[6]), .ZN(n4163) );
  INVD1BWP12T U2897 ( .I(r12[15]), .ZN(n4830) );
  ND2D1BWP12T U2898 ( .A1(n4764), .A2(n3137), .ZN(n4867) );
  ND2D1BWP12T U2899 ( .A1(n3138), .A2(n4867), .ZN(n4863) );
  ND2D1BWP12T U2900 ( .A1(n4678), .A2(n3129), .ZN(n3141) );
  OAI21D1BWP12T U2901 ( .A1(n3135), .A2(n4752), .B(n3141), .ZN(n3140) );
  ND2D1BWP12T U2902 ( .A1(n3123), .A2(n3141), .ZN(n3139) );
  NR2D1BWP12T U2903 ( .A1(n4752), .A2(n3135), .ZN(n3123) );
  ND2D1BWP12T U2904 ( .A1(n3129), .A2(n3137), .ZN(n4813) );
  OAI21D1BWP12T U2905 ( .A1(n3135), .A2(n3149), .B(n4813), .ZN(n4814) );
  ND2D1BWP12T U2906 ( .A1(n3130), .A2(n4813), .ZN(n4816) );
  ND2D1BWP12T U2907 ( .A1(n4678), .A2(n4759), .ZN(n4797) );
  OAI21D1BWP12T U2908 ( .A1(n3135), .A2(n4757), .B(n4797), .ZN(n4796) );
  ND2D1BWP12T U2909 ( .A1(n3131), .A2(n4797), .ZN(n4795) );
  NR2D1BWP12T U2910 ( .A1(n4757), .A2(n3135), .ZN(n3131) );
  INVD1BWP12T U2911 ( .I(r8[10]), .ZN(n4401) );
  INVD1BWP12T U2912 ( .I(r8[17]), .ZN(n4492) );
  INVD1BWP12T U2913 ( .I(r8[27]), .ZN(n4614) );
  INVD1BWP12T U2914 ( .I(r8[29]), .ZN(n4824) );
  ND2D1BWP12T U2915 ( .A1(n4759), .A2(n3137), .ZN(n4823) );
  ND2D1BWP12T U2916 ( .A1(n3136), .A2(n4823), .ZN(n4826) );
  ND2D1BWP12T U2917 ( .A1(n4753), .A2(n4758), .ZN(n4771) );
  ND2D1BWP12T U2918 ( .A1(n4754), .A2(n4771), .ZN(n4769) );
  ND2D1BWP12T U2919 ( .A1(n4753), .A2(n4763), .ZN(n4817) );
  OAI21D1BWP12T U2920 ( .A1(n4761), .A2(n3149), .B(n4817), .ZN(n4818) );
  ND2D1BWP12T U2921 ( .A1(n3148), .A2(n4817), .ZN(n4819) );
  NR2D1BWP12T U2922 ( .A1(n3149), .A2(n4761), .ZN(n3148) );
  ND2D1BWP12T U2923 ( .A1(n4764), .A2(n4758), .ZN(n4822) );
  OAI21D1BWP12T U2924 ( .A1(n4761), .A2(n4757), .B(n4822), .ZN(n4821) );
  ND2D1BWP12T U2925 ( .A1(n3152), .A2(n4822), .ZN(n4820) );
  NR2D1BWP12T U2926 ( .A1(n4757), .A2(n4761), .ZN(n3152) );
  ND2D1BWP12T U2927 ( .A1(n4764), .A2(n4763), .ZN(n4768) );
  ND2D1BWP12T U2928 ( .A1(n4765), .A2(n4768), .ZN(n4766) );
  INVD1BWP12T U2929 ( .I(r3[2]), .ZN(n4207) );
  INVD1BWP12T U2930 ( .I(r3[21]), .ZN(n3652) );
  INVD1BWP12T U2931 ( .I(r3[24]), .ZN(n3978) );
  ND2D1BWP12T U2932 ( .A1(n4758), .A2(n3129), .ZN(n4774) );
  ND2D1BWP12T U2933 ( .A1(n3127), .A2(n4774), .ZN(n4773) );
  ND2D1BWP12T U2934 ( .A1(n3126), .A2(n4774), .ZN(n4772) );
  INVD1BWP12T U2935 ( .I(r2[3]), .ZN(n3838) );
  INVD1BWP12T U2936 ( .I(r2[13]), .ZN(n4092) );
  INVD1BWP12T U2937 ( .I(r2[20]), .ZN(n4882) );
  INVD1BWP12T U2938 ( .I(r2[22]), .ZN(n4000) );
  INVD1BWP12T U2939 ( .I(r2[26]), .ZN(n3600) );
  ND2D1BWP12T U2940 ( .A1(n4763), .A2(n3129), .ZN(n4885) );
  ND2D1BWP12T U2941 ( .A1(n3127), .A2(n4885), .ZN(n4883) );
  ND2D1BWP12T U2942 ( .A1(n3126), .A2(n4885), .ZN(n4881) );
  INVD1BWP12T U2943 ( .I(r1[24]), .ZN(n4843) );
  INVD1BWP12T U2944 ( .I(r1[29]), .ZN(n4836) );
  ND2D1BWP12T U2945 ( .A1(n4759), .A2(n4758), .ZN(n4842) );
  ND2D1BWP12T U2946 ( .A1(n4760), .A2(n4842), .ZN(n4846) );
  INVD1BWP12T U2947 ( .I(write2_in[0]), .ZN(n4859) );
  INVD1BWP12T U2948 ( .I(write1_in[0]), .ZN(n4861) );
  INVD1BWP12T U2949 ( .I(write1_in[1]), .ZN(n4783) );
  INVD1BWP12T U2950 ( .I(write2_in[1]), .ZN(n4784) );
  INVD1BWP12T U2951 ( .I(write2_in[2]), .ZN(n4862) );
  INVD1BWP12T U2952 ( .I(write1_in[2]), .ZN(n4866) );
  INVD1BWP12T U2953 ( .I(write1_in[3]), .ZN(n4793) );
  INVD1BWP12T U2954 ( .I(write2_in[3]), .ZN(n4794) );
  INVD1BWP12T U2955 ( .I(write1_in[4]), .ZN(n4800) );
  INVD1BWP12T U2956 ( .I(write2_in[4]), .ZN(n4801) );
  INVD1BWP12T U2957 ( .I(r0[5]), .ZN(n4839) );
  INVD1BWP12T U2958 ( .I(write1_in[5]), .ZN(n4838) );
  INVD1BWP12T U2959 ( .I(write2_in[5]), .ZN(n4840) );
  INVD1BWP12T U2960 ( .I(write1_in[6]), .ZN(n4779) );
  INVD1BWP12T U2961 ( .I(write2_in[6]), .ZN(n4780) );
  INVD1BWP12T U2962 ( .I(write2_in[7]), .ZN(n4798) );
  INVD1BWP12T U2963 ( .I(write1_in[7]), .ZN(n4799) );
  INVD1BWP12T U2964 ( .I(write1_in[8]), .ZN(n4810) );
  INVD1BWP12T U2965 ( .I(write2_in[8]), .ZN(n4811) );
  INVD1BWP12T U2966 ( .I(r0[9]), .ZN(n4854) );
  INVD1BWP12T U2967 ( .I(write1_in[9]), .ZN(n4853) );
  INVD1BWP12T U2968 ( .I(write2_in[9]), .ZN(n4855) );
  INVD1BWP12T U2969 ( .I(write2_in[10]), .ZN(n4808) );
  INVD1BWP12T U2970 ( .I(write1_in[10]), .ZN(n4809) );
  INVD1BWP12T U2971 ( .I(write2_in[11]), .ZN(n4868) );
  INVD1BWP12T U2972 ( .I(write1_in[11]), .ZN(n4872) );
  INVD1BWP12T U2973 ( .I(write1_in[12]), .ZN(n4850) );
  INVD1BWP12T U2974 ( .I(write2_in[12]), .ZN(n4852) );
  INVD1BWP12T U2975 ( .I(write1_in[13]), .ZN(n4856) );
  INVD1BWP12T U2976 ( .I(write2_in[13]), .ZN(n4858) );
  INVD1BWP12T U2977 ( .I(write2_in[14]), .ZN(n4802) );
  INVD1BWP12T U2978 ( .I(write1_in[14]), .ZN(n4803) );
  INVD1BWP12T U2979 ( .I(r0[15]), .ZN(n4828) );
  INVD1BWP12T U2980 ( .I(write1_in[15]), .ZN(n4829) );
  INVD1BWP12T U2981 ( .I(write2_in[15]), .ZN(n4831) );
  INVD1BWP12T U2982 ( .I(r0[16]), .ZN(n4876) );
  INVD1BWP12T U2983 ( .I(write2_in[16]), .ZN(n4874) );
  INVD1BWP12T U2984 ( .I(write1_in[16]), .ZN(n4878) );
  INVD1BWP12T U2985 ( .I(write1_in[17]), .ZN(n4812) );
  INVD1BWP12T U2986 ( .I(write2_in[17]), .ZN(n4815) );
  INVD1BWP12T U2987 ( .I(write2_in[18]), .ZN(n4791) );
  INVD1BWP12T U2988 ( .I(write1_in[18]), .ZN(n4792) );
  INVD1BWP12T U2989 ( .I(write2_in[19]), .ZN(n4781) );
  INVD1BWP12T U2990 ( .I(write1_in[19]), .ZN(n4782) );
  INVD1BWP12T U2991 ( .I(write2_in[20]), .ZN(n4880) );
  INVD1BWP12T U2992 ( .I(write1_in[20]), .ZN(n4884) );
  INVD1BWP12T U2993 ( .I(write1_in[21]), .ZN(n4777) );
  INVD1BWP12T U2994 ( .I(write2_in[21]), .ZN(n4778) );
  INVD1BWP12T U2995 ( .I(write1_in[22]), .ZN(n4785) );
  INVD1BWP12T U2996 ( .I(write2_in[22]), .ZN(n4786) );
  INVD1BWP12T U2997 ( .I(r0[23]), .ZN(n4833) );
  INVD1BWP12T U2998 ( .I(write1_in[23]), .ZN(n4832) );
  INVD1BWP12T U2999 ( .I(write2_in[23]), .ZN(n4834) );
  INVD1BWP12T U3000 ( .I(write1_in[24]), .ZN(n4841) );
  INVD1BWP12T U3001 ( .I(write2_in[24]), .ZN(n4845) );
  INVD1BWP12T U3002 ( .I(write2_in[25]), .ZN(n4804) );
  INVD1BWP12T U3003 ( .I(write1_in[25]), .ZN(n4805) );
  INVD1BWP12T U3004 ( .I(write1_in[26]), .ZN(n4775) );
  INVD1BWP12T U3005 ( .I(write2_in[26]), .ZN(n4776) );
  INVD1BWP12T U3006 ( .I(write1_in[27]), .ZN(n4787) );
  INVD1BWP12T U3007 ( .I(write2_in[27]), .ZN(n4788) );
  INVD1BWP12T U3008 ( .I(write1_in[28]), .ZN(n4806) );
  INVD1BWP12T U3009 ( .I(write2_in[28]), .ZN(n4807) );
  INVD1BWP12T U3010 ( .I(write1_in[29]), .ZN(n4835) );
  INVD1BWP12T U3011 ( .I(write2_in[29]), .ZN(n4837) );
  INVD1BWP12T U3012 ( .I(write2_in[30]), .ZN(n4789) );
  INVD1BWP12T U3013 ( .I(write1_in[30]), .ZN(n4790) );
  INVD1BWP12T U3014 ( .I(r0[31]), .ZN(n4848) );
  ND2D1BWP12T U3015 ( .A1(n4759), .A2(n4763), .ZN(n4879) );
  ND2D1BWP12T U3016 ( .A1(n4755), .A2(n4879), .ZN(n4875) );
  INVD1BWP12T U3017 ( .I(write1_in[31]), .ZN(n4847) );
  INVD1BWP12T U3018 ( .I(write2_in[31]), .ZN(n4849) );
  OAI222D1BWP12T U3019 ( .A1(n4749), .A2(n4784), .B1(n4750), .B2(n3151), .C1(
        n4751), .C2(n4783), .ZN(n2170) );
  INVD1BWP12T U3020 ( .I(tmp1[1]), .ZN(n3151) );
  OAI222D1BWP12T U3021 ( .A1(n4751), .A2(n4799), .B1(n4750), .B2(n3153), .C1(
        n4749), .C2(n4798), .ZN(n2176) );
  INVD1BWP12T U3022 ( .I(tmp1[7]), .ZN(n3153) );
  INVD1BWP12T U3023 ( .I(tmp1[25]), .ZN(n4748) );
  OAI222D1BWP12T U3024 ( .A1(n4749), .A2(n4807), .B1(n4750), .B2(n3150), .C1(
        n4751), .C2(n4806), .ZN(n2197) );
  INVD1BWP12T U3025 ( .I(tmp1[28]), .ZN(n3150) );
  INVD1BWP12T U3026 ( .I(tmp1[30]), .ZN(n4747) );
  OAI222D1BWP12T U3027 ( .A1(n4873), .A2(n4866), .B1(n4871), .B2(n3850), .C1(
        n4869), .C2(n4862), .ZN(n2235) );
  OAI222D1BWP12T U3028 ( .A1(n4869), .A2(n4801), .B1(n4871), .B2(n4330), .C1(
        n4873), .C2(n4800), .ZN(n2237) );
  OAI222D1BWP12T U3029 ( .A1(n4869), .A2(n4811), .B1(n4871), .B2(n4377), .C1(
        n4873), .C2(n4810), .ZN(n2241) );
  OAI222D1BWP12T U3030 ( .A1(n4873), .A2(n4803), .B1(n4871), .B2(n4243), .C1(
        n4869), .C2(n4802), .ZN(n2247) );
  OAI222D1BWP12T U3031 ( .A1(n4873), .A2(n4792), .B1(n4871), .B2(n4504), .C1(
        n4869), .C2(n4791), .ZN(n2251) );
  OAI222D1BWP12T U3032 ( .A1(n4873), .A2(n4782), .B1(n4871), .B2(n4516), .C1(
        n4869), .C2(n4781), .ZN(n2252) );
  OAI222D1BWP12T U3033 ( .A1(n4869), .A2(n4776), .B1(n4871), .B2(n4602), .C1(
        n4873), .C2(n4775), .ZN(n2259) );
  OAI222D1BWP12T U3034 ( .A1(n4863), .A2(n4780), .B1(n4865), .B2(n4163), .C1(
        n4867), .C2(n4779), .ZN(n2271) );
  OAI222D1BWP12T U3035 ( .A1(n4823), .A2(n4809), .B1(n4825), .B2(n4401), .C1(
        n4826), .C2(n4808), .ZN(n2403) );
  OAI222D1BWP12T U3036 ( .A1(n4826), .A2(n4815), .B1(n4825), .B2(n4492), .C1(
        n4823), .C2(n4812), .ZN(n2410) );
  OAI222D1BWP12T U3037 ( .A1(n4826), .A2(n4788), .B1(n4825), .B2(n4614), .C1(
        n4823), .C2(n4787), .ZN(n2420) );
  OAI222D1BWP12T U3038 ( .A1(n4774), .A2(n4866), .B1(n4773), .B2(n4207), .C1(
        n4772), .C2(n4862), .ZN(n2555) );
  OAI222D1BWP12T U3039 ( .A1(n4772), .A2(n4778), .B1(n4773), .B2(n3652), .C1(
        n4774), .C2(n4777), .ZN(n2574) );
  OAI222D1BWP12T U3040 ( .A1(n4772), .A2(n4845), .B1(n4773), .B2(n3978), .C1(
        n4774), .C2(n4841), .ZN(n2577) );
  OAI222D1BWP12T U3041 ( .A1(n4881), .A2(n4794), .B1(n4883), .B2(n3838), .C1(
        n4885), .C2(n4793), .ZN(n2588) );
  OAI222D1BWP12T U3042 ( .A1(n4881), .A2(n4858), .B1(n4883), .B2(n4092), .C1(
        n4885), .C2(n4856), .ZN(n2598) );
  OAI222D1BWP12T U3043 ( .A1(n4881), .A2(n4786), .B1(n4883), .B2(n4000), .C1(
        n4885), .C2(n4785), .ZN(n2607) );
  OAI222D1BWP12T U3044 ( .A1(n4881), .A2(n4776), .B1(n4883), .B2(n3600), .C1(
        n4885), .C2(n4775), .ZN(n2611) );
  CKND0BWP12T U3045 ( .I(tmp1[0]), .ZN(n2681) );
  OAI222D0BWP12T U3046 ( .A1(n2681), .A2(n4750), .B1(n4749), .B2(n4859), .C1(
        n4861), .C2(n4751), .ZN(n2169) );
  CKND0BWP12T U3047 ( .I(tmp1[3]), .ZN(n2682) );
  OAI222D0BWP12T U3048 ( .A1(n2682), .A2(n4750), .B1(n4751), .B2(n4793), .C1(
        n4794), .C2(n4749), .ZN(n2172) );
  CKND0BWP12T U3049 ( .I(tmp1[4]), .ZN(n2683) );
  OAI222D0BWP12T U3050 ( .A1(n2683), .A2(n4750), .B1(n4751), .B2(n4800), .C1(
        n4801), .C2(n4749), .ZN(n2173) );
  CKND0BWP12T U3051 ( .I(tmp1[5]), .ZN(n2684) );
  OAI222D0BWP12T U3052 ( .A1(n2684), .A2(n4750), .B1(n4751), .B2(n4838), .C1(
        n4840), .C2(n4749), .ZN(n2174) );
  CKND0BWP12T U3053 ( .I(tmp1[6]), .ZN(n2685) );
  OAI222D0BWP12T U3054 ( .A1(n2685), .A2(n4750), .B1(n4751), .B2(n4779), .C1(
        n4780), .C2(n4749), .ZN(n2175) );
  CKND0BWP12T U3055 ( .I(tmp1[8]), .ZN(n2686) );
  OAI222D0BWP12T U3056 ( .A1(n2686), .A2(n4750), .B1(n4751), .B2(n4810), .C1(
        n4811), .C2(n4749), .ZN(n2177) );
  CKND0BWP12T U3057 ( .I(tmp1[10]), .ZN(n2687) );
  OAI222D0BWP12T U3058 ( .A1(n2687), .A2(n4750), .B1(n4749), .B2(n4808), .C1(
        n4809), .C2(n4751), .ZN(n2179) );
  CKND0BWP12T U3059 ( .I(tmp1[11]), .ZN(n2688) );
  OAI222D0BWP12T U3060 ( .A1(n2688), .A2(n4750), .B1(n4749), .B2(n4868), .C1(
        n4872), .C2(n4751), .ZN(n2180) );
  CKND0BWP12T U3061 ( .I(tmp1[12]), .ZN(n2689) );
  OAI222D0BWP12T U3062 ( .A1(n2689), .A2(n4750), .B1(n4751), .B2(n4850), .C1(
        n4852), .C2(n4749), .ZN(n2181) );
  CKND0BWP12T U3063 ( .I(tmp1[14]), .ZN(n2690) );
  OAI222D0BWP12T U3064 ( .A1(n2690), .A2(n4750), .B1(n4749), .B2(n4802), .C1(
        n4803), .C2(n4751), .ZN(n2183) );
  CKND0BWP12T U3065 ( .I(tmp1[16]), .ZN(n2691) );
  OAI222D0BWP12T U3066 ( .A1(n2691), .A2(n4750), .B1(n4749), .B2(n4874), .C1(
        n4878), .C2(n4751), .ZN(n2185) );
  CKND0BWP12T U3067 ( .I(tmp1[17]), .ZN(n2692) );
  OAI222D0BWP12T U3068 ( .A1(n2692), .A2(n4750), .B1(n4751), .B2(n4812), .C1(
        n4815), .C2(n4749), .ZN(n2186) );
  CKND0BWP12T U3069 ( .I(tmp1[18]), .ZN(n2693) );
  OAI222D0BWP12T U3070 ( .A1(n2693), .A2(n4750), .B1(n4749), .B2(n4791), .C1(
        n4792), .C2(n4751), .ZN(n2187) );
  CKND0BWP12T U3071 ( .I(tmp1[19]), .ZN(n2694) );
  OAI222D0BWP12T U3072 ( .A1(n2694), .A2(n4750), .B1(n4749), .B2(n4781), .C1(
        n4782), .C2(n4751), .ZN(n2188) );
  CKND0BWP12T U3073 ( .I(tmp1[20]), .ZN(n2695) );
  OAI222D0BWP12T U3074 ( .A1(n2695), .A2(n4750), .B1(n4749), .B2(n4880), .C1(
        n4884), .C2(n4751), .ZN(n2189) );
  CKND0BWP12T U3075 ( .I(tmp1[21]), .ZN(n2696) );
  OAI222D0BWP12T U3076 ( .A1(n2696), .A2(n4750), .B1(n4751), .B2(n4777), .C1(
        n4778), .C2(n4749), .ZN(n2190) );
  CKND0BWP12T U3077 ( .I(tmp1[22]), .ZN(n2697) );
  OAI222D0BWP12T U3078 ( .A1(n2697), .A2(n4750), .B1(n4751), .B2(n4785), .C1(
        n4786), .C2(n4749), .ZN(n2191) );
  CKND0BWP12T U3079 ( .I(tmp1[23]), .ZN(n2698) );
  OAI222D0BWP12T U3080 ( .A1(n2698), .A2(n4750), .B1(n4751), .B2(n4832), .C1(
        n4834), .C2(n4749), .ZN(n2192) );
  CKND0BWP12T U3081 ( .I(tmp1[27]), .ZN(n2699) );
  OAI222D0BWP12T U3082 ( .A1(n2699), .A2(n4750), .B1(n4751), .B2(n4787), .C1(
        n4788), .C2(n4749), .ZN(n2196) );
  CKND0BWP12T U3083 ( .I(tmp1[31]), .ZN(n2700) );
  OAI222D0BWP12T U3084 ( .A1(n2700), .A2(n4750), .B1(n4751), .B2(n4847), .C1(
        n4849), .C2(n4749), .ZN(n2200) );
  CKND0BWP12T U3085 ( .I(lr[1]), .ZN(n2701) );
  OAI222D0BWP12T U3086 ( .A1(n2701), .A2(n4871), .B1(n4873), .B2(n4783), .C1(
        n4784), .C2(n4869), .ZN(n2234) );
  CKND0BWP12T U3087 ( .I(lr[7]), .ZN(n2702) );
  OAI222D0BWP12T U3088 ( .A1(n2702), .A2(n4871), .B1(n4869), .B2(n4798), .C1(
        n4799), .C2(n4873), .ZN(n2240) );
  CKND0BWP12T U3089 ( .I(lr[25]), .ZN(n2703) );
  OAI222D0BWP12T U3090 ( .A1(n2703), .A2(n4871), .B1(n4869), .B2(n4804), .C1(
        n4805), .C2(n4873), .ZN(n2258) );
  CKND0BWP12T U3091 ( .I(lr[28]), .ZN(n2704) );
  OAI222D0BWP12T U3092 ( .A1(n2704), .A2(n4871), .B1(n4873), .B2(n4806), .C1(
        n4807), .C2(n4869), .ZN(n2261) );
  CKND0BWP12T U3093 ( .I(lr[30]), .ZN(n2705) );
  OAI222D0BWP12T U3094 ( .A1(n2705), .A2(n4871), .B1(n4869), .B2(n4789), .C1(
        n4790), .C2(n4873), .ZN(n2263) );
  CKND0BWP12T U3095 ( .I(tmp1[9]), .ZN(n2706) );
  OAI222D0BWP12T U3096 ( .A1(n2706), .A2(n4750), .B1(n4751), .B2(n4853), .C1(
        n4855), .C2(n4749), .ZN(n2178) );
  CKND0BWP12T U3097 ( .I(tmp1[13]), .ZN(n2707) );
  OAI222D0BWP12T U3098 ( .A1(n2707), .A2(n4750), .B1(n4751), .B2(n4856), .C1(
        n4858), .C2(n4749), .ZN(n2182) );
  CKND0BWP12T U3099 ( .I(tmp1[15]), .ZN(n2708) );
  OAI222D0BWP12T U3100 ( .A1(n2708), .A2(n4750), .B1(n4751), .B2(n4829), .C1(
        n4831), .C2(n4749), .ZN(n2184) );
  CKND0BWP12T U3101 ( .I(tmp1[24]), .ZN(n2709) );
  OAI222D0BWP12T U3102 ( .A1(n2709), .A2(n4750), .B1(n4751), .B2(n4841), .C1(
        n4845), .C2(n4749), .ZN(n2193) );
  CKND0BWP12T U3103 ( .I(tmp1[26]), .ZN(n2710) );
  OAI222D0BWP12T U3104 ( .A1(n2710), .A2(n4750), .B1(n4751), .B2(n4775), .C1(
        n4776), .C2(n4749), .ZN(n2195) );
  CKND0BWP12T U3105 ( .I(tmp1[29]), .ZN(n2711) );
  OAI222D0BWP12T U3106 ( .A1(n2711), .A2(n4750), .B1(n4751), .B2(n4835), .C1(
        n4837), .C2(n4749), .ZN(n2198) );
  CKND0BWP12T U3107 ( .I(lr[0]), .ZN(n2712) );
  OAI222D0BWP12T U3108 ( .A1(n2712), .A2(n4871), .B1(n4869), .B2(n4859), .C1(
        n4861), .C2(n4873), .ZN(n2233) );
  CKND0BWP12T U3109 ( .I(lr[3]), .ZN(n2713) );
  OAI222D0BWP12T U3110 ( .A1(n2713), .A2(n4871), .B1(n4873), .B2(n4793), .C1(
        n4794), .C2(n4869), .ZN(n2236) );
  CKND0BWP12T U3111 ( .I(lr[5]), .ZN(n2714) );
  OAI222D0BWP12T U3112 ( .A1(n2714), .A2(n4871), .B1(n4873), .B2(n4838), .C1(
        n4840), .C2(n4869), .ZN(n2238) );
  CKND0BWP12T U3113 ( .I(lr[6]), .ZN(n2715) );
  OAI222D0BWP12T U3114 ( .A1(n2715), .A2(n4871), .B1(n4873), .B2(n4779), .C1(
        n4780), .C2(n4869), .ZN(n2239) );
  CKND0BWP12T U3115 ( .I(lr[10]), .ZN(n2716) );
  OAI222D0BWP12T U3116 ( .A1(n2716), .A2(n4871), .B1(n4869), .B2(n4808), .C1(
        n4809), .C2(n4873), .ZN(n2243) );
  CKND0BWP12T U3117 ( .I(lr[16]), .ZN(n2717) );
  OAI222D0BWP12T U3118 ( .A1(n2717), .A2(n4871), .B1(n4869), .B2(n4874), .C1(
        n4878), .C2(n4873), .ZN(n2249) );
  CKND0BWP12T U3119 ( .I(lr[17]), .ZN(n2718) );
  OAI222D0BWP12T U3120 ( .A1(n2718), .A2(n4871), .B1(n4873), .B2(n4812), .C1(
        n4815), .C2(n4869), .ZN(n2250) );
  CKND0BWP12T U3121 ( .I(lr[20]), .ZN(n2719) );
  OAI222D0BWP12T U3122 ( .A1(n2719), .A2(n4871), .B1(n4869), .B2(n4880), .C1(
        n4884), .C2(n4873), .ZN(n2253) );
  CKND0BWP12T U3123 ( .I(lr[21]), .ZN(n2720) );
  OAI222D0BWP12T U3124 ( .A1(n2720), .A2(n4871), .B1(n4873), .B2(n4777), .C1(
        n4778), .C2(n4869), .ZN(n2254) );
  CKND0BWP12T U3125 ( .I(lr[22]), .ZN(n2721) );
  OAI222D0BWP12T U3126 ( .A1(n2721), .A2(n4871), .B1(n4873), .B2(n4785), .C1(
        n4786), .C2(n4869), .ZN(n2255) );
  CKND0BWP12T U3127 ( .I(lr[23]), .ZN(n2722) );
  OAI222D0BWP12T U3128 ( .A1(n2722), .A2(n4871), .B1(n4873), .B2(n4832), .C1(
        n4834), .C2(n4869), .ZN(n2256) );
  CKND0BWP12T U3129 ( .I(lr[27]), .ZN(n2723) );
  OAI222D0BWP12T U3130 ( .A1(n2723), .A2(n4871), .B1(n4873), .B2(n4787), .C1(
        n4788), .C2(n4869), .ZN(n2260) );
  CKND0BWP12T U3131 ( .I(lr[31]), .ZN(n2724) );
  OAI222D0BWP12T U3132 ( .A1(n2724), .A2(n4871), .B1(n4873), .B2(n4847), .C1(
        n4849), .C2(n4869), .ZN(n2264) );
  CKND0BWP12T U3133 ( .I(r12[1]), .ZN(n2725) );
  OAI222D0BWP12T U3134 ( .A1(n2725), .A2(n4865), .B1(n4867), .B2(n4783), .C1(
        n4784), .C2(n4863), .ZN(n2266) );
  CKND0BWP12T U3135 ( .I(r12[4]), .ZN(n2726) );
  OAI222D0BWP12T U3136 ( .A1(n2726), .A2(n4865), .B1(n4867), .B2(n4800), .C1(
        n4801), .C2(n4863), .ZN(n2269) );
  CKND0BWP12T U3137 ( .I(r12[7]), .ZN(n2727) );
  OAI222D0BWP12T U3138 ( .A1(n2727), .A2(n4865), .B1(n4863), .B2(n4798), .C1(
        n4799), .C2(n4867), .ZN(n2272) );
  CKND0BWP12T U3139 ( .I(r12[8]), .ZN(n2728) );
  OAI222D0BWP12T U3140 ( .A1(n2728), .A2(n4865), .B1(n4867), .B2(n4810), .C1(
        n4811), .C2(n4863), .ZN(n2273) );
  CKND0BWP12T U3141 ( .I(r12[11]), .ZN(n2729) );
  OAI222D0BWP12T U3142 ( .A1(n2729), .A2(n4865), .B1(n4863), .B2(n4868), .C1(
        n4872), .C2(n4867), .ZN(n2276) );
  CKND0BWP12T U3143 ( .I(r12[12]), .ZN(n2730) );
  OAI222D0BWP12T U3144 ( .A1(n2730), .A2(n4865), .B1(n4867), .B2(n4850), .C1(
        n4852), .C2(n4863), .ZN(n2277) );
  CKND0BWP12T U3145 ( .I(r12[14]), .ZN(n2731) );
  OAI222D0BWP12T U3146 ( .A1(n2731), .A2(n4865), .B1(n4863), .B2(n4802), .C1(
        n4803), .C2(n4867), .ZN(n2279) );
  CKND0BWP12T U3147 ( .I(r12[18]), .ZN(n2732) );
  OAI222D0BWP12T U3148 ( .A1(n2732), .A2(n4865), .B1(n4863), .B2(n4791), .C1(
        n4792), .C2(n4867), .ZN(n2283) );
  CKND0BWP12T U3149 ( .I(r12[19]), .ZN(n2733) );
  OAI222D0BWP12T U3150 ( .A1(n2733), .A2(n4865), .B1(n4863), .B2(n4781), .C1(
        n4782), .C2(n4867), .ZN(n2284) );
  CKND0BWP12T U3151 ( .I(r12[25]), .ZN(n2734) );
  OAI222D0BWP12T U3152 ( .A1(n2734), .A2(n4865), .B1(n4863), .B2(n4804), .C1(
        n4805), .C2(n4867), .ZN(n2290) );
  CKND0BWP12T U3153 ( .I(r12[28]), .ZN(n2735) );
  OAI222D0BWP12T U3154 ( .A1(n2735), .A2(n4865), .B1(n4867), .B2(n4806), .C1(
        n4807), .C2(n4863), .ZN(n2293) );
  CKND0BWP12T U3155 ( .I(r12[30]), .ZN(n2736) );
  OAI222D0BWP12T U3156 ( .A1(n2736), .A2(n4865), .B1(n4863), .B2(n4789), .C1(
        n4790), .C2(n4867), .ZN(n2295) );
  CKND0BWP12T U3157 ( .I(tmp1[2]), .ZN(n2737) );
  OAI222D0BWP12T U3158 ( .A1(n2737), .A2(n4750), .B1(n4749), .B2(n4862), .C1(
        n4866), .C2(n4751), .ZN(n2171) );
  CKND0BWP12T U3159 ( .I(lr[15]), .ZN(n2738) );
  OAI222D0BWP12T U3160 ( .A1(n2738), .A2(n4871), .B1(n4873), .B2(n4829), .C1(
        n4831), .C2(n4869), .ZN(n2248) );
  CKND0BWP12T U3161 ( .I(lr[24]), .ZN(n2739) );
  OAI222D0BWP12T U3162 ( .A1(n2739), .A2(n4871), .B1(n4873), .B2(n4841), .C1(
        n4845), .C2(n4869), .ZN(n2257) );
  CKND0BWP12T U3163 ( .I(lr[29]), .ZN(n2740) );
  OAI222D0BWP12T U3164 ( .A1(n2740), .A2(n4871), .B1(n4873), .B2(n4835), .C1(
        n4837), .C2(n4869), .ZN(n2262) );
  CKND0BWP12T U3165 ( .I(r12[3]), .ZN(n2741) );
  OAI222D0BWP12T U3166 ( .A1(n2741), .A2(n4865), .B1(n4867), .B2(n4793), .C1(
        n4794), .C2(n4863), .ZN(n2268) );
  CKND0BWP12T U3167 ( .I(r12[5]), .ZN(n2742) );
  OAI222D0BWP12T U3168 ( .A1(n2742), .A2(n4865), .B1(n4867), .B2(n4838), .C1(
        n4840), .C2(n4863), .ZN(n2270) );
  CKND0BWP12T U3169 ( .I(r12[9]), .ZN(n2743) );
  OAI222D0BWP12T U3170 ( .A1(n2743), .A2(n4865), .B1(n4867), .B2(n4853), .C1(
        n4855), .C2(n4863), .ZN(n2274) );
  CKND0BWP12T U3171 ( .I(r12[10]), .ZN(n2744) );
  OAI222D0BWP12T U3172 ( .A1(n2744), .A2(n4865), .B1(n4863), .B2(n4808), .C1(
        n4809), .C2(n4867), .ZN(n2275) );
  CKND0BWP12T U3173 ( .I(r12[13]), .ZN(n2745) );
  OAI222D0BWP12T U3174 ( .A1(n2745), .A2(n4865), .B1(n4867), .B2(n4856), .C1(
        n4858), .C2(n4863), .ZN(n2278) );
  CKND0BWP12T U3175 ( .I(r12[16]), .ZN(n2746) );
  OAI222D0BWP12T U3176 ( .A1(n2746), .A2(n4865), .B1(n4863), .B2(n4874), .C1(
        n4878), .C2(n4867), .ZN(n2281) );
  CKND0BWP12T U3177 ( .I(r12[17]), .ZN(n2747) );
  OAI222D0BWP12T U3178 ( .A1(n2747), .A2(n4865), .B1(n4867), .B2(n4812), .C1(
        n4815), .C2(n4863), .ZN(n2282) );
  CKND0BWP12T U3179 ( .I(r12[20]), .ZN(n2748) );
  OAI222D0BWP12T U3180 ( .A1(n2748), .A2(n4865), .B1(n4863), .B2(n4880), .C1(
        n4884), .C2(n4867), .ZN(n2285) );
  CKND0BWP12T U3181 ( .I(r12[21]), .ZN(n2749) );
  OAI222D0BWP12T U3182 ( .A1(n2749), .A2(n4865), .B1(n4867), .B2(n4777), .C1(
        n4778), .C2(n4863), .ZN(n2286) );
  CKND0BWP12T U3183 ( .I(r12[22]), .ZN(n2750) );
  OAI222D0BWP12T U3184 ( .A1(n2750), .A2(n4865), .B1(n4867), .B2(n4785), .C1(
        n4786), .C2(n4863), .ZN(n2287) );
  CKND0BWP12T U3185 ( .I(r12[23]), .ZN(n2751) );
  OAI222D0BWP12T U3186 ( .A1(n2751), .A2(n4865), .B1(n4867), .B2(n4832), .C1(
        n4834), .C2(n4863), .ZN(n2288) );
  CKND0BWP12T U3187 ( .I(r12[26]), .ZN(n2752) );
  OAI222D0BWP12T U3188 ( .A1(n2752), .A2(n4865), .B1(n4867), .B2(n4775), .C1(
        n4776), .C2(n4863), .ZN(n2291) );
  CKND0BWP12T U3189 ( .I(r12[27]), .ZN(n2753) );
  OAI222D0BWP12T U3190 ( .A1(n2753), .A2(n4865), .B1(n4867), .B2(n4787), .C1(
        n4788), .C2(n4863), .ZN(n2292) );
  CKND0BWP12T U3191 ( .I(r12[31]), .ZN(n2754) );
  OAI222D0BWP12T U3192 ( .A1(n2754), .A2(n4865), .B1(n4867), .B2(n4847), .C1(
        n4849), .C2(n4863), .ZN(n2296) );
  CKND0BWP12T U3193 ( .I(r11[0]), .ZN(n2755) );
  OAI222D0BWP12T U3194 ( .A1(n2755), .A2(n3140), .B1(n4859), .B2(n3139), .C1(
        n4861), .C2(n3141), .ZN(n2297) );
  CKND0BWP12T U3195 ( .I(r11[1]), .ZN(n2756) );
  OAI222D0BWP12T U3196 ( .A1(n2756), .A2(n3140), .B1(n4783), .B2(n3141), .C1(
        n4784), .C2(n3139), .ZN(n2298) );
  CKND0BWP12T U3197 ( .I(r11[4]), .ZN(n2757) );
  OAI222D0BWP12T U3198 ( .A1(n2757), .A2(n3140), .B1(n4800), .B2(n3141), .C1(
        n4801), .C2(n3139), .ZN(n2301) );
  CKND0BWP12T U3199 ( .I(r11[6]), .ZN(n2758) );
  OAI222D0BWP12T U3200 ( .A1(n2758), .A2(n3140), .B1(n4779), .B2(n3141), .C1(
        n4780), .C2(n3139), .ZN(n2303) );
  CKND0BWP12T U3201 ( .I(r11[7]), .ZN(n2759) );
  OAI222D0BWP12T U3202 ( .A1(n2759), .A2(n3140), .B1(n4798), .B2(n3139), .C1(
        n4799), .C2(n3141), .ZN(n2304) );
  CKND0BWP12T U3203 ( .I(r11[8]), .ZN(n2760) );
  OAI222D0BWP12T U3204 ( .A1(n2760), .A2(n3140), .B1(n4810), .B2(n3141), .C1(
        n4811), .C2(n3139), .ZN(n2305) );
  CKND0BWP12T U3205 ( .I(r11[11]), .ZN(n2761) );
  OAI222D0BWP12T U3206 ( .A1(n2761), .A2(n3140), .B1(n4868), .B2(n3139), .C1(
        n4872), .C2(n3141), .ZN(n2308) );
  CKND0BWP12T U3207 ( .I(r11[12]), .ZN(n2762) );
  OAI222D0BWP12T U3208 ( .A1(n2762), .A2(n3140), .B1(n4850), .B2(n3141), .C1(
        n4852), .C2(n3139), .ZN(n2309) );
  CKND0BWP12T U3209 ( .I(r11[14]), .ZN(n2763) );
  OAI222D0BWP12T U3210 ( .A1(n2763), .A2(n3140), .B1(n4802), .B2(n3139), .C1(
        n4803), .C2(n3141), .ZN(n2311) );
  CKND0BWP12T U3211 ( .I(r11[18]), .ZN(n2764) );
  OAI222D0BWP12T U3212 ( .A1(n2764), .A2(n3140), .B1(n4791), .B2(n3139), .C1(
        n4792), .C2(n3141), .ZN(n2315) );
  CKND0BWP12T U3213 ( .I(r11[19]), .ZN(n2765) );
  OAI222D0BWP12T U3214 ( .A1(n2765), .A2(n3140), .B1(n4781), .B2(n3139), .C1(
        n4782), .C2(n3141), .ZN(n2316) );
  CKND0BWP12T U3215 ( .I(r11[25]), .ZN(n2766) );
  OAI222D0BWP12T U3216 ( .A1(n2766), .A2(n3140), .B1(n4804), .B2(n3139), .C1(
        n4805), .C2(n3141), .ZN(n2322) );
  CKND0BWP12T U3217 ( .I(r11[28]), .ZN(n2767) );
  OAI222D0BWP12T U3218 ( .A1(n2767), .A2(n3140), .B1(n4806), .B2(n3141), .C1(
        n4807), .C2(n3139), .ZN(n2325) );
  CKND0BWP12T U3219 ( .I(r11[30]), .ZN(n2768) );
  OAI222D0BWP12T U3220 ( .A1(n2768), .A2(n3140), .B1(n4789), .B2(n3139), .C1(
        n4790), .C2(n3141), .ZN(n2327) );
  CKND0BWP12T U3221 ( .I(r12[24]), .ZN(n2769) );
  OAI222D0BWP12T U3222 ( .A1(n2769), .A2(n4865), .B1(n4867), .B2(n4841), .C1(
        n4845), .C2(n4863), .ZN(n2289) );
  CKND0BWP12T U3223 ( .I(r12[29]), .ZN(n2770) );
  OAI222D0BWP12T U3224 ( .A1(n2770), .A2(n4865), .B1(n4867), .B2(n4835), .C1(
        n4837), .C2(n4863), .ZN(n2294) );
  CKND0BWP12T U3225 ( .I(r11[2]), .ZN(n2771) );
  OAI222D0BWP12T U3226 ( .A1(n2771), .A2(n3140), .B1(n4862), .B2(n3139), .C1(
        n4866), .C2(n3141), .ZN(n2299) );
  CKND0BWP12T U3227 ( .I(r11[3]), .ZN(n2772) );
  OAI222D0BWP12T U3228 ( .A1(n2772), .A2(n3140), .B1(n4793), .B2(n3141), .C1(
        n4794), .C2(n3139), .ZN(n2300) );
  CKND0BWP12T U3229 ( .I(r11[5]), .ZN(n2773) );
  OAI222D0BWP12T U3230 ( .A1(n2773), .A2(n3140), .B1(n4838), .B2(n3141), .C1(
        n4840), .C2(n3139), .ZN(n2302) );
  CKND0BWP12T U3231 ( .I(r11[9]), .ZN(n2774) );
  OAI222D0BWP12T U3232 ( .A1(n2774), .A2(n3140), .B1(n4853), .B2(n3141), .C1(
        n4855), .C2(n3139), .ZN(n2306) );
  CKND0BWP12T U3233 ( .I(r11[10]), .ZN(n2775) );
  OAI222D0BWP12T U3234 ( .A1(n2775), .A2(n3140), .B1(n4808), .B2(n3139), .C1(
        n4809), .C2(n3141), .ZN(n2307) );
  CKND0BWP12T U3235 ( .I(r11[13]), .ZN(n2776) );
  OAI222D0BWP12T U3236 ( .A1(n2776), .A2(n3140), .B1(n4856), .B2(n3141), .C1(
        n4858), .C2(n3139), .ZN(n2310) );
  CKND0BWP12T U3237 ( .I(r11[15]), .ZN(n2777) );
  OAI222D0BWP12T U3238 ( .A1(n2777), .A2(n3140), .B1(n4829), .B2(n3141), .C1(
        n4831), .C2(n3139), .ZN(n2312) );
  CKND0BWP12T U3239 ( .I(r11[16]), .ZN(n2778) );
  OAI222D0BWP12T U3240 ( .A1(n2778), .A2(n3140), .B1(n4874), .B2(n3139), .C1(
        n4878), .C2(n3141), .ZN(n2313) );
  CKND0BWP12T U3241 ( .I(r11[17]), .ZN(n2779) );
  OAI222D0BWP12T U3242 ( .A1(n2779), .A2(n3140), .B1(n4812), .B2(n3141), .C1(
        n4815), .C2(n3139), .ZN(n2314) );
  CKND0BWP12T U3243 ( .I(r11[20]), .ZN(n2780) );
  OAI222D0BWP12T U3244 ( .A1(n2780), .A2(n3140), .B1(n4880), .B2(n3139), .C1(
        n4884), .C2(n3141), .ZN(n2317) );
  CKND0BWP12T U3245 ( .I(r11[21]), .ZN(n2781) );
  OAI222D0BWP12T U3246 ( .A1(n2781), .A2(n3140), .B1(n4777), .B2(n3141), .C1(
        n4778), .C2(n3139), .ZN(n2318) );
  CKND0BWP12T U3247 ( .I(r11[22]), .ZN(n2782) );
  OAI222D0BWP12T U3248 ( .A1(n2782), .A2(n3140), .B1(n4785), .B2(n3141), .C1(
        n4786), .C2(n3139), .ZN(n2319) );
  CKND0BWP12T U3249 ( .I(r11[23]), .ZN(n2783) );
  OAI222D0BWP12T U3250 ( .A1(n2783), .A2(n3140), .B1(n4832), .B2(n3141), .C1(
        n4834), .C2(n3139), .ZN(n2320) );
  CKND0BWP12T U3251 ( .I(r11[26]), .ZN(n2784) );
  OAI222D0BWP12T U3252 ( .A1(n2784), .A2(n3140), .B1(n4775), .B2(n3141), .C1(
        n4776), .C2(n3139), .ZN(n2323) );
  CKND0BWP12T U3253 ( .I(r11[27]), .ZN(n2785) );
  OAI222D0BWP12T U3254 ( .A1(n2785), .A2(n3140), .B1(n4787), .B2(n3141), .C1(
        n4788), .C2(n3139), .ZN(n2324) );
  CKND0BWP12T U3255 ( .I(r11[31]), .ZN(n2786) );
  OAI222D0BWP12T U3256 ( .A1(n2786), .A2(n3140), .B1(n4847), .B2(n3141), .C1(
        n4849), .C2(n3139), .ZN(n2328) );
  CKND0BWP12T U3257 ( .I(r10[0]), .ZN(n2787) );
  OAI222D0BWP12T U3258 ( .A1(n2787), .A2(n4814), .B1(n4816), .B2(n4859), .C1(
        n4861), .C2(n4813), .ZN(n2329) );
  CKND0BWP12T U3259 ( .I(r10[1]), .ZN(n2788) );
  OAI222D0BWP12T U3260 ( .A1(n2788), .A2(n4814), .B1(n4813), .B2(n4783), .C1(
        n4784), .C2(n4816), .ZN(n2330) );
  CKND0BWP12T U3261 ( .I(r10[4]), .ZN(n2789) );
  OAI222D0BWP12T U3262 ( .A1(n2789), .A2(n4814), .B1(n4813), .B2(n4800), .C1(
        n4801), .C2(n4816), .ZN(n2333) );
  CKND0BWP12T U3263 ( .I(r10[6]), .ZN(n2790) );
  OAI222D0BWP12T U3264 ( .A1(n2790), .A2(n4814), .B1(n4813), .B2(n4779), .C1(
        n4780), .C2(n4816), .ZN(n2335) );
  CKND0BWP12T U3265 ( .I(r10[7]), .ZN(n2791) );
  OAI222D0BWP12T U3266 ( .A1(n2791), .A2(n4814), .B1(n4816), .B2(n4798), .C1(
        n4799), .C2(n4813), .ZN(n2336) );
  CKND0BWP12T U3267 ( .I(r10[8]), .ZN(n2792) );
  OAI222D0BWP12T U3268 ( .A1(n2792), .A2(n4814), .B1(n4813), .B2(n4810), .C1(
        n4811), .C2(n4816), .ZN(n2337) );
  CKND0BWP12T U3269 ( .I(r10[11]), .ZN(n2793) );
  OAI222D0BWP12T U3270 ( .A1(n2793), .A2(n4814), .B1(n4816), .B2(n4868), .C1(
        n4872), .C2(n4813), .ZN(n2340) );
  CKND0BWP12T U3271 ( .I(r10[12]), .ZN(n2794) );
  OAI222D0BWP12T U3272 ( .A1(n2794), .A2(n4814), .B1(n4813), .B2(n4850), .C1(
        n4852), .C2(n4816), .ZN(n2341) );
  CKND0BWP12T U3273 ( .I(r10[14]), .ZN(n2795) );
  OAI222D0BWP12T U3274 ( .A1(n2795), .A2(n4814), .B1(n4816), .B2(n4802), .C1(
        n4803), .C2(n4813), .ZN(n2343) );
  CKND0BWP12T U3275 ( .I(r10[18]), .ZN(n2796) );
  OAI222D0BWP12T U3276 ( .A1(n2796), .A2(n4814), .B1(n4816), .B2(n4791), .C1(
        n4792), .C2(n4813), .ZN(n2347) );
  CKND0BWP12T U3277 ( .I(r10[19]), .ZN(n2797) );
  OAI222D0BWP12T U3278 ( .A1(n2797), .A2(n4814), .B1(n4816), .B2(n4781), .C1(
        n4782), .C2(n4813), .ZN(n2348) );
  CKND0BWP12T U3279 ( .I(r10[25]), .ZN(n2798) );
  OAI222D0BWP12T U3280 ( .A1(n2798), .A2(n4814), .B1(n4816), .B2(n4804), .C1(
        n4805), .C2(n4813), .ZN(n2354) );
  CKND0BWP12T U3281 ( .I(r10[28]), .ZN(n2799) );
  OAI222D0BWP12T U3282 ( .A1(n2799), .A2(n4814), .B1(n4813), .B2(n4806), .C1(
        n4807), .C2(n4816), .ZN(n2357) );
  CKND0BWP12T U3283 ( .I(r10[30]), .ZN(n2800) );
  OAI222D0BWP12T U3284 ( .A1(n2800), .A2(n4814), .B1(n4816), .B2(n4789), .C1(
        n4790), .C2(n4813), .ZN(n2359) );
  CKND0BWP12T U3285 ( .I(r11[24]), .ZN(n2801) );
  OAI222D0BWP12T U3286 ( .A1(n2801), .A2(n3140), .B1(n4841), .B2(n3141), .C1(
        n4845), .C2(n3139), .ZN(n2321) );
  CKND0BWP12T U3287 ( .I(r11[29]), .ZN(n2802) );
  OAI222D0BWP12T U3288 ( .A1(n2802), .A2(n3140), .B1(n4835), .B2(n3141), .C1(
        n4837), .C2(n3139), .ZN(n2326) );
  CKND0BWP12T U3289 ( .I(r10[2]), .ZN(n2803) );
  OAI222D0BWP12T U3290 ( .A1(n2803), .A2(n4814), .B1(n4816), .B2(n4862), .C1(
        n4866), .C2(n4813), .ZN(n2331) );
  CKND0BWP12T U3291 ( .I(r10[3]), .ZN(n2804) );
  OAI222D0BWP12T U3292 ( .A1(n2804), .A2(n4814), .B1(n4813), .B2(n4793), .C1(
        n4794), .C2(n4816), .ZN(n2332) );
  CKND0BWP12T U3293 ( .I(r10[5]), .ZN(n2805) );
  OAI222D0BWP12T U3294 ( .A1(n2805), .A2(n4814), .B1(n4813), .B2(n4838), .C1(
        n4840), .C2(n4816), .ZN(n2334) );
  CKND0BWP12T U3295 ( .I(r10[9]), .ZN(n2806) );
  OAI222D0BWP12T U3296 ( .A1(n2806), .A2(n4814), .B1(n4813), .B2(n4853), .C1(
        n4855), .C2(n4816), .ZN(n2338) );
  CKND0BWP12T U3297 ( .I(r10[10]), .ZN(n2807) );
  OAI222D0BWP12T U3298 ( .A1(n2807), .A2(n4814), .B1(n4816), .B2(n4808), .C1(
        n4809), .C2(n4813), .ZN(n2339) );
  CKND0BWP12T U3299 ( .I(r10[13]), .ZN(n2808) );
  OAI222D0BWP12T U3300 ( .A1(n2808), .A2(n4814), .B1(n4813), .B2(n4856), .C1(
        n4858), .C2(n4816), .ZN(n2342) );
  CKND0BWP12T U3301 ( .I(r10[15]), .ZN(n2809) );
  OAI222D0BWP12T U3302 ( .A1(n2809), .A2(n4814), .B1(n4813), .B2(n4829), .C1(
        n4831), .C2(n4816), .ZN(n2344) );
  CKND0BWP12T U3303 ( .I(r10[16]), .ZN(n2810) );
  OAI222D0BWP12T U3304 ( .A1(n2810), .A2(n4814), .B1(n4816), .B2(n4874), .C1(
        n4878), .C2(n4813), .ZN(n2345) );
  CKND0BWP12T U3305 ( .I(r10[17]), .ZN(n2811) );
  OAI222D0BWP12T U3306 ( .A1(n2811), .A2(n4814), .B1(n4813), .B2(n4812), .C1(
        n4815), .C2(n4816), .ZN(n2346) );
  CKND0BWP12T U3307 ( .I(r10[20]), .ZN(n2812) );
  OAI222D0BWP12T U3308 ( .A1(n2812), .A2(n4814), .B1(n4816), .B2(n4880), .C1(
        n4884), .C2(n4813), .ZN(n2349) );
  CKND0BWP12T U3309 ( .I(r10[21]), .ZN(n2813) );
  OAI222D0BWP12T U3310 ( .A1(n2813), .A2(n4814), .B1(n4813), .B2(n4777), .C1(
        n4778), .C2(n4816), .ZN(n2350) );
  CKND0BWP12T U3311 ( .I(r10[22]), .ZN(n2814) );
  OAI222D0BWP12T U3312 ( .A1(n2814), .A2(n4814), .B1(n4813), .B2(n4785), .C1(
        n4786), .C2(n4816), .ZN(n2351) );
  CKND0BWP12T U3313 ( .I(r10[23]), .ZN(n2815) );
  OAI222D0BWP12T U3314 ( .A1(n2815), .A2(n4814), .B1(n4813), .B2(n4832), .C1(
        n4834), .C2(n4816), .ZN(n2352) );
  CKND0BWP12T U3315 ( .I(r10[26]), .ZN(n2816) );
  OAI222D0BWP12T U3316 ( .A1(n2816), .A2(n4814), .B1(n4813), .B2(n4775), .C1(
        n4776), .C2(n4816), .ZN(n2355) );
  CKND0BWP12T U3317 ( .I(r10[27]), .ZN(n2817) );
  OAI222D0BWP12T U3318 ( .A1(n2817), .A2(n4814), .B1(n4813), .B2(n4787), .C1(
        n4788), .C2(n4816), .ZN(n2356) );
  CKND0BWP12T U3319 ( .I(r10[31]), .ZN(n2818) );
  OAI222D0BWP12T U3320 ( .A1(n2818), .A2(n4814), .B1(n4813), .B2(n4847), .C1(
        n4849), .C2(n4816), .ZN(n2360) );
  CKND0BWP12T U3321 ( .I(r9[0]), .ZN(n2819) );
  OAI222D0BWP12T U3322 ( .A1(n2819), .A2(n4796), .B1(n4795), .B2(n4859), .C1(
        n4861), .C2(n4797), .ZN(n2361) );
  CKND0BWP12T U3323 ( .I(r9[1]), .ZN(n2820) );
  OAI222D0BWP12T U3324 ( .A1(n2820), .A2(n4796), .B1(n4797), .B2(n4783), .C1(
        n4784), .C2(n4795), .ZN(n2362) );
  CKND0BWP12T U3325 ( .I(r9[4]), .ZN(n2821) );
  OAI222D0BWP12T U3326 ( .A1(n2821), .A2(n4796), .B1(n4797), .B2(n4800), .C1(
        n4801), .C2(n4795), .ZN(n2365) );
  CKND0BWP12T U3327 ( .I(r9[6]), .ZN(n2822) );
  OAI222D0BWP12T U3328 ( .A1(n2822), .A2(n4796), .B1(n4797), .B2(n4779), .C1(
        n4780), .C2(n4795), .ZN(n2367) );
  CKND0BWP12T U3329 ( .I(r9[7]), .ZN(n2823) );
  OAI222D0BWP12T U3330 ( .A1(n2823), .A2(n4796), .B1(n4795), .B2(n4798), .C1(
        n4799), .C2(n4797), .ZN(n2368) );
  CKND0BWP12T U3331 ( .I(r9[8]), .ZN(n2824) );
  OAI222D0BWP12T U3332 ( .A1(n2824), .A2(n4796), .B1(n4797), .B2(n4810), .C1(
        n4811), .C2(n4795), .ZN(n2369) );
  CKND0BWP12T U3333 ( .I(r9[11]), .ZN(n2825) );
  OAI222D0BWP12T U3334 ( .A1(n2825), .A2(n4796), .B1(n4795), .B2(n4868), .C1(
        n4872), .C2(n4797), .ZN(n2372) );
  CKND0BWP12T U3335 ( .I(r9[12]), .ZN(n2826) );
  OAI222D0BWP12T U3336 ( .A1(n2826), .A2(n4796), .B1(n4797), .B2(n4850), .C1(
        n4852), .C2(n4795), .ZN(n2373) );
  CKND0BWP12T U3337 ( .I(r9[14]), .ZN(n2827) );
  OAI222D0BWP12T U3338 ( .A1(n2827), .A2(n4796), .B1(n4795), .B2(n4802), .C1(
        n4803), .C2(n4797), .ZN(n2375) );
  CKND0BWP12T U3339 ( .I(r9[18]), .ZN(n2828) );
  OAI222D0BWP12T U3340 ( .A1(n2828), .A2(n4796), .B1(n4795), .B2(n4791), .C1(
        n4792), .C2(n4797), .ZN(n2379) );
  CKND0BWP12T U3341 ( .I(r9[19]), .ZN(n2829) );
  OAI222D0BWP12T U3342 ( .A1(n2829), .A2(n4796), .B1(n4795), .B2(n4781), .C1(
        n4782), .C2(n4797), .ZN(n2380) );
  CKND0BWP12T U3343 ( .I(r9[25]), .ZN(n2830) );
  OAI222D0BWP12T U3344 ( .A1(n2830), .A2(n4796), .B1(n4795), .B2(n4804), .C1(
        n4805), .C2(n4797), .ZN(n2386) );
  CKND0BWP12T U3345 ( .I(r9[28]), .ZN(n2831) );
  OAI222D0BWP12T U3346 ( .A1(n2831), .A2(n4796), .B1(n4797), .B2(n4806), .C1(
        n4807), .C2(n4795), .ZN(n2389) );
  CKND0BWP12T U3347 ( .I(r9[30]), .ZN(n2832) );
  OAI222D0BWP12T U3348 ( .A1(n2832), .A2(n4796), .B1(n4795), .B2(n4789), .C1(
        n4790), .C2(n4797), .ZN(n2391) );
  CKND0BWP12T U3349 ( .I(r10[24]), .ZN(n2833) );
  OAI222D0BWP12T U3350 ( .A1(n2833), .A2(n4814), .B1(n4813), .B2(n4841), .C1(
        n4845), .C2(n4816), .ZN(n2353) );
  CKND0BWP12T U3351 ( .I(r10[29]), .ZN(n2834) );
  OAI222D0BWP12T U3352 ( .A1(n2834), .A2(n4814), .B1(n4813), .B2(n4835), .C1(
        n4837), .C2(n4816), .ZN(n2358) );
  CKND0BWP12T U3353 ( .I(r9[2]), .ZN(n2835) );
  OAI222D0BWP12T U3354 ( .A1(n2835), .A2(n4796), .B1(n4795), .B2(n4862), .C1(
        n4866), .C2(n4797), .ZN(n2363) );
  CKND0BWP12T U3355 ( .I(r9[3]), .ZN(n2836) );
  OAI222D0BWP12T U3356 ( .A1(n2836), .A2(n4796), .B1(n4797), .B2(n4793), .C1(
        n4794), .C2(n4795), .ZN(n2364) );
  CKND0BWP12T U3357 ( .I(r9[5]), .ZN(n2837) );
  OAI222D0BWP12T U3358 ( .A1(n2837), .A2(n4796), .B1(n4797), .B2(n4838), .C1(
        n4840), .C2(n4795), .ZN(n2366) );
  CKND0BWP12T U3359 ( .I(r9[9]), .ZN(n2838) );
  OAI222D0BWP12T U3360 ( .A1(n2838), .A2(n4796), .B1(n4797), .B2(n4853), .C1(
        n4855), .C2(n4795), .ZN(n2370) );
  CKND0BWP12T U3361 ( .I(r9[10]), .ZN(n2839) );
  OAI222D0BWP12T U3362 ( .A1(n2839), .A2(n4796), .B1(n4795), .B2(n4808), .C1(
        n4809), .C2(n4797), .ZN(n2371) );
  CKND0BWP12T U3363 ( .I(r9[13]), .ZN(n2840) );
  OAI222D0BWP12T U3364 ( .A1(n2840), .A2(n4796), .B1(n4797), .B2(n4856), .C1(
        n4858), .C2(n4795), .ZN(n2374) );
  CKND0BWP12T U3365 ( .I(r9[15]), .ZN(n2841) );
  OAI222D0BWP12T U3366 ( .A1(n2841), .A2(n4796), .B1(n4797), .B2(n4829), .C1(
        n4831), .C2(n4795), .ZN(n2376) );
  CKND0BWP12T U3367 ( .I(r9[16]), .ZN(n2842) );
  OAI222D0BWP12T U3368 ( .A1(n2842), .A2(n4796), .B1(n4795), .B2(n4874), .C1(
        n4878), .C2(n4797), .ZN(n2377) );
  CKND0BWP12T U3369 ( .I(r9[17]), .ZN(n2843) );
  OAI222D0BWP12T U3370 ( .A1(n2843), .A2(n4796), .B1(n4797), .B2(n4812), .C1(
        n4815), .C2(n4795), .ZN(n2378) );
  CKND0BWP12T U3371 ( .I(r9[20]), .ZN(n2844) );
  OAI222D0BWP12T U3372 ( .A1(n2844), .A2(n4796), .B1(n4795), .B2(n4880), .C1(
        n4884), .C2(n4797), .ZN(n2381) );
  CKND0BWP12T U3373 ( .I(r9[21]), .ZN(n2845) );
  OAI222D0BWP12T U3374 ( .A1(n2845), .A2(n4796), .B1(n4797), .B2(n4777), .C1(
        n4778), .C2(n4795), .ZN(n2382) );
  CKND0BWP12T U3375 ( .I(r9[22]), .ZN(n2846) );
  OAI222D0BWP12T U3376 ( .A1(n2846), .A2(n4796), .B1(n4797), .B2(n4785), .C1(
        n4786), .C2(n4795), .ZN(n2383) );
  CKND0BWP12T U3377 ( .I(r9[23]), .ZN(n2847) );
  OAI222D0BWP12T U3378 ( .A1(n2847), .A2(n4796), .B1(n4797), .B2(n4832), .C1(
        n4834), .C2(n4795), .ZN(n2384) );
  CKND0BWP12T U3379 ( .I(r9[26]), .ZN(n2848) );
  OAI222D0BWP12T U3380 ( .A1(n2848), .A2(n4796), .B1(n4797), .B2(n4775), .C1(
        n4776), .C2(n4795), .ZN(n2387) );
  CKND0BWP12T U3381 ( .I(r9[27]), .ZN(n2849) );
  OAI222D0BWP12T U3382 ( .A1(n2849), .A2(n4796), .B1(n4797), .B2(n4787), .C1(
        n4788), .C2(n4795), .ZN(n2388) );
  CKND0BWP12T U3383 ( .I(r9[31]), .ZN(n2850) );
  OAI222D0BWP12T U3384 ( .A1(n2850), .A2(n4796), .B1(n4797), .B2(n4847), .C1(
        n4849), .C2(n4795), .ZN(n2392) );
  CKND0BWP12T U3385 ( .I(r8[0]), .ZN(n2851) );
  OAI222D0BWP12T U3386 ( .A1(n2851), .A2(n4825), .B1(n4826), .B2(n4859), .C1(
        n4861), .C2(n4823), .ZN(n2393) );
  CKND0BWP12T U3387 ( .I(r8[1]), .ZN(n2852) );
  OAI222D0BWP12T U3388 ( .A1(n2852), .A2(n4825), .B1(n4823), .B2(n4783), .C1(
        n4784), .C2(n4826), .ZN(n2394) );
  CKND0BWP12T U3389 ( .I(r8[4]), .ZN(n2853) );
  OAI222D0BWP12T U3390 ( .A1(n2853), .A2(n4825), .B1(n4823), .B2(n4800), .C1(
        n4801), .C2(n4826), .ZN(n2397) );
  CKND0BWP12T U3391 ( .I(r8[6]), .ZN(n2854) );
  OAI222D0BWP12T U3392 ( .A1(n2854), .A2(n4825), .B1(n4823), .B2(n4779), .C1(
        n4780), .C2(n4826), .ZN(n2399) );
  CKND0BWP12T U3393 ( .I(r8[7]), .ZN(n2855) );
  OAI222D0BWP12T U3394 ( .A1(n2855), .A2(n4825), .B1(n4826), .B2(n4798), .C1(
        n4799), .C2(n4823), .ZN(n2400) );
  CKND0BWP12T U3395 ( .I(r8[8]), .ZN(n2856) );
  OAI222D0BWP12T U3396 ( .A1(n2856), .A2(n4825), .B1(n4823), .B2(n4810), .C1(
        n4811), .C2(n4826), .ZN(n2401) );
  CKND0BWP12T U3397 ( .I(r8[11]), .ZN(n2857) );
  OAI222D0BWP12T U3398 ( .A1(n2857), .A2(n4825), .B1(n4826), .B2(n4868), .C1(
        n4872), .C2(n4823), .ZN(n2404) );
  CKND0BWP12T U3399 ( .I(r8[12]), .ZN(n2858) );
  OAI222D0BWP12T U3400 ( .A1(n2858), .A2(n4825), .B1(n4823), .B2(n4850), .C1(
        n4852), .C2(n4826), .ZN(n2405) );
  CKND0BWP12T U3401 ( .I(r8[14]), .ZN(n2859) );
  OAI222D0BWP12T U3402 ( .A1(n2859), .A2(n4825), .B1(n4826), .B2(n4802), .C1(
        n4803), .C2(n4823), .ZN(n2407) );
  CKND0BWP12T U3403 ( .I(r8[18]), .ZN(n2860) );
  OAI222D0BWP12T U3404 ( .A1(n2860), .A2(n4825), .B1(n4826), .B2(n4791), .C1(
        n4792), .C2(n4823), .ZN(n2411) );
  CKND0BWP12T U3405 ( .I(r8[19]), .ZN(n2861) );
  OAI222D0BWP12T U3406 ( .A1(n2861), .A2(n4825), .B1(n4826), .B2(n4781), .C1(
        n4782), .C2(n4823), .ZN(n2412) );
  CKND0BWP12T U3407 ( .I(r8[25]), .ZN(n2862) );
  OAI222D0BWP12T U3408 ( .A1(n2862), .A2(n4825), .B1(n4826), .B2(n4804), .C1(
        n4805), .C2(n4823), .ZN(n2418) );
  CKND0BWP12T U3409 ( .I(r8[28]), .ZN(n2863) );
  OAI222D0BWP12T U3410 ( .A1(n2863), .A2(n4825), .B1(n4823), .B2(n4806), .C1(
        n4807), .C2(n4826), .ZN(n2421) );
  CKND0BWP12T U3411 ( .I(r8[30]), .ZN(n2864) );
  OAI222D0BWP12T U3412 ( .A1(n2864), .A2(n4825), .B1(n4826), .B2(n4789), .C1(
        n4790), .C2(n4823), .ZN(n2423) );
  CKND0BWP12T U3413 ( .I(r9[24]), .ZN(n2865) );
  OAI222D0BWP12T U3414 ( .A1(n2865), .A2(n4796), .B1(n4797), .B2(n4841), .C1(
        n4845), .C2(n4795), .ZN(n2385) );
  CKND0BWP12T U3415 ( .I(r9[29]), .ZN(n2866) );
  OAI222D0BWP12T U3416 ( .A1(n2866), .A2(n4796), .B1(n4797), .B2(n4835), .C1(
        n4837), .C2(n4795), .ZN(n2390) );
  CKND0BWP12T U3417 ( .I(r8[2]), .ZN(n2867) );
  OAI222D0BWP12T U3418 ( .A1(n2867), .A2(n4825), .B1(n4826), .B2(n4862), .C1(
        n4866), .C2(n4823), .ZN(n2395) );
  CKND0BWP12T U3419 ( .I(r8[3]), .ZN(n2868) );
  OAI222D0BWP12T U3420 ( .A1(n2868), .A2(n4825), .B1(n4823), .B2(n4793), .C1(
        n4794), .C2(n4826), .ZN(n2396) );
  CKND0BWP12T U3421 ( .I(r8[5]), .ZN(n2869) );
  OAI222D0BWP12T U3422 ( .A1(n2869), .A2(n4825), .B1(n4823), .B2(n4838), .C1(
        n4840), .C2(n4826), .ZN(n2398) );
  CKND0BWP12T U3423 ( .I(r8[9]), .ZN(n2870) );
  OAI222D0BWP12T U3424 ( .A1(n2870), .A2(n4825), .B1(n4823), .B2(n4853), .C1(
        n4855), .C2(n4826), .ZN(n2402) );
  CKND0BWP12T U3425 ( .I(r8[13]), .ZN(n2871) );
  OAI222D0BWP12T U3426 ( .A1(n2871), .A2(n4825), .B1(n4823), .B2(n4856), .C1(
        n4858), .C2(n4826), .ZN(n2406) );
  CKND0BWP12T U3427 ( .I(r8[15]), .ZN(n2872) );
  OAI222D0BWP12T U3428 ( .A1(n2872), .A2(n4825), .B1(n4823), .B2(n4829), .C1(
        n4831), .C2(n4826), .ZN(n2408) );
  CKND0BWP12T U3429 ( .I(r8[16]), .ZN(n2873) );
  OAI222D0BWP12T U3430 ( .A1(n2873), .A2(n4825), .B1(n4826), .B2(n4874), .C1(
        n4878), .C2(n4823), .ZN(n2409) );
  CKND0BWP12T U3431 ( .I(r8[20]), .ZN(n2874) );
  OAI222D0BWP12T U3432 ( .A1(n2874), .A2(n4825), .B1(n4826), .B2(n4880), .C1(
        n4884), .C2(n4823), .ZN(n2413) );
  CKND0BWP12T U3433 ( .I(r8[21]), .ZN(n2875) );
  OAI222D0BWP12T U3434 ( .A1(n2875), .A2(n4825), .B1(n4823), .B2(n4777), .C1(
        n4778), .C2(n4826), .ZN(n2414) );
  CKND0BWP12T U3435 ( .I(r8[22]), .ZN(n2876) );
  OAI222D0BWP12T U3436 ( .A1(n2876), .A2(n4825), .B1(n4823), .B2(n4785), .C1(
        n4786), .C2(n4826), .ZN(n2415) );
  CKND0BWP12T U3437 ( .I(r8[23]), .ZN(n2877) );
  OAI222D0BWP12T U3438 ( .A1(n2877), .A2(n4825), .B1(n4823), .B2(n4832), .C1(
        n4834), .C2(n4826), .ZN(n2416) );
  CKND0BWP12T U3439 ( .I(r8[26]), .ZN(n2878) );
  OAI222D0BWP12T U3440 ( .A1(n2878), .A2(n4825), .B1(n4823), .B2(n4775), .C1(
        n4776), .C2(n4826), .ZN(n2419) );
  CKND0BWP12T U3441 ( .I(r8[31]), .ZN(n2879) );
  OAI222D0BWP12T U3442 ( .A1(n2879), .A2(n4825), .B1(n4823), .B2(n4847), .C1(
        n4849), .C2(n4826), .ZN(n2424) );
  CKND0BWP12T U3443 ( .I(r7[0]), .ZN(n2880) );
  OAI222D0BWP12T U3444 ( .A1(n2880), .A2(n4770), .B1(n4859), .B2(n4769), .C1(
        n4861), .C2(n4771), .ZN(n2425) );
  CKND0BWP12T U3445 ( .I(r7[1]), .ZN(n2881) );
  OAI222D0BWP12T U3446 ( .A1(n2881), .A2(n4770), .B1(n4783), .B2(n4771), .C1(
        n4784), .C2(n4769), .ZN(n2426) );
  CKND0BWP12T U3447 ( .I(r7[4]), .ZN(n2882) );
  OAI222D0BWP12T U3448 ( .A1(n2882), .A2(n4770), .B1(n4800), .B2(n4771), .C1(
        n4801), .C2(n4769), .ZN(n2429) );
  CKND0BWP12T U3449 ( .I(r7[6]), .ZN(n2883) );
  OAI222D0BWP12T U3450 ( .A1(n2883), .A2(n4770), .B1(n4779), .B2(n4771), .C1(
        n4780), .C2(n4769), .ZN(n2431) );
  CKND0BWP12T U3451 ( .I(r7[7]), .ZN(n2884) );
  OAI222D0BWP12T U3452 ( .A1(n2884), .A2(n4770), .B1(n4798), .B2(n4769), .C1(
        n4799), .C2(n4771), .ZN(n2432) );
  CKND0BWP12T U3453 ( .I(r7[8]), .ZN(n2885) );
  OAI222D0BWP12T U3454 ( .A1(n2885), .A2(n4770), .B1(n4810), .B2(n4771), .C1(
        n4811), .C2(n4769), .ZN(n2433) );
  CKND0BWP12T U3455 ( .I(r7[10]), .ZN(n2886) );
  OAI222D0BWP12T U3456 ( .A1(n2886), .A2(n4770), .B1(n4808), .B2(n4769), .C1(
        n4809), .C2(n4771), .ZN(n2435) );
  CKND0BWP12T U3457 ( .I(r7[11]), .ZN(n2887) );
  OAI222D0BWP12T U3458 ( .A1(n2887), .A2(n4770), .B1(n4868), .B2(n4769), .C1(
        n4872), .C2(n4771), .ZN(n2436) );
  CKND0BWP12T U3459 ( .I(r7[12]), .ZN(n2888) );
  OAI222D0BWP12T U3460 ( .A1(n2888), .A2(n4770), .B1(n4850), .B2(n4771), .C1(
        n4852), .C2(n4769), .ZN(n2437) );
  CKND0BWP12T U3461 ( .I(r7[14]), .ZN(n2889) );
  OAI222D0BWP12T U3462 ( .A1(n2889), .A2(n4770), .B1(n4802), .B2(n4769), .C1(
        n4803), .C2(n4771), .ZN(n2439) );
  CKND0BWP12T U3463 ( .I(r7[17]), .ZN(n2890) );
  OAI222D0BWP12T U3464 ( .A1(n2890), .A2(n4770), .B1(n4812), .B2(n4771), .C1(
        n4815), .C2(n4769), .ZN(n2442) );
  CKND0BWP12T U3465 ( .I(r7[18]), .ZN(n2891) );
  OAI222D0BWP12T U3466 ( .A1(n2891), .A2(n4770), .B1(n4791), .B2(n4769), .C1(
        n4792), .C2(n4771), .ZN(n2443) );
  CKND0BWP12T U3467 ( .I(r7[19]), .ZN(n2892) );
  OAI222D0BWP12T U3468 ( .A1(n2892), .A2(n4770), .B1(n4781), .B2(n4769), .C1(
        n4782), .C2(n4771), .ZN(n2444) );
  CKND0BWP12T U3469 ( .I(r7[25]), .ZN(n2893) );
  OAI222D0BWP12T U3470 ( .A1(n2893), .A2(n4770), .B1(n4804), .B2(n4769), .C1(
        n4805), .C2(n4771), .ZN(n2450) );
  CKND0BWP12T U3471 ( .I(r7[27]), .ZN(n2894) );
  OAI222D0BWP12T U3472 ( .A1(n2894), .A2(n4770), .B1(n4787), .B2(n4771), .C1(
        n4788), .C2(n4769), .ZN(n2452) );
  CKND0BWP12T U3473 ( .I(r7[28]), .ZN(n2895) );
  OAI222D0BWP12T U3474 ( .A1(n2895), .A2(n4770), .B1(n4806), .B2(n4771), .C1(
        n4807), .C2(n4769), .ZN(n2453) );
  CKND0BWP12T U3475 ( .I(r7[30]), .ZN(n2896) );
  OAI222D0BWP12T U3476 ( .A1(n2896), .A2(n4770), .B1(n4789), .B2(n4769), .C1(
        n4790), .C2(n4771), .ZN(n2455) );
  CKND0BWP12T U3477 ( .I(r8[24]), .ZN(n2897) );
  OAI222D0BWP12T U3478 ( .A1(n2897), .A2(n4825), .B1(n4823), .B2(n4841), .C1(
        n4845), .C2(n4826), .ZN(n2417) );
  CKND0BWP12T U3479 ( .I(r7[2]), .ZN(n2898) );
  OAI222D0BWP12T U3480 ( .A1(n2898), .A2(n4770), .B1(n4862), .B2(n4769), .C1(
        n4866), .C2(n4771), .ZN(n2427) );
  CKND0BWP12T U3481 ( .I(r7[3]), .ZN(n2899) );
  OAI222D0BWP12T U3482 ( .A1(n2899), .A2(n4770), .B1(n4793), .B2(n4771), .C1(
        n4794), .C2(n4769), .ZN(n2428) );
  CKND0BWP12T U3483 ( .I(r7[5]), .ZN(n2900) );
  OAI222D0BWP12T U3484 ( .A1(n2900), .A2(n4770), .B1(n4838), .B2(n4771), .C1(
        n4840), .C2(n4769), .ZN(n2430) );
  CKND0BWP12T U3485 ( .I(r7[9]), .ZN(n2901) );
  OAI222D0BWP12T U3486 ( .A1(n2901), .A2(n4770), .B1(n4853), .B2(n4771), .C1(
        n4855), .C2(n4769), .ZN(n2434) );
  CKND0BWP12T U3487 ( .I(r7[13]), .ZN(n2902) );
  OAI222D0BWP12T U3488 ( .A1(n2902), .A2(n4770), .B1(n4856), .B2(n4771), .C1(
        n4858), .C2(n4769), .ZN(n2438) );
  CKND0BWP12T U3489 ( .I(r7[15]), .ZN(n2903) );
  OAI222D0BWP12T U3490 ( .A1(n2903), .A2(n4770), .B1(n4829), .B2(n4771), .C1(
        n4831), .C2(n4769), .ZN(n2440) );
  CKND0BWP12T U3491 ( .I(r7[16]), .ZN(n2904) );
  OAI222D0BWP12T U3492 ( .A1(n2904), .A2(n4770), .B1(n4874), .B2(n4769), .C1(
        n4878), .C2(n4771), .ZN(n2441) );
  CKND0BWP12T U3493 ( .I(r7[20]), .ZN(n2905) );
  OAI222D0BWP12T U3494 ( .A1(n2905), .A2(n4770), .B1(n4880), .B2(n4769), .C1(
        n4884), .C2(n4771), .ZN(n2445) );
  CKND0BWP12T U3495 ( .I(r7[21]), .ZN(n2906) );
  OAI222D0BWP12T U3496 ( .A1(n2906), .A2(n4770), .B1(n4777), .B2(n4771), .C1(
        n4778), .C2(n4769), .ZN(n2446) );
  CKND0BWP12T U3497 ( .I(r7[22]), .ZN(n2907) );
  OAI222D0BWP12T U3498 ( .A1(n2907), .A2(n4770), .B1(n4785), .B2(n4771), .C1(
        n4786), .C2(n4769), .ZN(n2447) );
  CKND0BWP12T U3499 ( .I(r7[23]), .ZN(n2908) );
  OAI222D0BWP12T U3500 ( .A1(n2908), .A2(n4770), .B1(n4832), .B2(n4771), .C1(
        n4834), .C2(n4769), .ZN(n2448) );
  CKND0BWP12T U3501 ( .I(r7[26]), .ZN(n2909) );
  OAI222D0BWP12T U3502 ( .A1(n2909), .A2(n4770), .B1(n4775), .B2(n4771), .C1(
        n4776), .C2(n4769), .ZN(n2451) );
  CKND0BWP12T U3503 ( .I(r7[29]), .ZN(n2910) );
  OAI222D0BWP12T U3504 ( .A1(n2910), .A2(n4770), .B1(n4835), .B2(n4771), .C1(
        n4837), .C2(n4769), .ZN(n2454) );
  CKND0BWP12T U3505 ( .I(r7[31]), .ZN(n2911) );
  OAI222D0BWP12T U3506 ( .A1(n2911), .A2(n4770), .B1(n4847), .B2(n4771), .C1(
        n4849), .C2(n4769), .ZN(n2456) );
  CKND0BWP12T U3507 ( .I(r6[0]), .ZN(n2912) );
  OAI222D0BWP12T U3508 ( .A1(n2912), .A2(n4818), .B1(n4819), .B2(n4859), .C1(
        n4861), .C2(n4817), .ZN(n2457) );
  CKND0BWP12T U3509 ( .I(r6[1]), .ZN(n2913) );
  OAI222D0BWP12T U3510 ( .A1(n2913), .A2(n4818), .B1(n4817), .B2(n4783), .C1(
        n4784), .C2(n4819), .ZN(n2458) );
  CKND0BWP12T U3511 ( .I(r6[4]), .ZN(n2914) );
  OAI222D0BWP12T U3512 ( .A1(n2914), .A2(n4818), .B1(n4817), .B2(n4800), .C1(
        n4801), .C2(n4819), .ZN(n2461) );
  CKND0BWP12T U3513 ( .I(r6[6]), .ZN(n2915) );
  OAI222D0BWP12T U3514 ( .A1(n2915), .A2(n4818), .B1(n4817), .B2(n4779), .C1(
        n4780), .C2(n4819), .ZN(n2463) );
  CKND0BWP12T U3515 ( .I(r6[7]), .ZN(n2916) );
  OAI222D0BWP12T U3516 ( .A1(n2916), .A2(n4818), .B1(n4819), .B2(n4798), .C1(
        n4799), .C2(n4817), .ZN(n2464) );
  CKND0BWP12T U3517 ( .I(r6[8]), .ZN(n2917) );
  OAI222D0BWP12T U3518 ( .A1(n2917), .A2(n4818), .B1(n4817), .B2(n4810), .C1(
        n4811), .C2(n4819), .ZN(n2465) );
  CKND0BWP12T U3519 ( .I(r6[10]), .ZN(n2918) );
  OAI222D0BWP12T U3520 ( .A1(n2918), .A2(n4818), .B1(n4819), .B2(n4808), .C1(
        n4809), .C2(n4817), .ZN(n2467) );
  CKND0BWP12T U3521 ( .I(r6[11]), .ZN(n2919) );
  OAI222D0BWP12T U3522 ( .A1(n2919), .A2(n4818), .B1(n4819), .B2(n4868), .C1(
        n4872), .C2(n4817), .ZN(n2468) );
  CKND0BWP12T U3523 ( .I(r6[12]), .ZN(n2920) );
  OAI222D0BWP12T U3524 ( .A1(n2920), .A2(n4818), .B1(n4817), .B2(n4850), .C1(
        n4852), .C2(n4819), .ZN(n2469) );
  CKND0BWP12T U3525 ( .I(r6[14]), .ZN(n2921) );
  OAI222D0BWP12T U3526 ( .A1(n2921), .A2(n4818), .B1(n4819), .B2(n4802), .C1(
        n4803), .C2(n4817), .ZN(n2471) );
  CKND0BWP12T U3527 ( .I(r6[17]), .ZN(n2922) );
  OAI222D0BWP12T U3528 ( .A1(n2922), .A2(n4818), .B1(n4817), .B2(n4812), .C1(
        n4815), .C2(n4819), .ZN(n2474) );
  CKND0BWP12T U3529 ( .I(r6[18]), .ZN(n2923) );
  OAI222D0BWP12T U3530 ( .A1(n2923), .A2(n4818), .B1(n4819), .B2(n4791), .C1(
        n4792), .C2(n4817), .ZN(n2475) );
  CKND0BWP12T U3531 ( .I(r6[19]), .ZN(n2924) );
  OAI222D0BWP12T U3532 ( .A1(n2924), .A2(n4818), .B1(n4819), .B2(n4781), .C1(
        n4782), .C2(n4817), .ZN(n2476) );
  CKND0BWP12T U3533 ( .I(r6[25]), .ZN(n2925) );
  OAI222D0BWP12T U3534 ( .A1(n2925), .A2(n4818), .B1(n4819), .B2(n4804), .C1(
        n4805), .C2(n4817), .ZN(n2482) );
  CKND0BWP12T U3535 ( .I(r6[27]), .ZN(n2926) );
  OAI222D0BWP12T U3536 ( .A1(n2926), .A2(n4818), .B1(n4817), .B2(n4787), .C1(
        n4788), .C2(n4819), .ZN(n2484) );
  CKND0BWP12T U3537 ( .I(r6[28]), .ZN(n2927) );
  OAI222D0BWP12T U3538 ( .A1(n2927), .A2(n4818), .B1(n4817), .B2(n4806), .C1(
        n4807), .C2(n4819), .ZN(n2485) );
  CKND0BWP12T U3539 ( .I(r6[30]), .ZN(n2928) );
  OAI222D0BWP12T U3540 ( .A1(n2928), .A2(n4818), .B1(n4819), .B2(n4789), .C1(
        n4790), .C2(n4817), .ZN(n2487) );
  CKND0BWP12T U3541 ( .I(r7[24]), .ZN(n2929) );
  OAI222D0BWP12T U3542 ( .A1(n2929), .A2(n4770), .B1(n4841), .B2(n4771), .C1(
        n4845), .C2(n4769), .ZN(n2449) );
  CKND0BWP12T U3543 ( .I(r6[2]), .ZN(n2930) );
  OAI222D0BWP12T U3544 ( .A1(n2930), .A2(n4818), .B1(n4819), .B2(n4862), .C1(
        n4866), .C2(n4817), .ZN(n2459) );
  CKND0BWP12T U3545 ( .I(r6[3]), .ZN(n2931) );
  OAI222D0BWP12T U3546 ( .A1(n2931), .A2(n4818), .B1(n4817), .B2(n4793), .C1(
        n4794), .C2(n4819), .ZN(n2460) );
  CKND0BWP12T U3547 ( .I(r6[5]), .ZN(n2932) );
  OAI222D0BWP12T U3548 ( .A1(n2932), .A2(n4818), .B1(n4817), .B2(n4838), .C1(
        n4840), .C2(n4819), .ZN(n2462) );
  CKND0BWP12T U3549 ( .I(r6[9]), .ZN(n2933) );
  OAI222D0BWP12T U3550 ( .A1(n2933), .A2(n4818), .B1(n4817), .B2(n4853), .C1(
        n4855), .C2(n4819), .ZN(n2466) );
  CKND0BWP12T U3551 ( .I(r6[13]), .ZN(n2934) );
  OAI222D0BWP12T U3552 ( .A1(n2934), .A2(n4818), .B1(n4817), .B2(n4856), .C1(
        n4858), .C2(n4819), .ZN(n2470) );
  CKND0BWP12T U3553 ( .I(r6[15]), .ZN(n2935) );
  OAI222D0BWP12T U3554 ( .A1(n2935), .A2(n4818), .B1(n4817), .B2(n4829), .C1(
        n4831), .C2(n4819), .ZN(n2472) );
  CKND0BWP12T U3555 ( .I(r6[16]), .ZN(n2936) );
  OAI222D0BWP12T U3556 ( .A1(n2936), .A2(n4818), .B1(n4819), .B2(n4874), .C1(
        n4878), .C2(n4817), .ZN(n2473) );
  CKND0BWP12T U3557 ( .I(r6[20]), .ZN(n2937) );
  OAI222D0BWP12T U3558 ( .A1(n2937), .A2(n4818), .B1(n4819), .B2(n4880), .C1(
        n4884), .C2(n4817), .ZN(n2477) );
  CKND0BWP12T U3559 ( .I(r6[21]), .ZN(n2938) );
  OAI222D0BWP12T U3560 ( .A1(n2938), .A2(n4818), .B1(n4817), .B2(n4777), .C1(
        n4778), .C2(n4819), .ZN(n2478) );
  CKND0BWP12T U3561 ( .I(r6[22]), .ZN(n2939) );
  OAI222D0BWP12T U3562 ( .A1(n2939), .A2(n4818), .B1(n4817), .B2(n4785), .C1(
        n4786), .C2(n4819), .ZN(n2479) );
  CKND0BWP12T U3563 ( .I(r6[23]), .ZN(n2940) );
  OAI222D0BWP12T U3564 ( .A1(n2940), .A2(n4818), .B1(n4817), .B2(n4832), .C1(
        n4834), .C2(n4819), .ZN(n2480) );
  CKND0BWP12T U3565 ( .I(r6[26]), .ZN(n2941) );
  OAI222D0BWP12T U3566 ( .A1(n2941), .A2(n4818), .B1(n4817), .B2(n4775), .C1(
        n4776), .C2(n4819), .ZN(n2483) );
  CKND0BWP12T U3567 ( .I(r6[29]), .ZN(n2942) );
  OAI222D0BWP12T U3568 ( .A1(n2942), .A2(n4818), .B1(n4817), .B2(n4835), .C1(
        n4837), .C2(n4819), .ZN(n2486) );
  CKND0BWP12T U3569 ( .I(r6[31]), .ZN(n2943) );
  OAI222D0BWP12T U3570 ( .A1(n2943), .A2(n4818), .B1(n4817), .B2(n4847), .C1(
        n4849), .C2(n4819), .ZN(n2488) );
  CKND0BWP12T U3571 ( .I(r5[0]), .ZN(n2944) );
  OAI222D0BWP12T U3572 ( .A1(n2944), .A2(n4821), .B1(n4820), .B2(n4859), .C1(
        n4861), .C2(n4822), .ZN(n2489) );
  CKND0BWP12T U3573 ( .I(r5[1]), .ZN(n2945) );
  OAI222D0BWP12T U3574 ( .A1(n2945), .A2(n4821), .B1(n4822), .B2(n4783), .C1(
        n4784), .C2(n4820), .ZN(n2490) );
  CKND0BWP12T U3575 ( .I(r5[4]), .ZN(n2946) );
  OAI222D0BWP12T U3576 ( .A1(n2946), .A2(n4821), .B1(n4822), .B2(n4800), .C1(
        n4801), .C2(n4820), .ZN(n2493) );
  CKND0BWP12T U3577 ( .I(r5[6]), .ZN(n2947) );
  OAI222D0BWP12T U3578 ( .A1(n2947), .A2(n4821), .B1(n4822), .B2(n4779), .C1(
        n4780), .C2(n4820), .ZN(n2495) );
  CKND0BWP12T U3579 ( .I(r5[7]), .ZN(n2948) );
  OAI222D0BWP12T U3580 ( .A1(n2948), .A2(n4821), .B1(n4820), .B2(n4798), .C1(
        n4799), .C2(n4822), .ZN(n2496) );
  CKND0BWP12T U3581 ( .I(r5[8]), .ZN(n2949) );
  OAI222D0BWP12T U3582 ( .A1(n2949), .A2(n4821), .B1(n4822), .B2(n4810), .C1(
        n4811), .C2(n4820), .ZN(n2497) );
  CKND0BWP12T U3583 ( .I(r5[10]), .ZN(n2950) );
  OAI222D0BWP12T U3584 ( .A1(n2950), .A2(n4821), .B1(n4820), .B2(n4808), .C1(
        n4809), .C2(n4822), .ZN(n2499) );
  CKND0BWP12T U3585 ( .I(r5[11]), .ZN(n2951) );
  OAI222D0BWP12T U3586 ( .A1(n2951), .A2(n4821), .B1(n4820), .B2(n4868), .C1(
        n4872), .C2(n4822), .ZN(n2500) );
  CKND0BWP12T U3587 ( .I(r5[12]), .ZN(n2952) );
  OAI222D0BWP12T U3588 ( .A1(n2952), .A2(n4821), .B1(n4822), .B2(n4850), .C1(
        n4852), .C2(n4820), .ZN(n2501) );
  CKND0BWP12T U3589 ( .I(r5[14]), .ZN(n2953) );
  OAI222D0BWP12T U3590 ( .A1(n2953), .A2(n4821), .B1(n4820), .B2(n4802), .C1(
        n4803), .C2(n4822), .ZN(n2503) );
  CKND0BWP12T U3591 ( .I(r5[17]), .ZN(n2954) );
  OAI222D0BWP12T U3592 ( .A1(n2954), .A2(n4821), .B1(n4822), .B2(n4812), .C1(
        n4815), .C2(n4820), .ZN(n2506) );
  CKND0BWP12T U3593 ( .I(r5[18]), .ZN(n2955) );
  OAI222D0BWP12T U3594 ( .A1(n2955), .A2(n4821), .B1(n4820), .B2(n4791), .C1(
        n4792), .C2(n4822), .ZN(n2507) );
  CKND0BWP12T U3595 ( .I(r5[19]), .ZN(n2956) );
  OAI222D0BWP12T U3596 ( .A1(n2956), .A2(n4821), .B1(n4820), .B2(n4781), .C1(
        n4782), .C2(n4822), .ZN(n2508) );
  CKND0BWP12T U3597 ( .I(r5[25]), .ZN(n2957) );
  OAI222D0BWP12T U3598 ( .A1(n2957), .A2(n4821), .B1(n4820), .B2(n4804), .C1(
        n4805), .C2(n4822), .ZN(n2514) );
  CKND0BWP12T U3599 ( .I(r5[27]), .ZN(n2958) );
  OAI222D0BWP12T U3600 ( .A1(n2958), .A2(n4821), .B1(n4822), .B2(n4787), .C1(
        n4788), .C2(n4820), .ZN(n2516) );
  CKND0BWP12T U3601 ( .I(r5[28]), .ZN(n2959) );
  OAI222D0BWP12T U3602 ( .A1(n2959), .A2(n4821), .B1(n4822), .B2(n4806), .C1(
        n4807), .C2(n4820), .ZN(n2517) );
  CKND0BWP12T U3603 ( .I(r5[30]), .ZN(n2960) );
  OAI222D0BWP12T U3604 ( .A1(n2960), .A2(n4821), .B1(n4820), .B2(n4789), .C1(
        n4790), .C2(n4822), .ZN(n2519) );
  CKND0BWP12T U3605 ( .I(r6[24]), .ZN(n2961) );
  OAI222D0BWP12T U3606 ( .A1(n2961), .A2(n4818), .B1(n4817), .B2(n4841), .C1(
        n4845), .C2(n4819), .ZN(n2481) );
  CKND0BWP12T U3607 ( .I(r5[2]), .ZN(n2962) );
  OAI222D0BWP12T U3608 ( .A1(n2962), .A2(n4821), .B1(n4820), .B2(n4862), .C1(
        n4866), .C2(n4822), .ZN(n2491) );
  CKND0BWP12T U3609 ( .I(r5[3]), .ZN(n2963) );
  OAI222D0BWP12T U3610 ( .A1(n2963), .A2(n4821), .B1(n4822), .B2(n4793), .C1(
        n4794), .C2(n4820), .ZN(n2492) );
  CKND0BWP12T U3611 ( .I(r5[5]), .ZN(n2964) );
  OAI222D0BWP12T U3612 ( .A1(n2964), .A2(n4821), .B1(n4822), .B2(n4838), .C1(
        n4840), .C2(n4820), .ZN(n2494) );
  CKND0BWP12T U3613 ( .I(r5[9]), .ZN(n2965) );
  OAI222D0BWP12T U3614 ( .A1(n2965), .A2(n4821), .B1(n4822), .B2(n4853), .C1(
        n4855), .C2(n4820), .ZN(n2498) );
  CKND0BWP12T U3615 ( .I(r5[13]), .ZN(n2966) );
  OAI222D0BWP12T U3616 ( .A1(n2966), .A2(n4821), .B1(n4822), .B2(n4856), .C1(
        n4858), .C2(n4820), .ZN(n2502) );
  CKND0BWP12T U3617 ( .I(r5[15]), .ZN(n2967) );
  OAI222D0BWP12T U3618 ( .A1(n2967), .A2(n4821), .B1(n4822), .B2(n4829), .C1(
        n4831), .C2(n4820), .ZN(n2504) );
  CKND0BWP12T U3619 ( .I(r5[16]), .ZN(n2968) );
  OAI222D0BWP12T U3620 ( .A1(n2968), .A2(n4821), .B1(n4820), .B2(n4874), .C1(
        n4878), .C2(n4822), .ZN(n2505) );
  CKND0BWP12T U3621 ( .I(r5[20]), .ZN(n2969) );
  OAI222D0BWP12T U3622 ( .A1(n2969), .A2(n4821), .B1(n4820), .B2(n4880), .C1(
        n4884), .C2(n4822), .ZN(n2509) );
  CKND0BWP12T U3623 ( .I(r5[21]), .ZN(n2970) );
  OAI222D0BWP12T U3624 ( .A1(n2970), .A2(n4821), .B1(n4822), .B2(n4777), .C1(
        n4778), .C2(n4820), .ZN(n2510) );
  CKND0BWP12T U3625 ( .I(r5[22]), .ZN(n2971) );
  OAI222D0BWP12T U3626 ( .A1(n2971), .A2(n4821), .B1(n4822), .B2(n4785), .C1(
        n4786), .C2(n4820), .ZN(n2511) );
  CKND0BWP12T U3627 ( .I(r5[23]), .ZN(n2972) );
  OAI222D0BWP12T U3628 ( .A1(n2972), .A2(n4821), .B1(n4822), .B2(n4832), .C1(
        n4834), .C2(n4820), .ZN(n2512) );
  CKND0BWP12T U3629 ( .I(r5[26]), .ZN(n2973) );
  OAI222D0BWP12T U3630 ( .A1(n2973), .A2(n4821), .B1(n4822), .B2(n4775), .C1(
        n4776), .C2(n4820), .ZN(n2515) );
  CKND0BWP12T U3631 ( .I(r5[29]), .ZN(n2974) );
  OAI222D0BWP12T U3632 ( .A1(n2974), .A2(n4821), .B1(n4822), .B2(n4835), .C1(
        n4837), .C2(n4820), .ZN(n2518) );
  CKND0BWP12T U3633 ( .I(r5[31]), .ZN(n2975) );
  OAI222D0BWP12T U3634 ( .A1(n2975), .A2(n4821), .B1(n4822), .B2(n4847), .C1(
        n4849), .C2(n4820), .ZN(n2520) );
  CKND0BWP12T U3635 ( .I(r4[0]), .ZN(n2976) );
  OAI222D0BWP12T U3636 ( .A1(n2976), .A2(n4767), .B1(n4766), .B2(n4859), .C1(
        n4861), .C2(n4768), .ZN(n2521) );
  CKND0BWP12T U3637 ( .I(r4[1]), .ZN(n2977) );
  OAI222D0BWP12T U3638 ( .A1(n2977), .A2(n4767), .B1(n4768), .B2(n4783), .C1(
        n4784), .C2(n4766), .ZN(n2522) );
  CKND0BWP12T U3639 ( .I(r4[4]), .ZN(n2978) );
  OAI222D0BWP12T U3640 ( .A1(n2978), .A2(n4767), .B1(n4768), .B2(n4800), .C1(
        n4801), .C2(n4766), .ZN(n2525) );
  CKND0BWP12T U3641 ( .I(r4[6]), .ZN(n2979) );
  OAI222D0BWP12T U3642 ( .A1(n2979), .A2(n4767), .B1(n4768), .B2(n4779), .C1(
        n4780), .C2(n4766), .ZN(n2527) );
  CKND0BWP12T U3643 ( .I(r4[7]), .ZN(n2980) );
  OAI222D0BWP12T U3644 ( .A1(n2980), .A2(n4767), .B1(n4766), .B2(n4798), .C1(
        n4799), .C2(n4768), .ZN(n2528) );
  CKND0BWP12T U3645 ( .I(r4[8]), .ZN(n2981) );
  OAI222D0BWP12T U3646 ( .A1(n2981), .A2(n4767), .B1(n4768), .B2(n4810), .C1(
        n4811), .C2(n4766), .ZN(n2529) );
  CKND0BWP12T U3647 ( .I(r4[10]), .ZN(n2982) );
  OAI222D0BWP12T U3648 ( .A1(n2982), .A2(n4767), .B1(n4766), .B2(n4808), .C1(
        n4809), .C2(n4768), .ZN(n2531) );
  CKND0BWP12T U3649 ( .I(r4[11]), .ZN(n2983) );
  OAI222D0BWP12T U3650 ( .A1(n2983), .A2(n4767), .B1(n4766), .B2(n4868), .C1(
        n4872), .C2(n4768), .ZN(n2532) );
  CKND0BWP12T U3651 ( .I(r4[12]), .ZN(n2984) );
  OAI222D0BWP12T U3652 ( .A1(n2984), .A2(n4767), .B1(n4768), .B2(n4850), .C1(
        n4852), .C2(n4766), .ZN(n2533) );
  CKND0BWP12T U3653 ( .I(r4[14]), .ZN(n2985) );
  OAI222D0BWP12T U3654 ( .A1(n2985), .A2(n4767), .B1(n4766), .B2(n4802), .C1(
        n4803), .C2(n4768), .ZN(n2535) );
  CKND0BWP12T U3655 ( .I(r4[17]), .ZN(n2986) );
  OAI222D0BWP12T U3656 ( .A1(n2986), .A2(n4767), .B1(n4768), .B2(n4812), .C1(
        n4815), .C2(n4766), .ZN(n2538) );
  CKND0BWP12T U3657 ( .I(r4[18]), .ZN(n2987) );
  OAI222D0BWP12T U3658 ( .A1(n2987), .A2(n4767), .B1(n4766), .B2(n4791), .C1(
        n4792), .C2(n4768), .ZN(n2539) );
  CKND0BWP12T U3659 ( .I(r4[19]), .ZN(n2988) );
  OAI222D0BWP12T U3660 ( .A1(n2988), .A2(n4767), .B1(n4766), .B2(n4781), .C1(
        n4782), .C2(n4768), .ZN(n2540) );
  CKND0BWP12T U3661 ( .I(r4[25]), .ZN(n2989) );
  OAI222D0BWP12T U3662 ( .A1(n2989), .A2(n4767), .B1(n4766), .B2(n4804), .C1(
        n4805), .C2(n4768), .ZN(n2546) );
  CKND0BWP12T U3663 ( .I(r4[27]), .ZN(n2990) );
  OAI222D0BWP12T U3664 ( .A1(n2990), .A2(n4767), .B1(n4768), .B2(n4787), .C1(
        n4788), .C2(n4766), .ZN(n2548) );
  CKND0BWP12T U3665 ( .I(r4[28]), .ZN(n2991) );
  OAI222D0BWP12T U3666 ( .A1(n2991), .A2(n4767), .B1(n4768), .B2(n4806), .C1(
        n4807), .C2(n4766), .ZN(n2549) );
  CKND0BWP12T U3667 ( .I(r4[30]), .ZN(n2992) );
  OAI222D0BWP12T U3668 ( .A1(n2992), .A2(n4767), .B1(n4766), .B2(n4789), .C1(
        n4790), .C2(n4768), .ZN(n2551) );
  CKND0BWP12T U3669 ( .I(r5[24]), .ZN(n2993) );
  OAI222D0BWP12T U3670 ( .A1(n2993), .A2(n4821), .B1(n4822), .B2(n4841), .C1(
        n4845), .C2(n4820), .ZN(n2513) );
  CKND0BWP12T U3671 ( .I(r4[2]), .ZN(n2994) );
  OAI222D0BWP12T U3672 ( .A1(n2994), .A2(n4767), .B1(n4766), .B2(n4862), .C1(
        n4866), .C2(n4768), .ZN(n2523) );
  CKND0BWP12T U3673 ( .I(r4[3]), .ZN(n2995) );
  OAI222D0BWP12T U3674 ( .A1(n2995), .A2(n4767), .B1(n4768), .B2(n4793), .C1(
        n4794), .C2(n4766), .ZN(n2524) );
  CKND0BWP12T U3675 ( .I(r4[5]), .ZN(n2996) );
  OAI222D0BWP12T U3676 ( .A1(n2996), .A2(n4767), .B1(n4768), .B2(n4838), .C1(
        n4840), .C2(n4766), .ZN(n2526) );
  CKND0BWP12T U3677 ( .I(r4[9]), .ZN(n2997) );
  OAI222D0BWP12T U3678 ( .A1(n2997), .A2(n4767), .B1(n4768), .B2(n4853), .C1(
        n4855), .C2(n4766), .ZN(n2530) );
  CKND0BWP12T U3679 ( .I(r4[13]), .ZN(n2998) );
  OAI222D0BWP12T U3680 ( .A1(n2998), .A2(n4767), .B1(n4768), .B2(n4856), .C1(
        n4858), .C2(n4766), .ZN(n2534) );
  CKND0BWP12T U3681 ( .I(r4[15]), .ZN(n2999) );
  OAI222D0BWP12T U3682 ( .A1(n2999), .A2(n4767), .B1(n4768), .B2(n4829), .C1(
        n4831), .C2(n4766), .ZN(n2536) );
  CKND0BWP12T U3683 ( .I(r4[16]), .ZN(n3000) );
  OAI222D0BWP12T U3684 ( .A1(n3000), .A2(n4767), .B1(n4766), .B2(n4874), .C1(
        n4878), .C2(n4768), .ZN(n2537) );
  CKND0BWP12T U3685 ( .I(r4[20]), .ZN(n3001) );
  OAI222D0BWP12T U3686 ( .A1(n3001), .A2(n4767), .B1(n4766), .B2(n4880), .C1(
        n4884), .C2(n4768), .ZN(n2541) );
  CKND0BWP12T U3687 ( .I(r4[21]), .ZN(n3002) );
  OAI222D0BWP12T U3688 ( .A1(n3002), .A2(n4767), .B1(n4768), .B2(n4777), .C1(
        n4778), .C2(n4766), .ZN(n2542) );
  CKND0BWP12T U3689 ( .I(r4[22]), .ZN(n3003) );
  OAI222D0BWP12T U3690 ( .A1(n3003), .A2(n4767), .B1(n4768), .B2(n4785), .C1(
        n4786), .C2(n4766), .ZN(n2543) );
  CKND0BWP12T U3691 ( .I(r4[23]), .ZN(n3004) );
  OAI222D0BWP12T U3692 ( .A1(n3004), .A2(n4767), .B1(n4768), .B2(n4832), .C1(
        n4834), .C2(n4766), .ZN(n2544) );
  CKND0BWP12T U3693 ( .I(r4[26]), .ZN(n3005) );
  OAI222D0BWP12T U3694 ( .A1(n3005), .A2(n4767), .B1(n4768), .B2(n4775), .C1(
        n4776), .C2(n4766), .ZN(n2547) );
  CKND0BWP12T U3695 ( .I(r4[29]), .ZN(n3006) );
  OAI222D0BWP12T U3696 ( .A1(n3006), .A2(n4767), .B1(n4768), .B2(n4835), .C1(
        n4837), .C2(n4766), .ZN(n2550) );
  CKND0BWP12T U3697 ( .I(r4[31]), .ZN(n3007) );
  OAI222D0BWP12T U3698 ( .A1(n3007), .A2(n4767), .B1(n4768), .B2(n4847), .C1(
        n4849), .C2(n4766), .ZN(n2552) );
  CKND0BWP12T U3699 ( .I(r3[0]), .ZN(n3008) );
  OAI222D0BWP12T U3700 ( .A1(n3008), .A2(n4773), .B1(n4772), .B2(n4859), .C1(
        n4861), .C2(n4774), .ZN(n2553) );
  CKND0BWP12T U3701 ( .I(r3[1]), .ZN(n3009) );
  OAI222D0BWP12T U3702 ( .A1(n3009), .A2(n4773), .B1(n4774), .B2(n4783), .C1(
        n4784), .C2(n4772), .ZN(n2554) );
  CKND0BWP12T U3703 ( .I(r3[4]), .ZN(n3010) );
  OAI222D0BWP12T U3704 ( .A1(n3010), .A2(n4773), .B1(n4774), .B2(n4800), .C1(
        n4801), .C2(n4772), .ZN(n2557) );
  CKND0BWP12T U3705 ( .I(r3[6]), .ZN(n3011) );
  OAI222D0BWP12T U3706 ( .A1(n3011), .A2(n4773), .B1(n4774), .B2(n4779), .C1(
        n4780), .C2(n4772), .ZN(n2559) );
  CKND0BWP12T U3707 ( .I(r3[7]), .ZN(n3012) );
  OAI222D0BWP12T U3708 ( .A1(n3012), .A2(n4773), .B1(n4772), .B2(n4798), .C1(
        n4799), .C2(n4774), .ZN(n2560) );
  CKND0BWP12T U3709 ( .I(r3[8]), .ZN(n3013) );
  OAI222D0BWP12T U3710 ( .A1(n3013), .A2(n4773), .B1(n4774), .B2(n4810), .C1(
        n4811), .C2(n4772), .ZN(n2561) );
  CKND0BWP12T U3711 ( .I(r3[10]), .ZN(n3014) );
  OAI222D0BWP12T U3712 ( .A1(n3014), .A2(n4773), .B1(n4772), .B2(n4808), .C1(
        n4809), .C2(n4774), .ZN(n2563) );
  CKND0BWP12T U3713 ( .I(r3[11]), .ZN(n3015) );
  OAI222D0BWP12T U3714 ( .A1(n3015), .A2(n4773), .B1(n4772), .B2(n4868), .C1(
        n4872), .C2(n4774), .ZN(n2564) );
  CKND0BWP12T U3715 ( .I(r3[12]), .ZN(n3016) );
  OAI222D0BWP12T U3716 ( .A1(n3016), .A2(n4773), .B1(n4774), .B2(n4850), .C1(
        n4852), .C2(n4772), .ZN(n2565) );
  CKND0BWP12T U3717 ( .I(r3[14]), .ZN(n3017) );
  OAI222D0BWP12T U3718 ( .A1(n3017), .A2(n4773), .B1(n4772), .B2(n4802), .C1(
        n4803), .C2(n4774), .ZN(n2567) );
  CKND0BWP12T U3719 ( .I(r3[17]), .ZN(n3018) );
  OAI222D0BWP12T U3720 ( .A1(n3018), .A2(n4773), .B1(n4774), .B2(n4812), .C1(
        n4815), .C2(n4772), .ZN(n2570) );
  CKND0BWP12T U3721 ( .I(r3[18]), .ZN(n3019) );
  OAI222D0BWP12T U3722 ( .A1(n3019), .A2(n4773), .B1(n4772), .B2(n4791), .C1(
        n4792), .C2(n4774), .ZN(n2571) );
  CKND0BWP12T U3723 ( .I(r3[19]), .ZN(n3020) );
  OAI222D0BWP12T U3724 ( .A1(n3020), .A2(n4773), .B1(n4772), .B2(n4781), .C1(
        n4782), .C2(n4774), .ZN(n2572) );
  CKND0BWP12T U3725 ( .I(r3[25]), .ZN(n3021) );
  OAI222D0BWP12T U3726 ( .A1(n3021), .A2(n4773), .B1(n4772), .B2(n4804), .C1(
        n4805), .C2(n4774), .ZN(n2578) );
  CKND0BWP12T U3727 ( .I(r3[27]), .ZN(n3022) );
  OAI222D0BWP12T U3728 ( .A1(n3022), .A2(n4773), .B1(n4774), .B2(n4787), .C1(
        n4788), .C2(n4772), .ZN(n2580) );
  CKND0BWP12T U3729 ( .I(r3[28]), .ZN(n3023) );
  OAI222D0BWP12T U3730 ( .A1(n3023), .A2(n4773), .B1(n4774), .B2(n4806), .C1(
        n4807), .C2(n4772), .ZN(n2581) );
  CKND0BWP12T U3731 ( .I(r3[30]), .ZN(n3024) );
  OAI222D0BWP12T U3732 ( .A1(n3024), .A2(n4773), .B1(n4772), .B2(n4789), .C1(
        n4790), .C2(n4774), .ZN(n2583) );
  CKND0BWP12T U3733 ( .I(r4[24]), .ZN(n3025) );
  OAI222D0BWP12T U3734 ( .A1(n3025), .A2(n4767), .B1(n4768), .B2(n4841), .C1(
        n4845), .C2(n4766), .ZN(n2545) );
  CKND0BWP12T U3735 ( .I(r3[3]), .ZN(n3026) );
  OAI222D0BWP12T U3736 ( .A1(n3026), .A2(n4773), .B1(n4774), .B2(n4793), .C1(
        n4794), .C2(n4772), .ZN(n2556) );
  CKND0BWP12T U3737 ( .I(r3[5]), .ZN(n3027) );
  OAI222D0BWP12T U3738 ( .A1(n3027), .A2(n4773), .B1(n4774), .B2(n4838), .C1(
        n4840), .C2(n4772), .ZN(n2558) );
  CKND0BWP12T U3739 ( .I(r3[9]), .ZN(n3028) );
  OAI222D0BWP12T U3740 ( .A1(n3028), .A2(n4773), .B1(n4774), .B2(n4853), .C1(
        n4855), .C2(n4772), .ZN(n2562) );
  CKND0BWP12T U3741 ( .I(r3[13]), .ZN(n3029) );
  OAI222D0BWP12T U3742 ( .A1(n3029), .A2(n4773), .B1(n4774), .B2(n4856), .C1(
        n4858), .C2(n4772), .ZN(n2566) );
  CKND0BWP12T U3743 ( .I(r3[15]), .ZN(n3030) );
  OAI222D0BWP12T U3744 ( .A1(n3030), .A2(n4773), .B1(n4774), .B2(n4829), .C1(
        n4831), .C2(n4772), .ZN(n2568) );
  CKND0BWP12T U3745 ( .I(r3[16]), .ZN(n3031) );
  OAI222D0BWP12T U3746 ( .A1(n3031), .A2(n4773), .B1(n4772), .B2(n4874), .C1(
        n4878), .C2(n4774), .ZN(n2569) );
  CKND0BWP12T U3747 ( .I(r3[20]), .ZN(n3032) );
  OAI222D0BWP12T U3748 ( .A1(n3032), .A2(n4773), .B1(n4772), .B2(n4880), .C1(
        n4884), .C2(n4774), .ZN(n2573) );
  CKND0BWP12T U3749 ( .I(r3[22]), .ZN(n3033) );
  OAI222D0BWP12T U3750 ( .A1(n3033), .A2(n4773), .B1(n4774), .B2(n4785), .C1(
        n4786), .C2(n4772), .ZN(n2575) );
  CKND0BWP12T U3751 ( .I(r3[23]), .ZN(n3034) );
  OAI222D0BWP12T U3752 ( .A1(n3034), .A2(n4773), .B1(n4774), .B2(n4832), .C1(
        n4834), .C2(n4772), .ZN(n2576) );
  CKND0BWP12T U3753 ( .I(r3[26]), .ZN(n3035) );
  OAI222D0BWP12T U3754 ( .A1(n3035), .A2(n4773), .B1(n4774), .B2(n4775), .C1(
        n4776), .C2(n4772), .ZN(n2579) );
  CKND0BWP12T U3755 ( .I(r3[29]), .ZN(n3036) );
  OAI222D0BWP12T U3756 ( .A1(n3036), .A2(n4773), .B1(n4774), .B2(n4835), .C1(
        n4837), .C2(n4772), .ZN(n2582) );
  CKND0BWP12T U3757 ( .I(r3[31]), .ZN(n3037) );
  OAI222D0BWP12T U3758 ( .A1(n3037), .A2(n4773), .B1(n4774), .B2(n4847), .C1(
        n4849), .C2(n4772), .ZN(n2584) );
  CKND0BWP12T U3759 ( .I(r2[0]), .ZN(n3038) );
  OAI222D0BWP12T U3760 ( .A1(n3038), .A2(n4883), .B1(n4881), .B2(n4859), .C1(
        n4861), .C2(n4885), .ZN(n2585) );
  CKND0BWP12T U3761 ( .I(r2[1]), .ZN(n3039) );
  OAI222D0BWP12T U3762 ( .A1(n3039), .A2(n4883), .B1(n4885), .B2(n4783), .C1(
        n4784), .C2(n4881), .ZN(n2586) );
  CKND0BWP12T U3763 ( .I(r2[2]), .ZN(n3040) );
  OAI222D0BWP12T U3764 ( .A1(n3040), .A2(n4883), .B1(n4881), .B2(n4862), .C1(
        n4866), .C2(n4885), .ZN(n2587) );
  CKND0BWP12T U3765 ( .I(r2[4]), .ZN(n3041) );
  OAI222D0BWP12T U3766 ( .A1(n3041), .A2(n4883), .B1(n4885), .B2(n4800), .C1(
        n4801), .C2(n4881), .ZN(n2589) );
  CKND0BWP12T U3767 ( .I(r2[6]), .ZN(n3042) );
  OAI222D0BWP12T U3768 ( .A1(n3042), .A2(n4883), .B1(n4885), .B2(n4779), .C1(
        n4780), .C2(n4881), .ZN(n2591) );
  CKND0BWP12T U3769 ( .I(r2[7]), .ZN(n3043) );
  OAI222D0BWP12T U3770 ( .A1(n3043), .A2(n4883), .B1(n4881), .B2(n4798), .C1(
        n4799), .C2(n4885), .ZN(n2592) );
  CKND0BWP12T U3771 ( .I(r2[8]), .ZN(n3044) );
  OAI222D0BWP12T U3772 ( .A1(n3044), .A2(n4883), .B1(n4885), .B2(n4810), .C1(
        n4811), .C2(n4881), .ZN(n2593) );
  CKND0BWP12T U3773 ( .I(r2[10]), .ZN(n3045) );
  OAI222D0BWP12T U3774 ( .A1(n3045), .A2(n4883), .B1(n4881), .B2(n4808), .C1(
        n4809), .C2(n4885), .ZN(n2595) );
  CKND0BWP12T U3775 ( .I(r2[11]), .ZN(n3046) );
  OAI222D0BWP12T U3776 ( .A1(n3046), .A2(n4883), .B1(n4881), .B2(n4868), .C1(
        n4872), .C2(n4885), .ZN(n2596) );
  CKND0BWP12T U3777 ( .I(r2[12]), .ZN(n3047) );
  OAI222D0BWP12T U3778 ( .A1(n3047), .A2(n4883), .B1(n4885), .B2(n4850), .C1(
        n4852), .C2(n4881), .ZN(n2597) );
  CKND0BWP12T U3779 ( .I(r2[14]), .ZN(n3048) );
  OAI222D0BWP12T U3780 ( .A1(n3048), .A2(n4883), .B1(n4881), .B2(n4802), .C1(
        n4803), .C2(n4885), .ZN(n2599) );
  CKND0BWP12T U3781 ( .I(r2[17]), .ZN(n3049) );
  OAI222D0BWP12T U3782 ( .A1(n3049), .A2(n4883), .B1(n4885), .B2(n4812), .C1(
        n4815), .C2(n4881), .ZN(n2602) );
  CKND0BWP12T U3783 ( .I(r2[18]), .ZN(n3050) );
  OAI222D0BWP12T U3784 ( .A1(n3050), .A2(n4883), .B1(n4881), .B2(n4791), .C1(
        n4792), .C2(n4885), .ZN(n2603) );
  CKND0BWP12T U3785 ( .I(r2[19]), .ZN(n3051) );
  OAI222D0BWP12T U3786 ( .A1(n3051), .A2(n4883), .B1(n4881), .B2(n4781), .C1(
        n4782), .C2(n4885), .ZN(n2604) );
  CKND0BWP12T U3787 ( .I(r2[21]), .ZN(n3052) );
  OAI222D0BWP12T U3788 ( .A1(n3052), .A2(n4883), .B1(n4885), .B2(n4777), .C1(
        n4778), .C2(n4881), .ZN(n2606) );
  CKND0BWP12T U3789 ( .I(r2[25]), .ZN(n3053) );
  OAI222D0BWP12T U3790 ( .A1(n3053), .A2(n4883), .B1(n4881), .B2(n4804), .C1(
        n4805), .C2(n4885), .ZN(n2610) );
  CKND0BWP12T U3791 ( .I(r2[27]), .ZN(n3054) );
  OAI222D0BWP12T U3792 ( .A1(n3054), .A2(n4883), .B1(n4885), .B2(n4787), .C1(
        n4788), .C2(n4881), .ZN(n2612) );
  CKND0BWP12T U3793 ( .I(r2[28]), .ZN(n3055) );
  OAI222D0BWP12T U3794 ( .A1(n3055), .A2(n4883), .B1(n4885), .B2(n4806), .C1(
        n4807), .C2(n4881), .ZN(n2613) );
  CKND0BWP12T U3795 ( .I(r2[30]), .ZN(n3056) );
  OAI222D0BWP12T U3796 ( .A1(n3056), .A2(n4883), .B1(n4881), .B2(n4789), .C1(
        n4790), .C2(n4885), .ZN(n2615) );
  CKND0BWP12T U3797 ( .I(r2[5]), .ZN(n3057) );
  OAI222D0BWP12T U3798 ( .A1(n3057), .A2(n4883), .B1(n4885), .B2(n4838), .C1(
        n4840), .C2(n4881), .ZN(n2590) );
  CKND0BWP12T U3799 ( .I(r2[9]), .ZN(n3058) );
  OAI222D0BWP12T U3800 ( .A1(n3058), .A2(n4883), .B1(n4885), .B2(n4853), .C1(
        n4855), .C2(n4881), .ZN(n2594) );
  CKND0BWP12T U3801 ( .I(r2[15]), .ZN(n3059) );
  OAI222D0BWP12T U3802 ( .A1(n3059), .A2(n4883), .B1(n4885), .B2(n4829), .C1(
        n4831), .C2(n4881), .ZN(n2600) );
  CKND0BWP12T U3803 ( .I(r2[16]), .ZN(n3060) );
  OAI222D0BWP12T U3804 ( .A1(n3060), .A2(n4883), .B1(n4881), .B2(n4874), .C1(
        n4878), .C2(n4885), .ZN(n2601) );
  CKND0BWP12T U3805 ( .I(r2[23]), .ZN(n3061) );
  OAI222D0BWP12T U3806 ( .A1(n3061), .A2(n4883), .B1(n4885), .B2(n4832), .C1(
        n4834), .C2(n4881), .ZN(n2608) );
  CKND0BWP12T U3807 ( .I(r2[24]), .ZN(n3062) );
  OAI222D0BWP12T U3808 ( .A1(n3062), .A2(n4883), .B1(n4885), .B2(n4841), .C1(
        n4845), .C2(n4881), .ZN(n2609) );
  CKND0BWP12T U3809 ( .I(r2[29]), .ZN(n3063) );
  OAI222D0BWP12T U3810 ( .A1(n3063), .A2(n4883), .B1(n4885), .B2(n4835), .C1(
        n4837), .C2(n4881), .ZN(n2614) );
  CKND0BWP12T U3811 ( .I(r2[31]), .ZN(n3064) );
  OAI222D0BWP12T U3812 ( .A1(n3064), .A2(n4883), .B1(n4885), .B2(n4847), .C1(
        n4849), .C2(n4881), .ZN(n2616) );
  CKND0BWP12T U3813 ( .I(r1[0]), .ZN(n3065) );
  OAI222D0BWP12T U3814 ( .A1(n3065), .A2(n4844), .B1(n4846), .B2(n4859), .C1(
        n4861), .C2(n4842), .ZN(n2617) );
  CKND0BWP12T U3815 ( .I(r1[1]), .ZN(n3066) );
  OAI222D0BWP12T U3816 ( .A1(n3066), .A2(n4844), .B1(n4842), .B2(n4783), .C1(
        n4784), .C2(n4846), .ZN(n2618) );
  CKND0BWP12T U3817 ( .I(r1[2]), .ZN(n3067) );
  OAI222D0BWP12T U3818 ( .A1(n3067), .A2(n4844), .B1(n4846), .B2(n4862), .C1(
        n4866), .C2(n4842), .ZN(n2619) );
  CKND0BWP12T U3819 ( .I(r1[3]), .ZN(n3068) );
  OAI222D0BWP12T U3820 ( .A1(n3068), .A2(n4844), .B1(n4842), .B2(n4793), .C1(
        n4794), .C2(n4846), .ZN(n2620) );
  CKND0BWP12T U3821 ( .I(r1[4]), .ZN(n3069) );
  OAI222D0BWP12T U3822 ( .A1(n3069), .A2(n4844), .B1(n4842), .B2(n4800), .C1(
        n4801), .C2(n4846), .ZN(n2621) );
  CKND0BWP12T U3823 ( .I(r1[6]), .ZN(n3070) );
  OAI222D0BWP12T U3824 ( .A1(n3070), .A2(n4844), .B1(n4842), .B2(n4779), .C1(
        n4780), .C2(n4846), .ZN(n2623) );
  CKND0BWP12T U3825 ( .I(r1[7]), .ZN(n3071) );
  OAI222D0BWP12T U3826 ( .A1(n3071), .A2(n4844), .B1(n4846), .B2(n4798), .C1(
        n4799), .C2(n4842), .ZN(n2624) );
  CKND0BWP12T U3827 ( .I(r1[8]), .ZN(n3072) );
  OAI222D0BWP12T U3828 ( .A1(n3072), .A2(n4844), .B1(n4842), .B2(n4810), .C1(
        n4811), .C2(n4846), .ZN(n2625) );
  CKND0BWP12T U3829 ( .I(r1[10]), .ZN(n3073) );
  OAI222D0BWP12T U3830 ( .A1(n3073), .A2(n4844), .B1(n4846), .B2(n4808), .C1(
        n4809), .C2(n4842), .ZN(n2627) );
  CKND0BWP12T U3831 ( .I(r1[11]), .ZN(n3074) );
  OAI222D0BWP12T U3832 ( .A1(n3074), .A2(n4844), .B1(n4846), .B2(n4868), .C1(
        n4872), .C2(n4842), .ZN(n2628) );
  CKND0BWP12T U3833 ( .I(r1[12]), .ZN(n3075) );
  OAI222D0BWP12T U3834 ( .A1(n3075), .A2(n4844), .B1(n4842), .B2(n4850), .C1(
        n4852), .C2(n4846), .ZN(n2629) );
  CKND0BWP12T U3835 ( .I(r1[13]), .ZN(n3076) );
  OAI222D0BWP12T U3836 ( .A1(n3076), .A2(n4844), .B1(n4842), .B2(n4856), .C1(
        n4858), .C2(n4846), .ZN(n2630) );
  CKND0BWP12T U3837 ( .I(r1[14]), .ZN(n3077) );
  OAI222D0BWP12T U3838 ( .A1(n3077), .A2(n4844), .B1(n4846), .B2(n4802), .C1(
        n4803), .C2(n4842), .ZN(n2631) );
  CKND0BWP12T U3839 ( .I(r1[17]), .ZN(n3078) );
  OAI222D0BWP12T U3840 ( .A1(n3078), .A2(n4844), .B1(n4842), .B2(n4812), .C1(
        n4815), .C2(n4846), .ZN(n2634) );
  CKND0BWP12T U3841 ( .I(r1[18]), .ZN(n3079) );
  OAI222D0BWP12T U3842 ( .A1(n3079), .A2(n4844), .B1(n4846), .B2(n4791), .C1(
        n4792), .C2(n4842), .ZN(n2635) );
  CKND0BWP12T U3843 ( .I(r1[19]), .ZN(n3080) );
  OAI222D0BWP12T U3844 ( .A1(n3080), .A2(n4844), .B1(n4846), .B2(n4781), .C1(
        n4782), .C2(n4842), .ZN(n2636) );
  CKND0BWP12T U3845 ( .I(r1[20]), .ZN(n3081) );
  OAI222D0BWP12T U3846 ( .A1(n3081), .A2(n4844), .B1(n4846), .B2(n4880), .C1(
        n4884), .C2(n4842), .ZN(n2637) );
  CKND0BWP12T U3847 ( .I(r1[21]), .ZN(n3082) );
  OAI222D0BWP12T U3848 ( .A1(n3082), .A2(n4844), .B1(n4842), .B2(n4777), .C1(
        n4778), .C2(n4846), .ZN(n2638) );
  CKND0BWP12T U3849 ( .I(r1[22]), .ZN(n3083) );
  OAI222D0BWP12T U3850 ( .A1(n3083), .A2(n4844), .B1(n4842), .B2(n4785), .C1(
        n4786), .C2(n4846), .ZN(n2639) );
  CKND0BWP12T U3851 ( .I(r1[25]), .ZN(n3084) );
  OAI222D0BWP12T U3852 ( .A1(n3084), .A2(n4844), .B1(n4846), .B2(n4804), .C1(
        n4805), .C2(n4842), .ZN(n2642) );
  CKND0BWP12T U3853 ( .I(r1[26]), .ZN(n3085) );
  OAI222D0BWP12T U3854 ( .A1(n3085), .A2(n4844), .B1(n4842), .B2(n4775), .C1(
        n4776), .C2(n4846), .ZN(n2643) );
  CKND0BWP12T U3855 ( .I(r1[27]), .ZN(n3086) );
  OAI222D0BWP12T U3856 ( .A1(n3086), .A2(n4844), .B1(n4842), .B2(n4787), .C1(
        n4788), .C2(n4846), .ZN(n2644) );
  CKND0BWP12T U3857 ( .I(r1[28]), .ZN(n3087) );
  OAI222D0BWP12T U3858 ( .A1(n3087), .A2(n4844), .B1(n4842), .B2(n4806), .C1(
        n4807), .C2(n4846), .ZN(n2645) );
  CKND0BWP12T U3859 ( .I(r1[30]), .ZN(n3088) );
  OAI222D0BWP12T U3860 ( .A1(n3088), .A2(n4844), .B1(n4846), .B2(n4789), .C1(
        n4790), .C2(n4842), .ZN(n2647) );
  AOI22D0BWP12T U3861 ( .A1(next_pc_in[31]), .A2(n4743), .B1(n4744), .B2(
        pc_out[31]), .ZN(n3089) );
  AOI22D0BWP12T U3862 ( .A1(n4741), .A2(write2_in[31]), .B1(write1_in[31]), 
        .B2(n4742), .ZN(n3090) );
  CKND2D0BWP12T U3863 ( .A1(n3089), .A2(n3090), .ZN(n2232) );
  CKND0BWP12T U3864 ( .I(r1[5]), .ZN(n3091) );
  OAI222D0BWP12T U3865 ( .A1(n3091), .A2(n4844), .B1(n4842), .B2(n4838), .C1(
        n4840), .C2(n4846), .ZN(n2622) );
  CKND0BWP12T U3866 ( .I(r1[9]), .ZN(n3092) );
  OAI222D0BWP12T U3867 ( .A1(n3092), .A2(n4844), .B1(n4842), .B2(n4853), .C1(
        n4855), .C2(n4846), .ZN(n2626) );
  CKND0BWP12T U3868 ( .I(r1[15]), .ZN(n3093) );
  OAI222D0BWP12T U3869 ( .A1(n3093), .A2(n4844), .B1(n4842), .B2(n4829), .C1(
        n4831), .C2(n4846), .ZN(n2632) );
  CKND0BWP12T U3870 ( .I(r1[16]), .ZN(n3094) );
  OAI222D0BWP12T U3871 ( .A1(n3094), .A2(n4844), .B1(n4846), .B2(n4874), .C1(
        n4878), .C2(n4842), .ZN(n2633) );
  CKND0BWP12T U3872 ( .I(r1[23]), .ZN(n3095) );
  OAI222D0BWP12T U3873 ( .A1(n3095), .A2(n4844), .B1(n4842), .B2(n4832), .C1(
        n4834), .C2(n4846), .ZN(n2640) );
  CKND0BWP12T U3874 ( .I(r1[31]), .ZN(n3096) );
  OAI222D0BWP12T U3875 ( .A1(n3096), .A2(n4844), .B1(n4842), .B2(n4847), .C1(
        n4849), .C2(n4846), .ZN(n2648) );
  CKND0BWP12T U3876 ( .I(r0[0]), .ZN(n3097) );
  OAI222D0BWP12T U3877 ( .A1(n3097), .A2(n4877), .B1(n4875), .B2(n4859), .C1(
        n4861), .C2(n4879), .ZN(n2649) );
  CKND0BWP12T U3878 ( .I(r0[1]), .ZN(n3098) );
  OAI222D0BWP12T U3879 ( .A1(n3098), .A2(n4877), .B1(n4879), .B2(n4783), .C1(
        n4784), .C2(n4875), .ZN(n2650) );
  CKND0BWP12T U3880 ( .I(r0[2]), .ZN(n3099) );
  OAI222D0BWP12T U3881 ( .A1(n3099), .A2(n4877), .B1(n4875), .B2(n4862), .C1(
        n4866), .C2(n4879), .ZN(n2651) );
  CKND0BWP12T U3882 ( .I(r0[3]), .ZN(n3100) );
  OAI222D0BWP12T U3883 ( .A1(n3100), .A2(n4877), .B1(n4879), .B2(n4793), .C1(
        n4794), .C2(n4875), .ZN(n2652) );
  CKND0BWP12T U3884 ( .I(r0[4]), .ZN(n3101) );
  OAI222D0BWP12T U3885 ( .A1(n3101), .A2(n4877), .B1(n4879), .B2(n4800), .C1(
        n4801), .C2(n4875), .ZN(n2653) );
  CKND0BWP12T U3886 ( .I(r0[6]), .ZN(n3102) );
  OAI222D0BWP12T U3887 ( .A1(n3102), .A2(n4877), .B1(n4879), .B2(n4779), .C1(
        n4780), .C2(n4875), .ZN(n2655) );
  CKND0BWP12T U3888 ( .I(r0[7]), .ZN(n3103) );
  OAI222D0BWP12T U3889 ( .A1(n3103), .A2(n4877), .B1(n4875), .B2(n4798), .C1(
        n4799), .C2(n4879), .ZN(n2656) );
  CKND0BWP12T U3890 ( .I(r0[8]), .ZN(n3104) );
  OAI222D0BWP12T U3891 ( .A1(n3104), .A2(n4877), .B1(n4879), .B2(n4810), .C1(
        n4811), .C2(n4875), .ZN(n2657) );
  CKND0BWP12T U3892 ( .I(r0[10]), .ZN(n3105) );
  OAI222D0BWP12T U3893 ( .A1(n3105), .A2(n4877), .B1(n4875), .B2(n4808), .C1(
        n4809), .C2(n4879), .ZN(n2659) );
  CKND0BWP12T U3894 ( .I(r0[11]), .ZN(n3106) );
  OAI222D0BWP12T U3895 ( .A1(n3106), .A2(n4877), .B1(n4875), .B2(n4868), .C1(
        n4872), .C2(n4879), .ZN(n2660) );
  CKND0BWP12T U3896 ( .I(r0[12]), .ZN(n3107) );
  OAI222D0BWP12T U3897 ( .A1(n3107), .A2(n4877), .B1(n4879), .B2(n4850), .C1(
        n4852), .C2(n4875), .ZN(n2661) );
  CKND0BWP12T U3898 ( .I(r0[13]), .ZN(n3108) );
  OAI222D0BWP12T U3899 ( .A1(n3108), .A2(n4877), .B1(n4879), .B2(n4856), .C1(
        n4858), .C2(n4875), .ZN(n2662) );
  CKND0BWP12T U3900 ( .I(r0[14]), .ZN(n3109) );
  OAI222D0BWP12T U3901 ( .A1(n3109), .A2(n4877), .B1(n4875), .B2(n4802), .C1(
        n4803), .C2(n4879), .ZN(n2663) );
  CKND0BWP12T U3902 ( .I(r0[17]), .ZN(n3110) );
  OAI222D0BWP12T U3903 ( .A1(n3110), .A2(n4877), .B1(n4879), .B2(n4812), .C1(
        n4815), .C2(n4875), .ZN(n2666) );
  CKND0BWP12T U3904 ( .I(r0[18]), .ZN(n3111) );
  OAI222D0BWP12T U3905 ( .A1(n3111), .A2(n4877), .B1(n4875), .B2(n4791), .C1(
        n4792), .C2(n4879), .ZN(n2667) );
  CKND0BWP12T U3906 ( .I(r0[19]), .ZN(n3112) );
  OAI222D0BWP12T U3907 ( .A1(n3112), .A2(n4877), .B1(n4875), .B2(n4781), .C1(
        n4782), .C2(n4879), .ZN(n2668) );
  CKND0BWP12T U3908 ( .I(r0[20]), .ZN(n3113) );
  OAI222D0BWP12T U3909 ( .A1(n3113), .A2(n4877), .B1(n4875), .B2(n4880), .C1(
        n4884), .C2(n4879), .ZN(n2669) );
  CKND0BWP12T U3910 ( .I(r0[21]), .ZN(n3114) );
  OAI222D0BWP12T U3911 ( .A1(n3114), .A2(n4877), .B1(n4879), .B2(n4777), .C1(
        n4778), .C2(n4875), .ZN(n2670) );
  CKND0BWP12T U3912 ( .I(r0[22]), .ZN(n3115) );
  OAI222D0BWP12T U3913 ( .A1(n3115), .A2(n4877), .B1(n4879), .B2(n4785), .C1(
        n4786), .C2(n4875), .ZN(n2671) );
  CKND0BWP12T U3914 ( .I(r0[24]), .ZN(n3116) );
  OAI222D0BWP12T U3915 ( .A1(n3116), .A2(n4877), .B1(n4879), .B2(n4841), .C1(
        n4845), .C2(n4875), .ZN(n2673) );
  CKND0BWP12T U3916 ( .I(r0[25]), .ZN(n3117) );
  OAI222D0BWP12T U3917 ( .A1(n3117), .A2(n4877), .B1(n4875), .B2(n4804), .C1(
        n4805), .C2(n4879), .ZN(n2674) );
  CKND0BWP12T U3918 ( .I(r0[26]), .ZN(n3118) );
  OAI222D0BWP12T U3919 ( .A1(n3118), .A2(n4877), .B1(n4879), .B2(n4775), .C1(
        n4776), .C2(n4875), .ZN(n2675) );
  CKND0BWP12T U3920 ( .I(r0[27]), .ZN(n3119) );
  OAI222D0BWP12T U3921 ( .A1(n3119), .A2(n4877), .B1(n4879), .B2(n4787), .C1(
        n4788), .C2(n4875), .ZN(n2676) );
  CKND0BWP12T U3922 ( .I(r0[28]), .ZN(n3120) );
  OAI222D0BWP12T U3923 ( .A1(n3120), .A2(n4877), .B1(n4879), .B2(n4806), .C1(
        n4807), .C2(n4875), .ZN(n2677) );
  CKND0BWP12T U3924 ( .I(r0[29]), .ZN(n3121) );
  OAI222D0BWP12T U3925 ( .A1(n3121), .A2(n4877), .B1(n4879), .B2(n4835), .C1(
        n4837), .C2(n4875), .ZN(n2678) );
  CKND0BWP12T U3926 ( .I(r0[30]), .ZN(n3122) );
  OAI222D0BWP12T U3927 ( .A1(n3122), .A2(n4877), .B1(n4875), .B2(n4789), .C1(
        n4790), .C2(n4879), .ZN(n2679) );
  IND2XD1BWP12T U3928 ( .A1(n3125), .B1(write1_sel[3]), .ZN(n3128) );
  INR2XD0BWP12T U3929 ( .A1(write1_sel[1]), .B1(write1_sel[2]), .ZN(n3129) );
  INVD0BWP12T U3930 ( .I(n3126), .ZN(n3127) );
  NR2XD0BWP12T U3931 ( .A1(n3149), .A2(n3135), .ZN(n3130) );
  NR2XD0BWP12T U3932 ( .A1(write1_sel[0]), .A2(n3128), .ZN(n3137) );
  AN2XD1BWP12T U3933 ( .A1(write1_sel[1]), .A2(write1_sel[2]), .Z(n4753) );
  IND2XD1BWP12T U3934 ( .A1(n3132), .B1(n4873), .ZN(n4871) );
  IND2XD1BWP12T U3935 ( .A1(n3136), .B1(n4823), .ZN(n4825) );
  IND2XD1BWP12T U3936 ( .A1(n3138), .B1(n4867), .ZN(n4865) );
  AN4D0BWP12T U3937 ( .A1(n3142), .A2(n4753), .A3(write1_sel[3]), .A4(
        write1_sel[4]), .Z(n3143) );
  AN2D1BWP12T U3938 ( .A1(n4678), .A2(n4764), .Z(n3157) );
  NR2D1BWP12T U3939 ( .A1(n4679), .A2(n4757), .ZN(n3154) );
  INR2D1BWP12T U3940 ( .A1(n3154), .B1(n3157), .ZN(n3156) );
  NR2D1BWP12T U3941 ( .A1(n3157), .A2(n3154), .ZN(n3155) );
  AO222D1BWP12T U3942 ( .A1(write1_in[5]), .A2(n3157), .B1(write2_in[5]), .B2(
        n3156), .C1(n3155), .C2(next_sp_in[5]), .Z(spin[5]) );
  AO222D1BWP12T U3943 ( .A1(write1_in[4]), .A2(n3157), .B1(write2_in[4]), .B2(
        n3156), .C1(n3155), .C2(next_sp_in[4]), .Z(spin[4]) );
  AO222D1BWP12T U3944 ( .A1(write1_in[31]), .A2(n3157), .B1(write2_in[31]), 
        .B2(n3156), .C1(n3155), .C2(next_sp_in[31]), .Z(spin[31]) );
  AO222D1BWP12T U3945 ( .A1(write2_in[30]), .A2(n3156), .B1(n3157), .B2(
        write1_in[30]), .C1(n3155), .C2(next_sp_in[30]), .Z(spin[30]) );
  AO222D1BWP12T U3946 ( .A1(write1_in[29]), .A2(n3157), .B1(write2_in[29]), 
        .B2(n3156), .C1(n3155), .C2(next_sp_in[29]), .Z(spin[29]) );
  AO222D1BWP12T U3947 ( .A1(write1_in[28]), .A2(n3157), .B1(write2_in[28]), 
        .B2(n3156), .C1(n3155), .C2(next_sp_in[28]), .Z(spin[28]) );
  AO222D1BWP12T U3948 ( .A1(write1_in[27]), .A2(n3157), .B1(write2_in[27]), 
        .B2(n3156), .C1(n3155), .C2(next_sp_in[27]), .Z(spin[27]) );
  AO222D1BWP12T U3949 ( .A1(write1_in[26]), .A2(n3157), .B1(write2_in[26]), 
        .B2(n3156), .C1(n3155), .C2(next_sp_in[26]), .Z(spin[26]) );
  AO222D1BWP12T U3950 ( .A1(write2_in[25]), .A2(n3156), .B1(n3157), .B2(
        write1_in[25]), .C1(n3155), .C2(next_sp_in[25]), .Z(spin[25]) );
  AO222D1BWP12T U3951 ( .A1(write1_in[24]), .A2(n3157), .B1(write2_in[24]), 
        .B2(n3156), .C1(n3155), .C2(next_sp_in[24]), .Z(spin[24]) );
  AO222D1BWP12T U3952 ( .A1(write1_in[23]), .A2(n3157), .B1(write2_in[23]), 
        .B2(n3156), .C1(n3155), .C2(next_sp_in[23]), .Z(spin[23]) );
  AO222D1BWP12T U3953 ( .A1(write1_in[22]), .A2(n3157), .B1(write2_in[22]), 
        .B2(n3156), .C1(n3155), .C2(next_sp_in[22]), .Z(spin[22]) );
  AO222D1BWP12T U3954 ( .A1(write1_in[21]), .A2(n3157), .B1(write2_in[21]), 
        .B2(n3156), .C1(n3155), .C2(next_sp_in[21]), .Z(spin[21]) );
  AO222D1BWP12T U3955 ( .A1(write2_in[20]), .A2(n3156), .B1(n3157), .B2(
        write1_in[20]), .C1(n3155), .C2(next_sp_in[20]), .Z(spin[20]) );
  AO222D1BWP12T U3956 ( .A1(write2_in[19]), .A2(n3156), .B1(n3157), .B2(
        write1_in[19]), .C1(n3155), .C2(next_sp_in[19]), .Z(spin[19]) );
  AO222D1BWP12T U3957 ( .A1(write2_in[18]), .A2(n3156), .B1(n3157), .B2(
        write1_in[18]), .C1(n3155), .C2(next_sp_in[18]), .Z(spin[18]) );
  AO222D1BWP12T U3958 ( .A1(write1_in[17]), .A2(n3157), .B1(write2_in[17]), 
        .B2(n3156), .C1(n3155), .C2(next_sp_in[17]), .Z(spin[17]) );
  AO222D1BWP12T U3959 ( .A1(write2_in[16]), .A2(n3156), .B1(n3157), .B2(
        write1_in[16]), .C1(n3155), .C2(next_sp_in[16]), .Z(spin[16]) );
  AO222D1BWP12T U3960 ( .A1(write1_in[15]), .A2(n3157), .B1(write2_in[15]), 
        .B2(n3156), .C1(n3155), .C2(next_sp_in[15]), .Z(spin[15]) );
  AO222D1BWP12T U3961 ( .A1(write2_in[14]), .A2(n3156), .B1(n3157), .B2(
        write1_in[14]), .C1(n3155), .C2(next_sp_in[14]), .Z(spin[14]) );
  AO222D1BWP12T U3962 ( .A1(write1_in[13]), .A2(n3157), .B1(write2_in[13]), 
        .B2(n3156), .C1(n3155), .C2(next_sp_in[13]), .Z(spin[13]) );
  AO222D1BWP12T U3963 ( .A1(write1_in[12]), .A2(n3157), .B1(write2_in[12]), 
        .B2(n3156), .C1(n3155), .C2(next_sp_in[12]), .Z(spin[12]) );
  AO222D1BWP12T U3964 ( .A1(write2_in[11]), .A2(n3156), .B1(n3157), .B2(
        write1_in[11]), .C1(n3155), .C2(next_sp_in[11]), .Z(spin[11]) );
  AO222D1BWP12T U3965 ( .A1(write2_in[10]), .A2(n3156), .B1(n3157), .B2(
        write1_in[10]), .C1(n3155), .C2(next_sp_in[10]), .Z(spin[10]) );
  AO222D1BWP12T U3966 ( .A1(write1_in[9]), .A2(n3157), .B1(write2_in[9]), .B2(
        n3156), .C1(n3155), .C2(next_sp_in[9]), .Z(spin[9]) );
  AO222D1BWP12T U3967 ( .A1(write1_in[8]), .A2(n3157), .B1(write2_in[8]), .B2(
        n3156), .C1(n3155), .C2(next_sp_in[8]), .Z(spin[8]) );
  AO222D1BWP12T U3968 ( .A1(write2_in[7]), .A2(n3156), .B1(n3157), .B2(
        write1_in[7]), .C1(n3155), .C2(next_sp_in[7]), .Z(spin[7]) );
  AO222D1BWP12T U3969 ( .A1(write1_in[6]), .A2(n3157), .B1(write2_in[6]), .B2(
        n3156), .C1(n3155), .C2(next_sp_in[6]), .Z(spin[6]) );
  AO222D1BWP12T U3970 ( .A1(write2_in[0]), .A2(n3156), .B1(n3157), .B2(
        write1_in[0]), .C1(n3155), .C2(next_sp_in[0]), .Z(spin[0]) );
  AO222D1BWP12T U3971 ( .A1(write2_in[2]), .A2(n3156), .B1(n3157), .B2(
        write1_in[2]), .C1(n3155), .C2(next_sp_in[2]), .Z(spin[2]) );
  AO222D1BWP12T U3972 ( .A1(write1_in[3]), .A2(n3157), .B1(write2_in[3]), .B2(
        n3156), .C1(n3155), .C2(next_sp_in[3]), .Z(spin[3]) );
  AO222D1BWP12T U3973 ( .A1(write1_in[1]), .A2(n3157), .B1(write2_in[1]), .B2(
        n3156), .C1(n3155), .C2(next_sp_in[1]), .Z(spin[1]) );
  INVD1BWP12T U3974 ( .I(readB_sel[0]), .ZN(n3161) );
  ND4D1BWP12T U3975 ( .A1(readB_sel[3]), .A2(readB_sel[4]), .A3(readB_sel[1]), 
        .A4(readB_sel[2]), .ZN(n3170) );
  NR2D1BWP12T U3976 ( .A1(n3161), .A2(n3170), .ZN(n4269) );
  NR2D1BWP12T U3977 ( .A1(readB_sel[3]), .A2(readB_sel[4]), .ZN(n3158) );
  ND2D1BWP12T U3978 ( .A1(readB_sel[0]), .A2(n3158), .ZN(n3164) );
  INVD1BWP12T U3979 ( .I(readB_sel[1]), .ZN(n3160) );
  ND2D1BWP12T U3980 ( .A1(readB_sel[2]), .A2(n3160), .ZN(n3167) );
  NR2D1BWP12T U3981 ( .A1(n3164), .A2(n3167), .ZN(n4256) );
  AOI22D1BWP12T U3982 ( .A1(n4269), .A2(immediate2_in[28]), .B1(n4256), .B2(
        r5[28]), .ZN(n3182) );
  INR2D1BWP12T U3983 ( .A1(readB_sel[3]), .B1(readB_sel[4]), .ZN(n3162) );
  ND2D1BWP12T U3984 ( .A1(readB_sel[0]), .A2(n3162), .ZN(n3165) );
  NR2D1BWP12T U3985 ( .A1(n3165), .A2(n3167), .ZN(n4266) );
  INVD1BWP12T U3986 ( .I(readB_sel[2]), .ZN(n3159) );
  ND2D1BWP12T U3987 ( .A1(readB_sel[1]), .A2(n3159), .ZN(n3166) );
  ND2D1BWP12T U3988 ( .A1(n3158), .A2(n3161), .ZN(n3169) );
  NR2D1BWP12T U3989 ( .A1(n3166), .A2(n3169), .ZN(n4268) );
  AOI22D1BWP12T U3990 ( .A1(n4266), .A2(sp_out[28]), .B1(n4268), .B2(r2[28]), 
        .ZN(n3181) );
  NR2D1BWP12T U3991 ( .A1(n3169), .A2(n3167), .ZN(n4265) );
  ND2D1BWP12T U3992 ( .A1(readB_sel[1]), .A2(readB_sel[2]), .ZN(n3168) );
  NR2D1BWP12T U3993 ( .A1(n3164), .A2(n3168), .ZN(n4259) );
  AOI22D1BWP12T U3994 ( .A1(n4265), .A2(r4[28]), .B1(n4259), .B2(r7[28]), .ZN(
        n3180) );
  NR2D1BWP12T U3995 ( .A1(n3165), .A2(n3166), .ZN(n4276) );
  NR2D1BWP12T U3996 ( .A1(n3165), .A2(n3168), .ZN(n3486) );
  INVD1BWP12T U3997 ( .I(n3486), .ZN(n4263) );
  INVD1BWP12T U3998 ( .I(pc_out[28]), .ZN(n4630) );
  ND2D1BWP12T U3999 ( .A1(n3160), .A2(n3159), .ZN(n3172) );
  NR2D1BWP12T U4000 ( .A1(n3172), .A2(n3169), .ZN(n4229) );
  ND2D1BWP12T U4001 ( .A1(n3162), .A2(n3161), .ZN(n3171) );
  NR2D1BWP12T U4002 ( .A1(n3168), .A2(n3171), .ZN(n4267) );
  INVD1BWP12T U4003 ( .I(n4267), .ZN(n3488) );
  AOI22D1BWP12T U4004 ( .A1(n4229), .A2(r0[28]), .B1(n4267), .B2(lr[28]), .ZN(
        n3163) );
  OAI21D1BWP12T U4005 ( .A1(n4263), .A2(n4630), .B(n3163), .ZN(n3178) );
  NR2D1BWP12T U4006 ( .A1(n3172), .A2(n3164), .ZN(n4255) );
  NR2D1BWP12T U4007 ( .A1(n3166), .A2(n3164), .ZN(n3462) );
  AOI22D1BWP12T U4008 ( .A1(n4255), .A2(r1[28]), .B1(n3462), .B2(r3[28]), .ZN(
        n3176) );
  NR2D1BWP12T U4009 ( .A1(n3165), .A2(n3172), .ZN(n4260) );
  NR2D1BWP12T U4010 ( .A1(n3166), .A2(n3171), .ZN(n4257) );
  AOI22D1BWP12T U4011 ( .A1(n4260), .A2(r9[28]), .B1(n4257), .B2(r10[28]), 
        .ZN(n3175) );
  NR2D1BWP12T U4012 ( .A1(n3167), .A2(n3171), .ZN(n4258) );
  NR2D1BWP12T U4013 ( .A1(n3169), .A2(n3168), .ZN(n4230) );
  AOI22D1BWP12T U4014 ( .A1(n4258), .A2(r12[28]), .B1(n4230), .B2(r6[28]), 
        .ZN(n3174) );
  NR2D1BWP12T U4015 ( .A1(readB_sel[0]), .A2(n3170), .ZN(n4254) );
  NR2D1BWP12T U4016 ( .A1(n3172), .A2(n3171), .ZN(n4264) );
  INVD1BWP12T U4017 ( .I(n4264), .ZN(n3475) );
  AOI22D1BWP12T U4018 ( .A1(n4254), .A2(tmp1[28]), .B1(n4264), .B2(r8[28]), 
        .ZN(n3173) );
  ND4D1BWP12T U4019 ( .A1(n3176), .A2(n3175), .A3(n3174), .A4(n3173), .ZN(
        n3177) );
  AOI211D1BWP12T U4020 ( .A1(n4276), .A2(r11[28]), .B(n3178), .C(n3177), .ZN(
        n3179) );
  ND4D1BWP12T U4021 ( .A1(n3182), .A2(n3181), .A3(n3180), .A4(n3179), .ZN(
        regB_out[28]) );
  INVD1BWP12T U4022 ( .I(readA_sel[2]), .ZN(n3183) );
  ND2D1BWP12T U4023 ( .A1(readA_sel[1]), .A2(n3183), .ZN(n3192) );
  NR2D1BWP12T U4024 ( .A1(readA_sel[3]), .A2(readA_sel[4]), .ZN(n3184) );
  INVD1BWP12T U4025 ( .I(readA_sel[0]), .ZN(n3187) );
  ND2D1BWP12T U4026 ( .A1(n3184), .A2(n3187), .ZN(n3195) );
  NR2D1BWP12T U4027 ( .A1(n3192), .A2(n3195), .ZN(n4674) );
  INVD1BWP12T U4028 ( .I(readA_sel[1]), .ZN(n3185) );
  ND2D1BWP12T U4029 ( .A1(n3183), .A2(n3185), .ZN(n3196) );
  ND2D1BWP12T U4030 ( .A1(readA_sel[0]), .A2(n3184), .ZN(n3191) );
  NR2D1BWP12T U4031 ( .A1(n3196), .A2(n3191), .ZN(n4615) );
  AOI22D1BWP12T U4032 ( .A1(r2[31]), .A2(n4674), .B1(r1[31]), .B2(n4615), .ZN(
        n3208) );
  ND2D1BWP12T U4033 ( .A1(readA_sel[2]), .A2(n3185), .ZN(n3197) );
  NR2D1BWP12T U4034 ( .A1(n3197), .A2(n3195), .ZN(n4663) );
  ND2D1BWP12T U4035 ( .A1(readA_sel[2]), .A2(readA_sel[1]), .ZN(n3189) );
  NR2D1BWP12T U4036 ( .A1(n3195), .A2(n3189), .ZN(n4667) );
  AOI22D1BWP12T U4037 ( .A1(r4[31]), .A2(n4663), .B1(r6[31]), .B2(n4667), .ZN(
        n3207) );
  NR2D1BWP12T U4038 ( .A1(n3191), .A2(n3189), .ZN(n4656) );
  ND4D1BWP12T U4039 ( .A1(readA_sel[2]), .A2(readA_sel[1]), .A3(readA_sel[3]), 
        .A4(readA_sel[4]), .ZN(n3193) );
  NR2D1BWP12T U4040 ( .A1(n3187), .A2(n3193), .ZN(n3186) );
  AOI22D1BWP12T U4041 ( .A1(r7[31]), .A2(n4656), .B1(n3186), .B2(
        immediate1_in[31]), .ZN(n3206) );
  INR2D1BWP12T U4042 ( .A1(readA_sel[3]), .B1(readA_sel[4]), .ZN(n3188) );
  ND2D1BWP12T U4043 ( .A1(n3188), .A2(n3187), .ZN(n3198) );
  OR2XD1BWP12T U4044 ( .A1(n3198), .A2(n3189), .Z(n4601) );
  INVD1BWP12T U4045 ( .I(pc_out[31]), .ZN(n4262) );
  ND2D1BWP12T U4046 ( .A1(readA_sel[0]), .A2(n3188), .ZN(n3194) );
  NR2D1BWP12T U4047 ( .A1(n3194), .A2(n3189), .ZN(n4658) );
  INVD1BWP12T U4048 ( .I(n4658), .ZN(n4641) );
  NR2D1BWP12T U4049 ( .A1(n3192), .A2(n3198), .ZN(n4665) );
  NR2D1BWP12T U4050 ( .A1(n3191), .A2(n3197), .ZN(n4664) );
  AOI22D1BWP12T U4051 ( .A1(r10[31]), .A2(n4665), .B1(r5[31]), .B2(n4664), 
        .ZN(n3190) );
  OAI21D1BWP12T U4052 ( .A1(n4262), .A2(n4641), .B(n3190), .ZN(n3204) );
  NR2D1BWP12T U4053 ( .A1(n3192), .A2(n3191), .ZN(n4589) );
  NR2D1BWP12T U4054 ( .A1(n3192), .A2(n3194), .ZN(n4659) );
  AOI22D1BWP12T U4055 ( .A1(r3[31]), .A2(n4589), .B1(r11[31]), .B2(n4659), 
        .ZN(n3202) );
  NR2D1BWP12T U4056 ( .A1(n3194), .A2(n3197), .ZN(n4655) );
  NR2D1BWP12T U4057 ( .A1(readA_sel[0]), .A2(n3193), .ZN(n4657) );
  AOI22D1BWP12T U4058 ( .A1(sp_out[31]), .A2(n4655), .B1(tmp1[31]), .B2(n4657), 
        .ZN(n3201) );
  NR2D1BWP12T U4059 ( .A1(n3196), .A2(n3194), .ZN(n4666) );
  NR2D1BWP12T U4060 ( .A1(n3196), .A2(n3195), .ZN(n4626) );
  AOI22D1BWP12T U4061 ( .A1(r9[31]), .A2(n4666), .B1(r0[31]), .B2(n4626), .ZN(
        n3200) );
  NR2D1BWP12T U4062 ( .A1(n3198), .A2(n3196), .ZN(n4627) );
  NR2D1BWP12T U4063 ( .A1(n3198), .A2(n3197), .ZN(n4654) );
  AOI22D1BWP12T U4064 ( .A1(r8[31]), .A2(n4627), .B1(r12[31]), .B2(n4654), 
        .ZN(n3199) );
  ND4D1BWP12T U4065 ( .A1(n3202), .A2(n3201), .A3(n3200), .A4(n3199), .ZN(
        n3203) );
  AOI211D1BWP12T U4066 ( .A1(lr[31]), .A2(n4653), .B(n3204), .C(n3203), .ZN(
        n3205) );
  ND4D1BWP12T U4067 ( .A1(n3208), .A2(n3207), .A3(n3206), .A4(n3205), .ZN(
        regA_out[31]) );
  AOI22D1BWP12T U4068 ( .A1(n3462), .A2(r3[23]), .B1(n4267), .B2(lr[23]), .ZN(
        n3219) );
  AOI22D1BWP12T U4069 ( .A1(n4258), .A2(r12[23]), .B1(n4265), .B2(r4[23]), 
        .ZN(n3218) );
  AOI22D1BWP12T U4070 ( .A1(n4266), .A2(sp_out[23]), .B1(n4264), .B2(r8[23]), 
        .ZN(n3217) );
  INVD1BWP12T U4071 ( .I(pc_out[23]), .ZN(n4564) );
  AOI22D1BWP12T U4072 ( .A1(n4254), .A2(tmp1[23]), .B1(n4256), .B2(r5[23]), 
        .ZN(n3209) );
  OAI21D1BWP12T U4073 ( .A1(n4263), .A2(n4564), .B(n3209), .ZN(n3215) );
  AOI22D1BWP12T U4074 ( .A1(n4269), .A2(immediate2_in[23]), .B1(n4230), .B2(
        r6[23]), .ZN(n3213) );
  AOI22D1BWP12T U4075 ( .A1(n4260), .A2(r9[23]), .B1(n4259), .B2(r7[23]), .ZN(
        n3212) );
  AOI22D1BWP12T U4076 ( .A1(n4255), .A2(r1[23]), .B1(n4268), .B2(r2[23]), .ZN(
        n3211) );
  AOI22D1BWP12T U4077 ( .A1(n4276), .A2(r11[23]), .B1(n4257), .B2(r10[23]), 
        .ZN(n3210) );
  ND4D1BWP12T U4078 ( .A1(n3213), .A2(n3212), .A3(n3211), .A4(n3210), .ZN(
        n3214) );
  AOI211D1BWP12T U4079 ( .A1(n4229), .A2(r0[23]), .B(n3215), .C(n3214), .ZN(
        n3216) );
  ND4D1BWP12T U4080 ( .A1(n3219), .A2(n3218), .A3(n3217), .A4(n3216), .ZN(
        regB_out[23]) );
  AOI22D1BWP12T U4081 ( .A1(n4257), .A2(r10[22]), .B1(n4265), .B2(r4[22]), 
        .ZN(n3230) );
  AOI22D1BWP12T U4082 ( .A1(n4276), .A2(r11[22]), .B1(n4264), .B2(r8[22]), 
        .ZN(n3229) );
  AOI22D1BWP12T U4083 ( .A1(n4269), .A2(immediate2_in[22]), .B1(n3462), .B2(
        r3[22]), .ZN(n3228) );
  INVD1BWP12T U4084 ( .I(pc_out[22]), .ZN(n4552) );
  AOI22D1BWP12T U4085 ( .A1(n4259), .A2(r7[22]), .B1(n4268), .B2(r2[22]), .ZN(
        n3220) );
  OAI21D1BWP12T U4086 ( .A1(n4263), .A2(n4552), .B(n3220), .ZN(n3226) );
  AOI22D1BWP12T U4087 ( .A1(n4260), .A2(r9[22]), .B1(n4255), .B2(r1[22]), .ZN(
        n3224) );
  AOI22D1BWP12T U4088 ( .A1(n4254), .A2(tmp1[22]), .B1(n4256), .B2(r5[22]), 
        .ZN(n3223) );
  AOI22D1BWP12T U4089 ( .A1(n4229), .A2(r0[22]), .B1(n4258), .B2(r12[22]), 
        .ZN(n3222) );
  AOI22D1BWP12T U4090 ( .A1(n4230), .A2(r6[22]), .B1(n4267), .B2(lr[22]), .ZN(
        n3221) );
  ND4D1BWP12T U4091 ( .A1(n3224), .A2(n3223), .A3(n3222), .A4(n3221), .ZN(
        n3225) );
  AOI211D1BWP12T U4092 ( .A1(n4266), .A2(sp_out[22]), .B(n3226), .C(n3225), 
        .ZN(n3227) );
  ND4D1BWP12T U4093 ( .A1(n3230), .A2(n3229), .A3(n3228), .A4(n3227), .ZN(
        regB_out[22]) );
  AOI22D1BWP12T U4094 ( .A1(n4254), .A2(tmp1[21]), .B1(n4258), .B2(r12[21]), 
        .ZN(n3241) );
  AOI22D1BWP12T U4095 ( .A1(n4229), .A2(r0[21]), .B1(n4268), .B2(r2[21]), .ZN(
        n3240) );
  AOI22D1BWP12T U4096 ( .A1(n4265), .A2(r4[21]), .B1(n4256), .B2(r5[21]), .ZN(
        n3239) );
  INVD1BWP12T U4097 ( .I(pc_out[21]), .ZN(n4541) );
  AOI22D1BWP12T U4098 ( .A1(n3462), .A2(r3[21]), .B1(n4267), .B2(lr[21]), .ZN(
        n3231) );
  OAI21D1BWP12T U4099 ( .A1(n4263), .A2(n4541), .B(n3231), .ZN(n3237) );
  AOI22D1BWP12T U4100 ( .A1(n4255), .A2(r1[21]), .B1(n4230), .B2(r6[21]), .ZN(
        n3235) );
  AOI22D1BWP12T U4101 ( .A1(n4276), .A2(r11[21]), .B1(n4266), .B2(sp_out[21]), 
        .ZN(n3234) );
  AOI22D1BWP12T U4102 ( .A1(n4264), .A2(r8[21]), .B1(n4259), .B2(r7[21]), .ZN(
        n3233) );
  AOI22D1BWP12T U4103 ( .A1(n4269), .A2(immediate2_in[21]), .B1(n4257), .B2(
        r10[21]), .ZN(n3232) );
  ND4D1BWP12T U4104 ( .A1(n3235), .A2(n3234), .A3(n3233), .A4(n3232), .ZN(
        n3236) );
  AOI211D1BWP12T U4105 ( .A1(n4260), .A2(r9[21]), .B(n3237), .C(n3236), .ZN(
        n3238) );
  ND4D1BWP12T U4106 ( .A1(n3241), .A2(n3240), .A3(n3239), .A4(n3238), .ZN(
        regB_out[21]) );
  AOI22D1BWP12T U4107 ( .A1(n4255), .A2(r1[20]), .B1(n4258), .B2(r12[20]), 
        .ZN(n3252) );
  AOI22D1BWP12T U4108 ( .A1(n4254), .A2(tmp1[20]), .B1(n4256), .B2(r5[20]), 
        .ZN(n3251) );
  AOI22D1BWP12T U4109 ( .A1(n4257), .A2(r10[20]), .B1(n4264), .B2(r8[20]), 
        .ZN(n3250) );
  INVD1BWP12T U4110 ( .I(pc_out[20]), .ZN(n4528) );
  AOI22D1BWP12T U4111 ( .A1(n4268), .A2(r2[20]), .B1(n4230), .B2(r6[20]), .ZN(
        n3242) );
  OAI21D1BWP12T U4112 ( .A1(n4263), .A2(n4528), .B(n3242), .ZN(n3248) );
  AOI22D1BWP12T U4113 ( .A1(n4265), .A2(r4[20]), .B1(n4259), .B2(r7[20]), .ZN(
        n3246) );
  AOI22D1BWP12T U4114 ( .A1(n4276), .A2(r11[20]), .B1(n4269), .B2(
        immediate2_in[20]), .ZN(n3245) );
  AOI22D1BWP12T U4115 ( .A1(n4229), .A2(r0[20]), .B1(n3462), .B2(r3[20]), .ZN(
        n3244) );
  AOI22D1BWP12T U4116 ( .A1(n4260), .A2(r9[20]), .B1(n4267), .B2(lr[20]), .ZN(
        n3243) );
  ND4D1BWP12T U4117 ( .A1(n3246), .A2(n3245), .A3(n3244), .A4(n3243), .ZN(
        n3247) );
  AOI211D1BWP12T U4118 ( .A1(n4266), .A2(sp_out[20]), .B(n3248), .C(n3247), 
        .ZN(n3249) );
  ND4D1BWP12T U4119 ( .A1(n3252), .A2(n3251), .A3(n3250), .A4(n3249), .ZN(
        regB_out[20]) );
  AOI22D1BWP12T U4120 ( .A1(n4256), .A2(r5[19]), .B1(n4230), .B2(r6[19]), .ZN(
        n3263) );
  AOI22D1BWP12T U4121 ( .A1(n4254), .A2(tmp1[19]), .B1(n4259), .B2(r7[19]), 
        .ZN(n3262) );
  AOI22D1BWP12T U4122 ( .A1(n3486), .A2(pc_out[19]), .B1(n4266), .B2(
        sp_out[19]), .ZN(n3254) );
  AOI22D1BWP12T U4123 ( .A1(n4268), .A2(r2[19]), .B1(n3462), .B2(r3[19]), .ZN(
        n3253) );
  OAI211D1BWP12T U4124 ( .A1(n3488), .A2(n4516), .B(n3254), .C(n3253), .ZN(
        n3260) );
  AOI22D1BWP12T U4125 ( .A1(n4255), .A2(r1[19]), .B1(n4229), .B2(r0[19]), .ZN(
        n3258) );
  AOI22D1BWP12T U4126 ( .A1(n4276), .A2(r11[19]), .B1(n4269), .B2(
        immediate2_in[19]), .ZN(n3257) );
  AOI22D1BWP12T U4127 ( .A1(n4257), .A2(r10[19]), .B1(n4264), .B2(r8[19]), 
        .ZN(n3256) );
  AOI22D1BWP12T U4128 ( .A1(n4260), .A2(r9[19]), .B1(n4258), .B2(r12[19]), 
        .ZN(n3255) );
  ND4D1BWP12T U4129 ( .A1(n3258), .A2(n3257), .A3(n3256), .A4(n3255), .ZN(
        n3259) );
  AOI211D1BWP12T U4130 ( .A1(n4265), .A2(r4[19]), .B(n3260), .C(n3259), .ZN(
        n3261) );
  ND3D1BWP12T U4131 ( .A1(n3263), .A2(n3262), .A3(n3261), .ZN(regB_out[19]) );
  AOI22D1BWP12T U4132 ( .A1(n4269), .A2(immediate2_in[18]), .B1(n4259), .B2(
        r7[18]), .ZN(n3274) );
  AOI22D1BWP12T U4133 ( .A1(n3486), .A2(pc_out[18]), .B1(n3462), .B2(r3[18]), 
        .ZN(n3273) );
  AOI22D1BWP12T U4134 ( .A1(n4258), .A2(r12[18]), .B1(n4230), .B2(r6[18]), 
        .ZN(n3272) );
  AOI22D1BWP12T U4135 ( .A1(n4229), .A2(r0[18]), .B1(n4254), .B2(tmp1[18]), 
        .ZN(n3264) );
  OAI21D1BWP12T U4136 ( .A1(n3488), .A2(n4504), .B(n3264), .ZN(n3270) );
  AOI22D1BWP12T U4137 ( .A1(n4265), .A2(r4[18]), .B1(n4256), .B2(r5[18]), .ZN(
        n3268) );
  AOI22D1BWP12T U4138 ( .A1(n4266), .A2(sp_out[18]), .B1(n4257), .B2(r10[18]), 
        .ZN(n3267) );
  AOI22D1BWP12T U4139 ( .A1(n4264), .A2(r8[18]), .B1(n4268), .B2(r2[18]), .ZN(
        n3266) );
  AOI22D1BWP12T U4140 ( .A1(n4276), .A2(r11[18]), .B1(n4260), .B2(r9[18]), 
        .ZN(n3265) );
  ND4D1BWP12T U4141 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(
        n3269) );
  AOI211D1BWP12T U4142 ( .A1(n4255), .A2(r1[18]), .B(n3270), .C(n3269), .ZN(
        n3271) );
  ND4D1BWP12T U4143 ( .A1(n3274), .A2(n3273), .A3(n3272), .A4(n3271), .ZN(
        regB_out[18]) );
  AOI22D1BWP12T U4144 ( .A1(n4254), .A2(tmp1[17]), .B1(n4267), .B2(lr[17]), 
        .ZN(n3285) );
  AOI22D1BWP12T U4145 ( .A1(n4255), .A2(r1[17]), .B1(n4268), .B2(r2[17]), .ZN(
        n3284) );
  AOI22D1BWP12T U4146 ( .A1(n4276), .A2(r11[17]), .B1(n4259), .B2(r7[17]), 
        .ZN(n3276) );
  AOI22D1BWP12T U4147 ( .A1(n3486), .A2(pc_out[17]), .B1(n4257), .B2(r10[17]), 
        .ZN(n3275) );
  OAI211D1BWP12T U4148 ( .A1(n3475), .A2(n4492), .B(n3276), .C(n3275), .ZN(
        n3282) );
  AOI22D1BWP12T U4149 ( .A1(n4229), .A2(r0[17]), .B1(n4265), .B2(r4[17]), .ZN(
        n3280) );
  AOI22D1BWP12T U4150 ( .A1(n4266), .A2(sp_out[17]), .B1(n4256), .B2(r5[17]), 
        .ZN(n3279) );
  AOI22D1BWP12T U4151 ( .A1(n3462), .A2(r3[17]), .B1(n4230), .B2(r6[17]), .ZN(
        n3278) );
  AOI22D1BWP12T U4152 ( .A1(n4269), .A2(immediate2_in[17]), .B1(n4258), .B2(
        r12[17]), .ZN(n3277) );
  ND4D1BWP12T U4153 ( .A1(n3280), .A2(n3279), .A3(n3278), .A4(n3277), .ZN(
        n3281) );
  AOI211D1BWP12T U4154 ( .A1(n4260), .A2(r9[17]), .B(n3282), .C(n3281), .ZN(
        n3283) );
  ND3D1BWP12T U4155 ( .A1(n3285), .A2(n3284), .A3(n3283), .ZN(regB_out[17]) );
  AOI22D1BWP12T U4156 ( .A1(n4266), .A2(sp_out[16]), .B1(n4268), .B2(r2[16]), 
        .ZN(n3296) );
  AOI22D1BWP12T U4157 ( .A1(n4260), .A2(r9[16]), .B1(n4229), .B2(r0[16]), .ZN(
        n3295) );
  AOI22D1BWP12T U4158 ( .A1(n4276), .A2(r11[16]), .B1(n4255), .B2(r1[16]), 
        .ZN(n3294) );
  INVD1BWP12T U4159 ( .I(pc_out[16]), .ZN(n4481) );
  AOI22D1BWP12T U4160 ( .A1(n4264), .A2(r8[16]), .B1(n3462), .B2(r3[16]), .ZN(
        n3286) );
  OAI21D1BWP12T U4161 ( .A1(n4263), .A2(n4481), .B(n3286), .ZN(n3292) );
  AOI22D1BWP12T U4162 ( .A1(n4257), .A2(r10[16]), .B1(n4267), .B2(lr[16]), 
        .ZN(n3290) );
  AOI22D1BWP12T U4163 ( .A1(n4269), .A2(immediate2_in[16]), .B1(n4256), .B2(
        r5[16]), .ZN(n3289) );
  AOI22D1BWP12T U4164 ( .A1(n4265), .A2(r4[16]), .B1(n4230), .B2(r6[16]), .ZN(
        n3288) );
  AOI22D1BWP12T U4165 ( .A1(n4254), .A2(tmp1[16]), .B1(n4259), .B2(r7[16]), 
        .ZN(n3287) );
  ND4D1BWP12T U4166 ( .A1(n3290), .A2(n3289), .A3(n3288), .A4(n3287), .ZN(
        n3291) );
  AOI211D1BWP12T U4167 ( .A1(n4258), .A2(r12[16]), .B(n3292), .C(n3291), .ZN(
        n3293) );
  ND4D1BWP12T U4168 ( .A1(n3296), .A2(n3295), .A3(n3294), .A4(n3293), .ZN(
        regB_out[16]) );
  AOI22D1BWP12T U4169 ( .A1(n4269), .A2(immediate2_in[15]), .B1(n4265), .B2(
        r4[15]), .ZN(n3307) );
  AOI22D1BWP12T U4170 ( .A1(n4276), .A2(r11[15]), .B1(n3462), .B2(r3[15]), 
        .ZN(n3306) );
  AOI22D1BWP12T U4171 ( .A1(n4264), .A2(r8[15]), .B1(n4267), .B2(lr[15]), .ZN(
        n3305) );
  AOI22D1BWP12T U4172 ( .A1(n4259), .A2(r7[15]), .B1(n4268), .B2(r2[15]), .ZN(
        n3297) );
  OAI21D1BWP12T U4173 ( .A1(n4263), .A2(n4886), .B(n3297), .ZN(n3303) );
  AOI22D1BWP12T U4174 ( .A1(n4260), .A2(r9[15]), .B1(n4230), .B2(r6[15]), .ZN(
        n3301) );
  AOI22D1BWP12T U4175 ( .A1(n4258), .A2(r12[15]), .B1(n4257), .B2(r10[15]), 
        .ZN(n3300) );
  AOI22D1BWP12T U4176 ( .A1(n4229), .A2(r0[15]), .B1(n4256), .B2(r5[15]), .ZN(
        n3299) );
  AOI22D1BWP12T U4177 ( .A1(n4255), .A2(r1[15]), .B1(n4254), .B2(tmp1[15]), 
        .ZN(n3298) );
  ND4D1BWP12T U4178 ( .A1(n3301), .A2(n3300), .A3(n3299), .A4(n3298), .ZN(
        n3302) );
  AOI211D1BWP12T U4179 ( .A1(n4266), .A2(sp_out[15]), .B(n3303), .C(n3302), 
        .ZN(n3304) );
  ND4D1BWP12T U4180 ( .A1(n3307), .A2(n3306), .A3(n3305), .A4(n3304), .ZN(
        regB_out[15]) );
  AOI22D1BWP12T U4181 ( .A1(n4229), .A2(r0[14]), .B1(n3486), .B2(pc_out[14]), 
        .ZN(n3318) );
  AOI22D1BWP12T U4182 ( .A1(n4257), .A2(r10[14]), .B1(n4264), .B2(r8[14]), 
        .ZN(n3317) );
  AOI22D1BWP12T U4183 ( .A1(n4276), .A2(r11[14]), .B1(n4268), .B2(r2[14]), 
        .ZN(n3316) );
  AOI22D1BWP12T U4184 ( .A1(n4255), .A2(r1[14]), .B1(n4259), .B2(r7[14]), .ZN(
        n3308) );
  OAI21D1BWP12T U4185 ( .A1(n3488), .A2(n4243), .B(n3308), .ZN(n3314) );
  AOI22D1BWP12T U4186 ( .A1(n4266), .A2(sp_out[14]), .B1(n4265), .B2(r4[14]), 
        .ZN(n3312) );
  AOI22D1BWP12T U4187 ( .A1(n4258), .A2(r12[14]), .B1(n4230), .B2(r6[14]), 
        .ZN(n3311) );
  AOI22D1BWP12T U4188 ( .A1(n4256), .A2(r5[14]), .B1(n3462), .B2(r3[14]), .ZN(
        n3310) );
  AOI22D1BWP12T U4189 ( .A1(n4269), .A2(immediate2_in[14]), .B1(n4254), .B2(
        tmp1[14]), .ZN(n3309) );
  ND4D1BWP12T U4190 ( .A1(n3312), .A2(n3311), .A3(n3310), .A4(n3309), .ZN(
        n3313) );
  AOI211D1BWP12T U4191 ( .A1(n4260), .A2(r9[14]), .B(n3314), .C(n3313), .ZN(
        n3315) );
  ND4D1BWP12T U4192 ( .A1(n3318), .A2(n3317), .A3(n3316), .A4(n3315), .ZN(
        regB_out[14]) );
  AOI22D1BWP12T U4193 ( .A1(n4255), .A2(r1[13]), .B1(n4230), .B2(r6[13]), .ZN(
        n3329) );
  AOI22D1BWP12T U4194 ( .A1(n4256), .A2(r5[13]), .B1(n4267), .B2(lr[13]), .ZN(
        n3328) );
  AOI22D1BWP12T U4195 ( .A1(n4229), .A2(r0[13]), .B1(n4265), .B2(r4[13]), .ZN(
        n3327) );
  INVD1BWP12T U4196 ( .I(pc_out[13]), .ZN(n4436) );
  AOI22D1BWP12T U4197 ( .A1(n4266), .A2(sp_out[13]), .B1(n4257), .B2(r10[13]), 
        .ZN(n3319) );
  OAI21D1BWP12T U4198 ( .A1(n4263), .A2(n4436), .B(n3319), .ZN(n3325) );
  AOI22D1BWP12T U4199 ( .A1(n4258), .A2(r12[13]), .B1(n4268), .B2(r2[13]), 
        .ZN(n3323) );
  AOI22D1BWP12T U4200 ( .A1(n4260), .A2(r9[13]), .B1(n4259), .B2(r7[13]), .ZN(
        n3322) );
  AOI22D1BWP12T U4201 ( .A1(n4276), .A2(r11[13]), .B1(n3462), .B2(r3[13]), 
        .ZN(n3321) );
  AOI22D1BWP12T U4202 ( .A1(n4254), .A2(tmp1[13]), .B1(n4264), .B2(r8[13]), 
        .ZN(n3320) );
  ND4D1BWP12T U4203 ( .A1(n3323), .A2(n3322), .A3(n3321), .A4(n3320), .ZN(
        n3324) );
  AOI211D1BWP12T U4204 ( .A1(n4269), .A2(immediate2_in[13]), .B(n3325), .C(
        n3324), .ZN(n3326) );
  ND4D1BWP12T U4205 ( .A1(n3329), .A2(n3328), .A3(n3327), .A4(n3326), .ZN(
        regB_out[13]) );
  AOI22D1BWP12T U4206 ( .A1(n4254), .A2(tmp1[12]), .B1(n3462), .B2(r3[12]), 
        .ZN(n3340) );
  AOI22D1BWP12T U4207 ( .A1(n4229), .A2(r0[12]), .B1(n4258), .B2(r12[12]), 
        .ZN(n3339) );
  INVD1BWP12T U4208 ( .I(pc_out[12]), .ZN(n4424) );
  AOI22D1BWP12T U4209 ( .A1(n4255), .A2(r1[12]), .B1(n4257), .B2(r10[12]), 
        .ZN(n3331) );
  AOI22D1BWP12T U4210 ( .A1(n4260), .A2(r9[12]), .B1(n4230), .B2(r6[12]), .ZN(
        n3330) );
  OAI211D1BWP12T U4211 ( .A1(n4263), .A2(n4424), .B(n3331), .C(n3330), .ZN(
        n3337) );
  AOI22D1BWP12T U4212 ( .A1(n4276), .A2(r11[12]), .B1(n4256), .B2(r5[12]), 
        .ZN(n3335) );
  AOI22D1BWP12T U4213 ( .A1(n4266), .A2(sp_out[12]), .B1(n4265), .B2(r4[12]), 
        .ZN(n3334) );
  AOI22D1BWP12T U4214 ( .A1(n4264), .A2(r8[12]), .B1(n4259), .B2(r7[12]), .ZN(
        n3333) );
  AOI22D1BWP12T U4215 ( .A1(n4269), .A2(immediate2_in[12]), .B1(n4267), .B2(
        lr[12]), .ZN(n3332) );
  ND4D1BWP12T U4216 ( .A1(n3335), .A2(n3334), .A3(n3333), .A4(n3332), .ZN(
        n3336) );
  AOI211D1BWP12T U4217 ( .A1(n4268), .A2(r2[12]), .B(n3337), .C(n3336), .ZN(
        n3338) );
  ND3D1BWP12T U4218 ( .A1(n3340), .A2(n3339), .A3(n3338), .ZN(regB_out[12]) );
  AOI22D1BWP12T U4219 ( .A1(n4276), .A2(r11[11]), .B1(n4259), .B2(r7[11]), 
        .ZN(n3351) );
  AOI22D1BWP12T U4220 ( .A1(n4266), .A2(sp_out[11]), .B1(n4265), .B2(r4[11]), 
        .ZN(n3350) );
  AOI22D1BWP12T U4221 ( .A1(n4254), .A2(tmp1[11]), .B1(n4256), .B2(r5[11]), 
        .ZN(n3349) );
  INVD1BWP12T U4222 ( .I(pc_out[11]), .ZN(n4412) );
  AOI22D1BWP12T U4223 ( .A1(n3462), .A2(r3[11]), .B1(n4230), .B2(r6[11]), .ZN(
        n3341) );
  OAI21D1BWP12T U4224 ( .A1(n4263), .A2(n4412), .B(n3341), .ZN(n3347) );
  AOI22D1BWP12T U4225 ( .A1(n4269), .A2(immediate2_in[11]), .B1(n4264), .B2(
        r8[11]), .ZN(n3345) );
  AOI22D1BWP12T U4226 ( .A1(n4260), .A2(r9[11]), .B1(n4229), .B2(r0[11]), .ZN(
        n3344) );
  AOI22D1BWP12T U4227 ( .A1(n4255), .A2(r1[11]), .B1(n4257), .B2(r10[11]), 
        .ZN(n3343) );
  AOI22D1BWP12T U4228 ( .A1(n4258), .A2(r12[11]), .B1(n4267), .B2(lr[11]), 
        .ZN(n3342) );
  ND4D1BWP12T U4229 ( .A1(n3345), .A2(n3344), .A3(n3343), .A4(n3342), .ZN(
        n3346) );
  AOI211D1BWP12T U4230 ( .A1(n4268), .A2(r2[11]), .B(n3347), .C(n3346), .ZN(
        n3348) );
  ND4D1BWP12T U4231 ( .A1(n3351), .A2(n3350), .A3(n3349), .A4(n3348), .ZN(
        regB_out[11]) );
  AOI22D1BWP12T U4232 ( .A1(n4257), .A2(r10[10]), .B1(n4259), .B2(r7[10]), 
        .ZN(n3362) );
  AOI22D1BWP12T U4233 ( .A1(n4276), .A2(r11[10]), .B1(n4256), .B2(r5[10]), 
        .ZN(n3361) );
  AOI22D1BWP12T U4234 ( .A1(n4255), .A2(r1[10]), .B1(n3486), .B2(pc_out[10]), 
        .ZN(n3353) );
  AOI22D1BWP12T U4235 ( .A1(n4268), .A2(r2[10]), .B1(n4267), .B2(lr[10]), .ZN(
        n3352) );
  OAI211D1BWP12T U4236 ( .A1(n3475), .A2(n4401), .B(n3353), .C(n3352), .ZN(
        n3359) );
  AOI22D1BWP12T U4237 ( .A1(n4260), .A2(r9[10]), .B1(n3462), .B2(r3[10]), .ZN(
        n3357) );
  AOI22D1BWP12T U4238 ( .A1(n4229), .A2(r0[10]), .B1(n4269), .B2(
        immediate2_in[10]), .ZN(n3356) );
  AOI22D1BWP12T U4239 ( .A1(n4254), .A2(tmp1[10]), .B1(n4258), .B2(r12[10]), 
        .ZN(n3355) );
  AOI22D1BWP12T U4240 ( .A1(n4266), .A2(sp_out[10]), .B1(n4230), .B2(r6[10]), 
        .ZN(n3354) );
  ND4D1BWP12T U4241 ( .A1(n3357), .A2(n3356), .A3(n3355), .A4(n3354), .ZN(
        n3358) );
  AOI211D1BWP12T U4242 ( .A1(n4265), .A2(r4[10]), .B(n3359), .C(n3358), .ZN(
        n3360) );
  ND3D1BWP12T U4243 ( .A1(n3362), .A2(n3361), .A3(n3360), .ZN(regB_out[10]) );
  AOI22D1BWP12T U4244 ( .A1(n4229), .A2(r0[9]), .B1(n4266), .B2(sp_out[9]), 
        .ZN(n3373) );
  AOI22D1BWP12T U4245 ( .A1(n4257), .A2(r10[9]), .B1(n3462), .B2(r3[9]), .ZN(
        n3372) );
  AOI22D1BWP12T U4246 ( .A1(n4269), .A2(immediate2_in[9]), .B1(n4264), .B2(
        r8[9]), .ZN(n3371) );
  INVD1BWP12T U4247 ( .I(pc_out[9]), .ZN(n3773) );
  AOI22D1BWP12T U4248 ( .A1(n4255), .A2(r1[9]), .B1(n4267), .B2(lr[9]), .ZN(
        n3363) );
  OAI21D1BWP12T U4249 ( .A1(n4263), .A2(n3773), .B(n3363), .ZN(n3369) );
  AOI22D1BWP12T U4250 ( .A1(n4260), .A2(r9[9]), .B1(n4259), .B2(r7[9]), .ZN(
        n3367) );
  AOI22D1BWP12T U4251 ( .A1(n4258), .A2(r12[9]), .B1(n4268), .B2(r2[9]), .ZN(
        n3366) );
  AOI22D1BWP12T U4252 ( .A1(n4265), .A2(r4[9]), .B1(n4256), .B2(r5[9]), .ZN(
        n3365) );
  AOI22D1BWP12T U4253 ( .A1(n4254), .A2(tmp1[9]), .B1(n4230), .B2(r6[9]), .ZN(
        n3364) );
  ND4D1BWP12T U4254 ( .A1(n3367), .A2(n3366), .A3(n3365), .A4(n3364), .ZN(
        n3368) );
  AOI211D1BWP12T U4255 ( .A1(n4276), .A2(r11[9]), .B(n3369), .C(n3368), .ZN(
        n3370) );
  ND4D1BWP12T U4256 ( .A1(n3373), .A2(n3372), .A3(n3371), .A4(n3370), .ZN(
        regB_out[9]) );
  AOI22D1BWP12T U4257 ( .A1(n4254), .A2(tmp1[8]), .B1(n3486), .B2(pc_out[8]), 
        .ZN(n3384) );
  AOI22D1BWP12T U4258 ( .A1(n4266), .A2(sp_out[8]), .B1(n4257), .B2(r10[8]), 
        .ZN(n3383) );
  AOI22D1BWP12T U4259 ( .A1(n4255), .A2(r1[8]), .B1(n4265), .B2(r4[8]), .ZN(
        n3382) );
  AOI22D1BWP12T U4260 ( .A1(n4229), .A2(r0[8]), .B1(n4264), .B2(r8[8]), .ZN(
        n3374) );
  OAI21D1BWP12T U4261 ( .A1(n3488), .A2(n4377), .B(n3374), .ZN(n3380) );
  AOI22D1BWP12T U4262 ( .A1(n4256), .A2(r5[8]), .B1(n4268), .B2(r2[8]), .ZN(
        n3378) );
  AOI22D1BWP12T U4263 ( .A1(n4259), .A2(r7[8]), .B1(n3462), .B2(r3[8]), .ZN(
        n3377) );
  AOI22D1BWP12T U4264 ( .A1(n4269), .A2(immediate2_in[8]), .B1(n4230), .B2(
        r6[8]), .ZN(n3376) );
  AOI22D1BWP12T U4265 ( .A1(n4260), .A2(r9[8]), .B1(n4258), .B2(r12[8]), .ZN(
        n3375) );
  ND4D1BWP12T U4266 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(
        n3379) );
  AOI211D1BWP12T U4267 ( .A1(n4276), .A2(r11[8]), .B(n3380), .C(n3379), .ZN(
        n3381) );
  ND4D1BWP12T U4268 ( .A1(n3384), .A2(n3383), .A3(n3382), .A4(n3381), .ZN(
        regB_out[8]) );
  AOI22D1BWP12T U4269 ( .A1(n4269), .A2(immediate2_in[7]), .B1(n4268), .B2(
        r2[7]), .ZN(n3395) );
  AOI22D1BWP12T U4270 ( .A1(n4230), .A2(r6[7]), .B1(n4267), .B2(lr[7]), .ZN(
        n3394) );
  AOI22D1BWP12T U4271 ( .A1(n4276), .A2(r11[7]), .B1(n4254), .B2(tmp1[7]), 
        .ZN(n3393) );
  INVD1BWP12T U4272 ( .I(pc_out[7]), .ZN(n4365) );
  AOI22D1BWP12T U4273 ( .A1(n4257), .A2(r10[7]), .B1(n4264), .B2(r8[7]), .ZN(
        n3385) );
  OAI21D1BWP12T U4274 ( .A1(n4263), .A2(n4365), .B(n3385), .ZN(n3391) );
  AOI22D1BWP12T U4275 ( .A1(n4260), .A2(r9[7]), .B1(n4265), .B2(r4[7]), .ZN(
        n3389) );
  AOI22D1BWP12T U4276 ( .A1(n4258), .A2(r12[7]), .B1(n4259), .B2(r7[7]), .ZN(
        n3388) );
  AOI22D1BWP12T U4277 ( .A1(n4229), .A2(r0[7]), .B1(n3462), .B2(r3[7]), .ZN(
        n3387) );
  AOI22D1BWP12T U4278 ( .A1(n4266), .A2(sp_out[7]), .B1(n4256), .B2(r5[7]), 
        .ZN(n3386) );
  ND4D1BWP12T U4279 ( .A1(n3389), .A2(n3388), .A3(n3387), .A4(n3386), .ZN(
        n3390) );
  AOI211D1BWP12T U4280 ( .A1(n4255), .A2(r1[7]), .B(n3391), .C(n3390), .ZN(
        n3392) );
  ND4D1BWP12T U4281 ( .A1(n3395), .A2(n3394), .A3(n3393), .A4(n3392), .ZN(
        regB_out[7]) );
  AOI22D1BWP12T U4282 ( .A1(n4269), .A2(immediate2_in[6]), .B1(n4268), .B2(
        r2[6]), .ZN(n3406) );
  AOI22D1BWP12T U4283 ( .A1(n4276), .A2(r11[6]), .B1(n4266), .B2(sp_out[6]), 
        .ZN(n3405) );
  AOI22D1BWP12T U4284 ( .A1(n4254), .A2(tmp1[6]), .B1(n4256), .B2(r5[6]), .ZN(
        n3404) );
  INVD1BWP12T U4285 ( .I(pc_out[6]), .ZN(n4353) );
  AOI22D1BWP12T U4286 ( .A1(n4259), .A2(r7[6]), .B1(n4230), .B2(r6[6]), .ZN(
        n3396) );
  OAI21D1BWP12T U4287 ( .A1(n4263), .A2(n4353), .B(n3396), .ZN(n3402) );
  AOI22D1BWP12T U4288 ( .A1(n4257), .A2(r10[6]), .B1(n4265), .B2(r4[6]), .ZN(
        n3400) );
  AOI22D1BWP12T U4289 ( .A1(n4260), .A2(r9[6]), .B1(n4258), .B2(r12[6]), .ZN(
        n3399) );
  AOI22D1BWP12T U4290 ( .A1(n4255), .A2(r1[6]), .B1(n3462), .B2(r3[6]), .ZN(
        n3398) );
  AOI22D1BWP12T U4291 ( .A1(n4229), .A2(r0[6]), .B1(n4267), .B2(lr[6]), .ZN(
        n3397) );
  ND4D1BWP12T U4292 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(
        n3401) );
  AOI211D1BWP12T U4293 ( .A1(n4264), .A2(r8[6]), .B(n3402), .C(n3401), .ZN(
        n3403) );
  ND4D1BWP12T U4294 ( .A1(n3406), .A2(n3405), .A3(n3404), .A4(n3403), .ZN(
        regB_out[6]) );
  AOI22D1BWP12T U4295 ( .A1(n4264), .A2(r8[5]), .B1(n4259), .B2(r7[5]), .ZN(
        n3417) );
  AOI22D1BWP12T U4296 ( .A1(n4266), .A2(sp_out[5]), .B1(n4256), .B2(r5[5]), 
        .ZN(n3416) );
  AOI22D1BWP12T U4297 ( .A1(n4269), .A2(immediate2_in[5]), .B1(n4254), .B2(
        tmp1[5]), .ZN(n3415) );
  INVD1BWP12T U4298 ( .I(pc_out[5]), .ZN(n4341) );
  AOI22D1BWP12T U4299 ( .A1(n4265), .A2(r4[5]), .B1(n4230), .B2(r6[5]), .ZN(
        n3407) );
  OAI21D1BWP12T U4300 ( .A1(n4263), .A2(n4341), .B(n3407), .ZN(n3413) );
  AOI22D1BWP12T U4301 ( .A1(n4276), .A2(r11[5]), .B1(n4229), .B2(r0[5]), .ZN(
        n3411) );
  AOI22D1BWP12T U4302 ( .A1(n4258), .A2(r12[5]), .B1(n4257), .B2(r10[5]), .ZN(
        n3410) );
  AOI22D1BWP12T U4303 ( .A1(n4260), .A2(r9[5]), .B1(n3462), .B2(r3[5]), .ZN(
        n3409) );
  AOI22D1BWP12T U4304 ( .A1(n4268), .A2(r2[5]), .B1(n4267), .B2(lr[5]), .ZN(
        n3408) );
  ND4D1BWP12T U4305 ( .A1(n3411), .A2(n3410), .A3(n3409), .A4(n3408), .ZN(
        n3412) );
  AOI211D1BWP12T U4306 ( .A1(n4255), .A2(r1[5]), .B(n3413), .C(n3412), .ZN(
        n3414) );
  ND4D1BWP12T U4307 ( .A1(n3417), .A2(n3416), .A3(n3415), .A4(n3414), .ZN(
        regB_out[5]) );
  AOI22D1BWP12T U4308 ( .A1(n4264), .A2(r8[4]), .B1(n4268), .B2(r2[4]), .ZN(
        n3428) );
  AOI22D1BWP12T U4309 ( .A1(n3486), .A2(pc_out[4]), .B1(n4257), .B2(r10[4]), 
        .ZN(n3427) );
  AOI22D1BWP12T U4310 ( .A1(n4276), .A2(r11[4]), .B1(n4256), .B2(r5[4]), .ZN(
        n3426) );
  AOI22D1BWP12T U4311 ( .A1(n4259), .A2(r7[4]), .B1(n3462), .B2(r3[4]), .ZN(
        n3418) );
  OAI21D1BWP12T U4312 ( .A1(n3488), .A2(n4330), .B(n3418), .ZN(n3424) );
  AOI22D1BWP12T U4313 ( .A1(n4255), .A2(r1[4]), .B1(n4269), .B2(
        immediate2_in[4]), .ZN(n3422) );
  AOI22D1BWP12T U4314 ( .A1(n4260), .A2(r9[4]), .B1(n4258), .B2(r12[4]), .ZN(
        n3421) );
  AOI22D1BWP12T U4315 ( .A1(n4229), .A2(r0[4]), .B1(n4230), .B2(r6[4]), .ZN(
        n3420) );
  AOI22D1BWP12T U4316 ( .A1(n4266), .A2(sp_out[4]), .B1(n4265), .B2(r4[4]), 
        .ZN(n3419) );
  ND4D1BWP12T U4317 ( .A1(n3422), .A2(n3421), .A3(n3420), .A4(n3419), .ZN(
        n3423) );
  AOI211D1BWP12T U4318 ( .A1(n4254), .A2(tmp1[4]), .B(n3424), .C(n3423), .ZN(
        n3425) );
  ND4D1BWP12T U4319 ( .A1(n3428), .A2(n3427), .A3(n3426), .A4(n3425), .ZN(
        regB_out[4]) );
  AOI22D1BWP12T U4320 ( .A1(n4258), .A2(r12[3]), .B1(n4256), .B2(r5[3]), .ZN(
        n3439) );
  AOI22D1BWP12T U4321 ( .A1(n4269), .A2(immediate2_in[3]), .B1(n4230), .B2(
        r6[3]), .ZN(n3438) );
  INVD1BWP12T U4322 ( .I(pc_out[3]), .ZN(n4317) );
  AOI22D1BWP12T U4323 ( .A1(n4260), .A2(r9[3]), .B1(n4255), .B2(r1[3]), .ZN(
        n3430) );
  AOI22D1BWP12T U4324 ( .A1(n4254), .A2(tmp1[3]), .B1(n4264), .B2(r8[3]), .ZN(
        n3429) );
  OAI211D1BWP12T U4325 ( .A1(n4263), .A2(n4317), .B(n3430), .C(n3429), .ZN(
        n3436) );
  AOI22D1BWP12T U4326 ( .A1(n4229), .A2(r0[3]), .B1(n3462), .B2(r3[3]), .ZN(
        n3434) );
  AOI22D1BWP12T U4327 ( .A1(n4266), .A2(sp_out[3]), .B1(n4267), .B2(lr[3]), 
        .ZN(n3433) );
  AOI22D1BWP12T U4328 ( .A1(n4276), .A2(r11[3]), .B1(n4257), .B2(r10[3]), .ZN(
        n3432) );
  AOI22D1BWP12T U4329 ( .A1(n4265), .A2(r4[3]), .B1(n4259), .B2(r7[3]), .ZN(
        n3431) );
  ND4D1BWP12T U4330 ( .A1(n3434), .A2(n3433), .A3(n3432), .A4(n3431), .ZN(
        n3435) );
  AOI211D1BWP12T U4331 ( .A1(n4268), .A2(r2[3]), .B(n3436), .C(n3435), .ZN(
        n3437) );
  ND3D1BWP12T U4332 ( .A1(n3439), .A2(n3438), .A3(n3437), .ZN(regB_out[3]) );
  AOI22D1BWP12T U4333 ( .A1(n4266), .A2(sp_out[2]), .B1(n4264), .B2(r8[2]), 
        .ZN(n3450) );
  AOI22D1BWP12T U4334 ( .A1(n4257), .A2(r10[2]), .B1(n4268), .B2(r2[2]), .ZN(
        n3449) );
  AOI22D1BWP12T U4335 ( .A1(n4255), .A2(r1[2]), .B1(n3486), .B2(pc_out[2]), 
        .ZN(n3441) );
  AOI22D1BWP12T U4336 ( .A1(n4265), .A2(r4[2]), .B1(n4259), .B2(r7[2]), .ZN(
        n3440) );
  OAI211D1BWP12T U4337 ( .A1(n3488), .A2(n3850), .B(n3441), .C(n3440), .ZN(
        n3447) );
  AOI22D1BWP12T U4338 ( .A1(n4260), .A2(r9[2]), .B1(n3462), .B2(r3[2]), .ZN(
        n3445) );
  AOI22D1BWP12T U4339 ( .A1(n4254), .A2(tmp1[2]), .B1(n4230), .B2(r6[2]), .ZN(
        n3444) );
  AOI22D1BWP12T U4340 ( .A1(n4276), .A2(r11[2]), .B1(n4269), .B2(
        immediate2_in[2]), .ZN(n3443) );
  AOI22D1BWP12T U4341 ( .A1(n4258), .A2(r12[2]), .B1(n4256), .B2(r5[2]), .ZN(
        n3442) );
  ND4D1BWP12T U4342 ( .A1(n3445), .A2(n3444), .A3(n3443), .A4(n3442), .ZN(
        n3446) );
  AOI211D1BWP12T U4343 ( .A1(n4229), .A2(r0[2]), .B(n3447), .C(n3446), .ZN(
        n3448) );
  ND3D1BWP12T U4344 ( .A1(n3450), .A2(n3449), .A3(n3448), .ZN(regB_out[2]) );
  AOI22D1BWP12T U4345 ( .A1(n4229), .A2(r0[1]), .B1(n4267), .B2(lr[1]), .ZN(
        n3461) );
  AOI22D1BWP12T U4346 ( .A1(n4254), .A2(tmp1[1]), .B1(n4268), .B2(r2[1]), .ZN(
        n3460) );
  AOI22D1BWP12T U4347 ( .A1(n4260), .A2(r9[1]), .B1(n4265), .B2(r4[1]), .ZN(
        n3459) );
  INVD1BWP12T U4348 ( .I(pc_out[1]), .ZN(n4293) );
  AOI22D1BWP12T U4349 ( .A1(n4257), .A2(r10[1]), .B1(n4264), .B2(r8[1]), .ZN(
        n3451) );
  OAI21D1BWP12T U4350 ( .A1(n4263), .A2(n4293), .B(n3451), .ZN(n3457) );
  AOI22D1BWP12T U4351 ( .A1(n4258), .A2(r12[1]), .B1(n3462), .B2(r3[1]), .ZN(
        n3455) );
  AOI22D1BWP12T U4352 ( .A1(n4255), .A2(r1[1]), .B1(n4259), .B2(r7[1]), .ZN(
        n3454) );
  AOI22D1BWP12T U4353 ( .A1(n4256), .A2(r5[1]), .B1(n4230), .B2(r6[1]), .ZN(
        n3453) );
  AOI22D1BWP12T U4354 ( .A1(n4269), .A2(immediate2_in[1]), .B1(n4266), .B2(
        sp_out[1]), .ZN(n3452) );
  ND4D1BWP12T U4355 ( .A1(n3455), .A2(n3454), .A3(n3453), .A4(n3452), .ZN(
        n3456) );
  AOI211D1BWP12T U4356 ( .A1(n4276), .A2(r11[1]), .B(n3457), .C(n3456), .ZN(
        n3458) );
  ND4D1BWP12T U4357 ( .A1(n3461), .A2(n3460), .A3(n3459), .A4(n3458), .ZN(
        regB_out[1]) );
  AOI22D1BWP12T U4358 ( .A1(r2[0]), .A2(n4268), .B1(r3[0]), .B2(n3462), .ZN(
        n3473) );
  AOI22D1BWP12T U4359 ( .A1(r6[0]), .A2(n4230), .B1(lr[0]), .B2(n4267), .ZN(
        n3472) );
  AOI22D1BWP12T U4360 ( .A1(r8[0]), .A2(n4264), .B1(r7[0]), .B2(n4259), .ZN(
        n3471) );
  INVD1BWP12T U4361 ( .I(pc_out[0]), .ZN(n4459) );
  AOI22D1BWP12T U4362 ( .A1(tmp1[0]), .A2(n4254), .B1(r12[0]), .B2(n4258), 
        .ZN(n3463) );
  OAI21D1BWP12T U4363 ( .A1(n4459), .A2(n4263), .B(n3463), .ZN(n3469) );
  AOI22D1BWP12T U4364 ( .A1(r1[0]), .A2(n4255), .B1(r0[0]), .B2(n4229), .ZN(
        n3467) );
  AOI22D1BWP12T U4365 ( .A1(r11[0]), .A2(n4276), .B1(r9[0]), .B2(n4260), .ZN(
        n3466) );
  AOI22D1BWP12T U4366 ( .A1(r4[0]), .A2(n4265), .B1(r5[0]), .B2(n4256), .ZN(
        n3465) );
  AOI22D1BWP12T U4367 ( .A1(sp_out[0]), .A2(n4266), .B1(r10[0]), .B2(n4257), 
        .ZN(n3464) );
  ND4D1BWP12T U4368 ( .A1(n3467), .A2(n3466), .A3(n3465), .A4(n3464), .ZN(
        n3468) );
  AOI211D1BWP12T U4369 ( .A1(n4269), .A2(immediate2_in[0]), .B(n3469), .C(
        n3468), .ZN(n3470) );
  ND4D1BWP12T U4370 ( .A1(n3473), .A2(n3472), .A3(n3471), .A4(n3470), .ZN(
        regB_out[0]) );
  AOI22D1BWP12T U4371 ( .A1(n4276), .A2(r11[27]), .B1(n4256), .B2(r5[27]), 
        .ZN(n3485) );
  AOI22D1BWP12T U4372 ( .A1(n3486), .A2(pc_out[27]), .B1(n4268), .B2(r2[27]), 
        .ZN(n3484) );
  AOI22D1BWP12T U4373 ( .A1(n4265), .A2(r4[27]), .B1(n3462), .B2(r3[27]), .ZN(
        n3483) );
  AOI22D1BWP12T U4374 ( .A1(n4257), .A2(r10[27]), .B1(n4230), .B2(r6[27]), 
        .ZN(n3474) );
  OAI21D1BWP12T U4375 ( .A1(n3475), .A2(n4614), .B(n3474), .ZN(n3481) );
  AOI22D1BWP12T U4376 ( .A1(n4229), .A2(r0[27]), .B1(n4267), .B2(lr[27]), .ZN(
        n3479) );
  AOI22D1BWP12T U4377 ( .A1(n4254), .A2(tmp1[27]), .B1(n4259), .B2(r7[27]), 
        .ZN(n3478) );
  AOI22D1BWP12T U4378 ( .A1(n4255), .A2(r1[27]), .B1(n4258), .B2(r12[27]), 
        .ZN(n3477) );
  AOI22D1BWP12T U4379 ( .A1(n4260), .A2(r9[27]), .B1(n4269), .B2(
        immediate2_in[27]), .ZN(n3476) );
  ND4D1BWP12T U4380 ( .A1(n3479), .A2(n3478), .A3(n3477), .A4(n3476), .ZN(
        n3480) );
  AOI211D1BWP12T U4381 ( .A1(n4266), .A2(sp_out[27]), .B(n3481), .C(n3480), 
        .ZN(n3482) );
  ND4D1BWP12T U4382 ( .A1(n3485), .A2(n3484), .A3(n3483), .A4(n3482), .ZN(
        regB_out[27]) );
  AOI22D1BWP12T U4383 ( .A1(n4260), .A2(r9[26]), .B1(n4269), .B2(
        immediate2_in[26]), .ZN(n3498) );
  AOI22D1BWP12T U4384 ( .A1(n3486), .A2(pc_out[26]), .B1(n4264), .B2(r8[26]), 
        .ZN(n3497) );
  AOI22D1BWP12T U4385 ( .A1(n4265), .A2(r4[26]), .B1(n4259), .B2(r7[26]), .ZN(
        n3496) );
  AOI22D1BWP12T U4386 ( .A1(n4229), .A2(r0[26]), .B1(n4258), .B2(r12[26]), 
        .ZN(n3487) );
  OAI21D1BWP12T U4387 ( .A1(n3488), .A2(n4602), .B(n3487), .ZN(n3494) );
  AOI22D1BWP12T U4388 ( .A1(n4254), .A2(tmp1[26]), .B1(n4266), .B2(sp_out[26]), 
        .ZN(n3492) );
  AOI22D1BWP12T U4389 ( .A1(n4256), .A2(r5[26]), .B1(n4230), .B2(r6[26]), .ZN(
        n3491) );
  AOI22D1BWP12T U4390 ( .A1(n4255), .A2(r1[26]), .B1(n3462), .B2(r3[26]), .ZN(
        n3490) );
  AOI22D1BWP12T U4391 ( .A1(n4257), .A2(r10[26]), .B1(n4268), .B2(r2[26]), 
        .ZN(n3489) );
  ND4D1BWP12T U4392 ( .A1(n3492), .A2(n3491), .A3(n3490), .A4(n3489), .ZN(
        n3493) );
  AOI211D1BWP12T U4393 ( .A1(n4276), .A2(r11[26]), .B(n3494), .C(n3493), .ZN(
        n3495) );
  ND4D1BWP12T U4394 ( .A1(n3498), .A2(n3497), .A3(n3496), .A4(n3495), .ZN(
        regB_out[26]) );
  AOI22D1BWP12T U4395 ( .A1(n4255), .A2(r1[25]), .B1(n4269), .B2(
        immediate2_in[25]), .ZN(n3509) );
  AOI22D1BWP12T U4396 ( .A1(n4258), .A2(r12[25]), .B1(n4256), .B2(r5[25]), 
        .ZN(n3508) );
  AOI22D1BWP12T U4397 ( .A1(n4229), .A2(r0[25]), .B1(n4266), .B2(sp_out[25]), 
        .ZN(n3507) );
  INVD1BWP12T U4398 ( .I(pc_out[25]), .ZN(n4588) );
  AOI22D1BWP12T U4399 ( .A1(n4264), .A2(r8[25]), .B1(n4230), .B2(r6[25]), .ZN(
        n3499) );
  OAI21D1BWP12T U4400 ( .A1(n4263), .A2(n4588), .B(n3499), .ZN(n3505) );
  AOI22D1BWP12T U4401 ( .A1(n4276), .A2(r11[25]), .B1(n4257), .B2(r10[25]), 
        .ZN(n3503) );
  AOI22D1BWP12T U4402 ( .A1(n4259), .A2(r7[25]), .B1(n4268), .B2(r2[25]), .ZN(
        n3502) );
  AOI22D1BWP12T U4403 ( .A1(n4260), .A2(r9[25]), .B1(n4254), .B2(tmp1[25]), 
        .ZN(n3501) );
  AOI22D1BWP12T U4404 ( .A1(n3462), .A2(r3[25]), .B1(n4267), .B2(lr[25]), .ZN(
        n3500) );
  ND4D1BWP12T U4405 ( .A1(n3503), .A2(n3502), .A3(n3501), .A4(n3500), .ZN(
        n3504) );
  AOI211D1BWP12T U4406 ( .A1(n4265), .A2(r4[25]), .B(n3505), .C(n3504), .ZN(
        n3506) );
  ND4D1BWP12T U4407 ( .A1(n3509), .A2(n3508), .A3(n3507), .A4(n3506), .ZN(
        regB_out[25]) );
  AOI22D1BWP12T U4408 ( .A1(n4255), .A2(r1[24]), .B1(n4265), .B2(r4[24]), .ZN(
        n3520) );
  AOI22D1BWP12T U4409 ( .A1(n4258), .A2(r12[24]), .B1(n4268), .B2(r2[24]), 
        .ZN(n3519) );
  AOI22D1BWP12T U4410 ( .A1(n4269), .A2(immediate2_in[24]), .B1(n4254), .B2(
        tmp1[24]), .ZN(n3518) );
  INVD1BWP12T U4411 ( .I(pc_out[24]), .ZN(n4576) );
  AOI22D1BWP12T U4412 ( .A1(n4230), .A2(r6[24]), .B1(n4267), .B2(lr[24]), .ZN(
        n3510) );
  OAI21D1BWP12T U4413 ( .A1(n4263), .A2(n4576), .B(n3510), .ZN(n3516) );
  AOI22D1BWP12T U4414 ( .A1(n4257), .A2(r10[24]), .B1(n4256), .B2(r5[24]), 
        .ZN(n3514) );
  AOI22D1BWP12T U4415 ( .A1(n4260), .A2(r9[24]), .B1(n4264), .B2(r8[24]), .ZN(
        n3513) );
  AOI22D1BWP12T U4416 ( .A1(n4276), .A2(r11[24]), .B1(n4229), .B2(r0[24]), 
        .ZN(n3512) );
  AOI22D1BWP12T U4417 ( .A1(n4266), .A2(sp_out[24]), .B1(n3462), .B2(r3[24]), 
        .ZN(n3511) );
  ND4D1BWP12T U4418 ( .A1(n3514), .A2(n3513), .A3(n3512), .A4(n3511), .ZN(
        n3515) );
  AOI211D1BWP12T U4419 ( .A1(n4259), .A2(r7[24]), .B(n3516), .C(n3515), .ZN(
        n3517) );
  ND4D1BWP12T U4420 ( .A1(n3520), .A2(n3519), .A3(n3518), .A4(n3517), .ZN(
        regB_out[24]) );
  ND2D1BWP12T U4421 ( .A1(readC_sel[1]), .A2(readC_sel[0]), .ZN(n3535) );
  INVD1BWP12T U4422 ( .I(readC_sel[4]), .ZN(n3892) );
  INVD1BWP12T U4423 ( .I(readC_sel[3]), .ZN(n3523) );
  INVD1BWP12T U4424 ( .I(readC_sel[2]), .ZN(n3525) );
  ND3D1BWP12T U4425 ( .A1(n3892), .A2(n3523), .A3(n3525), .ZN(n3536) );
  NR2D1BWP12T U4426 ( .A1(n3535), .A2(n3536), .ZN(n3880) );
  INVD1BWP12T U4427 ( .I(n3880), .ZN(n3853) );
  INVD1BWP12T U4428 ( .I(readC_sel[1]), .ZN(n3522) );
  INVD1BWP12T U4429 ( .I(readC_sel[0]), .ZN(n3521) );
  ND2D1BWP12T U4430 ( .A1(n3522), .A2(n3521), .ZN(n3537) );
  ND3D1BWP12T U4431 ( .A1(readC_sel[3]), .A2(readC_sel[2]), .A3(n3892), .ZN(
        n3534) );
  OR2XD1BWP12T U4432 ( .A1(n3537), .A2(n3534), .Z(n3851) );
  INVD1BWP12T U4433 ( .I(n3851), .ZN(n3884) );
  AOI22D1BWP12T U4434 ( .A1(r3[31]), .A2(n3880), .B1(r12[31]), .B2(n3884), 
        .ZN(n3543) );
  ND2D1BWP12T U4435 ( .A1(readC_sel[1]), .A2(n3521), .ZN(n3528) );
  NR2D1BWP12T U4436 ( .A1(n3528), .A2(n3536), .ZN(n3864) );
  NR2D1BWP12T U4437 ( .A1(n3528), .A2(n3534), .ZN(n3831) );
  INVD1BWP12T U4438 ( .I(n3831), .ZN(n3849) );
  AOI22D1BWP12T U4439 ( .A1(r2[31]), .A2(n3864), .B1(lr[31]), .B2(n3831), .ZN(
        n3542) );
  ND2D1BWP12T U4440 ( .A1(readC_sel[0]), .A2(n3522), .ZN(n3527) );
  NR2D1BWP12T U4441 ( .A1(n3527), .A2(n3534), .ZN(n3885) );
  NR2D1BWP12T U4442 ( .A1(n3527), .A2(n3536), .ZN(n3882) );
  INVD1BWP12T U4443 ( .I(n3882), .ZN(n3621) );
  AOI22D1BWP12T U4444 ( .A1(sp_out[31]), .A2(n3885), .B1(r1[31]), .B2(n3882), 
        .ZN(n3541) );
  ND2D1BWP12T U4445 ( .A1(readC_sel[2]), .A2(n3523), .ZN(n3526) );
  NR2D1BWP12T U4446 ( .A1(n3526), .A2(n3535), .ZN(n3524) );
  ND2D1BWP12T U4447 ( .A1(readC_sel[3]), .A2(n3525), .ZN(n3529) );
  NR2D1BWP12T U4448 ( .A1(n3529), .A2(n3535), .ZN(n3595) );
  AOI22D1BWP12T U4449 ( .A1(r7[31]), .A2(n3524), .B1(r11[31]), .B2(n3595), 
        .ZN(n3533) );
  NR2D1BWP12T U4450 ( .A1(n3537), .A2(n3529), .ZN(n3871) );
  NR2D1BWP12T U4451 ( .A1(n3526), .A2(n3527), .ZN(n3875) );
  AOI22D1BWP12T U4452 ( .A1(r8[31]), .A2(n3871), .B1(r5[31]), .B2(n3875), .ZN(
        n3532) );
  NR2D1BWP12T U4453 ( .A1(n3537), .A2(n3526), .ZN(n3832) );
  NR2D1BWP12T U4454 ( .A1(n3526), .A2(n3528), .ZN(n3873) );
  AOI22D1BWP12T U4455 ( .A1(r4[31]), .A2(n3832), .B1(r6[31]), .B2(n3873), .ZN(
        n3531) );
  NR2D1BWP12T U4456 ( .A1(n3529), .A2(n3527), .ZN(n3872) );
  NR2D1BWP12T U4457 ( .A1(n3529), .A2(n3528), .ZN(n3874) );
  AOI22D1BWP12T U4458 ( .A1(r9[31]), .A2(n3872), .B1(r10[31]), .B2(n3874), 
        .ZN(n3530) );
  ND4D1BWP12T U4459 ( .A1(n3533), .A2(n3532), .A3(n3531), .A4(n3530), .ZN(
        n3539) );
  NR2D1BWP12T U4460 ( .A1(n3535), .A2(n3534), .ZN(n3883) );
  INVD1BWP12T U4461 ( .I(n3883), .ZN(n3852) );
  OR2XD1BWP12T U4462 ( .A1(n3537), .A2(n3536), .Z(n3814) );
  OAI22D1BWP12T U4463 ( .A1(n4262), .A2(n3852), .B1(n4848), .B2(n3814), .ZN(
        n3538) );
  AOI21D1BWP12T U4464 ( .A1(n3892), .A2(n3539), .B(n3538), .ZN(n3540) );
  ND4D1BWP12T U4465 ( .A1(n3543), .A2(n3542), .A3(n3541), .A4(n3540), .ZN(
        regC_out[31]) );
  AOI22D1BWP12T U4466 ( .A1(n4229), .A2(r0[29]), .B1(n4266), .B2(sp_out[29]), 
        .ZN(n3554) );
  AOI22D1BWP12T U4467 ( .A1(n4260), .A2(r9[29]), .B1(n4265), .B2(r4[29]), .ZN(
        n3553) );
  AOI22D1BWP12T U4468 ( .A1(n4268), .A2(r2[29]), .B1(n3462), .B2(r3[29]), .ZN(
        n3552) );
  INVD1BWP12T U4469 ( .I(pc_out[29]), .ZN(n3925) );
  AOI22D1BWP12T U4470 ( .A1(n4254), .A2(tmp1[29]), .B1(n4256), .B2(r5[29]), 
        .ZN(n3544) );
  OAI21D1BWP12T U4471 ( .A1(n4263), .A2(n3925), .B(n3544), .ZN(n3550) );
  AOI22D1BWP12T U4472 ( .A1(n4276), .A2(r11[29]), .B1(n4230), .B2(r6[29]), 
        .ZN(n3548) );
  AOI22D1BWP12T U4473 ( .A1(n4258), .A2(r12[29]), .B1(n4257), .B2(r10[29]), 
        .ZN(n3547) );
  AOI22D1BWP12T U4474 ( .A1(n4264), .A2(r8[29]), .B1(n4267), .B2(lr[29]), .ZN(
        n3546) );
  AOI22D1BWP12T U4475 ( .A1(n4269), .A2(immediate2_in[29]), .B1(n4259), .B2(
        r7[29]), .ZN(n3545) );
  ND4D1BWP12T U4476 ( .A1(n3548), .A2(n3547), .A3(n3546), .A4(n3545), .ZN(
        n3549) );
  AOI211D1BWP12T U4477 ( .A1(n4255), .A2(r1[29]), .B(n3550), .C(n3549), .ZN(
        n3551) );
  ND4D1BWP12T U4478 ( .A1(n3554), .A2(n3553), .A3(n3552), .A4(n3551), .ZN(
        regB_out[29]) );
  AOI22D1BWP12T U4479 ( .A1(r10[30]), .A2(n3874), .B1(r6[30]), .B2(n3873), 
        .ZN(n3558) );
  AOI22D1BWP12T U4480 ( .A1(r11[30]), .A2(n3595), .B1(r8[30]), .B2(n3871), 
        .ZN(n3557) );
  AOI22D1BWP12T U4481 ( .A1(r9[30]), .A2(n3872), .B1(r4[30]), .B2(n3832), .ZN(
        n3556) );
  AOI22D1BWP12T U4482 ( .A1(r5[30]), .A2(n3875), .B1(r7[30]), .B2(n3524), .ZN(
        n3555) );
  ND4D1BWP12T U4483 ( .A1(n3558), .A2(n3557), .A3(n3556), .A4(n3555), .ZN(
        n3564) );
  AOI22D1BWP12T U4484 ( .A1(r1[30]), .A2(n3882), .B1(r12[30]), .B2(n3884), 
        .ZN(n3562) );
  INVD1BWP12T U4485 ( .I(n3814), .ZN(n3881) );
  AOI22D1BWP12T U4486 ( .A1(sp_out[30]), .A2(n3885), .B1(r0[30]), .B2(n3881), 
        .ZN(n3561) );
  INVD1BWP12T U4487 ( .I(n3864), .ZN(n3837) );
  AOI22D1BWP12T U4488 ( .A1(r2[30]), .A2(n3864), .B1(r3[30]), .B2(n3880), .ZN(
        n3560) );
  AOI22D1BWP12T U4489 ( .A1(lr[30]), .A2(n3831), .B1(pc_out[30]), .B2(n3883), 
        .ZN(n3559) );
  ND4D1BWP12T U4490 ( .A1(n3562), .A2(n3561), .A3(n3560), .A4(n3559), .ZN(
        n3563) );
  AO21D1BWP12T U4491 ( .A1(n3892), .A2(n3564), .B(n3563), .Z(regC_out[30]) );
  AOI22D1BWP12T U4492 ( .A1(r2[29]), .A2(n3864), .B1(r0[29]), .B2(n3881), .ZN(
        n3574) );
  AOI22D1BWP12T U4493 ( .A1(lr[29]), .A2(n3831), .B1(sp_out[29]), .B2(n3885), 
        .ZN(n3573) );
  AOI22D1BWP12T U4494 ( .A1(r12[29]), .A2(n3884), .B1(r3[29]), .B2(n3880), 
        .ZN(n3572) );
  AOI22D1BWP12T U4495 ( .A1(r10[29]), .A2(n3874), .B1(r7[29]), .B2(n3524), 
        .ZN(n3568) );
  AOI22D1BWP12T U4496 ( .A1(r11[29]), .A2(n3595), .B1(r5[29]), .B2(n3875), 
        .ZN(n3567) );
  AOI22D1BWP12T U4497 ( .A1(r6[29]), .A2(n3873), .B1(r8[29]), .B2(n3871), .ZN(
        n3566) );
  AOI22D1BWP12T U4498 ( .A1(r4[29]), .A2(n3832), .B1(r9[29]), .B2(n3872), .ZN(
        n3565) );
  ND4D1BWP12T U4499 ( .A1(n3568), .A2(n3567), .A3(n3566), .A4(n3565), .ZN(
        n3570) );
  OAI22D1BWP12T U4500 ( .A1(n4836), .A2(n3621), .B1(n3925), .B2(n3852), .ZN(
        n3569) );
  AOI21D1BWP12T U4501 ( .A1(n3892), .A2(n3570), .B(n3569), .ZN(n3571) );
  ND4D1BWP12T U4502 ( .A1(n3574), .A2(n3573), .A3(n3572), .A4(n3571), .ZN(
        regC_out[29]) );
  AOI22D1BWP12T U4503 ( .A1(r11[28]), .A2(n3595), .B1(r5[28]), .B2(n3875), 
        .ZN(n3578) );
  AOI22D1BWP12T U4504 ( .A1(r8[28]), .A2(n3871), .B1(r6[28]), .B2(n3873), .ZN(
        n3577) );
  AOI22D1BWP12T U4505 ( .A1(r9[28]), .A2(n3872), .B1(r7[28]), .B2(n3524), .ZN(
        n3576) );
  AOI22D1BWP12T U4506 ( .A1(r10[28]), .A2(n3874), .B1(r4[28]), .B2(n3832), 
        .ZN(n3575) );
  ND4D1BWP12T U4507 ( .A1(n3578), .A2(n3577), .A3(n3576), .A4(n3575), .ZN(
        n3584) );
  AOI22D1BWP12T U4508 ( .A1(r3[28]), .A2(n3880), .B1(sp_out[28]), .B2(n3885), 
        .ZN(n3582) );
  AOI22D1BWP12T U4509 ( .A1(lr[28]), .A2(n3831), .B1(r2[28]), .B2(n3864), .ZN(
        n3581) );
  AOI22D1BWP12T U4510 ( .A1(pc_out[28]), .A2(n3883), .B1(r12[28]), .B2(n3884), 
        .ZN(n3580) );
  AOI22D1BWP12T U4511 ( .A1(r1[28]), .A2(n3882), .B1(r0[28]), .B2(n3881), .ZN(
        n3579) );
  ND4D1BWP12T U4512 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(
        n3583) );
  AO21D1BWP12T U4513 ( .A1(n3892), .A2(n3584), .B(n3583), .Z(regC_out[28]) );
  AOI22D1BWP12T U4514 ( .A1(r8[27]), .A2(n3871), .B1(r9[27]), .B2(n3872), .ZN(
        n3588) );
  AOI22D1BWP12T U4515 ( .A1(r7[27]), .A2(n3524), .B1(r5[27]), .B2(n3875), .ZN(
        n3587) );
  AOI22D1BWP12T U4516 ( .A1(r10[27]), .A2(n3874), .B1(r4[27]), .B2(n3832), 
        .ZN(n3586) );
  AOI22D1BWP12T U4517 ( .A1(r6[27]), .A2(n3873), .B1(r11[27]), .B2(n3595), 
        .ZN(n3585) );
  ND4D1BWP12T U4518 ( .A1(n3588), .A2(n3587), .A3(n3586), .A4(n3585), .ZN(
        n3594) );
  AOI22D1BWP12T U4519 ( .A1(r1[27]), .A2(n3882), .B1(pc_out[27]), .B2(n3883), 
        .ZN(n3592) );
  AOI22D1BWP12T U4520 ( .A1(lr[27]), .A2(n3831), .B1(r0[27]), .B2(n3881), .ZN(
        n3591) );
  AOI22D1BWP12T U4521 ( .A1(sp_out[27]), .A2(n3885), .B1(r2[27]), .B2(n3864), 
        .ZN(n3590) );
  AOI22D1BWP12T U4522 ( .A1(r12[27]), .A2(n3884), .B1(r3[27]), .B2(n3880), 
        .ZN(n3589) );
  ND4D1BWP12T U4523 ( .A1(n3592), .A2(n3591), .A3(n3590), .A4(n3589), .ZN(
        n3593) );
  AO21D1BWP12T U4524 ( .A1(n3892), .A2(n3594), .B(n3593), .Z(regC_out[27]) );
  AOI22D1BWP12T U4525 ( .A1(sp_out[26]), .A2(n3885), .B1(r12[26]), .B2(n3884), 
        .ZN(n3606) );
  AOI22D1BWP12T U4526 ( .A1(r1[26]), .A2(n3882), .B1(pc_out[26]), .B2(n3883), 
        .ZN(n3605) );
  AOI22D1BWP12T U4527 ( .A1(r3[26]), .A2(n3880), .B1(r0[26]), .B2(n3881), .ZN(
        n3604) );
  AOI22D1BWP12T U4528 ( .A1(r6[26]), .A2(n3873), .B1(r8[26]), .B2(n3871), .ZN(
        n3599) );
  AOI22D1BWP12T U4529 ( .A1(r11[26]), .A2(n3595), .B1(r9[26]), .B2(n3872), 
        .ZN(n3598) );
  AOI22D1BWP12T U4530 ( .A1(r10[26]), .A2(n3874), .B1(r4[26]), .B2(n3832), 
        .ZN(n3597) );
  AOI22D1BWP12T U4531 ( .A1(r5[26]), .A2(n3875), .B1(r7[26]), .B2(n3524), .ZN(
        n3596) );
  ND4D1BWP12T U4532 ( .A1(n3599), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(
        n3602) );
  OAI22D1BWP12T U4533 ( .A1(n3600), .A2(n3837), .B1(n4602), .B2(n3849), .ZN(
        n3601) );
  AOI21D1BWP12T U4534 ( .A1(n3892), .A2(n3602), .B(n3601), .ZN(n3603) );
  ND4D1BWP12T U4535 ( .A1(n3606), .A2(n3605), .A3(n3604), .A4(n3603), .ZN(
        regC_out[26]) );
  AOI22D1BWP12T U4536 ( .A1(r6[25]), .A2(n3873), .B1(r9[25]), .B2(n3872), .ZN(
        n3610) );
  AOI22D1BWP12T U4537 ( .A1(r4[25]), .A2(n3832), .B1(r11[25]), .B2(n3595), 
        .ZN(n3609) );
  AOI22D1BWP12T U4538 ( .A1(r7[25]), .A2(n3524), .B1(r5[25]), .B2(n3875), .ZN(
        n3608) );
  AOI22D1BWP12T U4539 ( .A1(r8[25]), .A2(n3871), .B1(r10[25]), .B2(n3874), 
        .ZN(n3607) );
  ND4D1BWP12T U4540 ( .A1(n3610), .A2(n3609), .A3(n3608), .A4(n3607), .ZN(
        n3616) );
  AOI22D1BWP12T U4541 ( .A1(r2[25]), .A2(n3864), .B1(r0[25]), .B2(n3881), .ZN(
        n3614) );
  AOI22D1BWP12T U4542 ( .A1(r1[25]), .A2(n3882), .B1(r12[25]), .B2(n3884), 
        .ZN(n3613) );
  AOI22D1BWP12T U4543 ( .A1(pc_out[25]), .A2(n3883), .B1(r3[25]), .B2(n3880), 
        .ZN(n3612) );
  AOI22D1BWP12T U4544 ( .A1(lr[25]), .A2(n3831), .B1(sp_out[25]), .B2(n3885), 
        .ZN(n3611) );
  ND4D1BWP12T U4545 ( .A1(n3614), .A2(n3613), .A3(n3612), .A4(n3611), .ZN(
        n3615) );
  AO21D1BWP12T U4546 ( .A1(n3892), .A2(n3616), .B(n3615), .Z(regC_out[25]) );
  AOI22D1BWP12T U4547 ( .A1(r2[24]), .A2(n3864), .B1(r12[24]), .B2(n3884), 
        .ZN(n3627) );
  AOI22D1BWP12T U4548 ( .A1(pc_out[24]), .A2(n3883), .B1(sp_out[24]), .B2(
        n3885), .ZN(n3626) );
  AOI22D1BWP12T U4549 ( .A1(lr[24]), .A2(n3831), .B1(r0[24]), .B2(n3881), .ZN(
        n3625) );
  AOI22D1BWP12T U4550 ( .A1(r8[24]), .A2(n3871), .B1(r11[24]), .B2(n3595), 
        .ZN(n3620) );
  AOI22D1BWP12T U4551 ( .A1(r7[24]), .A2(n3524), .B1(r6[24]), .B2(n3873), .ZN(
        n3619) );
  AOI22D1BWP12T U4552 ( .A1(r5[24]), .A2(n3875), .B1(r4[24]), .B2(n3832), .ZN(
        n3618) );
  AOI22D1BWP12T U4553 ( .A1(r9[24]), .A2(n3872), .B1(r10[24]), .B2(n3874), 
        .ZN(n3617) );
  ND4D1BWP12T U4554 ( .A1(n3620), .A2(n3619), .A3(n3618), .A4(n3617), .ZN(
        n3623) );
  OAI22D1BWP12T U4555 ( .A1(n3978), .A2(n3853), .B1(n4843), .B2(n3621), .ZN(
        n3622) );
  AOI21D1BWP12T U4556 ( .A1(n3892), .A2(n3623), .B(n3622), .ZN(n3624) );
  ND4D1BWP12T U4557 ( .A1(n3627), .A2(n3626), .A3(n3625), .A4(n3624), .ZN(
        regC_out[24]) );
  AOI22D1BWP12T U4558 ( .A1(r1[23]), .A2(n3882), .B1(r12[23]), .B2(n3884), 
        .ZN(n3637) );
  AOI22D1BWP12T U4559 ( .A1(sp_out[23]), .A2(n3885), .B1(r3[23]), .B2(n3880), 
        .ZN(n3636) );
  AOI22D1BWP12T U4560 ( .A1(r2[23]), .A2(n3864), .B1(lr[23]), .B2(n3831), .ZN(
        n3635) );
  AOI22D1BWP12T U4561 ( .A1(r11[23]), .A2(n3595), .B1(r4[23]), .B2(n3832), 
        .ZN(n3631) );
  AOI22D1BWP12T U4562 ( .A1(r10[23]), .A2(n3874), .B1(r8[23]), .B2(n3871), 
        .ZN(n3630) );
  AOI22D1BWP12T U4563 ( .A1(r6[23]), .A2(n3873), .B1(r5[23]), .B2(n3875), .ZN(
        n3629) );
  AOI22D1BWP12T U4564 ( .A1(r7[23]), .A2(n3524), .B1(r9[23]), .B2(n3872), .ZN(
        n3628) );
  ND4D1BWP12T U4565 ( .A1(n3631), .A2(n3630), .A3(n3629), .A4(n3628), .ZN(
        n3633) );
  OAI22D1BWP12T U4566 ( .A1(n4564), .A2(n3852), .B1(n4833), .B2(n3814), .ZN(
        n3632) );
  AOI21D1BWP12T U4567 ( .A1(n3892), .A2(n3633), .B(n3632), .ZN(n3634) );
  ND4D1BWP12T U4568 ( .A1(n3637), .A2(n3636), .A3(n3635), .A4(n3634), .ZN(
        regC_out[23]) );
  AOI22D1BWP12T U4569 ( .A1(r6[22]), .A2(n3873), .B1(r4[22]), .B2(n3832), .ZN(
        n3641) );
  AOI22D1BWP12T U4570 ( .A1(r9[22]), .A2(n3872), .B1(r8[22]), .B2(n3871), .ZN(
        n3640) );
  AOI22D1BWP12T U4571 ( .A1(r5[22]), .A2(n3875), .B1(r11[22]), .B2(n3595), 
        .ZN(n3639) );
  AOI22D1BWP12T U4572 ( .A1(r7[22]), .A2(n3524), .B1(r10[22]), .B2(n3874), 
        .ZN(n3638) );
  ND4D1BWP12T U4573 ( .A1(n3641), .A2(n3640), .A3(n3639), .A4(n3638), .ZN(
        n3647) );
  AOI22D1BWP12T U4574 ( .A1(sp_out[22]), .A2(n3885), .B1(r3[22]), .B2(n3880), 
        .ZN(n3645) );
  AOI22D1BWP12T U4575 ( .A1(lr[22]), .A2(n3831), .B1(r12[22]), .B2(n3884), 
        .ZN(n3644) );
  AOI22D1BWP12T U4576 ( .A1(r2[22]), .A2(n3864), .B1(r0[22]), .B2(n3881), .ZN(
        n3643) );
  AOI22D1BWP12T U4577 ( .A1(r1[22]), .A2(n3882), .B1(pc_out[22]), .B2(n3883), 
        .ZN(n3642) );
  ND4D1BWP12T U4578 ( .A1(n3645), .A2(n3644), .A3(n3643), .A4(n3642), .ZN(
        n3646) );
  AO21D1BWP12T U4579 ( .A1(n3892), .A2(n3647), .B(n3646), .Z(regC_out[22]) );
  AOI22D1BWP12T U4580 ( .A1(lr[21]), .A2(n3831), .B1(r2[21]), .B2(n3864), .ZN(
        n3658) );
  AOI22D1BWP12T U4581 ( .A1(r12[21]), .A2(n3884), .B1(r0[21]), .B2(n3881), 
        .ZN(n3657) );
  AOI22D1BWP12T U4582 ( .A1(sp_out[21]), .A2(n3885), .B1(r1[21]), .B2(n3882), 
        .ZN(n3656) );
  AOI22D1BWP12T U4583 ( .A1(r6[21]), .A2(n3873), .B1(r7[21]), .B2(n3524), .ZN(
        n3651) );
  AOI22D1BWP12T U4584 ( .A1(r9[21]), .A2(n3872), .B1(r5[21]), .B2(n3875), .ZN(
        n3650) );
  AOI22D1BWP12T U4585 ( .A1(r10[21]), .A2(n3874), .B1(r4[21]), .B2(n3832), 
        .ZN(n3649) );
  AOI22D1BWP12T U4586 ( .A1(r11[21]), .A2(n3595), .B1(r8[21]), .B2(n3871), 
        .ZN(n3648) );
  ND4D1BWP12T U4587 ( .A1(n3651), .A2(n3650), .A3(n3649), .A4(n3648), .ZN(
        n3654) );
  OAI22D1BWP12T U4588 ( .A1(n4541), .A2(n3852), .B1(n3652), .B2(n3853), .ZN(
        n3653) );
  AOI21D1BWP12T U4589 ( .A1(n3892), .A2(n3654), .B(n3653), .ZN(n3655) );
  ND4D1BWP12T U4590 ( .A1(n3658), .A2(n3657), .A3(n3656), .A4(n3655), .ZN(
        regC_out[21]) );
  AOI22D1BWP12T U4591 ( .A1(r3[20]), .A2(n3880), .B1(r1[20]), .B2(n3882), .ZN(
        n3668) );
  AOI22D1BWP12T U4592 ( .A1(sp_out[20]), .A2(n3885), .B1(r12[20]), .B2(n3884), 
        .ZN(n3667) );
  AOI22D1BWP12T U4593 ( .A1(lr[20]), .A2(n3831), .B1(r0[20]), .B2(n3881), .ZN(
        n3666) );
  AOI22D1BWP12T U4594 ( .A1(r7[20]), .A2(n3524), .B1(r8[20]), .B2(n3871), .ZN(
        n3662) );
  AOI22D1BWP12T U4595 ( .A1(r4[20]), .A2(n3832), .B1(r9[20]), .B2(n3872), .ZN(
        n3661) );
  AOI22D1BWP12T U4596 ( .A1(r11[20]), .A2(n3595), .B1(r10[20]), .B2(n3874), 
        .ZN(n3660) );
  AOI22D1BWP12T U4597 ( .A1(r6[20]), .A2(n3873), .B1(r5[20]), .B2(n3875), .ZN(
        n3659) );
  ND4D1BWP12T U4598 ( .A1(n3662), .A2(n3661), .A3(n3660), .A4(n3659), .ZN(
        n3664) );
  OAI22D1BWP12T U4599 ( .A1(n4882), .A2(n3837), .B1(n4528), .B2(n3852), .ZN(
        n3663) );
  AOI21D1BWP12T U4600 ( .A1(n3892), .A2(n3664), .B(n3663), .ZN(n3665) );
  ND4D1BWP12T U4601 ( .A1(n3668), .A2(n3667), .A3(n3666), .A4(n3665), .ZN(
        regC_out[20]) );
  AOI22D1BWP12T U4602 ( .A1(r6[19]), .A2(n3873), .B1(r4[19]), .B2(n3832), .ZN(
        n3672) );
  AOI22D1BWP12T U4603 ( .A1(r7[19]), .A2(n3524), .B1(r10[19]), .B2(n3874), 
        .ZN(n3671) );
  AOI22D1BWP12T U4604 ( .A1(r5[19]), .A2(n3875), .B1(r11[19]), .B2(n3595), 
        .ZN(n3670) );
  AOI22D1BWP12T U4605 ( .A1(r9[19]), .A2(n3872), .B1(r8[19]), .B2(n3871), .ZN(
        n3669) );
  ND4D1BWP12T U4606 ( .A1(n3672), .A2(n3671), .A3(n3670), .A4(n3669), .ZN(
        n3678) );
  AOI22D1BWP12T U4607 ( .A1(r0[19]), .A2(n3881), .B1(r2[19]), .B2(n3864), .ZN(
        n3676) );
  AOI22D1BWP12T U4608 ( .A1(r12[19]), .A2(n3884), .B1(sp_out[19]), .B2(n3885), 
        .ZN(n3675) );
  AOI22D1BWP12T U4609 ( .A1(lr[19]), .A2(n3831), .B1(r3[19]), .B2(n3880), .ZN(
        n3674) );
  AOI22D1BWP12T U4610 ( .A1(r1[19]), .A2(n3882), .B1(pc_out[19]), .B2(n3883), 
        .ZN(n3673) );
  ND4D1BWP12T U4611 ( .A1(n3676), .A2(n3675), .A3(n3674), .A4(n3673), .ZN(
        n3677) );
  AO21D1BWP12T U4612 ( .A1(n3892), .A2(n3678), .B(n3677), .Z(regC_out[19]) );
  AOI22D1BWP12T U4613 ( .A1(r10[18]), .A2(n3874), .B1(r6[18]), .B2(n3873), 
        .ZN(n3682) );
  AOI22D1BWP12T U4614 ( .A1(r5[18]), .A2(n3875), .B1(r9[18]), .B2(n3872), .ZN(
        n3681) );
  AOI22D1BWP12T U4615 ( .A1(r11[18]), .A2(n3595), .B1(r8[18]), .B2(n3871), 
        .ZN(n3680) );
  AOI22D1BWP12T U4616 ( .A1(r4[18]), .A2(n3832), .B1(r7[18]), .B2(n3524), .ZN(
        n3679) );
  ND4D1BWP12T U4617 ( .A1(n3682), .A2(n3681), .A3(n3680), .A4(n3679), .ZN(
        n3688) );
  AOI22D1BWP12T U4618 ( .A1(r0[18]), .A2(n3881), .B1(sp_out[18]), .B2(n3885), 
        .ZN(n3686) );
  AOI22D1BWP12T U4619 ( .A1(r2[18]), .A2(n3864), .B1(r3[18]), .B2(n3880), .ZN(
        n3685) );
  AOI22D1BWP12T U4620 ( .A1(lr[18]), .A2(n3831), .B1(r1[18]), .B2(n3882), .ZN(
        n3684) );
  AOI22D1BWP12T U4621 ( .A1(r12[18]), .A2(n3884), .B1(pc_out[18]), .B2(n3883), 
        .ZN(n3683) );
  ND4D1BWP12T U4622 ( .A1(n3686), .A2(n3685), .A3(n3684), .A4(n3683), .ZN(
        n3687) );
  AO21D1BWP12T U4623 ( .A1(n3892), .A2(n3688), .B(n3687), .Z(regC_out[18]) );
  AOI22D1BWP12T U4624 ( .A1(r4[17]), .A2(n3832), .B1(r6[17]), .B2(n3873), .ZN(
        n3692) );
  AOI22D1BWP12T U4625 ( .A1(r5[17]), .A2(n3875), .B1(r9[17]), .B2(n3872), .ZN(
        n3691) );
  AOI22D1BWP12T U4626 ( .A1(r8[17]), .A2(n3871), .B1(r7[17]), .B2(n3524), .ZN(
        n3690) );
  AOI22D1BWP12T U4627 ( .A1(r11[17]), .A2(n3595), .B1(r10[17]), .B2(n3874), 
        .ZN(n3689) );
  ND4D1BWP12T U4628 ( .A1(n3692), .A2(n3691), .A3(n3690), .A4(n3689), .ZN(
        n3698) );
  AOI22D1BWP12T U4629 ( .A1(lr[17]), .A2(n3831), .B1(sp_out[17]), .B2(n3885), 
        .ZN(n3696) );
  AOI22D1BWP12T U4630 ( .A1(r0[17]), .A2(n3881), .B1(r3[17]), .B2(n3880), .ZN(
        n3695) );
  AOI22D1BWP12T U4631 ( .A1(r2[17]), .A2(n3864), .B1(r1[17]), .B2(n3882), .ZN(
        n3694) );
  AOI22D1BWP12T U4632 ( .A1(r12[17]), .A2(n3884), .B1(pc_out[17]), .B2(n3883), 
        .ZN(n3693) );
  ND4D1BWP12T U4633 ( .A1(n3696), .A2(n3695), .A3(n3694), .A4(n3693), .ZN(
        n3697) );
  AO21D1BWP12T U4634 ( .A1(n3892), .A2(n3698), .B(n3697), .Z(regC_out[17]) );
  AOI22D1BWP12T U4635 ( .A1(r12[16]), .A2(n3884), .B1(r1[16]), .B2(n3882), 
        .ZN(n3708) );
  AOI22D1BWP12T U4636 ( .A1(r3[16]), .A2(n3880), .B1(r2[16]), .B2(n3864), .ZN(
        n3707) );
  AOI22D1BWP12T U4637 ( .A1(lr[16]), .A2(n3831), .B1(sp_out[16]), .B2(n3885), 
        .ZN(n3706) );
  AOI22D1BWP12T U4638 ( .A1(r10[16]), .A2(n3874), .B1(r11[16]), .B2(n3595), 
        .ZN(n3702) );
  AOI22D1BWP12T U4639 ( .A1(r8[16]), .A2(n3871), .B1(r5[16]), .B2(n3875), .ZN(
        n3701) );
  AOI22D1BWP12T U4640 ( .A1(r7[16]), .A2(n3524), .B1(r9[16]), .B2(n3872), .ZN(
        n3700) );
  AOI22D1BWP12T U4641 ( .A1(r6[16]), .A2(n3873), .B1(r4[16]), .B2(n3832), .ZN(
        n3699) );
  ND4D1BWP12T U4642 ( .A1(n3702), .A2(n3701), .A3(n3700), .A4(n3699), .ZN(
        n3704) );
  OAI22D1BWP12T U4643 ( .A1(n4481), .A2(n3852), .B1(n4876), .B2(n3814), .ZN(
        n3703) );
  AOI21D1BWP12T U4644 ( .A1(n3892), .A2(n3704), .B(n3703), .ZN(n3705) );
  ND4D1BWP12T U4645 ( .A1(n3708), .A2(n3707), .A3(n3706), .A4(n3705), .ZN(
        regC_out[16]) );
  AOI22D1BWP12T U4646 ( .A1(r1[15]), .A2(n3882), .B1(r3[15]), .B2(n3880), .ZN(
        n3718) );
  AOI22D1BWP12T U4647 ( .A1(r12[15]), .A2(n3884), .B1(r2[15]), .B2(n3864), 
        .ZN(n3717) );
  AOI22D1BWP12T U4648 ( .A1(sp_out[15]), .A2(n3885), .B1(lr[15]), .B2(n3831), 
        .ZN(n3716) );
  AOI22D1BWP12T U4649 ( .A1(r9[15]), .A2(n3872), .B1(r8[15]), .B2(n3871), .ZN(
        n3712) );
  AOI22D1BWP12T U4650 ( .A1(r10[15]), .A2(n3874), .B1(r11[15]), .B2(n3595), 
        .ZN(n3711) );
  AOI22D1BWP12T U4651 ( .A1(r5[15]), .A2(n3875), .B1(r7[15]), .B2(n3524), .ZN(
        n3710) );
  AOI22D1BWP12T U4652 ( .A1(r6[15]), .A2(n3873), .B1(r4[15]), .B2(n3832), .ZN(
        n3709) );
  ND4D1BWP12T U4653 ( .A1(n3712), .A2(n3711), .A3(n3710), .A4(n3709), .ZN(
        n3714) );
  OAI22D1BWP12T U4654 ( .A1(n4828), .A2(n3814), .B1(n4886), .B2(n3852), .ZN(
        n3713) );
  AOI21D1BWP12T U4655 ( .A1(n3892), .A2(n3714), .B(n3713), .ZN(n3715) );
  ND4D1BWP12T U4656 ( .A1(n3718), .A2(n3717), .A3(n3716), .A4(n3715), .ZN(
        regC_out[15]) );
  AOI22D1BWP12T U4657 ( .A1(r11[14]), .A2(n3595), .B1(r10[14]), .B2(n3874), 
        .ZN(n3722) );
  AOI22D1BWP12T U4658 ( .A1(r4[14]), .A2(n3832), .B1(r8[14]), .B2(n3871), .ZN(
        n3721) );
  AOI22D1BWP12T U4659 ( .A1(r9[14]), .A2(n3872), .B1(r7[14]), .B2(n3524), .ZN(
        n3720) );
  AOI22D1BWP12T U4660 ( .A1(r6[14]), .A2(n3873), .B1(r5[14]), .B2(n3875), .ZN(
        n3719) );
  ND4D1BWP12T U4661 ( .A1(n3722), .A2(n3721), .A3(n3720), .A4(n3719), .ZN(
        n3728) );
  AOI22D1BWP12T U4662 ( .A1(r12[14]), .A2(n3884), .B1(r0[14]), .B2(n3881), 
        .ZN(n3726) );
  AOI22D1BWP12T U4663 ( .A1(r3[14]), .A2(n3880), .B1(pc_out[14]), .B2(n3883), 
        .ZN(n3725) );
  AOI22D1BWP12T U4664 ( .A1(sp_out[14]), .A2(n3885), .B1(r2[14]), .B2(n3864), 
        .ZN(n3724) );
  AOI22D1BWP12T U4665 ( .A1(r1[14]), .A2(n3882), .B1(lr[14]), .B2(n3831), .ZN(
        n3723) );
  ND4D1BWP12T U4666 ( .A1(n3726), .A2(n3725), .A3(n3724), .A4(n3723), .ZN(
        n3727) );
  AO21D1BWP12T U4667 ( .A1(n3892), .A2(n3728), .B(n3727), .Z(regC_out[14]) );
  AOI22D1BWP12T U4668 ( .A1(r12[13]), .A2(n3884), .B1(r0[13]), .B2(n3881), 
        .ZN(n3738) );
  AOI22D1BWP12T U4669 ( .A1(r2[13]), .A2(n3864), .B1(r1[13]), .B2(n3882), .ZN(
        n3737) );
  AOI22D1BWP12T U4670 ( .A1(sp_out[13]), .A2(n3885), .B1(r3[13]), .B2(n3880), 
        .ZN(n3736) );
  AOI22D1BWP12T U4671 ( .A1(r7[13]), .A2(n3524), .B1(r10[13]), .B2(n3874), 
        .ZN(n3732) );
  AOI22D1BWP12T U4672 ( .A1(r11[13]), .A2(n3595), .B1(r4[13]), .B2(n3832), 
        .ZN(n3731) );
  AOI22D1BWP12T U4673 ( .A1(r9[13]), .A2(n3872), .B1(r8[13]), .B2(n3871), .ZN(
        n3730) );
  AOI22D1BWP12T U4674 ( .A1(r6[13]), .A2(n3873), .B1(r5[13]), .B2(n3875), .ZN(
        n3729) );
  ND4D1BWP12T U4675 ( .A1(n3732), .A2(n3731), .A3(n3730), .A4(n3729), .ZN(
        n3734) );
  OAI22D1BWP12T U4676 ( .A1(n4436), .A2(n3852), .B1(n4857), .B2(n3849), .ZN(
        n3733) );
  AOI21D1BWP12T U4677 ( .A1(n3892), .A2(n3734), .B(n3733), .ZN(n3735) );
  ND4D1BWP12T U4678 ( .A1(n3738), .A2(n3737), .A3(n3736), .A4(n3735), .ZN(
        regC_out[13]) );
  AOI22D1BWP12T U4679 ( .A1(r3[12]), .A2(n3880), .B1(sp_out[12]), .B2(n3885), 
        .ZN(n3748) );
  AOI22D1BWP12T U4680 ( .A1(r0[12]), .A2(n3881), .B1(r1[12]), .B2(n3882), .ZN(
        n3747) );
  AOI22D1BWP12T U4681 ( .A1(r12[12]), .A2(n3884), .B1(r2[12]), .B2(n3864), 
        .ZN(n3746) );
  AOI22D1BWP12T U4682 ( .A1(r8[12]), .A2(n3871), .B1(r10[12]), .B2(n3874), 
        .ZN(n3742) );
  AOI22D1BWP12T U4683 ( .A1(r4[12]), .A2(n3832), .B1(r7[12]), .B2(n3524), .ZN(
        n3741) );
  AOI22D1BWP12T U4684 ( .A1(r5[12]), .A2(n3875), .B1(r11[12]), .B2(n3595), 
        .ZN(n3740) );
  AOI22D1BWP12T U4685 ( .A1(r6[12]), .A2(n3873), .B1(r9[12]), .B2(n3872), .ZN(
        n3739) );
  ND4D1BWP12T U4686 ( .A1(n3742), .A2(n3741), .A3(n3740), .A4(n3739), .ZN(
        n3744) );
  OAI22D1BWP12T U4687 ( .A1(n4851), .A2(n3849), .B1(n4424), .B2(n3852), .ZN(
        n3743) );
  AOI21D1BWP12T U4688 ( .A1(n3892), .A2(n3744), .B(n3743), .ZN(n3745) );
  ND4D1BWP12T U4689 ( .A1(n3748), .A2(n3747), .A3(n3746), .A4(n3745), .ZN(
        regC_out[12]) );
  AOI22D1BWP12T U4690 ( .A1(r9[11]), .A2(n3872), .B1(r5[11]), .B2(n3875), .ZN(
        n3752) );
  AOI22D1BWP12T U4691 ( .A1(r10[11]), .A2(n3874), .B1(r4[11]), .B2(n3832), 
        .ZN(n3751) );
  AOI22D1BWP12T U4692 ( .A1(r8[11]), .A2(n3871), .B1(r6[11]), .B2(n3873), .ZN(
        n3750) );
  AOI22D1BWP12T U4693 ( .A1(r11[11]), .A2(n3595), .B1(r7[11]), .B2(n3524), 
        .ZN(n3749) );
  ND4D1BWP12T U4694 ( .A1(n3752), .A2(n3751), .A3(n3750), .A4(n3749), .ZN(
        n3758) );
  AOI22D1BWP12T U4695 ( .A1(r2[11]), .A2(n3864), .B1(sp_out[11]), .B2(n3885), 
        .ZN(n3756) );
  AOI22D1BWP12T U4696 ( .A1(r3[11]), .A2(n3880), .B1(r12[11]), .B2(n3884), 
        .ZN(n3755) );
  AOI22D1BWP12T U4697 ( .A1(lr[11]), .A2(n3831), .B1(r1[11]), .B2(n3882), .ZN(
        n3754) );
  AOI22D1BWP12T U4698 ( .A1(r0[11]), .A2(n3881), .B1(pc_out[11]), .B2(n3883), 
        .ZN(n3753) );
  ND4D1BWP12T U4699 ( .A1(n3756), .A2(n3755), .A3(n3754), .A4(n3753), .ZN(
        n3757) );
  AO21D1BWP12T U4700 ( .A1(n3892), .A2(n3758), .B(n3757), .Z(regC_out[11]) );
  AOI22D1BWP12T U4701 ( .A1(r11[10]), .A2(n3595), .B1(r10[10]), .B2(n3874), 
        .ZN(n3762) );
  AOI22D1BWP12T U4702 ( .A1(r6[10]), .A2(n3873), .B1(r4[10]), .B2(n3832), .ZN(
        n3761) );
  AOI22D1BWP12T U4703 ( .A1(r9[10]), .A2(n3872), .B1(r8[10]), .B2(n3871), .ZN(
        n3760) );
  AOI22D1BWP12T U4704 ( .A1(r5[10]), .A2(n3875), .B1(r7[10]), .B2(n3524), .ZN(
        n3759) );
  ND4D1BWP12T U4705 ( .A1(n3762), .A2(n3761), .A3(n3760), .A4(n3759), .ZN(
        n3768) );
  AOI22D1BWP12T U4706 ( .A1(r3[10]), .A2(n3880), .B1(sp_out[10]), .B2(n3885), 
        .ZN(n3766) );
  AOI22D1BWP12T U4707 ( .A1(r0[10]), .A2(n3881), .B1(lr[10]), .B2(n3831), .ZN(
        n3765) );
  AOI22D1BWP12T U4708 ( .A1(pc_out[10]), .A2(n3883), .B1(r1[10]), .B2(n3882), 
        .ZN(n3764) );
  AOI22D1BWP12T U4709 ( .A1(r12[10]), .A2(n3884), .B1(r2[10]), .B2(n3864), 
        .ZN(n3763) );
  ND4D1BWP12T U4710 ( .A1(n3766), .A2(n3765), .A3(n3764), .A4(n3763), .ZN(
        n3767) );
  AO21D1BWP12T U4711 ( .A1(n3892), .A2(n3768), .B(n3767), .Z(regC_out[10]) );
  AOI22D1BWP12T U4712 ( .A1(lr[9]), .A2(n3831), .B1(sp_out[9]), .B2(n3885), 
        .ZN(n3779) );
  AOI22D1BWP12T U4713 ( .A1(r2[9]), .A2(n3864), .B1(r3[9]), .B2(n3880), .ZN(
        n3778) );
  AOI22D1BWP12T U4714 ( .A1(r12[9]), .A2(n3884), .B1(r1[9]), .B2(n3882), .ZN(
        n3777) );
  AOI22D1BWP12T U4715 ( .A1(r6[9]), .A2(n3873), .B1(r11[9]), .B2(n3595), .ZN(
        n3772) );
  AOI22D1BWP12T U4716 ( .A1(r4[9]), .A2(n3832), .B1(r8[9]), .B2(n3871), .ZN(
        n3771) );
  AOI22D1BWP12T U4717 ( .A1(r9[9]), .A2(n3872), .B1(r5[9]), .B2(n3875), .ZN(
        n3770) );
  AOI22D1BWP12T U4718 ( .A1(r7[9]), .A2(n3524), .B1(r10[9]), .B2(n3874), .ZN(
        n3769) );
  ND4D1BWP12T U4719 ( .A1(n3772), .A2(n3771), .A3(n3770), .A4(n3769), .ZN(
        n3775) );
  OAI22D1BWP12T U4720 ( .A1(n3773), .A2(n3852), .B1(n4854), .B2(n3814), .ZN(
        n3774) );
  AOI21D1BWP12T U4721 ( .A1(n3892), .A2(n3775), .B(n3774), .ZN(n3776) );
  ND4D1BWP12T U4722 ( .A1(n3779), .A2(n3778), .A3(n3777), .A4(n3776), .ZN(
        regC_out[9]) );
  AOI22D1BWP12T U4723 ( .A1(r11[8]), .A2(n3595), .B1(r7[8]), .B2(n3524), .ZN(
        n3783) );
  AOI22D1BWP12T U4724 ( .A1(r9[8]), .A2(n3872), .B1(r10[8]), .B2(n3874), .ZN(
        n3782) );
  AOI22D1BWP12T U4725 ( .A1(r8[8]), .A2(n3871), .B1(r6[8]), .B2(n3873), .ZN(
        n3781) );
  AOI22D1BWP12T U4726 ( .A1(r5[8]), .A2(n3875), .B1(r4[8]), .B2(n3832), .ZN(
        n3780) );
  ND4D1BWP12T U4727 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(
        n3789) );
  AOI22D1BWP12T U4728 ( .A1(r0[8]), .A2(n3881), .B1(r3[8]), .B2(n3880), .ZN(
        n3787) );
  AOI22D1BWP12T U4729 ( .A1(r2[8]), .A2(n3864), .B1(sp_out[8]), .B2(n3885), 
        .ZN(n3786) );
  AOI22D1BWP12T U4730 ( .A1(lr[8]), .A2(n3831), .B1(r1[8]), .B2(n3882), .ZN(
        n3785) );
  AOI22D1BWP12T U4731 ( .A1(r12[8]), .A2(n3884), .B1(pc_out[8]), .B2(n3883), 
        .ZN(n3784) );
  ND4D1BWP12T U4732 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(
        n3788) );
  AO21D1BWP12T U4733 ( .A1(n3892), .A2(n3789), .B(n3788), .Z(regC_out[8]) );
  AOI22D1BWP12T U4734 ( .A1(r8[7]), .A2(n3871), .B1(r11[7]), .B2(n3595), .ZN(
        n3793) );
  AOI22D1BWP12T U4735 ( .A1(r7[7]), .A2(n3524), .B1(r10[7]), .B2(n3874), .ZN(
        n3792) );
  AOI22D1BWP12T U4736 ( .A1(r4[7]), .A2(n3832), .B1(r6[7]), .B2(n3873), .ZN(
        n3791) );
  AOI22D1BWP12T U4737 ( .A1(r9[7]), .A2(n3872), .B1(r5[7]), .B2(n3875), .ZN(
        n3790) );
  ND4D1BWP12T U4738 ( .A1(n3793), .A2(n3792), .A3(n3791), .A4(n3790), .ZN(
        n3799) );
  AOI22D1BWP12T U4739 ( .A1(r0[7]), .A2(n3881), .B1(r1[7]), .B2(n3882), .ZN(
        n3797) );
  AOI22D1BWP12T U4740 ( .A1(r12[7]), .A2(n3884), .B1(r3[7]), .B2(n3880), .ZN(
        n3796) );
  AOI22D1BWP12T U4741 ( .A1(sp_out[7]), .A2(n3885), .B1(r2[7]), .B2(n3864), 
        .ZN(n3795) );
  AOI22D1BWP12T U4742 ( .A1(pc_out[7]), .A2(n3883), .B1(lr[7]), .B2(n3831), 
        .ZN(n3794) );
  ND4D1BWP12T U4743 ( .A1(n3797), .A2(n3796), .A3(n3795), .A4(n3794), .ZN(
        n3798) );
  AO21D1BWP12T U4744 ( .A1(n3892), .A2(n3799), .B(n3798), .Z(regC_out[7]) );
  AOI22D1BWP12T U4745 ( .A1(r3[6]), .A2(n3880), .B1(r1[6]), .B2(n3882), .ZN(
        n3809) );
  AOI22D1BWP12T U4746 ( .A1(r2[6]), .A2(n3864), .B1(sp_out[6]), .B2(n3885), 
        .ZN(n3808) );
  AOI22D1BWP12T U4747 ( .A1(r0[6]), .A2(n3881), .B1(lr[6]), .B2(n3831), .ZN(
        n3807) );
  AOI22D1BWP12T U4748 ( .A1(r5[6]), .A2(n3875), .B1(r11[6]), .B2(n3595), .ZN(
        n3803) );
  AOI22D1BWP12T U4749 ( .A1(r6[6]), .A2(n3873), .B1(r7[6]), .B2(n3524), .ZN(
        n3802) );
  AOI22D1BWP12T U4750 ( .A1(r4[6]), .A2(n3832), .B1(r8[6]), .B2(n3871), .ZN(
        n3801) );
  AOI22D1BWP12T U4751 ( .A1(r9[6]), .A2(n3872), .B1(r10[6]), .B2(n3874), .ZN(
        n3800) );
  ND4D1BWP12T U4752 ( .A1(n3803), .A2(n3802), .A3(n3801), .A4(n3800), .ZN(
        n3805) );
  OAI22D1BWP12T U4753 ( .A1(n4163), .A2(n3851), .B1(n4353), .B2(n3852), .ZN(
        n3804) );
  AOI21D1BWP12T U4754 ( .A1(n3892), .A2(n3805), .B(n3804), .ZN(n3806) );
  ND4D1BWP12T U4755 ( .A1(n3809), .A2(n3808), .A3(n3807), .A4(n3806), .ZN(
        regC_out[6]) );
  AOI22D1BWP12T U4756 ( .A1(r1[5]), .A2(n3882), .B1(r2[5]), .B2(n3864), .ZN(
        n3820) );
  AOI22D1BWP12T U4757 ( .A1(lr[5]), .A2(n3831), .B1(r3[5]), .B2(n3880), .ZN(
        n3819) );
  AOI22D1BWP12T U4758 ( .A1(r12[5]), .A2(n3884), .B1(sp_out[5]), .B2(n3885), 
        .ZN(n3818) );
  AOI22D1BWP12T U4759 ( .A1(r11[5]), .A2(n3595), .B1(r6[5]), .B2(n3873), .ZN(
        n3813) );
  AOI22D1BWP12T U4760 ( .A1(r4[5]), .A2(n3832), .B1(r9[5]), .B2(n3872), .ZN(
        n3812) );
  AOI22D1BWP12T U4761 ( .A1(r10[5]), .A2(n3874), .B1(r5[5]), .B2(n3875), .ZN(
        n3811) );
  AOI22D1BWP12T U4762 ( .A1(r8[5]), .A2(n3871), .B1(r7[5]), .B2(n3524), .ZN(
        n3810) );
  ND4D1BWP12T U4763 ( .A1(n3813), .A2(n3812), .A3(n3811), .A4(n3810), .ZN(
        n3816) );
  OAI22D1BWP12T U4764 ( .A1(n4839), .A2(n3814), .B1(n4341), .B2(n3852), .ZN(
        n3815) );
  AOI21D1BWP12T U4765 ( .A1(n3892), .A2(n3816), .B(n3815), .ZN(n3817) );
  ND4D1BWP12T U4766 ( .A1(n3820), .A2(n3819), .A3(n3818), .A4(n3817), .ZN(
        regC_out[5]) );
  AOI22D1BWP12T U4767 ( .A1(r8[4]), .A2(n3871), .B1(r10[4]), .B2(n3874), .ZN(
        n3824) );
  AOI22D1BWP12T U4768 ( .A1(r6[4]), .A2(n3873), .B1(r11[4]), .B2(n3595), .ZN(
        n3823) );
  AOI22D1BWP12T U4769 ( .A1(r4[4]), .A2(n3832), .B1(r7[4]), .B2(n3524), .ZN(
        n3822) );
  AOI22D1BWP12T U4770 ( .A1(r9[4]), .A2(n3872), .B1(r5[4]), .B2(n3875), .ZN(
        n3821) );
  ND4D1BWP12T U4771 ( .A1(n3824), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(
        n3830) );
  AOI22D1BWP12T U4772 ( .A1(r1[4]), .A2(n3882), .B1(r0[4]), .B2(n3881), .ZN(
        n3828) );
  AOI22D1BWP12T U4773 ( .A1(r12[4]), .A2(n3884), .B1(r2[4]), .B2(n3864), .ZN(
        n3827) );
  AOI22D1BWP12T U4774 ( .A1(r3[4]), .A2(n3880), .B1(pc_out[4]), .B2(n3883), 
        .ZN(n3826) );
  AOI22D1BWP12T U4775 ( .A1(sp_out[4]), .A2(n3885), .B1(lr[4]), .B2(n3831), 
        .ZN(n3825) );
  ND4D1BWP12T U4776 ( .A1(n3828), .A2(n3827), .A3(n3826), .A4(n3825), .ZN(
        n3829) );
  AO21D1BWP12T U4777 ( .A1(n3892), .A2(n3830), .B(n3829), .Z(regC_out[4]) );
  AOI22D1BWP12T U4778 ( .A1(sp_out[3]), .A2(n3885), .B1(r1[3]), .B2(n3882), 
        .ZN(n3844) );
  AOI22D1BWP12T U4779 ( .A1(lr[3]), .A2(n3831), .B1(r0[3]), .B2(n3881), .ZN(
        n3843) );
  AOI22D1BWP12T U4780 ( .A1(r12[3]), .A2(n3884), .B1(r3[3]), .B2(n3880), .ZN(
        n3842) );
  AOI22D1BWP12T U4781 ( .A1(r6[3]), .A2(n3873), .B1(r9[3]), .B2(n3872), .ZN(
        n3836) );
  AOI22D1BWP12T U4782 ( .A1(r5[3]), .A2(n3875), .B1(r4[3]), .B2(n3832), .ZN(
        n3835) );
  AOI22D1BWP12T U4783 ( .A1(r7[3]), .A2(n3524), .B1(r8[3]), .B2(n3871), .ZN(
        n3834) );
  AOI22D1BWP12T U4784 ( .A1(r10[3]), .A2(n3874), .B1(r11[3]), .B2(n3595), .ZN(
        n3833) );
  ND4D1BWP12T U4785 ( .A1(n3836), .A2(n3835), .A3(n3834), .A4(n3833), .ZN(
        n3840) );
  OAI22D1BWP12T U4786 ( .A1(n3838), .A2(n3837), .B1(n4317), .B2(n3852), .ZN(
        n3839) );
  AOI21D1BWP12T U4787 ( .A1(n3892), .A2(n3840), .B(n3839), .ZN(n3841) );
  ND4D1BWP12T U4788 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(
        regC_out[3]) );
  AOI22D1BWP12T U4789 ( .A1(sp_out[2]), .A2(n3885), .B1(r1[2]), .B2(n3882), 
        .ZN(n3859) );
  AOI22D1BWP12T U4790 ( .A1(r2[2]), .A2(n3864), .B1(r0[2]), .B2(n3881), .ZN(
        n3858) );
  AOI22D1BWP12T U4791 ( .A1(r10[2]), .A2(n3874), .B1(r5[2]), .B2(n3875), .ZN(
        n3848) );
  AOI22D1BWP12T U4792 ( .A1(r6[2]), .A2(n3873), .B1(r4[2]), .B2(n3832), .ZN(
        n3847) );
  AOI22D1BWP12T U4793 ( .A1(r9[2]), .A2(n3872), .B1(r11[2]), .B2(n3595), .ZN(
        n3846) );
  AOI22D1BWP12T U4794 ( .A1(r8[2]), .A2(n3871), .B1(r7[2]), .B2(n3524), .ZN(
        n3845) );
  ND4D1BWP12T U4795 ( .A1(n3848), .A2(n3847), .A3(n3846), .A4(n3845), .ZN(
        n3856) );
  OAI22D1BWP12T U4796 ( .A1(n4864), .A2(n3851), .B1(n3850), .B2(n3849), .ZN(
        n3855) );
  INVD1BWP12T U4797 ( .I(pc_out[2]), .ZN(n4305) );
  OAI22D1BWP12T U4798 ( .A1(n4207), .A2(n3853), .B1(n4305), .B2(n3852), .ZN(
        n3854) );
  AOI211D1BWP12T U4799 ( .A1(n3892), .A2(n3856), .B(n3855), .C(n3854), .ZN(
        n3857) );
  ND3D1BWP12T U4800 ( .A1(n3859), .A2(n3858), .A3(n3857), .ZN(regC_out[2]) );
  AOI22D1BWP12T U4801 ( .A1(r10[1]), .A2(n3874), .B1(r8[1]), .B2(n3871), .ZN(
        n3863) );
  AOI22D1BWP12T U4802 ( .A1(r7[1]), .A2(n3524), .B1(r6[1]), .B2(n3873), .ZN(
        n3862) );
  AOI22D1BWP12T U4803 ( .A1(r4[1]), .A2(n3832), .B1(r9[1]), .B2(n3872), .ZN(
        n3861) );
  AOI22D1BWP12T U4804 ( .A1(r5[1]), .A2(n3875), .B1(r11[1]), .B2(n3595), .ZN(
        n3860) );
  ND4D1BWP12T U4805 ( .A1(n3863), .A2(n3862), .A3(n3861), .A4(n3860), .ZN(
        n3870) );
  AOI22D1BWP12T U4806 ( .A1(r0[1]), .A2(n3881), .B1(r2[1]), .B2(n3864), .ZN(
        n3868) );
  AOI22D1BWP12T U4807 ( .A1(r1[1]), .A2(n3882), .B1(lr[1]), .B2(n3831), .ZN(
        n3867) );
  AOI22D1BWP12T U4808 ( .A1(r3[1]), .A2(n3880), .B1(sp_out[1]), .B2(n3885), 
        .ZN(n3866) );
  AOI22D1BWP12T U4809 ( .A1(r12[1]), .A2(n3884), .B1(pc_out[1]), .B2(n3883), 
        .ZN(n3865) );
  ND4D1BWP12T U4810 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(
        n3869) );
  AO21D1BWP12T U4811 ( .A1(n3892), .A2(n3870), .B(n3869), .Z(regC_out[1]) );
  AOI22D1BWP12T U4812 ( .A1(r4[0]), .A2(n3832), .B1(r8[0]), .B2(n3871), .ZN(
        n3879) );
  AOI22D1BWP12T U4813 ( .A1(r9[0]), .A2(n3872), .B1(r7[0]), .B2(n3524), .ZN(
        n3878) );
  AOI22D1BWP12T U4814 ( .A1(r10[0]), .A2(n3874), .B1(r6[0]), .B2(n3873), .ZN(
        n3877) );
  AOI22D1BWP12T U4815 ( .A1(r11[0]), .A2(n3595), .B1(r5[0]), .B2(n3875), .ZN(
        n3876) );
  ND4D1BWP12T U4816 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(
        n3891) );
  AOI22D1BWP12T U4817 ( .A1(r2[0]), .A2(n3864), .B1(r3[0]), .B2(n3880), .ZN(
        n3889) );
  AOI22D1BWP12T U4818 ( .A1(r1[0]), .A2(n3882), .B1(r0[0]), .B2(n3881), .ZN(
        n3888) );
  AOI22D1BWP12T U4819 ( .A1(r12[0]), .A2(n3884), .B1(pc_out[0]), .B2(n3883), 
        .ZN(n3887) );
  AOI22D1BWP12T U4820 ( .A1(sp_out[0]), .A2(n3885), .B1(lr[0]), .B2(n3831), 
        .ZN(n3886) );
  ND4D1BWP12T U4821 ( .A1(n3889), .A2(n3888), .A3(n3887), .A4(n3886), .ZN(
        n3890) );
  AO21D1BWP12T U4822 ( .A1(n3892), .A2(n3891), .B(n3890), .Z(regC_out[0]) );
  INVD1BWP12T U4823 ( .I(readD_sel[4]), .ZN(n4463) );
  IND2D1BWP12T U4824 ( .A1(readD_sel[3]), .B1(readD_sel[2]), .ZN(n3893) );
  OR2XD1BWP12T U4825 ( .A1(readD_sel[0]), .A2(readD_sel[1]), .Z(n3900) );
  NR2D1BWP12T U4826 ( .A1(n3893), .A2(n3900), .ZN(n3942) );
  IND2D1BWP12T U4827 ( .A1(readD_sel[2]), .B1(readD_sel[3]), .ZN(n3894) );
  NR2D1BWP12T U4828 ( .A1(n3900), .A2(n3894), .ZN(n4452) );
  AOI22D1BWP12T U4829 ( .A1(r4[31]), .A2(n3942), .B1(r8[31]), .B2(n4452), .ZN(
        n3898) );
  IND2D1BWP12T U4830 ( .A1(readD_sel[1]), .B1(readD_sel[0]), .ZN(n3899) );
  NR2D1BWP12T U4831 ( .A1(n3894), .A2(n3899), .ZN(n4218) );
  IND2D1BWP12T U4832 ( .A1(readD_sel[0]), .B1(readD_sel[1]), .ZN(n3904) );
  NR2D1BWP12T U4833 ( .A1(n3904), .A2(n3893), .ZN(n4451) );
  AOI22D1BWP12T U4834 ( .A1(r9[31]), .A2(n4218), .B1(r6[31]), .B2(n4451), .ZN(
        n3897) );
  ND2D1BWP12T U4835 ( .A1(readD_sel[0]), .A2(readD_sel[1]), .ZN(n3902) );
  NR2D1BWP12T U4836 ( .A1(n3894), .A2(n3902), .ZN(n3953) );
  NR2D1BWP12T U4837 ( .A1(n3893), .A2(n3899), .ZN(n4453) );
  AOI22D1BWP12T U4838 ( .A1(r11[31]), .A2(n3953), .B1(r5[31]), .B2(n4453), 
        .ZN(n3896) );
  NR2D1BWP12T U4839 ( .A1(n3893), .A2(n3902), .ZN(n3985) );
  NR2D1BWP12T U4840 ( .A1(n3904), .A2(n3894), .ZN(n4217) );
  AOI22D1BWP12T U4841 ( .A1(r7[31]), .A2(n3985), .B1(r10[31]), .B2(n4217), 
        .ZN(n3895) );
  ND4D1BWP12T U4842 ( .A1(n3898), .A2(n3897), .A3(n3896), .A4(n3895), .ZN(
        n3910) );
  ND3D1BWP12T U4843 ( .A1(readD_sel[2]), .A2(readD_sel[3]), .A3(n4463), .ZN(
        n3901) );
  NR2D1BWP12T U4844 ( .A1(n3904), .A2(n3901), .ZN(n4447) );
  INVD1BWP12T U4845 ( .I(n4447), .ZN(n4184) );
  OR3XD1BWP12T U4846 ( .A1(readD_sel[4]), .A2(readD_sel[2]), .A3(readD_sel[3]), 
        .Z(n3903) );
  NR2D1BWP12T U4847 ( .A1(n3899), .A2(n3903), .ZN(n4450) );
  AOI22D1BWP12T U4848 ( .A1(lr[31]), .A2(n4447), .B1(r1[31]), .B2(n4450), .ZN(
        n3908) );
  NR2D1BWP12T U4849 ( .A1(n3899), .A2(n3901), .ZN(n4449) );
  NR2D1BWP12T U4850 ( .A1(n3902), .A2(n3903), .ZN(n4214) );
  INVD1BWP12T U4851 ( .I(n4214), .ZN(n4206) );
  AOI22D1BWP12T U4852 ( .A1(sp_out[31]), .A2(n4449), .B1(r3[31]), .B2(n4214), 
        .ZN(n3907) );
  NR2D1BWP12T U4853 ( .A1(n3900), .A2(n3903), .ZN(n4448) );
  OR2XD1BWP12T U4854 ( .A1(n3900), .A2(n3901), .Z(n4460) );
  INVD1BWP12T U4855 ( .I(n4460), .ZN(n4215) );
  AOI22D1BWP12T U4856 ( .A1(r0[31]), .A2(n4448), .B1(r12[31]), .B2(n4215), 
        .ZN(n3906) );
  NR2D1BWP12T U4857 ( .A1(n3902), .A2(n3901), .ZN(n4195) );
  NR2D1BWP12T U4858 ( .A1(n3904), .A2(n3903), .ZN(n4216) );
  INVD1BWP12T U4859 ( .I(n4216), .ZN(n4091) );
  AOI22D1BWP12T U4860 ( .A1(pc_out[31]), .A2(n4195), .B1(r2[31]), .B2(n4216), 
        .ZN(n3905) );
  ND4D1BWP12T U4861 ( .A1(n3908), .A2(n3907), .A3(n3906), .A4(n3905), .ZN(
        n3909) );
  AO21D1BWP12T U4862 ( .A1(n4463), .A2(n3910), .B(n3909), .Z(regD_out[31]) );
  AOI22D1BWP12T U4863 ( .A1(r4[30]), .A2(n3942), .B1(r10[30]), .B2(n4217), 
        .ZN(n3914) );
  AOI22D1BWP12T U4864 ( .A1(r11[30]), .A2(n3953), .B1(r8[30]), .B2(n4452), 
        .ZN(n3913) );
  AOI22D1BWP12T U4865 ( .A1(r9[30]), .A2(n4218), .B1(r6[30]), .B2(n4451), .ZN(
        n3912) );
  AOI22D1BWP12T U4866 ( .A1(r5[30]), .A2(n4453), .B1(r7[30]), .B2(n3985), .ZN(
        n3911) );
  ND4D1BWP12T U4867 ( .A1(n3914), .A2(n3913), .A3(n3912), .A4(n3911), .ZN(
        n3920) );
  AOI22D1BWP12T U4868 ( .A1(r12[30]), .A2(n4215), .B1(sp_out[30]), .B2(n4449), 
        .ZN(n3918) );
  AOI22D1BWP12T U4869 ( .A1(r1[30]), .A2(n4450), .B1(r2[30]), .B2(n4216), .ZN(
        n3917) );
  AOI22D1BWP12T U4870 ( .A1(lr[30]), .A2(n4447), .B1(r3[30]), .B2(n4214), .ZN(
        n3916) );
  AOI22D1BWP12T U4871 ( .A1(pc_out[30]), .A2(n4195), .B1(r0[30]), .B2(n4448), 
        .ZN(n3915) );
  ND4D1BWP12T U4872 ( .A1(n3918), .A2(n3917), .A3(n3916), .A4(n3915), .ZN(
        n3919) );
  AO21D1BWP12T U4873 ( .A1(n4463), .A2(n3920), .B(n3919), .Z(regD_out[30]) );
  AOI22D1BWP12T U4874 ( .A1(r3[29]), .A2(n4214), .B1(r0[29]), .B2(n4448), .ZN(
        n3931) );
  AOI22D1BWP12T U4875 ( .A1(lr[29]), .A2(n4447), .B1(r2[29]), .B2(n4216), .ZN(
        n3930) );
  AOI22D1BWP12T U4876 ( .A1(r12[29]), .A2(n4215), .B1(r1[29]), .B2(n4450), 
        .ZN(n3929) );
  AOI22D1BWP12T U4877 ( .A1(r11[29]), .A2(n3953), .B1(r7[29]), .B2(n3985), 
        .ZN(n3924) );
  AOI22D1BWP12T U4878 ( .A1(r8[29]), .A2(n4452), .B1(r4[29]), .B2(n3942), .ZN(
        n3923) );
  AOI22D1BWP12T U4879 ( .A1(r6[29]), .A2(n4451), .B1(r9[29]), .B2(n4218), .ZN(
        n3922) );
  AOI22D1BWP12T U4880 ( .A1(r10[29]), .A2(n4217), .B1(r5[29]), .B2(n4453), 
        .ZN(n3921) );
  ND4D1BWP12T U4881 ( .A1(n3924), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(
        n3927) );
  INVD1BWP12T U4882 ( .I(n4195), .ZN(n4458) );
  MOAI22D0BWP12T U4883 ( .A1(n3925), .A2(n4458), .B1(sp_out[29]), .B2(n4449), 
        .ZN(n3926) );
  AOI21D1BWP12T U4884 ( .A1(n4463), .A2(n3927), .B(n3926), .ZN(n3928) );
  ND4D1BWP12T U4885 ( .A1(n3931), .A2(n3930), .A3(n3929), .A4(n3928), .ZN(
        regD_out[29]) );
  AOI22D1BWP12T U4886 ( .A1(r6[28]), .A2(n4451), .B1(r5[28]), .B2(n4453), .ZN(
        n3935) );
  AOI22D1BWP12T U4887 ( .A1(r11[28]), .A2(n3953), .B1(r8[28]), .B2(n4452), 
        .ZN(n3934) );
  AOI22D1BWP12T U4888 ( .A1(r10[28]), .A2(n4217), .B1(r9[28]), .B2(n4218), 
        .ZN(n3933) );
  AOI22D1BWP12T U4889 ( .A1(r4[28]), .A2(n3942), .B1(r7[28]), .B2(n3985), .ZN(
        n3932) );
  ND4D1BWP12T U4890 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(
        n3941) );
  AOI22D1BWP12T U4891 ( .A1(lr[28]), .A2(n4447), .B1(r12[28]), .B2(n4215), 
        .ZN(n3939) );
  AOI22D1BWP12T U4892 ( .A1(r1[28]), .A2(n4450), .B1(r2[28]), .B2(n4216), .ZN(
        n3938) );
  AOI22D1BWP12T U4893 ( .A1(r3[28]), .A2(n4214), .B1(pc_out[28]), .B2(n4195), 
        .ZN(n3937) );
  AOI22D1BWP12T U4894 ( .A1(r0[28]), .A2(n4448), .B1(sp_out[28]), .B2(n4449), 
        .ZN(n3936) );
  ND4D1BWP12T U4895 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(
        n3940) );
  AO21D1BWP12T U4896 ( .A1(n4463), .A2(n3941), .B(n3940), .Z(regD_out[28]) );
  AOI22D1BWP12T U4897 ( .A1(r8[27]), .A2(n4452), .B1(r5[27]), .B2(n4453), .ZN(
        n3946) );
  AOI22D1BWP12T U4898 ( .A1(r6[27]), .A2(n4451), .B1(r7[27]), .B2(n3985), .ZN(
        n3945) );
  AOI22D1BWP12T U4899 ( .A1(r4[27]), .A2(n3942), .B1(r11[27]), .B2(n3953), 
        .ZN(n3944) );
  AOI22D1BWP12T U4900 ( .A1(r10[27]), .A2(n4217), .B1(r9[27]), .B2(n4218), 
        .ZN(n3943) );
  ND4D1BWP12T U4901 ( .A1(n3946), .A2(n3945), .A3(n3944), .A4(n3943), .ZN(
        n3952) );
  AOI22D1BWP12T U4902 ( .A1(sp_out[27]), .A2(n4449), .B1(r2[27]), .B2(n4216), 
        .ZN(n3950) );
  AOI22D1BWP12T U4903 ( .A1(lr[27]), .A2(n4447), .B1(r1[27]), .B2(n4450), .ZN(
        n3949) );
  AOI22D1BWP12T U4904 ( .A1(r12[27]), .A2(n4215), .B1(pc_out[27]), .B2(n4195), 
        .ZN(n3948) );
  AOI22D1BWP12T U4905 ( .A1(r0[27]), .A2(n4448), .B1(r3[27]), .B2(n4214), .ZN(
        n3947) );
  ND4D1BWP12T U4906 ( .A1(n3950), .A2(n3949), .A3(n3948), .A4(n3947), .ZN(
        n3951) );
  AO21D1BWP12T U4907 ( .A1(n4463), .A2(n3952), .B(n3951), .Z(regD_out[27]) );
  AOI22D1BWP12T U4908 ( .A1(r11[26]), .A2(n3953), .B1(r9[26]), .B2(n4218), 
        .ZN(n3957) );
  AOI22D1BWP12T U4909 ( .A1(r5[26]), .A2(n4453), .B1(r6[26]), .B2(n4451), .ZN(
        n3956) );
  AOI22D1BWP12T U4910 ( .A1(r7[26]), .A2(n3985), .B1(r4[26]), .B2(n3942), .ZN(
        n3955) );
  AOI22D1BWP12T U4911 ( .A1(r10[26]), .A2(n4217), .B1(r8[26]), .B2(n4452), 
        .ZN(n3954) );
  ND4D1BWP12T U4912 ( .A1(n3957), .A2(n3956), .A3(n3955), .A4(n3954), .ZN(
        n3963) );
  AOI22D1BWP12T U4913 ( .A1(r2[26]), .A2(n4216), .B1(r12[26]), .B2(n4215), 
        .ZN(n3961) );
  AOI22D1BWP12T U4914 ( .A1(sp_out[26]), .A2(n4449), .B1(r3[26]), .B2(n4214), 
        .ZN(n3960) );
  AOI22D1BWP12T U4915 ( .A1(r1[26]), .A2(n4450), .B1(pc_out[26]), .B2(n4195), 
        .ZN(n3959) );
  AOI22D1BWP12T U4916 ( .A1(r0[26]), .A2(n4448), .B1(lr[26]), .B2(n4447), .ZN(
        n3958) );
  ND4D1BWP12T U4917 ( .A1(n3961), .A2(n3960), .A3(n3959), .A4(n3958), .ZN(
        n3962) );
  AO21D1BWP12T U4918 ( .A1(n4463), .A2(n3963), .B(n3962), .Z(regD_out[26]) );
  AOI22D1BWP12T U4919 ( .A1(r10[25]), .A2(n4217), .B1(r5[25]), .B2(n4453), 
        .ZN(n3967) );
  AOI22D1BWP12T U4920 ( .A1(r6[25]), .A2(n4451), .B1(r7[25]), .B2(n3985), .ZN(
        n3966) );
  AOI22D1BWP12T U4921 ( .A1(r4[25]), .A2(n3942), .B1(r9[25]), .B2(n4218), .ZN(
        n3965) );
  AOI22D1BWP12T U4922 ( .A1(r8[25]), .A2(n4452), .B1(r11[25]), .B2(n3953), 
        .ZN(n3964) );
  ND4D1BWP12T U4923 ( .A1(n3967), .A2(n3966), .A3(n3965), .A4(n3964), .ZN(
        n3973) );
  AOI22D1BWP12T U4924 ( .A1(r2[25]), .A2(n4216), .B1(r1[25]), .B2(n4450), .ZN(
        n3971) );
  AOI22D1BWP12T U4925 ( .A1(lr[25]), .A2(n4447), .B1(r3[25]), .B2(n4214), .ZN(
        n3970) );
  AOI22D1BWP12T U4926 ( .A1(r0[25]), .A2(n4448), .B1(r12[25]), .B2(n4215), 
        .ZN(n3969) );
  AOI22D1BWP12T U4927 ( .A1(pc_out[25]), .A2(n4195), .B1(sp_out[25]), .B2(
        n4449), .ZN(n3968) );
  ND4D1BWP12T U4928 ( .A1(n3971), .A2(n3970), .A3(n3969), .A4(n3968), .ZN(
        n3972) );
  AO21D1BWP12T U4929 ( .A1(n4463), .A2(n3973), .B(n3972), .Z(regD_out[25]) );
  AOI22D1BWP12T U4930 ( .A1(r2[24]), .A2(n4216), .B1(r12[24]), .B2(n4215), 
        .ZN(n3984) );
  AOI22D1BWP12T U4931 ( .A1(lr[24]), .A2(n4447), .B1(r1[24]), .B2(n4450), .ZN(
        n3983) );
  AOI22D1BWP12T U4932 ( .A1(sp_out[24]), .A2(n4449), .B1(r0[24]), .B2(n4448), 
        .ZN(n3982) );
  AOI22D1BWP12T U4933 ( .A1(r5[24]), .A2(n4453), .B1(r6[24]), .B2(n4451), .ZN(
        n3977) );
  AOI22D1BWP12T U4934 ( .A1(r7[24]), .A2(n3985), .B1(r4[24]), .B2(n3942), .ZN(
        n3976) );
  AOI22D1BWP12T U4935 ( .A1(r8[24]), .A2(n4452), .B1(r10[24]), .B2(n4217), 
        .ZN(n3975) );
  AOI22D1BWP12T U4936 ( .A1(r9[24]), .A2(n4218), .B1(r11[24]), .B2(n3953), 
        .ZN(n3974) );
  ND4D1BWP12T U4937 ( .A1(n3977), .A2(n3976), .A3(n3975), .A4(n3974), .ZN(
        n3980) );
  OAI22D1BWP12T U4938 ( .A1(n4576), .A2(n4458), .B1(n3978), .B2(n4206), .ZN(
        n3979) );
  AOI21D1BWP12T U4939 ( .A1(n4463), .A2(n3980), .B(n3979), .ZN(n3981) );
  ND4D1BWP12T U4940 ( .A1(n3984), .A2(n3983), .A3(n3982), .A4(n3981), .ZN(
        regD_out[24]) );
  AOI22D1BWP12T U4941 ( .A1(r6[23]), .A2(n4451), .B1(r11[23]), .B2(n3953), 
        .ZN(n3989) );
  AOI22D1BWP12T U4942 ( .A1(r9[23]), .A2(n4218), .B1(r4[23]), .B2(n3942), .ZN(
        n3988) );
  AOI22D1BWP12T U4943 ( .A1(r10[23]), .A2(n4217), .B1(r5[23]), .B2(n4453), 
        .ZN(n3987) );
  AOI22D1BWP12T U4944 ( .A1(r7[23]), .A2(n3985), .B1(r8[23]), .B2(n4452), .ZN(
        n3986) );
  ND4D1BWP12T U4945 ( .A1(n3989), .A2(n3988), .A3(n3987), .A4(n3986), .ZN(
        n3995) );
  AOI22D1BWP12T U4946 ( .A1(r1[23]), .A2(n4450), .B1(r3[23]), .B2(n4214), .ZN(
        n3993) );
  AOI22D1BWP12T U4947 ( .A1(sp_out[23]), .A2(n4449), .B1(lr[23]), .B2(n4447), 
        .ZN(n3992) );
  AOI22D1BWP12T U4948 ( .A1(r0[23]), .A2(n4448), .B1(r12[23]), .B2(n4215), 
        .ZN(n3991) );
  AOI22D1BWP12T U4949 ( .A1(r2[23]), .A2(n4216), .B1(pc_out[23]), .B2(n4195), 
        .ZN(n3990) );
  ND4D1BWP12T U4950 ( .A1(n3993), .A2(n3992), .A3(n3991), .A4(n3990), .ZN(
        n3994) );
  AO21D1BWP12T U4951 ( .A1(n4463), .A2(n3995), .B(n3994), .Z(regD_out[23]) );
  AOI22D1BWP12T U4952 ( .A1(r0[22]), .A2(n4448), .B1(r12[22]), .B2(n4215), 
        .ZN(n4006) );
  AOI22D1BWP12T U4953 ( .A1(lr[22]), .A2(n4447), .B1(r3[22]), .B2(n4214), .ZN(
        n4005) );
  AOI22D1BWP12T U4954 ( .A1(r1[22]), .A2(n4450), .B1(sp_out[22]), .B2(n4449), 
        .ZN(n4004) );
  AOI22D1BWP12T U4955 ( .A1(r5[22]), .A2(n4453), .B1(r11[22]), .B2(n3953), 
        .ZN(n3999) );
  AOI22D1BWP12T U4956 ( .A1(r4[22]), .A2(n3942), .B1(r10[22]), .B2(n4217), 
        .ZN(n3998) );
  AOI22D1BWP12T U4957 ( .A1(r9[22]), .A2(n4218), .B1(r8[22]), .B2(n4452), .ZN(
        n3997) );
  AOI22D1BWP12T U4958 ( .A1(r7[22]), .A2(n3985), .B1(r6[22]), .B2(n4451), .ZN(
        n3996) );
  ND4D1BWP12T U4959 ( .A1(n3999), .A2(n3998), .A3(n3997), .A4(n3996), .ZN(
        n4002) );
  OAI22D1BWP12T U4960 ( .A1(n4552), .A2(n4458), .B1(n4000), .B2(n4091), .ZN(
        n4001) );
  AOI21D1BWP12T U4961 ( .A1(n4463), .A2(n4002), .B(n4001), .ZN(n4003) );
  ND4D1BWP12T U4962 ( .A1(n4006), .A2(n4005), .A3(n4004), .A4(n4003), .ZN(
        regD_out[22]) );
  AOI22D1BWP12T U4963 ( .A1(r9[21]), .A2(n4218), .B1(r5[21]), .B2(n4453), .ZN(
        n4010) );
  AOI22D1BWP12T U4964 ( .A1(r11[21]), .A2(n3953), .B1(r7[21]), .B2(n3985), 
        .ZN(n4009) );
  AOI22D1BWP12T U4965 ( .A1(r6[21]), .A2(n4451), .B1(r4[21]), .B2(n3942), .ZN(
        n4008) );
  AOI22D1BWP12T U4966 ( .A1(r10[21]), .A2(n4217), .B1(r8[21]), .B2(n4452), 
        .ZN(n4007) );
  ND4D1BWP12T U4967 ( .A1(n4010), .A2(n4009), .A3(n4008), .A4(n4007), .ZN(
        n4016) );
  AOI22D1BWP12T U4968 ( .A1(sp_out[21]), .A2(n4449), .B1(r0[21]), .B2(n4448), 
        .ZN(n4014) );
  AOI22D1BWP12T U4969 ( .A1(r1[21]), .A2(n4450), .B1(r12[21]), .B2(n4215), 
        .ZN(n4013) );
  AOI22D1BWP12T U4970 ( .A1(r3[21]), .A2(n4214), .B1(r2[21]), .B2(n4216), .ZN(
        n4012) );
  AOI22D1BWP12T U4971 ( .A1(pc_out[21]), .A2(n4195), .B1(lr[21]), .B2(n4447), 
        .ZN(n4011) );
  ND4D1BWP12T U4972 ( .A1(n4014), .A2(n4013), .A3(n4012), .A4(n4011), .ZN(
        n4015) );
  AO21D1BWP12T U4973 ( .A1(n4463), .A2(n4016), .B(n4015), .Z(regD_out[21]) );
  AOI22D1BWP12T U4974 ( .A1(r9[20]), .A2(n4218), .B1(r6[20]), .B2(n4451), .ZN(
        n4020) );
  AOI22D1BWP12T U4975 ( .A1(r11[20]), .A2(n3953), .B1(r7[20]), .B2(n3985), 
        .ZN(n4019) );
  AOI22D1BWP12T U4976 ( .A1(r8[20]), .A2(n4452), .B1(r10[20]), .B2(n4217), 
        .ZN(n4018) );
  AOI22D1BWP12T U4977 ( .A1(r4[20]), .A2(n3942), .B1(r5[20]), .B2(n4453), .ZN(
        n4017) );
  ND4D1BWP12T U4978 ( .A1(n4020), .A2(n4019), .A3(n4018), .A4(n4017), .ZN(
        n4026) );
  AOI22D1BWP12T U4979 ( .A1(lr[20]), .A2(n4447), .B1(r1[20]), .B2(n4450), .ZN(
        n4024) );
  AOI22D1BWP12T U4980 ( .A1(r3[20]), .A2(n4214), .B1(r12[20]), .B2(n4215), 
        .ZN(n4023) );
  AOI22D1BWP12T U4981 ( .A1(r0[20]), .A2(n4448), .B1(r2[20]), .B2(n4216), .ZN(
        n4022) );
  AOI22D1BWP12T U4982 ( .A1(sp_out[20]), .A2(n4449), .B1(pc_out[20]), .B2(
        n4195), .ZN(n4021) );
  ND4D1BWP12T U4983 ( .A1(n4024), .A2(n4023), .A3(n4022), .A4(n4021), .ZN(
        n4025) );
  AO21D1BWP12T U4984 ( .A1(n4463), .A2(n4026), .B(n4025), .Z(regD_out[20]) );
  AOI22D1BWP12T U4985 ( .A1(r7[19]), .A2(n3985), .B1(r4[19]), .B2(n3942), .ZN(
        n4030) );
  AOI22D1BWP12T U4986 ( .A1(r5[19]), .A2(n4453), .B1(r8[19]), .B2(n4452), .ZN(
        n4029) );
  AOI22D1BWP12T U4987 ( .A1(r6[19]), .A2(n4451), .B1(r9[19]), .B2(n4218), .ZN(
        n4028) );
  AOI22D1BWP12T U4988 ( .A1(r11[19]), .A2(n3953), .B1(r10[19]), .B2(n4217), 
        .ZN(n4027) );
  ND4D1BWP12T U4989 ( .A1(n4030), .A2(n4029), .A3(n4028), .A4(n4027), .ZN(
        n4036) );
  AOI22D1BWP12T U4990 ( .A1(sp_out[19]), .A2(n4449), .B1(r2[19]), .B2(n4216), 
        .ZN(n4034) );
  AOI22D1BWP12T U4991 ( .A1(r0[19]), .A2(n4448), .B1(r1[19]), .B2(n4450), .ZN(
        n4033) );
  AOI22D1BWP12T U4992 ( .A1(r12[19]), .A2(n4215), .B1(lr[19]), .B2(n4447), 
        .ZN(n4032) );
  AOI22D1BWP12T U4993 ( .A1(pc_out[19]), .A2(n4195), .B1(r3[19]), .B2(n4214), 
        .ZN(n4031) );
  ND4D1BWP12T U4994 ( .A1(n4034), .A2(n4033), .A3(n4032), .A4(n4031), .ZN(
        n4035) );
  AO21D1BWP12T U4995 ( .A1(n4463), .A2(n4036), .B(n4035), .Z(regD_out[19]) );
  AOI22D1BWP12T U4996 ( .A1(r0[18]), .A2(n4448), .B1(sp_out[18]), .B2(n4449), 
        .ZN(n4046) );
  AOI22D1BWP12T U4997 ( .A1(r1[18]), .A2(n4450), .B1(r12[18]), .B2(n4215), 
        .ZN(n4045) );
  AOI22D1BWP12T U4998 ( .A1(r2[18]), .A2(n4216), .B1(r3[18]), .B2(n4214), .ZN(
        n4044) );
  AOI22D1BWP12T U4999 ( .A1(r4[18]), .A2(n3942), .B1(r8[18]), .B2(n4452), .ZN(
        n4040) );
  AOI22D1BWP12T U5000 ( .A1(r10[18]), .A2(n4217), .B1(r9[18]), .B2(n4218), 
        .ZN(n4039) );
  AOI22D1BWP12T U5001 ( .A1(r5[18]), .A2(n4453), .B1(r11[18]), .B2(n3953), 
        .ZN(n4038) );
  AOI22D1BWP12T U5002 ( .A1(r6[18]), .A2(n4451), .B1(r7[18]), .B2(n3985), .ZN(
        n4037) );
  ND4D1BWP12T U5003 ( .A1(n4040), .A2(n4039), .A3(n4038), .A4(n4037), .ZN(
        n4042) );
  MOAI22D0BWP12T U5004 ( .A1(n4504), .A2(n4184), .B1(pc_out[18]), .B2(n4195), 
        .ZN(n4041) );
  AOI21D1BWP12T U5005 ( .A1(n4463), .A2(n4042), .B(n4041), .ZN(n4043) );
  ND4D1BWP12T U5006 ( .A1(n4046), .A2(n4045), .A3(n4044), .A4(n4043), .ZN(
        regD_out[18]) );
  AOI22D1BWP12T U5007 ( .A1(r6[17]), .A2(n4451), .B1(r8[17]), .B2(n4452), .ZN(
        n4050) );
  AOI22D1BWP12T U5008 ( .A1(r5[17]), .A2(n4453), .B1(r11[17]), .B2(n3953), 
        .ZN(n4049) );
  AOI22D1BWP12T U5009 ( .A1(r4[17]), .A2(n3942), .B1(r9[17]), .B2(n4218), .ZN(
        n4048) );
  AOI22D1BWP12T U5010 ( .A1(r7[17]), .A2(n3985), .B1(r10[17]), .B2(n4217), 
        .ZN(n4047) );
  ND4D1BWP12T U5011 ( .A1(n4050), .A2(n4049), .A3(n4048), .A4(n4047), .ZN(
        n4056) );
  AOI22D1BWP12T U5012 ( .A1(r12[17]), .A2(n4215), .B1(pc_out[17]), .B2(n4195), 
        .ZN(n4054) );
  AOI22D1BWP12T U5013 ( .A1(lr[17]), .A2(n4447), .B1(sp_out[17]), .B2(n4449), 
        .ZN(n4053) );
  AOI22D1BWP12T U5014 ( .A1(r2[17]), .A2(n4216), .B1(r3[17]), .B2(n4214), .ZN(
        n4052) );
  AOI22D1BWP12T U5015 ( .A1(r1[17]), .A2(n4450), .B1(r0[17]), .B2(n4448), .ZN(
        n4051) );
  ND4D1BWP12T U5016 ( .A1(n4054), .A2(n4053), .A3(n4052), .A4(n4051), .ZN(
        n4055) );
  AO21D1BWP12T U5017 ( .A1(n4463), .A2(n4056), .B(n4055), .Z(regD_out[17]) );
  AOI22D1BWP12T U5018 ( .A1(r8[16]), .A2(n4452), .B1(r7[16]), .B2(n3985), .ZN(
        n4060) );
  AOI22D1BWP12T U5019 ( .A1(r11[16]), .A2(n3953), .B1(r9[16]), .B2(n4218), 
        .ZN(n4059) );
  AOI22D1BWP12T U5020 ( .A1(r10[16]), .A2(n4217), .B1(r4[16]), .B2(n3942), 
        .ZN(n4058) );
  AOI22D1BWP12T U5021 ( .A1(r5[16]), .A2(n4453), .B1(r6[16]), .B2(n4451), .ZN(
        n4057) );
  ND4D1BWP12T U5022 ( .A1(n4060), .A2(n4059), .A3(n4058), .A4(n4057), .ZN(
        n4066) );
  AOI22D1BWP12T U5023 ( .A1(lr[16]), .A2(n4447), .B1(r1[16]), .B2(n4450), .ZN(
        n4064) );
  AOI22D1BWP12T U5024 ( .A1(r12[16]), .A2(n4215), .B1(sp_out[16]), .B2(n4449), 
        .ZN(n4063) );
  AOI22D1BWP12T U5025 ( .A1(pc_out[16]), .A2(n4195), .B1(r2[16]), .B2(n4216), 
        .ZN(n4062) );
  AOI22D1BWP12T U5026 ( .A1(r3[16]), .A2(n4214), .B1(r0[16]), .B2(n4448), .ZN(
        n4061) );
  ND4D1BWP12T U5027 ( .A1(n4064), .A2(n4063), .A3(n4062), .A4(n4061), .ZN(
        n4065) );
  AO21D1BWP12T U5028 ( .A1(n4463), .A2(n4066), .B(n4065), .Z(regD_out[16]) );
  AOI22D1BWP12T U5029 ( .A1(r0[15]), .A2(n4448), .B1(lr[15]), .B2(n4447), .ZN(
        n4076) );
  AOI22D1BWP12T U5030 ( .A1(sp_out[15]), .A2(n4449), .B1(r3[15]), .B2(n4214), 
        .ZN(n4075) );
  AOI22D1BWP12T U5031 ( .A1(r1[15]), .A2(n4450), .B1(r2[15]), .B2(n4216), .ZN(
        n4074) );
  AOI22D1BWP12T U5032 ( .A1(r10[15]), .A2(n4217), .B1(r5[15]), .B2(n4453), 
        .ZN(n4070) );
  AOI22D1BWP12T U5033 ( .A1(r6[15]), .A2(n4451), .B1(r4[15]), .B2(n3942), .ZN(
        n4069) );
  AOI22D1BWP12T U5034 ( .A1(r8[15]), .A2(n4452), .B1(r11[15]), .B2(n3953), 
        .ZN(n4068) );
  AOI22D1BWP12T U5035 ( .A1(r9[15]), .A2(n4218), .B1(r7[15]), .B2(n3985), .ZN(
        n4067) );
  ND4D1BWP12T U5036 ( .A1(n4070), .A2(n4069), .A3(n4068), .A4(n4067), .ZN(
        n4072) );
  OAI22D1BWP12T U5037 ( .A1(n4830), .A2(n4460), .B1(n4886), .B2(n4458), .ZN(
        n4071) );
  AOI21D1BWP12T U5038 ( .A1(n4463), .A2(n4072), .B(n4071), .ZN(n4073) );
  ND4D1BWP12T U5039 ( .A1(n4076), .A2(n4075), .A3(n4074), .A4(n4073), .ZN(
        regD_out[15]) );
  AOI22D1BWP12T U5040 ( .A1(r6[14]), .A2(n4451), .B1(r10[14]), .B2(n4217), 
        .ZN(n4080) );
  AOI22D1BWP12T U5041 ( .A1(r4[14]), .A2(n3942), .B1(r7[14]), .B2(n3985), .ZN(
        n4079) );
  AOI22D1BWP12T U5042 ( .A1(r5[14]), .A2(n4453), .B1(r9[14]), .B2(n4218), .ZN(
        n4078) );
  AOI22D1BWP12T U5043 ( .A1(r11[14]), .A2(n3953), .B1(r8[14]), .B2(n4452), 
        .ZN(n4077) );
  ND4D1BWP12T U5044 ( .A1(n4080), .A2(n4079), .A3(n4078), .A4(n4077), .ZN(
        n4086) );
  AOI22D1BWP12T U5045 ( .A1(r1[14]), .A2(n4450), .B1(pc_out[14]), .B2(n4195), 
        .ZN(n4084) );
  AOI22D1BWP12T U5046 ( .A1(r12[14]), .A2(n4215), .B1(sp_out[14]), .B2(n4449), 
        .ZN(n4083) );
  AOI22D1BWP12T U5047 ( .A1(lr[14]), .A2(n4447), .B1(r2[14]), .B2(n4216), .ZN(
        n4082) );
  AOI22D1BWP12T U5048 ( .A1(r3[14]), .A2(n4214), .B1(r0[14]), .B2(n4448), .ZN(
        n4081) );
  ND4D1BWP12T U5049 ( .A1(n4084), .A2(n4083), .A3(n4082), .A4(n4081), .ZN(
        n4085) );
  AO21D1BWP12T U5050 ( .A1(n4463), .A2(n4086), .B(n4085), .Z(regD_out[14]) );
  AOI22D1BWP12T U5051 ( .A1(sp_out[13]), .A2(n4449), .B1(lr[13]), .B2(n4447), 
        .ZN(n4098) );
  AOI22D1BWP12T U5052 ( .A1(r12[13]), .A2(n4215), .B1(r0[13]), .B2(n4448), 
        .ZN(n4097) );
  AOI22D1BWP12T U5053 ( .A1(r3[13]), .A2(n4214), .B1(r1[13]), .B2(n4450), .ZN(
        n4096) );
  AOI22D1BWP12T U5054 ( .A1(r11[13]), .A2(n3953), .B1(r6[13]), .B2(n4451), 
        .ZN(n4090) );
  AOI22D1BWP12T U5055 ( .A1(r7[13]), .A2(n3985), .B1(r10[13]), .B2(n4217), 
        .ZN(n4089) );
  AOI22D1BWP12T U5056 ( .A1(r9[13]), .A2(n4218), .B1(r4[13]), .B2(n3942), .ZN(
        n4088) );
  AOI22D1BWP12T U5057 ( .A1(r8[13]), .A2(n4452), .B1(r5[13]), .B2(n4453), .ZN(
        n4087) );
  ND4D1BWP12T U5058 ( .A1(n4090), .A2(n4089), .A3(n4088), .A4(n4087), .ZN(
        n4094) );
  OAI22D1BWP12T U5059 ( .A1(n4092), .A2(n4091), .B1(n4436), .B2(n4458), .ZN(
        n4093) );
  AOI21D1BWP12T U5060 ( .A1(n4463), .A2(n4094), .B(n4093), .ZN(n4095) );
  ND4D1BWP12T U5061 ( .A1(n4098), .A2(n4097), .A3(n4096), .A4(n4095), .ZN(
        regD_out[13]) );
  AOI22D1BWP12T U5062 ( .A1(r11[12]), .A2(n3953), .B1(r7[12]), .B2(n3985), 
        .ZN(n4102) );
  AOI22D1BWP12T U5063 ( .A1(r4[12]), .A2(n3942), .B1(r10[12]), .B2(n4217), 
        .ZN(n4101) );
  AOI22D1BWP12T U5064 ( .A1(r5[12]), .A2(n4453), .B1(r9[12]), .B2(n4218), .ZN(
        n4100) );
  AOI22D1BWP12T U5065 ( .A1(r8[12]), .A2(n4452), .B1(r6[12]), .B2(n4451), .ZN(
        n4099) );
  ND4D1BWP12T U5066 ( .A1(n4102), .A2(n4101), .A3(n4100), .A4(n4099), .ZN(
        n4108) );
  AOI22D1BWP12T U5067 ( .A1(r3[12]), .A2(n4214), .B1(r1[12]), .B2(n4450), .ZN(
        n4106) );
  AOI22D1BWP12T U5068 ( .A1(sp_out[12]), .A2(n4449), .B1(lr[12]), .B2(n4447), 
        .ZN(n4105) );
  AOI22D1BWP12T U5069 ( .A1(r0[12]), .A2(n4448), .B1(r12[12]), .B2(n4215), 
        .ZN(n4104) );
  AOI22D1BWP12T U5070 ( .A1(r2[12]), .A2(n4216), .B1(pc_out[12]), .B2(n4195), 
        .ZN(n4103) );
  ND4D1BWP12T U5071 ( .A1(n4106), .A2(n4105), .A3(n4104), .A4(n4103), .ZN(
        n4107) );
  AO21D1BWP12T U5072 ( .A1(n4463), .A2(n4108), .B(n4107), .Z(regD_out[12]) );
  AOI22D1BWP12T U5073 ( .A1(r3[11]), .A2(n4214), .B1(r1[11]), .B2(n4450), .ZN(
        n4118) );
  AOI22D1BWP12T U5074 ( .A1(r0[11]), .A2(n4448), .B1(r2[11]), .B2(n4216), .ZN(
        n4117) );
  AOI22D1BWP12T U5075 ( .A1(r12[11]), .A2(n4215), .B1(sp_out[11]), .B2(n4449), 
        .ZN(n4116) );
  AOI22D1BWP12T U5076 ( .A1(r8[11]), .A2(n4452), .B1(r11[11]), .B2(n3953), 
        .ZN(n4112) );
  AOI22D1BWP12T U5077 ( .A1(r9[11]), .A2(n4218), .B1(r5[11]), .B2(n4453), .ZN(
        n4111) );
  AOI22D1BWP12T U5078 ( .A1(r6[11]), .A2(n4451), .B1(r4[11]), .B2(n3942), .ZN(
        n4110) );
  AOI22D1BWP12T U5079 ( .A1(r10[11]), .A2(n4217), .B1(r7[11]), .B2(n3985), 
        .ZN(n4109) );
  ND4D1BWP12T U5080 ( .A1(n4112), .A2(n4111), .A3(n4110), .A4(n4109), .ZN(
        n4114) );
  OAI22D1BWP12T U5081 ( .A1(n4412), .A2(n4458), .B1(n4870), .B2(n4184), .ZN(
        n4113) );
  AOI21D1BWP12T U5082 ( .A1(n4463), .A2(n4114), .B(n4113), .ZN(n4115) );
  ND4D1BWP12T U5083 ( .A1(n4118), .A2(n4117), .A3(n4116), .A4(n4115), .ZN(
        regD_out[11]) );
  AOI22D1BWP12T U5084 ( .A1(r10[10]), .A2(n4217), .B1(r6[10]), .B2(n4451), 
        .ZN(n4122) );
  AOI22D1BWP12T U5085 ( .A1(r11[10]), .A2(n3953), .B1(r8[10]), .B2(n4452), 
        .ZN(n4121) );
  AOI22D1BWP12T U5086 ( .A1(r5[10]), .A2(n4453), .B1(r7[10]), .B2(n3985), .ZN(
        n4120) );
  AOI22D1BWP12T U5087 ( .A1(r9[10]), .A2(n4218), .B1(r4[10]), .B2(n3942), .ZN(
        n4119) );
  ND4D1BWP12T U5088 ( .A1(n4122), .A2(n4121), .A3(n4120), .A4(n4119), .ZN(
        n4128) );
  AOI22D1BWP12T U5089 ( .A1(r0[10]), .A2(n4448), .B1(r1[10]), .B2(n4450), .ZN(
        n4126) );
  AOI22D1BWP12T U5090 ( .A1(r2[10]), .A2(n4216), .B1(lr[10]), .B2(n4447), .ZN(
        n4125) );
  AOI22D1BWP12T U5091 ( .A1(r3[10]), .A2(n4214), .B1(pc_out[10]), .B2(n4195), 
        .ZN(n4124) );
  AOI22D1BWP12T U5092 ( .A1(sp_out[10]), .A2(n4449), .B1(r12[10]), .B2(n4215), 
        .ZN(n4123) );
  ND4D1BWP12T U5093 ( .A1(n4126), .A2(n4125), .A3(n4124), .A4(n4123), .ZN(
        n4127) );
  AO21D1BWP12T U5094 ( .A1(n4463), .A2(n4128), .B(n4127), .Z(regD_out[10]) );
  AOI22D1BWP12T U5095 ( .A1(r7[9]), .A2(n3985), .B1(r10[9]), .B2(n4217), .ZN(
        n4132) );
  AOI22D1BWP12T U5096 ( .A1(r6[9]), .A2(n4451), .B1(r11[9]), .B2(n3953), .ZN(
        n4131) );
  AOI22D1BWP12T U5097 ( .A1(r9[9]), .A2(n4218), .B1(r5[9]), .B2(n4453), .ZN(
        n4130) );
  AOI22D1BWP12T U5098 ( .A1(r4[9]), .A2(n3942), .B1(r8[9]), .B2(n4452), .ZN(
        n4129) );
  ND4D1BWP12T U5099 ( .A1(n4132), .A2(n4131), .A3(n4130), .A4(n4129), .ZN(
        n4138) );
  AOI22D1BWP12T U5100 ( .A1(r12[9]), .A2(n4215), .B1(r3[9]), .B2(n4214), .ZN(
        n4136) );
  AOI22D1BWP12T U5101 ( .A1(sp_out[9]), .A2(n4449), .B1(r0[9]), .B2(n4448), 
        .ZN(n4135) );
  AOI22D1BWP12T U5102 ( .A1(r2[9]), .A2(n4216), .B1(lr[9]), .B2(n4447), .ZN(
        n4134) );
  AOI22D1BWP12T U5103 ( .A1(pc_out[9]), .A2(n4195), .B1(r1[9]), .B2(n4450), 
        .ZN(n4133) );
  ND4D1BWP12T U5104 ( .A1(n4136), .A2(n4135), .A3(n4134), .A4(n4133), .ZN(
        n4137) );
  AO21D1BWP12T U5105 ( .A1(n4463), .A2(n4138), .B(n4137), .Z(regD_out[9]) );
  AOI22D1BWP12T U5106 ( .A1(r6[8]), .A2(n4451), .B1(r10[8]), .B2(n4217), .ZN(
        n4142) );
  AOI22D1BWP12T U5107 ( .A1(r8[8]), .A2(n4452), .B1(r7[8]), .B2(n3985), .ZN(
        n4141) );
  AOI22D1BWP12T U5108 ( .A1(r11[8]), .A2(n3953), .B1(r9[8]), .B2(n4218), .ZN(
        n4140) );
  AOI22D1BWP12T U5109 ( .A1(r5[8]), .A2(n4453), .B1(r4[8]), .B2(n3942), .ZN(
        n4139) );
  ND4D1BWP12T U5110 ( .A1(n4142), .A2(n4141), .A3(n4140), .A4(n4139), .ZN(
        n4148) );
  AOI22D1BWP12T U5111 ( .A1(pc_out[8]), .A2(n4195), .B1(sp_out[8]), .B2(n4449), 
        .ZN(n4146) );
  AOI22D1BWP12T U5112 ( .A1(r0[8]), .A2(n4448), .B1(r1[8]), .B2(n4450), .ZN(
        n4145) );
  AOI22D1BWP12T U5113 ( .A1(r2[8]), .A2(n4216), .B1(r12[8]), .B2(n4215), .ZN(
        n4144) );
  AOI22D1BWP12T U5114 ( .A1(lr[8]), .A2(n4447), .B1(r3[8]), .B2(n4214), .ZN(
        n4143) );
  ND4D1BWP12T U5115 ( .A1(n4146), .A2(n4145), .A3(n4144), .A4(n4143), .ZN(
        n4147) );
  AO21D1BWP12T U5116 ( .A1(n4463), .A2(n4148), .B(n4147), .Z(regD_out[8]) );
  AOI22D1BWP12T U5117 ( .A1(r5[7]), .A2(n4453), .B1(r11[7]), .B2(n3953), .ZN(
        n4152) );
  AOI22D1BWP12T U5118 ( .A1(r7[7]), .A2(n3985), .B1(r10[7]), .B2(n4217), .ZN(
        n4151) );
  AOI22D1BWP12T U5119 ( .A1(r4[7]), .A2(n3942), .B1(r8[7]), .B2(n4452), .ZN(
        n4150) );
  AOI22D1BWP12T U5120 ( .A1(r9[7]), .A2(n4218), .B1(r6[7]), .B2(n4451), .ZN(
        n4149) );
  ND4D1BWP12T U5121 ( .A1(n4152), .A2(n4151), .A3(n4150), .A4(n4149), .ZN(
        n4158) );
  AOI22D1BWP12T U5122 ( .A1(sp_out[7]), .A2(n4449), .B1(r3[7]), .B2(n4214), 
        .ZN(n4156) );
  AOI22D1BWP12T U5123 ( .A1(r1[7]), .A2(n4450), .B1(lr[7]), .B2(n4447), .ZN(
        n4155) );
  AOI22D1BWP12T U5124 ( .A1(pc_out[7]), .A2(n4195), .B1(r2[7]), .B2(n4216), 
        .ZN(n4154) );
  AOI22D1BWP12T U5125 ( .A1(r12[7]), .A2(n4215), .B1(r0[7]), .B2(n4448), .ZN(
        n4153) );
  ND4D1BWP12T U5126 ( .A1(n4156), .A2(n4155), .A3(n4154), .A4(n4153), .ZN(
        n4157) );
  AO21D1BWP12T U5127 ( .A1(n4463), .A2(n4158), .B(n4157), .Z(regD_out[7]) );
  AOI22D1BWP12T U5128 ( .A1(r0[6]), .A2(n4448), .B1(r1[6]), .B2(n4450), .ZN(
        n4169) );
  AOI22D1BWP12T U5129 ( .A1(lr[6]), .A2(n4447), .B1(r3[6]), .B2(n4214), .ZN(
        n4168) );
  AOI22D1BWP12T U5130 ( .A1(r2[6]), .A2(n4216), .B1(sp_out[6]), .B2(n4449), 
        .ZN(n4167) );
  AOI22D1BWP12T U5131 ( .A1(r4[6]), .A2(n3942), .B1(r8[6]), .B2(n4452), .ZN(
        n4162) );
  AOI22D1BWP12T U5132 ( .A1(r7[6]), .A2(n3985), .B1(r11[6]), .B2(n3953), .ZN(
        n4161) );
  AOI22D1BWP12T U5133 ( .A1(r9[6]), .A2(n4218), .B1(r5[6]), .B2(n4453), .ZN(
        n4160) );
  AOI22D1BWP12T U5134 ( .A1(r10[6]), .A2(n4217), .B1(r6[6]), .B2(n4451), .ZN(
        n4159) );
  ND4D1BWP12T U5135 ( .A1(n4162), .A2(n4161), .A3(n4160), .A4(n4159), .ZN(
        n4165) );
  OAI22D1BWP12T U5136 ( .A1(n4163), .A2(n4460), .B1(n4353), .B2(n4458), .ZN(
        n4164) );
  AOI21D1BWP12T U5137 ( .A1(n4463), .A2(n4165), .B(n4164), .ZN(n4166) );
  ND4D1BWP12T U5138 ( .A1(n4169), .A2(n4168), .A3(n4167), .A4(n4166), .ZN(
        regD_out[6]) );
  AOI22D1BWP12T U5139 ( .A1(r6[5]), .A2(n4451), .B1(r9[5]), .B2(n4218), .ZN(
        n4173) );
  AOI22D1BWP12T U5140 ( .A1(r8[5]), .A2(n4452), .B1(r7[5]), .B2(n3985), .ZN(
        n4172) );
  AOI22D1BWP12T U5141 ( .A1(r11[5]), .A2(n3953), .B1(r5[5]), .B2(n4453), .ZN(
        n4171) );
  AOI22D1BWP12T U5142 ( .A1(r10[5]), .A2(n4217), .B1(r4[5]), .B2(n3942), .ZN(
        n4170) );
  ND4D1BWP12T U5143 ( .A1(n4173), .A2(n4172), .A3(n4171), .A4(n4170), .ZN(
        n4179) );
  AOI22D1BWP12T U5144 ( .A1(r1[5]), .A2(n4450), .B1(r2[5]), .B2(n4216), .ZN(
        n4177) );
  AOI22D1BWP12T U5145 ( .A1(r0[5]), .A2(n4448), .B1(r3[5]), .B2(n4214), .ZN(
        n4176) );
  AOI22D1BWP12T U5146 ( .A1(pc_out[5]), .A2(n4195), .B1(lr[5]), .B2(n4447), 
        .ZN(n4175) );
  AOI22D1BWP12T U5147 ( .A1(r12[5]), .A2(n4215), .B1(sp_out[5]), .B2(n4449), 
        .ZN(n4174) );
  ND4D1BWP12T U5148 ( .A1(n4177), .A2(n4176), .A3(n4175), .A4(n4174), .ZN(
        n4178) );
  AO21D1BWP12T U5149 ( .A1(n4463), .A2(n4179), .B(n4178), .Z(regD_out[5]) );
  AOI22D1BWP12T U5150 ( .A1(r1[4]), .A2(n4450), .B1(r3[4]), .B2(n4214), .ZN(
        n4190) );
  AOI22D1BWP12T U5151 ( .A1(sp_out[4]), .A2(n4449), .B1(r2[4]), .B2(n4216), 
        .ZN(n4189) );
  AOI22D1BWP12T U5152 ( .A1(r12[4]), .A2(n4215), .B1(r0[4]), .B2(n4448), .ZN(
        n4188) );
  AOI22D1BWP12T U5153 ( .A1(r7[4]), .A2(n3985), .B1(r10[4]), .B2(n4217), .ZN(
        n4183) );
  AOI22D1BWP12T U5154 ( .A1(r4[4]), .A2(n3942), .B1(r5[4]), .B2(n4453), .ZN(
        n4182) );
  AOI22D1BWP12T U5155 ( .A1(r9[4]), .A2(n4218), .B1(r8[4]), .B2(n4452), .ZN(
        n4181) );
  AOI22D1BWP12T U5156 ( .A1(r6[4]), .A2(n4451), .B1(r11[4]), .B2(n3953), .ZN(
        n4180) );
  ND4D1BWP12T U5157 ( .A1(n4183), .A2(n4182), .A3(n4181), .A4(n4180), .ZN(
        n4186) );
  MOAI22D0BWP12T U5158 ( .A1(n4330), .A2(n4184), .B1(pc_out[4]), .B2(n4195), 
        .ZN(n4185) );
  AOI21D1BWP12T U5159 ( .A1(n4463), .A2(n4186), .B(n4185), .ZN(n4187) );
  ND4D1BWP12T U5160 ( .A1(n4190), .A2(n4189), .A3(n4188), .A4(n4187), .ZN(
        regD_out[4]) );
  AOI22D1BWP12T U5161 ( .A1(r7[3]), .A2(n3985), .B1(r10[3]), .B2(n4217), .ZN(
        n4194) );
  AOI22D1BWP12T U5162 ( .A1(r4[3]), .A2(n3942), .B1(r8[3]), .B2(n4452), .ZN(
        n4193) );
  AOI22D1BWP12T U5163 ( .A1(r5[3]), .A2(n4453), .B1(r9[3]), .B2(n4218), .ZN(
        n4192) );
  AOI22D1BWP12T U5164 ( .A1(r6[3]), .A2(n4451), .B1(r11[3]), .B2(n3953), .ZN(
        n4191) );
  ND4D1BWP12T U5165 ( .A1(n4194), .A2(n4193), .A3(n4192), .A4(n4191), .ZN(
        n4201) );
  AOI22D1BWP12T U5166 ( .A1(r12[3]), .A2(n4215), .B1(sp_out[3]), .B2(n4449), 
        .ZN(n4199) );
  AOI22D1BWP12T U5167 ( .A1(lr[3]), .A2(n4447), .B1(r1[3]), .B2(n4450), .ZN(
        n4198) );
  AOI22D1BWP12T U5168 ( .A1(r2[3]), .A2(n4216), .B1(pc_out[3]), .B2(n4195), 
        .ZN(n4197) );
  AOI22D1BWP12T U5169 ( .A1(r3[3]), .A2(n4214), .B1(r0[3]), .B2(n4448), .ZN(
        n4196) );
  ND4D1BWP12T U5170 ( .A1(n4199), .A2(n4198), .A3(n4197), .A4(n4196), .ZN(
        n4200) );
  AO21D1BWP12T U5171 ( .A1(n4463), .A2(n4201), .B(n4200), .Z(regD_out[3]) );
  AOI22D1BWP12T U5172 ( .A1(r0[2]), .A2(n4448), .B1(r1[2]), .B2(n4450), .ZN(
        n4213) );
  AOI22D1BWP12T U5173 ( .A1(sp_out[2]), .A2(n4449), .B1(lr[2]), .B2(n4447), 
        .ZN(n4212) );
  AOI22D1BWP12T U5174 ( .A1(r2[2]), .A2(n4216), .B1(r12[2]), .B2(n4215), .ZN(
        n4211) );
  AOI22D1BWP12T U5175 ( .A1(r8[2]), .A2(n4452), .B1(r11[2]), .B2(n3953), .ZN(
        n4205) );
  AOI22D1BWP12T U5176 ( .A1(r10[2]), .A2(n4217), .B1(r7[2]), .B2(n3985), .ZN(
        n4204) );
  AOI22D1BWP12T U5177 ( .A1(r9[2]), .A2(n4218), .B1(r4[2]), .B2(n3942), .ZN(
        n4203) );
  AOI22D1BWP12T U5178 ( .A1(r6[2]), .A2(n4451), .B1(r5[2]), .B2(n4453), .ZN(
        n4202) );
  ND4D1BWP12T U5179 ( .A1(n4205), .A2(n4204), .A3(n4203), .A4(n4202), .ZN(
        n4209) );
  OAI22D1BWP12T U5180 ( .A1(n4207), .A2(n4206), .B1(n4305), .B2(n4458), .ZN(
        n4208) );
  AOI21D1BWP12T U5181 ( .A1(n4463), .A2(n4209), .B(n4208), .ZN(n4210) );
  ND4D1BWP12T U5182 ( .A1(n4213), .A2(n4212), .A3(n4211), .A4(n4210), .ZN(
        regD_out[2]) );
  AOI22D1BWP12T U5183 ( .A1(r12[1]), .A2(n4215), .B1(r3[1]), .B2(n4214), .ZN(
        n4228) );
  AOI22D1BWP12T U5184 ( .A1(lr[1]), .A2(n4447), .B1(r2[1]), .B2(n4216), .ZN(
        n4227) );
  AOI22D1BWP12T U5185 ( .A1(r1[1]), .A2(n4450), .B1(r0[1]), .B2(n4448), .ZN(
        n4226) );
  AOI22D1BWP12T U5186 ( .A1(r5[1]), .A2(n4453), .B1(r8[1]), .B2(n4452), .ZN(
        n4222) );
  AOI22D1BWP12T U5187 ( .A1(r7[1]), .A2(n3985), .B1(r4[1]), .B2(n3942), .ZN(
        n4221) );
  AOI22D1BWP12T U5188 ( .A1(r11[1]), .A2(n3953), .B1(r10[1]), .B2(n4217), .ZN(
        n4220) );
  AOI22D1BWP12T U5189 ( .A1(r6[1]), .A2(n4451), .B1(r9[1]), .B2(n4218), .ZN(
        n4219) );
  ND4D1BWP12T U5190 ( .A1(n4222), .A2(n4221), .A3(n4220), .A4(n4219), .ZN(
        n4224) );
  MOAI22D0BWP12T U5191 ( .A1(n4293), .A2(n4458), .B1(sp_out[1]), .B2(n4449), 
        .ZN(n4223) );
  AOI21D1BWP12T U5192 ( .A1(n4463), .A2(n4224), .B(n4223), .ZN(n4225) );
  ND4D1BWP12T U5193 ( .A1(n4228), .A2(n4227), .A3(n4226), .A4(n4225), .ZN(
        regD_out[1]) );
  AOI22D1BWP12T U5194 ( .A1(n4229), .A2(r0[30]), .B1(n4254), .B2(tmp1[30]), 
        .ZN(n4241) );
  AOI22D1BWP12T U5195 ( .A1(n4264), .A2(r8[30]), .B1(n3462), .B2(r3[30]), .ZN(
        n4240) );
  AOI22D1BWP12T U5196 ( .A1(n4257), .A2(r10[30]), .B1(n4230), .B2(r6[30]), 
        .ZN(n4239) );
  INVD1BWP12T U5197 ( .I(pc_out[30]), .ZN(n4642) );
  AOI22D1BWP12T U5198 ( .A1(n4266), .A2(sp_out[30]), .B1(n4259), .B2(r7[30]), 
        .ZN(n4231) );
  OAI21D1BWP12T U5199 ( .A1(n4263), .A2(n4642), .B(n4231), .ZN(n4237) );
  AOI22D1BWP12T U5200 ( .A1(n4260), .A2(r9[30]), .B1(n4265), .B2(r4[30]), .ZN(
        n4235) );
  AOI22D1BWP12T U5201 ( .A1(n4255), .A2(r1[30]), .B1(n4256), .B2(r5[30]), .ZN(
        n4234) );
  AOI22D1BWP12T U5202 ( .A1(n4258), .A2(r12[30]), .B1(n4267), .B2(lr[30]), 
        .ZN(n4233) );
  AOI22D1BWP12T U5203 ( .A1(n4269), .A2(immediate2_in[30]), .B1(n4268), .B2(
        r2[30]), .ZN(n4232) );
  ND4D1BWP12T U5204 ( .A1(n4235), .A2(n4234), .A3(n4233), .A4(n4232), .ZN(
        n4236) );
  AOI211D1BWP12T U5205 ( .A1(n4276), .A2(r11[30]), .B(n4237), .C(n4236), .ZN(
        n4238) );
  ND4D1BWP12T U5206 ( .A1(n4241), .A2(n4240), .A3(n4239), .A4(n4238), .ZN(
        regB_out[30]) );
  AOI22D1BWP12T U5207 ( .A1(r6[14]), .A2(n4667), .B1(n3186), .B2(
        immediate1_in[14]), .ZN(n4253) );
  AOI22D1BWP12T U5208 ( .A1(r5[14]), .A2(n4664), .B1(r11[14]), .B2(n4659), 
        .ZN(n4252) );
  AOI22D1BWP12T U5209 ( .A1(r4[14]), .A2(n4663), .B1(r9[14]), .B2(n4666), .ZN(
        n4251) );
  AOI22D1BWP12T U5210 ( .A1(r1[14]), .A2(n4615), .B1(r7[14]), .B2(n4656), .ZN(
        n4242) );
  OAI21D1BWP12T U5211 ( .A1(n4243), .A2(n4601), .B(n4242), .ZN(n4249) );
  AOI22D1BWP12T U5212 ( .A1(r12[14]), .A2(n4654), .B1(pc_out[14]), .B2(n4658), 
        .ZN(n4247) );
  AOI22D1BWP12T U5213 ( .A1(tmp1[14]), .A2(n4657), .B1(r10[14]), .B2(n4665), 
        .ZN(n4246) );
  AOI22D1BWP12T U5214 ( .A1(sp_out[14]), .A2(n4655), .B1(r8[14]), .B2(n4627), 
        .ZN(n4245) );
  AOI22D1BWP12T U5215 ( .A1(r2[14]), .A2(n4674), .B1(r0[14]), .B2(n4626), .ZN(
        n4244) );
  ND4D1BWP12T U5216 ( .A1(n4247), .A2(n4246), .A3(n4245), .A4(n4244), .ZN(
        n4248) );
  AOI211D1BWP12T U5217 ( .A1(r3[14]), .A2(n4589), .B(n4249), .C(n4248), .ZN(
        n4250) );
  ND4D1BWP12T U5218 ( .A1(n4253), .A2(n4252), .A3(n4251), .A4(n4250), .ZN(
        regA_out[14]) );
  AOI22D1BWP12T U5219 ( .A1(n4255), .A2(r1[31]), .B1(n4254), .B2(tmp1[31]), 
        .ZN(n4280) );
  AOI22D1BWP12T U5220 ( .A1(n4256), .A2(r5[31]), .B1(n4230), .B2(r6[31]), .ZN(
        n4279) );
  AOI22D1BWP12T U5221 ( .A1(n4258), .A2(r12[31]), .B1(n4257), .B2(r10[31]), 
        .ZN(n4278) );
  AOI22D1BWP12T U5222 ( .A1(n4260), .A2(r9[31]), .B1(n4259), .B2(r7[31]), .ZN(
        n4261) );
  OAI21D1BWP12T U5223 ( .A1(n4263), .A2(n4262), .B(n4261), .ZN(n4275) );
  AOI22D1BWP12T U5224 ( .A1(n4264), .A2(r8[31]), .B1(n3462), .B2(r3[31]), .ZN(
        n4273) );
  AOI22D1BWP12T U5225 ( .A1(n4266), .A2(sp_out[31]), .B1(n4265), .B2(r4[31]), 
        .ZN(n4272) );
  AOI22D1BWP12T U5226 ( .A1(n4229), .A2(r0[31]), .B1(n4267), .B2(lr[31]), .ZN(
        n4271) );
  AOI22D1BWP12T U5227 ( .A1(n4269), .A2(immediate2_in[31]), .B1(n4268), .B2(
        r2[31]), .ZN(n4270) );
  ND4D1BWP12T U5228 ( .A1(n4273), .A2(n4272), .A3(n4271), .A4(n4270), .ZN(
        n4274) );
  AOI211D1BWP12T U5229 ( .A1(n4276), .A2(r11[31]), .B(n4275), .C(n4274), .ZN(
        n4277) );
  ND4D1BWP12T U5230 ( .A1(n4280), .A2(n4279), .A3(n4278), .A4(n4277), .ZN(
        regB_out[31]) );
  AOI22D1BWP12T U5231 ( .A1(lr[0]), .A2(n4653), .B1(n3186), .B2(
        immediate1_in[0]), .ZN(n4291) );
  AOI22D1BWP12T U5232 ( .A1(r11[0]), .A2(n4659), .B1(r3[0]), .B2(n4589), .ZN(
        n4290) );
  AOI22D1BWP12T U5233 ( .A1(r0[0]), .A2(n4626), .B1(tmp1[0]), .B2(n4657), .ZN(
        n4289) );
  AOI22D1BWP12T U5234 ( .A1(sp_out[0]), .A2(n4655), .B1(r7[0]), .B2(n4656), 
        .ZN(n4281) );
  OAI21D1BWP12T U5235 ( .A1(n4459), .A2(n4641), .B(n4281), .ZN(n4287) );
  AOI22D1BWP12T U5236 ( .A1(r1[0]), .A2(n4615), .B1(r5[0]), .B2(n4664), .ZN(
        n4285) );
  AOI22D1BWP12T U5237 ( .A1(r9[0]), .A2(n4666), .B1(r10[0]), .B2(n4665), .ZN(
        n4284) );
  AOI22D1BWP12T U5238 ( .A1(r2[0]), .A2(n4674), .B1(r6[0]), .B2(n4667), .ZN(
        n4283) );
  INVD1BWP12T U5239 ( .I(n4627), .ZN(n4662) );
  AOI22D1BWP12T U5240 ( .A1(r4[0]), .A2(n4663), .B1(r8[0]), .B2(n4627), .ZN(
        n4282) );
  ND4D1BWP12T U5241 ( .A1(n4285), .A2(n4284), .A3(n4283), .A4(n4282), .ZN(
        n4286) );
  AOI211D1BWP12T U5242 ( .A1(r12[0]), .A2(n4654), .B(n4287), .C(n4286), .ZN(
        n4288) );
  ND4D1BWP12T U5243 ( .A1(n4291), .A2(n4290), .A3(n4289), .A4(n4288), .ZN(
        regA_out[0]) );
  AOI22D1BWP12T U5244 ( .A1(r8[1]), .A2(n4627), .B1(n3186), .B2(
        immediate1_in[1]), .ZN(n4303) );
  AOI22D1BWP12T U5245 ( .A1(r4[1]), .A2(n4663), .B1(tmp1[1]), .B2(n4657), .ZN(
        n4302) );
  AOI22D1BWP12T U5246 ( .A1(r9[1]), .A2(n4666), .B1(lr[1]), .B2(n4653), .ZN(
        n4301) );
  AOI22D1BWP12T U5247 ( .A1(r3[1]), .A2(n4589), .B1(r2[1]), .B2(n4674), .ZN(
        n4292) );
  OAI21D1BWP12T U5248 ( .A1(n4293), .A2(n4641), .B(n4292), .ZN(n4299) );
  AOI22D1BWP12T U5249 ( .A1(r1[1]), .A2(n4615), .B1(r0[1]), .B2(n4626), .ZN(
        n4297) );
  AOI22D1BWP12T U5250 ( .A1(r7[1]), .A2(n4656), .B1(r10[1]), .B2(n4665), .ZN(
        n4296) );
  AOI22D1BWP12T U5251 ( .A1(sp_out[1]), .A2(n4655), .B1(r5[1]), .B2(n4664), 
        .ZN(n4295) );
  AOI22D1BWP12T U5252 ( .A1(r6[1]), .A2(n4667), .B1(r11[1]), .B2(n4659), .ZN(
        n4294) );
  ND4D1BWP12T U5253 ( .A1(n4297), .A2(n4296), .A3(n4295), .A4(n4294), .ZN(
        n4298) );
  AOI211D1BWP12T U5254 ( .A1(r12[1]), .A2(n4654), .B(n4299), .C(n4298), .ZN(
        n4300) );
  ND4D1BWP12T U5255 ( .A1(n4303), .A2(n4302), .A3(n4301), .A4(n4300), .ZN(
        regA_out[1]) );
  AOI22D1BWP12T U5256 ( .A1(r2[2]), .A2(n4674), .B1(lr[2]), .B2(n4653), .ZN(
        n4315) );
  AOI22D1BWP12T U5257 ( .A1(r6[2]), .A2(n4667), .B1(r5[2]), .B2(n4664), .ZN(
        n4314) );
  AOI22D1BWP12T U5258 ( .A1(r8[2]), .A2(n4627), .B1(r9[2]), .B2(n4666), .ZN(
        n4313) );
  AOI22D1BWP12T U5259 ( .A1(r12[2]), .A2(n4654), .B1(r7[2]), .B2(n4656), .ZN(
        n4304) );
  OAI21D1BWP12T U5260 ( .A1(n4305), .A2(n4641), .B(n4304), .ZN(n4311) );
  AOI22D1BWP12T U5261 ( .A1(r11[2]), .A2(n4659), .B1(r1[2]), .B2(n4615), .ZN(
        n4309) );
  AOI22D1BWP12T U5262 ( .A1(tmp1[2]), .A2(n4657), .B1(r4[2]), .B2(n4663), .ZN(
        n4308) );
  AOI22D1BWP12T U5263 ( .A1(r10[2]), .A2(n4665), .B1(r0[2]), .B2(n4626), .ZN(
        n4307) );
  AOI22D1BWP12T U5264 ( .A1(r3[2]), .A2(n4589), .B1(n3186), .B2(
        immediate1_in[2]), .ZN(n4306) );
  ND4D1BWP12T U5265 ( .A1(n4309), .A2(n4308), .A3(n4307), .A4(n4306), .ZN(
        n4310) );
  AOI211D1BWP12T U5266 ( .A1(sp_out[2]), .A2(n4655), .B(n4311), .C(n4310), 
        .ZN(n4312) );
  ND4D1BWP12T U5267 ( .A1(n4315), .A2(n4314), .A3(n4313), .A4(n4312), .ZN(
        regA_out[2]) );
  AOI22D1BWP12T U5268 ( .A1(r5[3]), .A2(n4664), .B1(r8[3]), .B2(n4627), .ZN(
        n4327) );
  AOI22D1BWP12T U5269 ( .A1(r6[3]), .A2(n4667), .B1(r1[3]), .B2(n4615), .ZN(
        n4326) );
  AOI22D1BWP12T U5270 ( .A1(r12[3]), .A2(n4654), .B1(tmp1[3]), .B2(n4657), 
        .ZN(n4325) );
  AOI22D1BWP12T U5271 ( .A1(r7[3]), .A2(n4656), .B1(r4[3]), .B2(n4663), .ZN(
        n4316) );
  OAI21D1BWP12T U5272 ( .A1(n4317), .A2(n4641), .B(n4316), .ZN(n4323) );
  AOI22D1BWP12T U5273 ( .A1(r0[3]), .A2(n4626), .B1(r11[3]), .B2(n4659), .ZN(
        n4321) );
  AOI22D1BWP12T U5274 ( .A1(r10[3]), .A2(n4665), .B1(r9[3]), .B2(n4666), .ZN(
        n4320) );
  AOI22D1BWP12T U5275 ( .A1(lr[3]), .A2(n4653), .B1(r2[3]), .B2(n4674), .ZN(
        n4319) );
  AOI22D1BWP12T U5276 ( .A1(sp_out[3]), .A2(n4655), .B1(n3186), .B2(
        immediate1_in[3]), .ZN(n4318) );
  ND4D1BWP12T U5277 ( .A1(n4321), .A2(n4320), .A3(n4319), .A4(n4318), .ZN(
        n4322) );
  AOI211D1BWP12T U5278 ( .A1(r3[3]), .A2(n4589), .B(n4323), .C(n4322), .ZN(
        n4324) );
  ND4D1BWP12T U5279 ( .A1(n4327), .A2(n4326), .A3(n4325), .A4(n4324), .ZN(
        regA_out[3]) );
  AOI22D1BWP12T U5280 ( .A1(r6[4]), .A2(n4667), .B1(r8[4]), .B2(n4627), .ZN(
        n4339) );
  AOI22D1BWP12T U5281 ( .A1(r12[4]), .A2(n4654), .B1(r3[4]), .B2(n4589), .ZN(
        n4338) );
  AOI22D1BWP12T U5282 ( .A1(r1[4]), .A2(n4615), .B1(tmp1[4]), .B2(n4657), .ZN(
        n4329) );
  AOI22D1BWP12T U5283 ( .A1(r0[4]), .A2(n4626), .B1(r5[4]), .B2(n4664), .ZN(
        n4328) );
  OAI211D1BWP12T U5284 ( .A1(n4330), .A2(n4601), .B(n4329), .C(n4328), .ZN(
        n4336) );
  AOI22D1BWP12T U5285 ( .A1(r11[4]), .A2(n4659), .B1(pc_out[4]), .B2(n4658), 
        .ZN(n4334) );
  AOI22D1BWP12T U5286 ( .A1(r2[4]), .A2(n4674), .B1(n3186), .B2(
        immediate1_in[4]), .ZN(n4333) );
  AOI22D1BWP12T U5287 ( .A1(r4[4]), .A2(n4663), .B1(r10[4]), .B2(n4665), .ZN(
        n4332) );
  AOI22D1BWP12T U5288 ( .A1(r9[4]), .A2(n4666), .B1(sp_out[4]), .B2(n4655), 
        .ZN(n4331) );
  ND4D1BWP12T U5289 ( .A1(n4334), .A2(n4333), .A3(n4332), .A4(n4331), .ZN(
        n4335) );
  AOI211D1BWP12T U5290 ( .A1(r7[4]), .A2(n4656), .B(n4336), .C(n4335), .ZN(
        n4337) );
  ND3D1BWP12T U5291 ( .A1(n4339), .A2(n4338), .A3(n4337), .ZN(regA_out[4]) );
  AOI22D1BWP12T U5292 ( .A1(r11[5]), .A2(n4659), .B1(r5[5]), .B2(n4664), .ZN(
        n4351) );
  AOI22D1BWP12T U5293 ( .A1(r0[5]), .A2(n4626), .B1(r3[5]), .B2(n4589), .ZN(
        n4350) );
  AOI22D1BWP12T U5294 ( .A1(r7[5]), .A2(n4656), .B1(sp_out[5]), .B2(n4655), 
        .ZN(n4349) );
  AOI22D1BWP12T U5295 ( .A1(r4[5]), .A2(n4663), .B1(r2[5]), .B2(n4674), .ZN(
        n4340) );
  OAI21D1BWP12T U5296 ( .A1(n4341), .A2(n4641), .B(n4340), .ZN(n4347) );
  AOI22D1BWP12T U5297 ( .A1(r10[5]), .A2(n4665), .B1(r1[5]), .B2(n4615), .ZN(
        n4345) );
  AOI22D1BWP12T U5298 ( .A1(lr[5]), .A2(n4653), .B1(tmp1[5]), .B2(n4657), .ZN(
        n4344) );
  AOI22D1BWP12T U5299 ( .A1(r8[5]), .A2(n4627), .B1(n3186), .B2(
        immediate1_in[5]), .ZN(n4343) );
  AOI22D1BWP12T U5300 ( .A1(r12[5]), .A2(n4654), .B1(r9[5]), .B2(n4666), .ZN(
        n4342) );
  ND4D1BWP12T U5301 ( .A1(n4345), .A2(n4344), .A3(n4343), .A4(n4342), .ZN(
        n4346) );
  AOI211D1BWP12T U5302 ( .A1(r6[5]), .A2(n4667), .B(n4347), .C(n4346), .ZN(
        n4348) );
  ND4D1BWP12T U5303 ( .A1(n4351), .A2(n4350), .A3(n4349), .A4(n4348), .ZN(
        regA_out[5]) );
  AOI22D1BWP12T U5304 ( .A1(sp_out[6]), .A2(n4655), .B1(r11[6]), .B2(n4659), 
        .ZN(n4363) );
  AOI22D1BWP12T U5305 ( .A1(r12[6]), .A2(n4654), .B1(r10[6]), .B2(n4665), .ZN(
        n4362) );
  AOI22D1BWP12T U5306 ( .A1(r8[6]), .A2(n4627), .B1(r7[6]), .B2(n4656), .ZN(
        n4361) );
  AOI22D1BWP12T U5307 ( .A1(r5[6]), .A2(n4664), .B1(n3186), .B2(
        immediate1_in[6]), .ZN(n4352) );
  OAI21D1BWP12T U5308 ( .A1(n4353), .A2(n4641), .B(n4352), .ZN(n4359) );
  AOI22D1BWP12T U5309 ( .A1(r4[6]), .A2(n4663), .B1(r6[6]), .B2(n4667), .ZN(
        n4357) );
  AOI22D1BWP12T U5310 ( .A1(lr[6]), .A2(n4653), .B1(r2[6]), .B2(n4674), .ZN(
        n4356) );
  AOI22D1BWP12T U5311 ( .A1(r9[6]), .A2(n4666), .B1(r1[6]), .B2(n4615), .ZN(
        n4355) );
  AOI22D1BWP12T U5312 ( .A1(r3[6]), .A2(n4589), .B1(tmp1[6]), .B2(n4657), .ZN(
        n4354) );
  ND4D1BWP12T U5313 ( .A1(n4357), .A2(n4356), .A3(n4355), .A4(n4354), .ZN(
        n4358) );
  AOI211D1BWP12T U5314 ( .A1(r0[6]), .A2(n4626), .B(n4359), .C(n4358), .ZN(
        n4360) );
  ND4D1BWP12T U5315 ( .A1(n4363), .A2(n4362), .A3(n4361), .A4(n4360), .ZN(
        regA_out[6]) );
  AOI22D1BWP12T U5316 ( .A1(r12[7]), .A2(n4654), .B1(r3[7]), .B2(n4589), .ZN(
        n4375) );
  AOI22D1BWP12T U5317 ( .A1(r4[7]), .A2(n4663), .B1(r6[7]), .B2(n4667), .ZN(
        n4374) );
  AOI22D1BWP12T U5318 ( .A1(r9[7]), .A2(n4666), .B1(r10[7]), .B2(n4665), .ZN(
        n4373) );
  AOI22D1BWP12T U5319 ( .A1(tmp1[7]), .A2(n4657), .B1(n3186), .B2(
        immediate1_in[7]), .ZN(n4364) );
  OAI21D1BWP12T U5320 ( .A1(n4365), .A2(n4641), .B(n4364), .ZN(n4371) );
  AOI22D1BWP12T U5321 ( .A1(r7[7]), .A2(n4656), .B1(sp_out[7]), .B2(n4655), 
        .ZN(n4369) );
  AOI22D1BWP12T U5322 ( .A1(r0[7]), .A2(n4626), .B1(r11[7]), .B2(n4659), .ZN(
        n4368) );
  AOI22D1BWP12T U5323 ( .A1(r5[7]), .A2(n4664), .B1(r2[7]), .B2(n4674), .ZN(
        n4367) );
  AOI22D1BWP12T U5324 ( .A1(r8[7]), .A2(n4627), .B1(lr[7]), .B2(n4653), .ZN(
        n4366) );
  ND4D1BWP12T U5325 ( .A1(n4369), .A2(n4368), .A3(n4367), .A4(n4366), .ZN(
        n4370) );
  AOI211D1BWP12T U5326 ( .A1(r1[7]), .A2(n4615), .B(n4371), .C(n4370), .ZN(
        n4372) );
  ND4D1BWP12T U5327 ( .A1(n4375), .A2(n4374), .A3(n4373), .A4(n4372), .ZN(
        regA_out[7]) );
  AOI22D1BWP12T U5328 ( .A1(r5[8]), .A2(n4664), .B1(r9[8]), .B2(n4666), .ZN(
        n4387) );
  AOI22D1BWP12T U5329 ( .A1(r0[8]), .A2(n4626), .B1(r2[8]), .B2(n4674), .ZN(
        n4386) );
  AOI22D1BWP12T U5330 ( .A1(r11[8]), .A2(n4659), .B1(n3186), .B2(
        immediate1_in[8]), .ZN(n4385) );
  AOI22D1BWP12T U5331 ( .A1(r4[8]), .A2(n4663), .B1(tmp1[8]), .B2(n4657), .ZN(
        n4376) );
  OAI21D1BWP12T U5332 ( .A1(n4377), .A2(n4601), .B(n4376), .ZN(n4383) );
  AOI22D1BWP12T U5333 ( .A1(r12[8]), .A2(n4654), .B1(r10[8]), .B2(n4665), .ZN(
        n4381) );
  AOI22D1BWP12T U5334 ( .A1(r8[8]), .A2(n4627), .B1(r6[8]), .B2(n4667), .ZN(
        n4380) );
  AOI22D1BWP12T U5335 ( .A1(r1[8]), .A2(n4615), .B1(sp_out[8]), .B2(n4655), 
        .ZN(n4379) );
  AOI22D1BWP12T U5336 ( .A1(r3[8]), .A2(n4589), .B1(pc_out[8]), .B2(n4658), 
        .ZN(n4378) );
  ND4D1BWP12T U5337 ( .A1(n4381), .A2(n4380), .A3(n4379), .A4(n4378), .ZN(
        n4382) );
  AOI211D1BWP12T U5338 ( .A1(r7[8]), .A2(n4656), .B(n4383), .C(n4382), .ZN(
        n4384) );
  ND4D1BWP12T U5339 ( .A1(n4387), .A2(n4386), .A3(n4385), .A4(n4384), .ZN(
        regA_out[8]) );
  AOI22D1BWP12T U5340 ( .A1(r4[9]), .A2(n4663), .B1(pc_out[9]), .B2(n4658), 
        .ZN(n4398) );
  AOI22D1BWP12T U5341 ( .A1(r12[9]), .A2(n4654), .B1(r9[9]), .B2(n4666), .ZN(
        n4397) );
  AOI22D1BWP12T U5342 ( .A1(r8[9]), .A2(n4627), .B1(sp_out[9]), .B2(n4655), 
        .ZN(n4396) );
  AOI22D1BWP12T U5343 ( .A1(tmp1[9]), .A2(n4657), .B1(r11[9]), .B2(n4659), 
        .ZN(n4388) );
  OAI21D1BWP12T U5344 ( .A1(n4827), .A2(n4601), .B(n4388), .ZN(n4394) );
  AOI22D1BWP12T U5345 ( .A1(r5[9]), .A2(n4664), .B1(r1[9]), .B2(n4615), .ZN(
        n4392) );
  AOI22D1BWP12T U5346 ( .A1(r2[9]), .A2(n4674), .B1(n3186), .B2(
        immediate1_in[9]), .ZN(n4391) );
  AOI22D1BWP12T U5347 ( .A1(r7[9]), .A2(n4656), .B1(r0[9]), .B2(n4626), .ZN(
        n4390) );
  AOI22D1BWP12T U5348 ( .A1(r3[9]), .A2(n4589), .B1(r10[9]), .B2(n4665), .ZN(
        n4389) );
  ND4D1BWP12T U5349 ( .A1(n4392), .A2(n4391), .A3(n4390), .A4(n4389), .ZN(
        n4393) );
  AOI211D1BWP12T U5350 ( .A1(r6[9]), .A2(n4667), .B(n4394), .C(n4393), .ZN(
        n4395) );
  ND4D1BWP12T U5351 ( .A1(n4398), .A2(n4397), .A3(n4396), .A4(n4395), .ZN(
        regA_out[9]) );
  AOI22D1BWP12T U5352 ( .A1(r3[10]), .A2(n4589), .B1(n3186), .B2(
        immediate1_in[10]), .ZN(n4410) );
  AOI22D1BWP12T U5353 ( .A1(r10[10]), .A2(n4665), .B1(r12[10]), .B2(n4654), 
        .ZN(n4409) );
  AOI22D1BWP12T U5354 ( .A1(r11[10]), .A2(n4659), .B1(r4[10]), .B2(n4663), 
        .ZN(n4400) );
  AOI22D1BWP12T U5355 ( .A1(r9[10]), .A2(n4666), .B1(r1[10]), .B2(n4615), .ZN(
        n4399) );
  OAI211D1BWP12T U5356 ( .A1(n4401), .A2(n4662), .B(n4400), .C(n4399), .ZN(
        n4407) );
  AOI22D1BWP12T U5357 ( .A1(r7[10]), .A2(n4656), .B1(r6[10]), .B2(n4667), .ZN(
        n4405) );
  AOI22D1BWP12T U5358 ( .A1(r5[10]), .A2(n4664), .B1(tmp1[10]), .B2(n4657), 
        .ZN(n4404) );
  AOI22D1BWP12T U5359 ( .A1(r0[10]), .A2(n4626), .B1(sp_out[10]), .B2(n4655), 
        .ZN(n4403) );
  AOI22D1BWP12T U5360 ( .A1(pc_out[10]), .A2(n4658), .B1(lr[10]), .B2(n4653), 
        .ZN(n4402) );
  ND4D1BWP12T U5361 ( .A1(n4405), .A2(n4404), .A3(n4403), .A4(n4402), .ZN(
        n4406) );
  AOI211D1BWP12T U5362 ( .A1(r2[10]), .A2(n4674), .B(n4407), .C(n4406), .ZN(
        n4408) );
  ND3D1BWP12T U5363 ( .A1(n4410), .A2(n4409), .A3(n4408), .ZN(regA_out[10]) );
  AOI22D1BWP12T U5364 ( .A1(r10[11]), .A2(n4665), .B1(r7[11]), .B2(n4656), 
        .ZN(n4422) );
  AOI22D1BWP12T U5365 ( .A1(lr[11]), .A2(n4653), .B1(r4[11]), .B2(n4663), .ZN(
        n4421) );
  AOI22D1BWP12T U5366 ( .A1(r9[11]), .A2(n4666), .B1(r6[11]), .B2(n4667), .ZN(
        n4420) );
  AOI22D1BWP12T U5367 ( .A1(r12[11]), .A2(n4654), .B1(r5[11]), .B2(n4664), 
        .ZN(n4411) );
  OAI21D1BWP12T U5368 ( .A1(n4412), .A2(n4641), .B(n4411), .ZN(n4418) );
  AOI22D1BWP12T U5369 ( .A1(r0[11]), .A2(n4626), .B1(r3[11]), .B2(n4589), .ZN(
        n4416) );
  AOI22D1BWP12T U5370 ( .A1(r11[11]), .A2(n4659), .B1(n3186), .B2(
        immediate1_in[11]), .ZN(n4415) );
  AOI22D1BWP12T U5371 ( .A1(r1[11]), .A2(n4615), .B1(sp_out[11]), .B2(n4655), 
        .ZN(n4414) );
  AOI22D1BWP12T U5372 ( .A1(r8[11]), .A2(n4627), .B1(tmp1[11]), .B2(n4657), 
        .ZN(n4413) );
  ND4D1BWP12T U5373 ( .A1(n4416), .A2(n4415), .A3(n4414), .A4(n4413), .ZN(
        n4417) );
  AOI211D1BWP12T U5374 ( .A1(r2[11]), .A2(n4674), .B(n4418), .C(n4417), .ZN(
        n4419) );
  ND4D1BWP12T U5375 ( .A1(n4422), .A2(n4421), .A3(n4420), .A4(n4419), .ZN(
        regA_out[11]) );
  AOI22D1BWP12T U5376 ( .A1(r2[12]), .A2(n4674), .B1(r6[12]), .B2(n4667), .ZN(
        n4434) );
  AOI22D1BWP12T U5377 ( .A1(r0[12]), .A2(n4626), .B1(r3[12]), .B2(n4589), .ZN(
        n4433) );
  AOI22D1BWP12T U5378 ( .A1(r4[12]), .A2(n4663), .B1(r7[12]), .B2(n4656), .ZN(
        n4432) );
  AOI22D1BWP12T U5379 ( .A1(lr[12]), .A2(n4653), .B1(r1[12]), .B2(n4615), .ZN(
        n4423) );
  OAI21D1BWP12T U5380 ( .A1(n4424), .A2(n4641), .B(n4423), .ZN(n4430) );
  AOI22D1BWP12T U5381 ( .A1(r12[12]), .A2(n4654), .B1(r10[12]), .B2(n4665), 
        .ZN(n4428) );
  AOI22D1BWP12T U5382 ( .A1(sp_out[12]), .A2(n4655), .B1(r5[12]), .B2(n4664), 
        .ZN(n4427) );
  AOI22D1BWP12T U5383 ( .A1(r11[12]), .A2(n4659), .B1(r8[12]), .B2(n4627), 
        .ZN(n4426) );
  AOI22D1BWP12T U5384 ( .A1(r9[12]), .A2(n4666), .B1(n3186), .B2(
        immediate1_in[12]), .ZN(n4425) );
  ND4D1BWP12T U5385 ( .A1(n4428), .A2(n4427), .A3(n4426), .A4(n4425), .ZN(
        n4429) );
  AOI211D1BWP12T U5386 ( .A1(tmp1[12]), .A2(n4657), .B(n4430), .C(n4429), .ZN(
        n4431) );
  ND4D1BWP12T U5387 ( .A1(n4434), .A2(n4433), .A3(n4432), .A4(n4431), .ZN(
        regA_out[12]) );
  AOI22D1BWP12T U5388 ( .A1(r9[13]), .A2(n4666), .B1(r6[13]), .B2(n4667), .ZN(
        n4446) );
  AOI22D1BWP12T U5389 ( .A1(r12[13]), .A2(n4654), .B1(r2[13]), .B2(n4674), 
        .ZN(n4445) );
  AOI22D1BWP12T U5390 ( .A1(r7[13]), .A2(n4656), .B1(sp_out[13]), .B2(n4655), 
        .ZN(n4444) );
  AOI22D1BWP12T U5391 ( .A1(r0[13]), .A2(n4626), .B1(r1[13]), .B2(n4615), .ZN(
        n4435) );
  OAI21D1BWP12T U5392 ( .A1(n4436), .A2(n4641), .B(n4435), .ZN(n4442) );
  AOI22D1BWP12T U5393 ( .A1(r10[13]), .A2(n4665), .B1(tmp1[13]), .B2(n4657), 
        .ZN(n4440) );
  AOI22D1BWP12T U5394 ( .A1(r5[13]), .A2(n4664), .B1(n3186), .B2(
        immediate1_in[13]), .ZN(n4439) );
  AOI22D1BWP12T U5395 ( .A1(r8[13]), .A2(n4627), .B1(r11[13]), .B2(n4659), 
        .ZN(n4438) );
  AOI22D1BWP12T U5396 ( .A1(r4[13]), .A2(n4663), .B1(lr[13]), .B2(n4653), .ZN(
        n4437) );
  ND4D1BWP12T U5397 ( .A1(n4440), .A2(n4439), .A3(n4438), .A4(n4437), .ZN(
        n4441) );
  AOI211D1BWP12T U5398 ( .A1(r3[13]), .A2(n4589), .B(n4442), .C(n4441), .ZN(
        n4443) );
  ND4D1BWP12T U5399 ( .A1(n4446), .A2(n4445), .A3(n4444), .A4(n4443), .ZN(
        regA_out[13]) );
  AOI22D1BWP12T U5400 ( .A1(r3[0]), .A2(n4214), .B1(lr[0]), .B2(n4447), .ZN(
        n4467) );
  AOI22D1BWP12T U5401 ( .A1(r0[0]), .A2(n4448), .B1(r2[0]), .B2(n4216), .ZN(
        n4466) );
  AOI22D1BWP12T U5402 ( .A1(r1[0]), .A2(n4450), .B1(sp_out[0]), .B2(n4449), 
        .ZN(n4465) );
  AOI22D1BWP12T U5403 ( .A1(r8[0]), .A2(n4452), .B1(r6[0]), .B2(n4451), .ZN(
        n4457) );
  AOI22D1BWP12T U5404 ( .A1(r11[0]), .A2(n3953), .B1(r4[0]), .B2(n3942), .ZN(
        n4456) );
  AOI22D1BWP12T U5405 ( .A1(r9[0]), .A2(n4218), .B1(r7[0]), .B2(n3985), .ZN(
        n4455) );
  AOI22D1BWP12T U5406 ( .A1(r10[0]), .A2(n4217), .B1(r5[0]), .B2(n4453), .ZN(
        n4454) );
  ND4D1BWP12T U5407 ( .A1(n4457), .A2(n4456), .A3(n4455), .A4(n4454), .ZN(
        n4462) );
  OAI22D1BWP12T U5408 ( .A1(n4860), .A2(n4460), .B1(n4459), .B2(n4458), .ZN(
        n4461) );
  AOI21D1BWP12T U5409 ( .A1(n4463), .A2(n4462), .B(n4461), .ZN(n4464) );
  ND4D1BWP12T U5410 ( .A1(n4467), .A2(n4466), .A3(n4465), .A4(n4464), .ZN(
        regD_out[0]) );
  AOI22D1BWP12T U5411 ( .A1(r12[15]), .A2(n4654), .B1(r3[15]), .B2(n4589), 
        .ZN(n4478) );
  AOI22D1BWP12T U5412 ( .A1(r0[15]), .A2(n4626), .B1(sp_out[15]), .B2(n4655), 
        .ZN(n4477) );
  AOI22D1BWP12T U5413 ( .A1(lr[15]), .A2(n4653), .B1(r4[15]), .B2(n4663), .ZN(
        n4476) );
  AOI22D1BWP12T U5414 ( .A1(r9[15]), .A2(n4666), .B1(r8[15]), .B2(n4627), .ZN(
        n4468) );
  OAI21D1BWP12T U5415 ( .A1(n4886), .A2(n4641), .B(n4468), .ZN(n4474) );
  AOI22D1BWP12T U5416 ( .A1(r11[15]), .A2(n4659), .B1(n3186), .B2(
        immediate1_in[15]), .ZN(n4472) );
  AOI22D1BWP12T U5417 ( .A1(tmp1[15]), .A2(n4657), .B1(r5[15]), .B2(n4664), 
        .ZN(n4471) );
  AOI22D1BWP12T U5418 ( .A1(r6[15]), .A2(n4667), .B1(r1[15]), .B2(n4615), .ZN(
        n4470) );
  AOI22D1BWP12T U5419 ( .A1(r7[15]), .A2(n4656), .B1(r2[15]), .B2(n4674), .ZN(
        n4469) );
  ND4D1BWP12T U5420 ( .A1(n4472), .A2(n4471), .A3(n4470), .A4(n4469), .ZN(
        n4473) );
  AOI211D1BWP12T U5421 ( .A1(r10[15]), .A2(n4665), .B(n4474), .C(n4473), .ZN(
        n4475) );
  ND4D1BWP12T U5422 ( .A1(n4478), .A2(n4477), .A3(n4476), .A4(n4475), .ZN(
        regA_out[15]) );
  AOI22D1BWP12T U5423 ( .A1(r3[16]), .A2(n4589), .B1(r9[16]), .B2(n4666), .ZN(
        n4490) );
  AOI22D1BWP12T U5424 ( .A1(r11[16]), .A2(n4659), .B1(r2[16]), .B2(n4674), 
        .ZN(n4489) );
  AOI22D1BWP12T U5425 ( .A1(r5[16]), .A2(n4664), .B1(tmp1[16]), .B2(n4657), 
        .ZN(n4480) );
  AOI22D1BWP12T U5426 ( .A1(r8[16]), .A2(n4627), .B1(r12[16]), .B2(n4654), 
        .ZN(n4479) );
  OAI211D1BWP12T U5427 ( .A1(n4481), .A2(n4641), .B(n4480), .C(n4479), .ZN(
        n4487) );
  AOI22D1BWP12T U5428 ( .A1(lr[16]), .A2(n4653), .B1(r6[16]), .B2(n4667), .ZN(
        n4485) );
  AOI22D1BWP12T U5429 ( .A1(sp_out[16]), .A2(n4655), .B1(r0[16]), .B2(n4626), 
        .ZN(n4484) );
  AOI22D1BWP12T U5430 ( .A1(r7[16]), .A2(n4656), .B1(r1[16]), .B2(n4615), .ZN(
        n4483) );
  AOI22D1BWP12T U5431 ( .A1(r10[16]), .A2(n4665), .B1(n3186), .B2(
        immediate1_in[16]), .ZN(n4482) );
  ND4D1BWP12T U5432 ( .A1(n4485), .A2(n4484), .A3(n4483), .A4(n4482), .ZN(
        n4486) );
  AOI211D1BWP12T U5433 ( .A1(r4[16]), .A2(n4663), .B(n4487), .C(n4486), .ZN(
        n4488) );
  ND3D1BWP12T U5434 ( .A1(n4490), .A2(n4489), .A3(n4488), .ZN(regA_out[16]) );
  AOI22D1BWP12T U5435 ( .A1(r6[17]), .A2(n4667), .B1(r7[17]), .B2(n4656), .ZN(
        n4502) );
  AOI22D1BWP12T U5436 ( .A1(r2[17]), .A2(n4674), .B1(pc_out[17]), .B2(n4658), 
        .ZN(n4501) );
  AOI22D1BWP12T U5437 ( .A1(r1[17]), .A2(n4615), .B1(sp_out[17]), .B2(n4655), 
        .ZN(n4500) );
  AOI22D1BWP12T U5438 ( .A1(r0[17]), .A2(n4626), .B1(n3186), .B2(
        immediate1_in[17]), .ZN(n4491) );
  OAI21D1BWP12T U5439 ( .A1(n4492), .A2(n4662), .B(n4491), .ZN(n4498) );
  AOI22D1BWP12T U5440 ( .A1(r12[17]), .A2(n4654), .B1(r9[17]), .B2(n4666), 
        .ZN(n4496) );
  AOI22D1BWP12T U5441 ( .A1(r4[17]), .A2(n4663), .B1(r11[17]), .B2(n4659), 
        .ZN(n4495) );
  AOI22D1BWP12T U5442 ( .A1(tmp1[17]), .A2(n4657), .B1(r5[17]), .B2(n4664), 
        .ZN(n4494) );
  AOI22D1BWP12T U5443 ( .A1(r3[17]), .A2(n4589), .B1(r10[17]), .B2(n4665), 
        .ZN(n4493) );
  ND4D1BWP12T U5444 ( .A1(n4496), .A2(n4495), .A3(n4494), .A4(n4493), .ZN(
        n4497) );
  AOI211D1BWP12T U5445 ( .A1(lr[17]), .A2(n4653), .B(n4498), .C(n4497), .ZN(
        n4499) );
  ND4D1BWP12T U5446 ( .A1(n4502), .A2(n4501), .A3(n4500), .A4(n4499), .ZN(
        regA_out[17]) );
  AOI22D1BWP12T U5447 ( .A1(r9[18]), .A2(n4666), .B1(r7[18]), .B2(n4656), .ZN(
        n4514) );
  AOI22D1BWP12T U5448 ( .A1(r12[18]), .A2(n4654), .B1(pc_out[18]), .B2(n4658), 
        .ZN(n4513) );
  AOI22D1BWP12T U5449 ( .A1(r1[18]), .A2(n4615), .B1(sp_out[18]), .B2(n4655), 
        .ZN(n4512) );
  AOI22D1BWP12T U5450 ( .A1(r5[18]), .A2(n4664), .B1(r2[18]), .B2(n4674), .ZN(
        n4503) );
  OAI21D1BWP12T U5451 ( .A1(n4504), .A2(n4601), .B(n4503), .ZN(n4510) );
  AOI22D1BWP12T U5452 ( .A1(r10[18]), .A2(n4665), .B1(r11[18]), .B2(n4659), 
        .ZN(n4508) );
  AOI22D1BWP12T U5453 ( .A1(r8[18]), .A2(n4627), .B1(n3186), .B2(
        immediate1_in[18]), .ZN(n4507) );
  AOI22D1BWP12T U5454 ( .A1(r0[18]), .A2(n4626), .B1(r4[18]), .B2(n4663), .ZN(
        n4506) );
  AOI22D1BWP12T U5455 ( .A1(r6[18]), .A2(n4667), .B1(r3[18]), .B2(n4589), .ZN(
        n4505) );
  ND4D1BWP12T U5456 ( .A1(n4508), .A2(n4507), .A3(n4506), .A4(n4505), .ZN(
        n4509) );
  AOI211D1BWP12T U5457 ( .A1(tmp1[18]), .A2(n4657), .B(n4510), .C(n4509), .ZN(
        n4511) );
  ND4D1BWP12T U5458 ( .A1(n4514), .A2(n4513), .A3(n4512), .A4(n4511), .ZN(
        regA_out[18]) );
  AOI22D1BWP12T U5459 ( .A1(r6[19]), .A2(n4667), .B1(sp_out[19]), .B2(n4655), 
        .ZN(n4526) );
  AOI22D1BWP12T U5460 ( .A1(r7[19]), .A2(n4656), .B1(r2[19]), .B2(n4674), .ZN(
        n4525) );
  AOI22D1BWP12T U5461 ( .A1(r9[19]), .A2(n4666), .B1(r8[19]), .B2(n4627), .ZN(
        n4524) );
  AOI22D1BWP12T U5462 ( .A1(r4[19]), .A2(n4663), .B1(n3186), .B2(
        immediate1_in[19]), .ZN(n4515) );
  OAI21D1BWP12T U5463 ( .A1(n4516), .A2(n4601), .B(n4515), .ZN(n4522) );
  AOI22D1BWP12T U5464 ( .A1(r0[19]), .A2(n4626), .B1(r12[19]), .B2(n4654), 
        .ZN(n4520) );
  AOI22D1BWP12T U5465 ( .A1(r11[19]), .A2(n4659), .B1(r1[19]), .B2(n4615), 
        .ZN(n4519) );
  AOI22D1BWP12T U5466 ( .A1(r5[19]), .A2(n4664), .B1(r3[19]), .B2(n4589), .ZN(
        n4518) );
  AOI22D1BWP12T U5467 ( .A1(r10[19]), .A2(n4665), .B1(pc_out[19]), .B2(n4658), 
        .ZN(n4517) );
  ND4D1BWP12T U5468 ( .A1(n4520), .A2(n4519), .A3(n4518), .A4(n4517), .ZN(
        n4521) );
  AOI211D1BWP12T U5469 ( .A1(tmp1[19]), .A2(n4657), .B(n4522), .C(n4521), .ZN(
        n4523) );
  ND4D1BWP12T U5470 ( .A1(n4526), .A2(n4525), .A3(n4524), .A4(n4523), .ZN(
        regA_out[19]) );
  AOI22D1BWP12T U5471 ( .A1(lr[20]), .A2(n4653), .B1(r0[20]), .B2(n4626), .ZN(
        n4538) );
  AOI22D1BWP12T U5472 ( .A1(r6[20]), .A2(n4667), .B1(r5[20]), .B2(n4664), .ZN(
        n4537) );
  AOI22D1BWP12T U5473 ( .A1(r3[20]), .A2(n4589), .B1(n3186), .B2(
        immediate1_in[20]), .ZN(n4536) );
  AOI22D1BWP12T U5474 ( .A1(sp_out[20]), .A2(n4655), .B1(r10[20]), .B2(n4665), 
        .ZN(n4527) );
  OAI21D1BWP12T U5475 ( .A1(n4528), .A2(n4641), .B(n4527), .ZN(n4534) );
  AOI22D1BWP12T U5476 ( .A1(r9[20]), .A2(n4666), .B1(r8[20]), .B2(n4627), .ZN(
        n4532) );
  AOI22D1BWP12T U5477 ( .A1(r7[20]), .A2(n4656), .B1(tmp1[20]), .B2(n4657), 
        .ZN(n4531) );
  AOI22D1BWP12T U5478 ( .A1(r2[20]), .A2(n4674), .B1(r1[20]), .B2(n4615), .ZN(
        n4530) );
  AOI22D1BWP12T U5479 ( .A1(r11[20]), .A2(n4659), .B1(r12[20]), .B2(n4654), 
        .ZN(n4529) );
  ND4D1BWP12T U5480 ( .A1(n4532), .A2(n4531), .A3(n4530), .A4(n4529), .ZN(
        n4533) );
  AOI211D1BWP12T U5481 ( .A1(r4[20]), .A2(n4663), .B(n4534), .C(n4533), .ZN(
        n4535) );
  ND4D1BWP12T U5482 ( .A1(n4538), .A2(n4537), .A3(n4536), .A4(n4535), .ZN(
        regA_out[20]) );
  AOI22D1BWP12T U5483 ( .A1(r7[21]), .A2(n4656), .B1(r12[21]), .B2(n4654), 
        .ZN(n4550) );
  AOI22D1BWP12T U5484 ( .A1(r10[21]), .A2(n4665), .B1(r8[21]), .B2(n4627), 
        .ZN(n4549) );
  AOI22D1BWP12T U5485 ( .A1(r6[21]), .A2(n4667), .B1(r9[21]), .B2(n4666), .ZN(
        n4540) );
  AOI22D1BWP12T U5486 ( .A1(r1[21]), .A2(n4615), .B1(tmp1[21]), .B2(n4657), 
        .ZN(n4539) );
  OAI211D1BWP12T U5487 ( .A1(n4541), .A2(n4641), .B(n4540), .C(n4539), .ZN(
        n4547) );
  AOI22D1BWP12T U5488 ( .A1(sp_out[21]), .A2(n4655), .B1(lr[21]), .B2(n4653), 
        .ZN(n4545) );
  AOI22D1BWP12T U5489 ( .A1(r3[21]), .A2(n4589), .B1(r5[21]), .B2(n4664), .ZN(
        n4544) );
  AOI22D1BWP12T U5490 ( .A1(r2[21]), .A2(n4674), .B1(n3186), .B2(
        immediate1_in[21]), .ZN(n4543) );
  AOI22D1BWP12T U5491 ( .A1(r11[21]), .A2(n4659), .B1(r4[21]), .B2(n4663), 
        .ZN(n4542) );
  ND4D1BWP12T U5492 ( .A1(n4545), .A2(n4544), .A3(n4543), .A4(n4542), .ZN(
        n4546) );
  AOI211D1BWP12T U5493 ( .A1(r0[21]), .A2(n4626), .B(n4547), .C(n4546), .ZN(
        n4548) );
  ND3D1BWP12T U5494 ( .A1(n4550), .A2(n4549), .A3(n4548), .ZN(regA_out[21]) );
  AOI22D1BWP12T U5495 ( .A1(lr[22]), .A2(n4653), .B1(r6[22]), .B2(n4667), .ZN(
        n4562) );
  AOI22D1BWP12T U5496 ( .A1(r1[22]), .A2(n4615), .B1(r8[22]), .B2(n4627), .ZN(
        n4561) );
  AOI22D1BWP12T U5497 ( .A1(sp_out[22]), .A2(n4655), .B1(r2[22]), .B2(n4674), 
        .ZN(n4560) );
  AOI22D1BWP12T U5498 ( .A1(r0[22]), .A2(n4626), .B1(r3[22]), .B2(n4589), .ZN(
        n4551) );
  OAI21D1BWP12T U5499 ( .A1(n4552), .A2(n4641), .B(n4551), .ZN(n4558) );
  AOI22D1BWP12T U5500 ( .A1(r7[22]), .A2(n4656), .B1(n3186), .B2(
        immediate1_in[22]), .ZN(n4556) );
  AOI22D1BWP12T U5501 ( .A1(r10[22]), .A2(n4665), .B1(r11[22]), .B2(n4659), 
        .ZN(n4555) );
  AOI22D1BWP12T U5502 ( .A1(r9[22]), .A2(n4666), .B1(r4[22]), .B2(n4663), .ZN(
        n4554) );
  AOI22D1BWP12T U5503 ( .A1(tmp1[22]), .A2(n4657), .B1(r12[22]), .B2(n4654), 
        .ZN(n4553) );
  ND4D1BWP12T U5504 ( .A1(n4556), .A2(n4555), .A3(n4554), .A4(n4553), .ZN(
        n4557) );
  AOI211D1BWP12T U5505 ( .A1(r5[22]), .A2(n4664), .B(n4558), .C(n4557), .ZN(
        n4559) );
  ND4D1BWP12T U5506 ( .A1(n4562), .A2(n4561), .A3(n4560), .A4(n4559), .ZN(
        regA_out[22]) );
  AOI22D1BWP12T U5507 ( .A1(r5[23]), .A2(n4664), .B1(n3186), .B2(
        immediate1_in[23]), .ZN(n4574) );
  AOI22D1BWP12T U5508 ( .A1(r9[23]), .A2(n4666), .B1(r4[23]), .B2(n4663), .ZN(
        n4573) );
  AOI22D1BWP12T U5509 ( .A1(r11[23]), .A2(n4659), .B1(r1[23]), .B2(n4615), 
        .ZN(n4572) );
  AOI22D1BWP12T U5510 ( .A1(lr[23]), .A2(n4653), .B1(r12[23]), .B2(n4654), 
        .ZN(n4563) );
  OAI21D1BWP12T U5511 ( .A1(n4564), .A2(n4641), .B(n4563), .ZN(n4570) );
  AOI22D1BWP12T U5512 ( .A1(r10[23]), .A2(n4665), .B1(r0[23]), .B2(n4626), 
        .ZN(n4568) );
  AOI22D1BWP12T U5513 ( .A1(r2[23]), .A2(n4674), .B1(sp_out[23]), .B2(n4655), 
        .ZN(n4567) );
  AOI22D1BWP12T U5514 ( .A1(r6[23]), .A2(n4667), .B1(r3[23]), .B2(n4589), .ZN(
        n4566) );
  AOI22D1BWP12T U5515 ( .A1(tmp1[23]), .A2(n4657), .B1(r8[23]), .B2(n4627), 
        .ZN(n4565) );
  ND4D1BWP12T U5516 ( .A1(n4568), .A2(n4567), .A3(n4566), .A4(n4565), .ZN(
        n4569) );
  AOI211D1BWP12T U5517 ( .A1(r7[23]), .A2(n4656), .B(n4570), .C(n4569), .ZN(
        n4571) );
  ND4D1BWP12T U5518 ( .A1(n4574), .A2(n4573), .A3(n4572), .A4(n4571), .ZN(
        regA_out[23]) );
  AOI22D1BWP12T U5519 ( .A1(r10[24]), .A2(n4665), .B1(r2[24]), .B2(n4674), 
        .ZN(n4586) );
  AOI22D1BWP12T U5520 ( .A1(r9[24]), .A2(n4666), .B1(r7[24]), .B2(n4656), .ZN(
        n4585) );
  AOI22D1BWP12T U5521 ( .A1(r3[24]), .A2(n4589), .B1(sp_out[24]), .B2(n4655), 
        .ZN(n4584) );
  AOI22D1BWP12T U5522 ( .A1(r1[24]), .A2(n4615), .B1(n3186), .B2(
        immediate1_in[24]), .ZN(n4575) );
  OAI21D1BWP12T U5523 ( .A1(n4576), .A2(n4641), .B(n4575), .ZN(n4582) );
  AOI22D1BWP12T U5524 ( .A1(r11[24]), .A2(n4659), .B1(tmp1[24]), .B2(n4657), 
        .ZN(n4580) );
  AOI22D1BWP12T U5525 ( .A1(r5[24]), .A2(n4664), .B1(r4[24]), .B2(n4663), .ZN(
        n4579) );
  AOI22D1BWP12T U5526 ( .A1(r8[24]), .A2(n4627), .B1(r6[24]), .B2(n4667), .ZN(
        n4578) );
  AOI22D1BWP12T U5527 ( .A1(lr[24]), .A2(n4653), .B1(r12[24]), .B2(n4654), 
        .ZN(n4577) );
  ND4D1BWP12T U5528 ( .A1(n4580), .A2(n4579), .A3(n4578), .A4(n4577), .ZN(
        n4581) );
  AOI211D1BWP12T U5529 ( .A1(r0[24]), .A2(n4626), .B(n4582), .C(n4581), .ZN(
        n4583) );
  ND4D1BWP12T U5530 ( .A1(n4586), .A2(n4585), .A3(n4584), .A4(n4583), .ZN(
        regA_out[24]) );
  AOI22D1BWP12T U5531 ( .A1(tmp1[25]), .A2(n4657), .B1(r0[25]), .B2(n4626), 
        .ZN(n4599) );
  AOI22D1BWP12T U5532 ( .A1(r2[25]), .A2(n4674), .B1(r7[25]), .B2(n4656), .ZN(
        n4598) );
  AOI22D1BWP12T U5533 ( .A1(sp_out[25]), .A2(n4655), .B1(r1[25]), .B2(n4615), 
        .ZN(n4597) );
  AOI22D1BWP12T U5534 ( .A1(lr[25]), .A2(n4653), .B1(r12[25]), .B2(n4654), 
        .ZN(n4587) );
  OAI21D1BWP12T U5535 ( .A1(n4588), .A2(n4641), .B(n4587), .ZN(n4595) );
  AOI22D1BWP12T U5536 ( .A1(r8[25]), .A2(n4627), .B1(r6[25]), .B2(n4667), .ZN(
        n4593) );
  AOI22D1BWP12T U5537 ( .A1(r3[25]), .A2(n4589), .B1(r5[25]), .B2(n4664), .ZN(
        n4592) );
  AOI22D1BWP12T U5538 ( .A1(r11[25]), .A2(n4659), .B1(r9[25]), .B2(n4666), 
        .ZN(n4591) );
  AOI22D1BWP12T U5539 ( .A1(r10[25]), .A2(n4665), .B1(n3186), .B2(
        immediate1_in[25]), .ZN(n4590) );
  ND4D1BWP12T U5540 ( .A1(n4593), .A2(n4592), .A3(n4591), .A4(n4590), .ZN(
        n4594) );
  AOI211D1BWP12T U5541 ( .A1(r4[25]), .A2(n4663), .B(n4595), .C(n4594), .ZN(
        n4596) );
  ND4D1BWP12T U5542 ( .A1(n4599), .A2(n4598), .A3(n4597), .A4(n4596), .ZN(
        regA_out[25]) );
  AOI22D1BWP12T U5543 ( .A1(r11[26]), .A2(n4659), .B1(pc_out[26]), .B2(n4658), 
        .ZN(n4612) );
  AOI22D1BWP12T U5544 ( .A1(r5[26]), .A2(n4664), .B1(r2[26]), .B2(n4674), .ZN(
        n4611) );
  AOI22D1BWP12T U5545 ( .A1(r4[26]), .A2(n4663), .B1(r8[26]), .B2(n4627), .ZN(
        n4610) );
  AOI22D1BWP12T U5546 ( .A1(tmp1[26]), .A2(n4657), .B1(r9[26]), .B2(n4666), 
        .ZN(n4600) );
  OAI21D1BWP12T U5547 ( .A1(n4602), .A2(n4601), .B(n4600), .ZN(n4608) );
  AOI22D1BWP12T U5548 ( .A1(r1[26]), .A2(n4615), .B1(r0[26]), .B2(n4626), .ZN(
        n4606) );
  AOI22D1BWP12T U5549 ( .A1(r12[26]), .A2(n4654), .B1(r7[26]), .B2(n4656), 
        .ZN(n4605) );
  AOI22D1BWP12T U5550 ( .A1(sp_out[26]), .A2(n4655), .B1(n3186), .B2(
        immediate1_in[26]), .ZN(n4604) );
  AOI22D1BWP12T U5551 ( .A1(r10[26]), .A2(n4665), .B1(r3[26]), .B2(n4589), 
        .ZN(n4603) );
  ND4D1BWP12T U5552 ( .A1(n4606), .A2(n4605), .A3(n4604), .A4(n4603), .ZN(
        n4607) );
  AOI211D1BWP12T U5553 ( .A1(r6[26]), .A2(n4667), .B(n4608), .C(n4607), .ZN(
        n4609) );
  ND4D1BWP12T U5554 ( .A1(n4612), .A2(n4611), .A3(n4610), .A4(n4609), .ZN(
        regA_out[26]) );
  AOI22D1BWP12T U5555 ( .A1(r4[27]), .A2(n4663), .B1(n3186), .B2(
        immediate1_in[27]), .ZN(n4625) );
  AOI22D1BWP12T U5556 ( .A1(lr[27]), .A2(n4653), .B1(r12[27]), .B2(n4654), 
        .ZN(n4624) );
  AOI22D1BWP12T U5557 ( .A1(r6[27]), .A2(n4667), .B1(tmp1[27]), .B2(n4657), 
        .ZN(n4623) );
  AOI22D1BWP12T U5558 ( .A1(r0[27]), .A2(n4626), .B1(pc_out[27]), .B2(n4658), 
        .ZN(n4613) );
  OAI21D1BWP12T U5559 ( .A1(n4614), .A2(n4662), .B(n4613), .ZN(n4621) );
  AOI22D1BWP12T U5560 ( .A1(r7[27]), .A2(n4656), .B1(r9[27]), .B2(n4666), .ZN(
        n4619) );
  AOI22D1BWP12T U5561 ( .A1(sp_out[27]), .A2(n4655), .B1(r3[27]), .B2(n4589), 
        .ZN(n4618) );
  AOI22D1BWP12T U5562 ( .A1(r5[27]), .A2(n4664), .B1(r2[27]), .B2(n4674), .ZN(
        n4617) );
  AOI22D1BWP12T U5563 ( .A1(r1[27]), .A2(n4615), .B1(r11[27]), .B2(n4659), 
        .ZN(n4616) );
  ND4D1BWP12T U5564 ( .A1(n4619), .A2(n4618), .A3(n4617), .A4(n4616), .ZN(
        n4620) );
  AOI211D1BWP12T U5565 ( .A1(r10[27]), .A2(n4665), .B(n4621), .C(n4620), .ZN(
        n4622) );
  ND4D1BWP12T U5566 ( .A1(n4625), .A2(n4624), .A3(n4623), .A4(n4622), .ZN(
        regA_out[27]) );
  AOI22D1BWP12T U5567 ( .A1(r0[28]), .A2(n4626), .B1(tmp1[28]), .B2(n4657), 
        .ZN(n4639) );
  AOI22D1BWP12T U5568 ( .A1(lr[28]), .A2(n4653), .B1(r8[28]), .B2(n4627), .ZN(
        n4638) );
  AOI22D1BWP12T U5569 ( .A1(r9[28]), .A2(n4666), .B1(r1[28]), .B2(n4615), .ZN(
        n4629) );
  AOI22D1BWP12T U5570 ( .A1(r3[28]), .A2(n4589), .B1(r6[28]), .B2(n4667), .ZN(
        n4628) );
  OAI211D1BWP12T U5571 ( .A1(n4630), .A2(n4641), .B(n4629), .C(n4628), .ZN(
        n4636) );
  AOI22D1BWP12T U5572 ( .A1(r7[28]), .A2(n4656), .B1(r2[28]), .B2(n4674), .ZN(
        n4634) );
  AOI22D1BWP12T U5573 ( .A1(r11[28]), .A2(n4659), .B1(r5[28]), .B2(n4664), 
        .ZN(n4633) );
  AOI22D1BWP12T U5574 ( .A1(r4[28]), .A2(n4663), .B1(sp_out[28]), .B2(n4655), 
        .ZN(n4632) );
  AOI22D1BWP12T U5575 ( .A1(r12[28]), .A2(n4654), .B1(n3186), .B2(
        immediate1_in[28]), .ZN(n4631) );
  ND4D1BWP12T U5576 ( .A1(n4634), .A2(n4633), .A3(n4632), .A4(n4631), .ZN(
        n4635) );
  AOI211D1BWP12T U5577 ( .A1(r10[28]), .A2(n4665), .B(n4636), .C(n4635), .ZN(
        n4637) );
  ND3D1BWP12T U5578 ( .A1(n4639), .A2(n4638), .A3(n4637), .ZN(regA_out[28]) );
  AOI22D1BWP12T U5579 ( .A1(r12[30]), .A2(n4654), .B1(r3[30]), .B2(n4589), 
        .ZN(n4652) );
  AOI22D1BWP12T U5580 ( .A1(tmp1[30]), .A2(n4657), .B1(r0[30]), .B2(n4626), 
        .ZN(n4651) );
  AOI22D1BWP12T U5581 ( .A1(r5[30]), .A2(n4664), .B1(r2[30]), .B2(n4674), .ZN(
        n4650) );
  AOI22D1BWP12T U5582 ( .A1(r10[30]), .A2(n4665), .B1(n3186), .B2(
        immediate1_in[30]), .ZN(n4640) );
  OAI21D1BWP12T U5583 ( .A1(n4642), .A2(n4641), .B(n4640), .ZN(n4648) );
  AOI22D1BWP12T U5584 ( .A1(r1[30]), .A2(n4615), .B1(r7[30]), .B2(n4656), .ZN(
        n4646) );
  AOI22D1BWP12T U5585 ( .A1(r6[30]), .A2(n4667), .B1(r8[30]), .B2(n4627), .ZN(
        n4645) );
  AOI22D1BWP12T U5586 ( .A1(r9[30]), .A2(n4666), .B1(sp_out[30]), .B2(n4655), 
        .ZN(n4644) );
  AOI22D1BWP12T U5587 ( .A1(lr[30]), .A2(n4653), .B1(r11[30]), .B2(n4659), 
        .ZN(n4643) );
  ND4D1BWP12T U5588 ( .A1(n4646), .A2(n4645), .A3(n4644), .A4(n4643), .ZN(
        n4647) );
  AOI211D1BWP12T U5589 ( .A1(r4[30]), .A2(n4663), .B(n4648), .C(n4647), .ZN(
        n4649) );
  ND4D1BWP12T U5590 ( .A1(n4652), .A2(n4651), .A3(n4650), .A4(n4649), .ZN(
        regA_out[30]) );
  AOI22D1BWP12T U5591 ( .A1(r12[29]), .A2(n4654), .B1(lr[29]), .B2(n4653), 
        .ZN(n4677) );
  AOI22D1BWP12T U5592 ( .A1(sp_out[29]), .A2(n4655), .B1(r0[29]), .B2(n4626), 
        .ZN(n4676) );
  AOI22D1BWP12T U5593 ( .A1(tmp1[29]), .A2(n4657), .B1(r7[29]), .B2(n4656), 
        .ZN(n4661) );
  AOI22D1BWP12T U5594 ( .A1(r11[29]), .A2(n4659), .B1(pc_out[29]), .B2(n4658), 
        .ZN(n4660) );
  OAI211D1BWP12T U5595 ( .A1(n4824), .A2(n4662), .B(n4661), .C(n4660), .ZN(
        n4673) );
  AOI22D1BWP12T U5596 ( .A1(r5[29]), .A2(n4664), .B1(r4[29]), .B2(n4663), .ZN(
        n4671) );
  AOI22D1BWP12T U5597 ( .A1(r10[29]), .A2(n4665), .B1(r1[29]), .B2(n4615), 
        .ZN(n4670) );
  AOI22D1BWP12T U5598 ( .A1(r9[29]), .A2(n4666), .B1(n3186), .B2(
        immediate1_in[29]), .ZN(n4669) );
  AOI22D1BWP12T U5599 ( .A1(r6[29]), .A2(n4667), .B1(r3[29]), .B2(n4589), .ZN(
        n4668) );
  ND4D1BWP12T U5600 ( .A1(n4671), .A2(n4670), .A3(n4669), .A4(n4668), .ZN(
        n4672) );
  AOI211D1BWP12T U5601 ( .A1(r2[29]), .A2(n4674), .B(n4673), .C(n4672), .ZN(
        n4675) );
  ND3D1BWP12T U5602 ( .A1(n4677), .A2(n4676), .A3(n4675), .ZN(regA_out[29]) );
  TPND2D0BWP12T U5603 ( .A1(n4753), .A2(n4678), .ZN(n4681) );
  OR2XD0BWP12T U5604 ( .A1(n4752), .A2(n4679), .Z(n4682) );
  ND2D1BWP12T U5605 ( .A1(n4681), .A2(n4682), .ZN(n4680) );
  AOI22D1BWP12T U5606 ( .A1(pc_out[15]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[15]), .ZN(n4887) );
  AOI22D1BWP12T U5607 ( .A1(n4742), .A2(write1_in[15]), .B1(n4741), .B2(
        write2_in[15]), .ZN(n4888) );
  AOI22D1BWP12T U5608 ( .A1(n4742), .A2(write1_in[6]), .B1(n4741), .B2(
        write2_in[6]), .ZN(n4684) );
  AOI22D1BWP12T U5609 ( .A1(pc_out[6]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[6]), .ZN(n4683) );
  ND2D1BWP12T U5610 ( .A1(n4684), .A2(n4683), .ZN(n2207) );
  AOI22D1BWP12T U5611 ( .A1(n4742), .A2(write1_in[13]), .B1(n4741), .B2(
        write2_in[13]), .ZN(n4686) );
  AOI22D1BWP12T U5612 ( .A1(pc_out[13]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[13]), .ZN(n4685) );
  ND2D1BWP12T U5613 ( .A1(n4686), .A2(n4685), .ZN(n2214) );
  AOI22D1BWP12T U5614 ( .A1(n4742), .A2(write1_in[2]), .B1(n4741), .B2(
        write2_in[2]), .ZN(n4688) );
  AOI22D1BWP12T U5615 ( .A1(pc_out[2]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[2]), .ZN(n4687) );
  ND2D1BWP12T U5616 ( .A1(n4688), .A2(n4687), .ZN(n2203) );
  AOI22D1BWP12T U5617 ( .A1(n4742), .A2(write1_in[20]), .B1(n4741), .B2(
        write2_in[20]), .ZN(n4690) );
  AOI22D1BWP12T U5618 ( .A1(pc_out[20]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[20]), .ZN(n4689) );
  ND2D1BWP12T U5619 ( .A1(n4690), .A2(n4689), .ZN(n2221) );
  AOI22D1BWP12T U5620 ( .A1(n4742), .A2(write1_in[0]), .B1(n4741), .B2(
        write2_in[0]), .ZN(n4692) );
  AOI22D1BWP12T U5621 ( .A1(pc_out[0]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[0]), .ZN(n4691) );
  ND2D1BWP12T U5622 ( .A1(n4692), .A2(n4691), .ZN(n2201) );
  AOI22D1BWP12T U5623 ( .A1(n4742), .A2(write1_in[22]), .B1(n4741), .B2(
        write2_in[22]), .ZN(n4694) );
  AOI22D1BWP12T U5624 ( .A1(pc_out[22]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[22]), .ZN(n4693) );
  ND2D1BWP12T U5625 ( .A1(n4694), .A2(n4693), .ZN(n2223) );
  AOI22D1BWP12T U5626 ( .A1(n4742), .A2(write1_in[23]), .B1(n4741), .B2(
        write2_in[23]), .ZN(n4696) );
  AOI22D1BWP12T U5627 ( .A1(pc_out[23]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[23]), .ZN(n4695) );
  ND2D1BWP12T U5628 ( .A1(n4696), .A2(n4695), .ZN(n2224) );
  AOI22D1BWP12T U5629 ( .A1(n4742), .A2(write1_in[12]), .B1(n4741), .B2(
        write2_in[12]), .ZN(n4698) );
  AOI22D1BWP12T U5630 ( .A1(pc_out[12]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[12]), .ZN(n4697) );
  ND2D1BWP12T U5631 ( .A1(n4698), .A2(n4697), .ZN(n2213) );
  AOI22D1BWP12T U5632 ( .A1(n4742), .A2(write1_in[11]), .B1(n4741), .B2(
        write2_in[11]), .ZN(n4700) );
  AOI22D1BWP12T U5633 ( .A1(pc_out[11]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[11]), .ZN(n4699) );
  ND2D1BWP12T U5634 ( .A1(n4700), .A2(n4699), .ZN(n2212) );
  AOI22D1BWP12T U5635 ( .A1(n4742), .A2(write1_in[1]), .B1(n4741), .B2(
        write2_in[1]), .ZN(n4702) );
  AOI22D1BWP12T U5636 ( .A1(pc_out[1]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[1]), .ZN(n4701) );
  ND2D1BWP12T U5637 ( .A1(n4702), .A2(n4701), .ZN(n2202) );
  AOI22D1BWP12T U5638 ( .A1(n4742), .A2(write1_in[29]), .B1(n4741), .B2(
        write2_in[29]), .ZN(n4704) );
  AOI22D1BWP12T U5639 ( .A1(pc_out[29]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[29]), .ZN(n4703) );
  ND2D1BWP12T U5640 ( .A1(n4704), .A2(n4703), .ZN(n2230) );
  AOI22D1BWP12T U5641 ( .A1(n4742), .A2(write1_in[3]), .B1(n4741), .B2(
        write2_in[3]), .ZN(n4706) );
  AOI22D1BWP12T U5642 ( .A1(pc_out[3]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[3]), .ZN(n4705) );
  ND2D1BWP12T U5643 ( .A1(n4706), .A2(n4705), .ZN(n2204) );
  AOI22D1BWP12T U5644 ( .A1(n4742), .A2(write1_in[24]), .B1(n4741), .B2(
        write2_in[24]), .ZN(n4708) );
  AOI22D1BWP12T U5645 ( .A1(pc_out[24]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[24]), .ZN(n4707) );
  ND2D1BWP12T U5646 ( .A1(n4708), .A2(n4707), .ZN(n2225) );
  AOI22D1BWP12T U5647 ( .A1(n4742), .A2(write1_in[21]), .B1(n4741), .B2(
        write2_in[21]), .ZN(n4710) );
  AOI22D1BWP12T U5648 ( .A1(pc_out[21]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[21]), .ZN(n4709) );
  ND2D1BWP12T U5649 ( .A1(n4710), .A2(n4709), .ZN(n2222) );
  AOI22D1BWP12T U5650 ( .A1(n4742), .A2(write1_in[16]), .B1(n4741), .B2(
        write2_in[16]), .ZN(n4712) );
  AOI22D1BWP12T U5651 ( .A1(pc_out[16]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[16]), .ZN(n4711) );
  ND2D1BWP12T U5652 ( .A1(n4712), .A2(n4711), .ZN(n2217) );
  AOI22D1BWP12T U5653 ( .A1(n4742), .A2(write1_in[5]), .B1(n4741), .B2(
        write2_in[5]), .ZN(n4714) );
  AOI22D1BWP12T U5654 ( .A1(pc_out[5]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[5]), .ZN(n4713) );
  ND2D1BWP12T U5655 ( .A1(n4714), .A2(n4713), .ZN(n2206) );
  AOI22D1BWP12T U5656 ( .A1(n4742), .A2(write1_in[28]), .B1(n4741), .B2(
        write2_in[28]), .ZN(n4716) );
  AOI22D1BWP12T U5657 ( .A1(pc_out[28]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[28]), .ZN(n4715) );
  ND2D1BWP12T U5658 ( .A1(n4716), .A2(n4715), .ZN(n2229) );
  AOI22D1BWP12T U5659 ( .A1(n4742), .A2(write1_in[9]), .B1(n4741), .B2(
        write2_in[9]), .ZN(n4718) );
  AOI22D1BWP12T U5660 ( .A1(pc_out[9]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[9]), .ZN(n4717) );
  ND2D1BWP12T U5661 ( .A1(n4718), .A2(n4717), .ZN(n2210) );
  AOI22D1BWP12T U5662 ( .A1(n4742), .A2(write1_in[30]), .B1(n4741), .B2(
        write2_in[30]), .ZN(n4720) );
  AOI22D1BWP12T U5663 ( .A1(pc_out[30]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[30]), .ZN(n4719) );
  ND2D1BWP12T U5664 ( .A1(n4720), .A2(n4719), .ZN(n2231) );
  AOI22D1BWP12T U5665 ( .A1(n4742), .A2(write1_in[7]), .B1(n4741), .B2(
        write2_in[7]), .ZN(n4722) );
  AOI22D1BWP12T U5666 ( .A1(pc_out[7]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[7]), .ZN(n4721) );
  ND2D1BWP12T U5667 ( .A1(n4722), .A2(n4721), .ZN(n2208) );
  AOI22D1BWP12T U5668 ( .A1(n4742), .A2(write1_in[25]), .B1(n4741), .B2(
        write2_in[25]), .ZN(n4724) );
  AOI22D1BWP12T U5669 ( .A1(pc_out[25]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[25]), .ZN(n4723) );
  ND2D1BWP12T U5670 ( .A1(n4724), .A2(n4723), .ZN(n2226) );
  AOI22D1BWP12T U5671 ( .A1(n4742), .A2(write1_in[14]), .B1(n4741), .B2(
        write2_in[14]), .ZN(n4726) );
  AOI22D1BWP12T U5672 ( .A1(pc_out[14]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[14]), .ZN(n4725) );
  ND2D1BWP12T U5673 ( .A1(n4726), .A2(n4725), .ZN(n2215) );
  AOI22D1BWP12T U5674 ( .A1(n4742), .A2(write1_in[8]), .B1(n4741), .B2(
        write2_in[8]), .ZN(n4728) );
  AOI22D1BWP12T U5675 ( .A1(pc_out[8]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[8]), .ZN(n4727) );
  ND2D1BWP12T U5676 ( .A1(n4728), .A2(n4727), .ZN(n2209) );
  AOI22D1BWP12T U5677 ( .A1(n4742), .A2(write1_in[26]), .B1(n4741), .B2(
        write2_in[26]), .ZN(n4730) );
  AOI22D1BWP12T U5678 ( .A1(pc_out[26]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[26]), .ZN(n4729) );
  ND2D1BWP12T U5679 ( .A1(n4730), .A2(n4729), .ZN(n2227) );
  AOI22D1BWP12T U5680 ( .A1(n4742), .A2(write1_in[17]), .B1(n4741), .B2(
        write2_in[17]), .ZN(n4732) );
  AOI22D1BWP12T U5681 ( .A1(pc_out[17]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[17]), .ZN(n4731) );
  ND2D1BWP12T U5682 ( .A1(n4732), .A2(n4731), .ZN(n2218) );
  AOI22D1BWP12T U5683 ( .A1(n4742), .A2(write1_in[10]), .B1(n4741), .B2(
        write2_in[10]), .ZN(n4734) );
  AOI22D1BWP12T U5684 ( .A1(pc_out[10]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[10]), .ZN(n4733) );
  ND2D1BWP12T U5685 ( .A1(n4734), .A2(n4733), .ZN(n2211) );
  AOI22D1BWP12T U5686 ( .A1(n4742), .A2(write1_in[27]), .B1(n4741), .B2(
        write2_in[27]), .ZN(n4736) );
  AOI22D1BWP12T U5687 ( .A1(pc_out[27]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[27]), .ZN(n4735) );
  ND2D1BWP12T U5688 ( .A1(n4736), .A2(n4735), .ZN(n2228) );
  AOI22D1BWP12T U5689 ( .A1(n4742), .A2(write1_in[19]), .B1(n4741), .B2(
        write2_in[19]), .ZN(n4738) );
  AOI22D1BWP12T U5690 ( .A1(pc_out[19]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[19]), .ZN(n4737) );
  ND2D1BWP12T U5691 ( .A1(n4738), .A2(n4737), .ZN(n2220) );
  AOI22D1BWP12T U5692 ( .A1(n4742), .A2(write1_in[18]), .B1(n4741), .B2(
        write2_in[18]), .ZN(n4740) );
  AOI22D1BWP12T U5693 ( .A1(pc_out[18]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[18]), .ZN(n4739) );
  ND2D1BWP12T U5694 ( .A1(n4740), .A2(n4739), .ZN(n2219) );
  AOI22D1BWP12T U5695 ( .A1(n4742), .A2(write1_in[4]), .B1(n4741), .B2(
        write2_in[4]), .ZN(n4746) );
  AOI22D1BWP12T U5696 ( .A1(pc_out[4]), .A2(n4744), .B1(n4743), .B2(
        next_pc_in[4]), .ZN(n4745) );
  ND2D1BWP12T U5697 ( .A1(n4746), .A2(n4745), .ZN(n2205) );
  OAI222D1BWP12T U5698 ( .A1(n4751), .A2(n4790), .B1(n4750), .B2(n4747), .C1(
        n4749), .C2(n4789), .ZN(n2199) );
  OAI222D1BWP12T U5699 ( .A1(n4751), .A2(n4805), .B1(n4750), .B2(n4748), .C1(
        n4749), .C2(n4804), .ZN(n2194) );
  IND2XD1BWP12T U5700 ( .A1(n4754), .B1(n4771), .ZN(n4770) );
  IND2XD1BWP12T U5701 ( .A1(n4755), .B1(n4879), .ZN(n4877) );
  IND2XD1BWP12T U5702 ( .A1(n4760), .B1(n4842), .ZN(n4844) );
  IND2XD1BWP12T U5703 ( .A1(n4765), .B1(n4768), .ZN(n4767) );
  OAI222D1BWP12T U5704 ( .A1(n4826), .A2(n4837), .B1(n4825), .B2(n4824), .C1(
        n4823), .C2(n4835), .ZN(n2422) );
  OAI222D1BWP12T U5705 ( .A1(n4869), .A2(n4855), .B1(n4871), .B2(n4827), .C1(
        n4873), .C2(n4853), .ZN(n2242) );
  OAI222D1BWP12T U5706 ( .A1(n4875), .A2(n4831), .B1(n4877), .B2(n4828), .C1(
        n4879), .C2(n4829), .ZN(n2664) );
  OAI222D1BWP12T U5707 ( .A1(n4863), .A2(n4831), .B1(n4865), .B2(n4830), .C1(
        n4867), .C2(n4829), .ZN(n2280) );
  OAI222D1BWP12T U5708 ( .A1(n4875), .A2(n4834), .B1(n4877), .B2(n4833), .C1(
        n4879), .C2(n4832), .ZN(n2672) );
  OAI222D1BWP12T U5709 ( .A1(n4846), .A2(n4837), .B1(n4844), .B2(n4836), .C1(
        n4842), .C2(n4835), .ZN(n2646) );
  OAI222D1BWP12T U5710 ( .A1(n4875), .A2(n4840), .B1(n4877), .B2(n4839), .C1(
        n4879), .C2(n4838), .ZN(n2654) );
  OAI222D1BWP12T U5711 ( .A1(n4846), .A2(n4845), .B1(n4844), .B2(n4843), .C1(
        n4842), .C2(n4841), .ZN(n2641) );
  OAI222D1BWP12T U5712 ( .A1(n4875), .A2(n4849), .B1(n4877), .B2(n4848), .C1(
        n4879), .C2(n4847), .ZN(n2680) );
  OAI222D1BWP12T U5713 ( .A1(n4869), .A2(n4852), .B1(n4871), .B2(n4851), .C1(
        n4873), .C2(n4850), .ZN(n2245) );
  OAI222D1BWP12T U5714 ( .A1(n4875), .A2(n4855), .B1(n4877), .B2(n4854), .C1(
        n4879), .C2(n4853), .ZN(n2658) );
  OAI222D1BWP12T U5715 ( .A1(n4869), .A2(n4858), .B1(n4871), .B2(n4857), .C1(
        n4873), .C2(n4856), .ZN(n2246) );
  OAI222D1BWP12T U5716 ( .A1(n4867), .A2(n4861), .B1(n4865), .B2(n4860), .C1(
        n4863), .C2(n4859), .ZN(n2265) );
  OAI222D1BWP12T U5717 ( .A1(n4867), .A2(n4866), .B1(n4865), .B2(n4864), .C1(
        n4863), .C2(n4862), .ZN(n2267) );
  OAI222D1BWP12T U5718 ( .A1(n4873), .A2(n4872), .B1(n4871), .B2(n4870), .C1(
        n4869), .C2(n4868), .ZN(n2244) );
  OAI222D1BWP12T U5719 ( .A1(n4879), .A2(n4878), .B1(n4877), .B2(n4876), .C1(
        n4875), .C2(n4874), .ZN(n2665) );
  OAI222D1BWP12T U5720 ( .A1(n4885), .A2(n4884), .B1(n4883), .B2(n4882), .C1(
        n4881), .C2(n4880), .ZN(n2605) );
endmodule

