
module register_file ( readA_sel, readB_sel, readC_sel, readD_sel, write1_sel, 
        write2_sel, write1_en, write2_en, write1_in, write2_in, immediate1_in, 
        immediate2_in, next_pc_in, next_cpsr_in, next_sp_in, next_pc_en, clk, 
        regA_out, regB_out, regC_out, regD_out, pc_out, cpsr_out, sp_out );
  input [4:0] readA_sel;
  input [4:0] readB_sel;
  input [4:0] readC_sel;
  input [4:0] readD_sel;
  input [4:0] write1_sel;
  input [4:0] write2_sel;
  input [31:0] write1_in;
  input [31:0] write2_in;
  input [31:0] immediate1_in;
  input [31:0] immediate2_in;
  input [31:0] next_pc_in;
  input [3:0] next_cpsr_in;
  input [31:0] next_sp_in;
  input [31:0] next_pc_en;
  output [31:0] regA_out;
  output [31:0] regB_out;
  output [31:0] regC_out;
  output [31:0] regD_out;
  output [31:0] pc_out;
  output [3:0] cpsr_out;
  output [31:0] sp_out;
  input write1_en, write2_en, clk;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242,
         N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253,
         N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264,
         N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374,
         N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385,
         N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396,
         N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440,
         N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451,
         N452, N453, N454, N455, N456, pc_write_select, N457, N458, N459, N460,
         N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471,
         N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482,
         N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493,
         N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, N504,
         N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515,
         N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526,
         N527, N528, N529, N530, N531, N532, N533, N534, N535, N536, N537,
         N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, N548,
         N549, N550, N551, N552, N553, N554, N555, N556, N557, N558, N559,
         N560, N561, N562, N563, N564, N565, N566, N567, N568, N569, N570,
         N571, N572, N573, N574, N575, N576, N577, N578, N579, N580, N581,
         N582, N583, N584, N585, N586, N587, N588, N589, N590, N591, N592,
         N593, N594, N595, N596, N597, N598, N599, N600, N601, N602, N603,
         N604, N605, N606, N607, N608, N609, N610, N611, N612;
  wire   [31:0] r0;
  wire   [31:0] r1;
  wire   [31:0] r2;
  wire   [31:0] r3;
  wire   [31:0] r4;
  wire   [31:0] r5;
  wire   [31:0] r6;
  wire   [31:0] r7;
  wire   [31:0] r8;
  wire   [31:0] r9;
  wire   [31:0] r10;
  wire   [31:0] r11;
  wire   [31:0] r12;
  wire   [31:0] lr;
  wire   [31:0] tmp1;
  wire   [31:0] r0in;
  wire   [31:0] r1in;
  wire   [31:0] r2in;
  wire   [31:0] r3in;
  wire   [31:0] r4in;
  wire   [31:0] r5in;
  wire   [31:0] r6in;
  wire   [31:0] r7in;
  wire   [31:0] r8in;
  wire   [31:0] r9in;
  wire   [31:0] r10in;
  wire   [31:0] r11in;
  wire   [31:0] r12in;
  wire   [31:0] spin;
  wire   [31:0] lrin;
  wire   [31:0] pc_write_in;
  wire   [31:0] pcin;
  wire   [31:0] tmp1in;

  GTECH_AND2 C9 ( .A(N93), .B(N151), .Z(N95) );
  GTECH_AND2 C10 ( .A(N153), .B(N155), .Z(N96) );
  GTECH_AND2 C11 ( .A(N95), .B(N96), .Z(N97) );
  GTECH_AND2 C12 ( .A(N97), .B(N94), .Z(N98) );
  GTECH_OR2 C14 ( .A(readA_sel[4]), .B(readA_sel[3]), .Z(N99) );
  GTECH_OR2 C15 ( .A(readA_sel[2]), .B(readA_sel[1]), .Z(N100) );
  GTECH_OR2 C16 ( .A(N99), .B(N100), .Z(N101) );
  GTECH_OR2 C17 ( .A(N101), .B(N94), .Z(N102) );
  GTECH_OR2 C21 ( .A(readA_sel[2]), .B(N155), .Z(N104) );
  GTECH_OR2 C22 ( .A(N99), .B(N104), .Z(N105) );
  GTECH_OR2 C23 ( .A(N105), .B(readA_sel[0]), .Z(N106) );
  GTECH_OR2 C30 ( .A(N105), .B(N94), .Z(N108) );
  GTECH_OR2 C34 ( .A(N153), .B(readA_sel[1]), .Z(N110) );
  GTECH_OR2 C35 ( .A(N99), .B(N110), .Z(N111) );
  GTECH_OR2 C36 ( .A(N111), .B(readA_sel[0]), .Z(N112) );
  GTECH_OR2 C43 ( .A(N111), .B(N94), .Z(N114) );
  GTECH_OR2 C48 ( .A(N153), .B(N155), .Z(N116) );
  GTECH_OR2 C49 ( .A(N99), .B(N116), .Z(N117) );
  GTECH_OR2 C50 ( .A(N117), .B(readA_sel[0]), .Z(N118) );
  GTECH_OR2 C58 ( .A(N117), .B(N94), .Z(N120) );
  GTECH_OR2 C61 ( .A(readA_sel[4]), .B(N151), .Z(N122) );
  GTECH_OR2 C63 ( .A(N122), .B(N100), .Z(N123) );
  GTECH_OR2 C64 ( .A(N123), .B(readA_sel[0]), .Z(N124) );
  GTECH_OR2 C71 ( .A(N123), .B(N94), .Z(N126) );
  GTECH_OR2 C77 ( .A(N122), .B(N104), .Z(N128) );
  GTECH_OR2 C78 ( .A(N128), .B(readA_sel[0]), .Z(N129) );
  GTECH_OR2 C86 ( .A(N128), .B(N94), .Z(N131) );
  GTECH_OR2 C92 ( .A(N122), .B(N110), .Z(N133) );
  GTECH_OR2 C93 ( .A(N133), .B(readA_sel[0]), .Z(N134) );
  GTECH_OR2 C101 ( .A(N133), .B(N94), .Z(N136) );
  GTECH_OR2 C108 ( .A(N122), .B(N116), .Z(N138) );
  GTECH_OR2 C109 ( .A(N138), .B(readA_sel[0]), .Z(N139) );
  GTECH_OR2 C118 ( .A(N138), .B(N94), .Z(N141) );
  GTECH_OR2 C124 ( .A(N93), .B(N151), .Z(N143) );
  GTECH_OR2 C126 ( .A(N143), .B(N116), .Z(N144) );
  GTECH_OR2 C127 ( .A(N144), .B(readA_sel[0]), .Z(N145) );
  GTECH_AND2 C129 ( .A(readA_sel[4]), .B(readA_sel[3]), .Z(N147) );
  GTECH_AND2 C130 ( .A(readA_sel[2]), .B(readA_sel[1]), .Z(N148) );
  GTECH_AND2 C131 ( .A(N147), .B(N148), .Z(N149) );
  GTECH_AND2 C132 ( .A(N149), .B(readA_sel[0]), .Z(N150) );
  GTECH_AND2 C134 ( .A(readA_sel[4]), .B(N151), .Z(N152) );
  GTECH_AND2 C136 ( .A(readA_sel[4]), .B(N153), .Z(N154) );
  GTECH_AND2 C138 ( .A(readA_sel[4]), .B(N155), .Z(N156) );
  GTECH_AND2 C215 ( .A(N158), .B(N216), .Z(N160) );
  GTECH_AND2 C216 ( .A(N218), .B(N220), .Z(N161) );
  GTECH_AND2 C217 ( .A(N160), .B(N161), .Z(N162) );
  GTECH_AND2 C218 ( .A(N162), .B(N159), .Z(N163) );
  GTECH_OR2 C220 ( .A(readB_sel[4]), .B(readB_sel[3]), .Z(N164) );
  GTECH_OR2 C221 ( .A(readB_sel[2]), .B(readB_sel[1]), .Z(N165) );
  GTECH_OR2 C222 ( .A(N164), .B(N165), .Z(N166) );
  GTECH_OR2 C223 ( .A(N166), .B(N159), .Z(N167) );
  GTECH_OR2 C227 ( .A(readB_sel[2]), .B(N220), .Z(N169) );
  GTECH_OR2 C228 ( .A(N164), .B(N169), .Z(N170) );
  GTECH_OR2 C229 ( .A(N170), .B(readB_sel[0]), .Z(N171) );
  GTECH_OR2 C236 ( .A(N170), .B(N159), .Z(N173) );
  GTECH_OR2 C240 ( .A(N218), .B(readB_sel[1]), .Z(N175) );
  GTECH_OR2 C241 ( .A(N164), .B(N175), .Z(N176) );
  GTECH_OR2 C242 ( .A(N176), .B(readB_sel[0]), .Z(N177) );
  GTECH_OR2 C249 ( .A(N176), .B(N159), .Z(N179) );
  GTECH_OR2 C254 ( .A(N218), .B(N220), .Z(N181) );
  GTECH_OR2 C255 ( .A(N164), .B(N181), .Z(N182) );
  GTECH_OR2 C256 ( .A(N182), .B(readB_sel[0]), .Z(N183) );
  GTECH_OR2 C264 ( .A(N182), .B(N159), .Z(N185) );
  GTECH_OR2 C267 ( .A(readB_sel[4]), .B(N216), .Z(N187) );
  GTECH_OR2 C269 ( .A(N187), .B(N165), .Z(N188) );
  GTECH_OR2 C270 ( .A(N188), .B(readB_sel[0]), .Z(N189) );
  GTECH_OR2 C277 ( .A(N188), .B(N159), .Z(N191) );
  GTECH_OR2 C283 ( .A(N187), .B(N169), .Z(N193) );
  GTECH_OR2 C284 ( .A(N193), .B(readB_sel[0]), .Z(N194) );
  GTECH_OR2 C292 ( .A(N193), .B(N159), .Z(N196) );
  GTECH_OR2 C298 ( .A(N187), .B(N175), .Z(N198) );
  GTECH_OR2 C299 ( .A(N198), .B(readB_sel[0]), .Z(N199) );
  GTECH_OR2 C307 ( .A(N198), .B(N159), .Z(N201) );
  GTECH_OR2 C314 ( .A(N187), .B(N181), .Z(N203) );
  GTECH_OR2 C315 ( .A(N203), .B(readB_sel[0]), .Z(N204) );
  GTECH_OR2 C324 ( .A(N203), .B(N159), .Z(N206) );
  GTECH_OR2 C330 ( .A(N158), .B(N216), .Z(N208) );
  GTECH_OR2 C332 ( .A(N208), .B(N181), .Z(N209) );
  GTECH_OR2 C333 ( .A(N209), .B(readB_sel[0]), .Z(N210) );
  GTECH_AND2 C335 ( .A(readB_sel[4]), .B(readB_sel[3]), .Z(N212) );
  GTECH_AND2 C336 ( .A(readB_sel[2]), .B(readB_sel[1]), .Z(N213) );
  GTECH_AND2 C337 ( .A(N212), .B(N213), .Z(N214) );
  GTECH_AND2 C338 ( .A(N214), .B(readB_sel[0]), .Z(N215) );
  GTECH_AND2 C340 ( .A(readB_sel[4]), .B(N216), .Z(N217) );
  GTECH_AND2 C342 ( .A(readB_sel[4]), .B(N218), .Z(N219) );
  GTECH_AND2 C344 ( .A(readB_sel[4]), .B(N220), .Z(N221) );
  GTECH_AND2 C424 ( .A(N224), .B(N225), .Z(N228) );
  GTECH_AND2 C425 ( .A(N226), .B(N227), .Z(N229) );
  GTECH_AND2 C426 ( .A(N228), .B(N229), .Z(N230) );
  GTECH_OR2 C428 ( .A(readC_sel[3]), .B(readC_sel[2]), .Z(N231) );
  GTECH_OR2 C429 ( .A(readC_sel[1]), .B(N227), .Z(N232) );
  GTECH_OR2 C430 ( .A(N231), .B(N232), .Z(N233) );
  GTECH_OR2 C434 ( .A(N226), .B(readC_sel[0]), .Z(N235) );
  GTECH_OR2 C435 ( .A(N231), .B(N235), .Z(N236) );
  GTECH_OR2 C440 ( .A(N226), .B(N227), .Z(N238) );
  GTECH_OR2 C441 ( .A(N231), .B(N238), .Z(N239) );
  GTECH_OR2 C444 ( .A(readC_sel[3]), .B(N225), .Z(N241) );
  GTECH_OR2 C445 ( .A(readC_sel[1]), .B(readC_sel[0]), .Z(N242) );
  GTECH_OR2 C446 ( .A(N241), .B(N242), .Z(N243) );
  GTECH_OR2 C452 ( .A(N241), .B(N232), .Z(N245) );
  GTECH_OR2 C458 ( .A(N241), .B(N235), .Z(N247) );
  GTECH_OR2 C465 ( .A(N241), .B(N238), .Z(N249) );
  GTECH_OR2 C468 ( .A(N224), .B(readC_sel[2]), .Z(N251) );
  GTECH_OR2 C470 ( .A(N251), .B(N242), .Z(N252) );
  GTECH_OR2 C476 ( .A(N251), .B(N232), .Z(N254) );
  GTECH_OR2 C482 ( .A(N251), .B(N235), .Z(N256) );
  GTECH_OR2 C489 ( .A(N251), .B(N238), .Z(N258) );
  GTECH_OR2 C493 ( .A(N224), .B(N225), .Z(N260) );
  GTECH_OR2 C495 ( .A(N260), .B(N242), .Z(N261) );
  GTECH_OR2 C502 ( .A(N260), .B(N232), .Z(N263) );
  GTECH_OR2 C509 ( .A(N260), .B(N235), .Z(N265) );
  GTECH_AND2 C511 ( .A(readC_sel[3]), .B(readC_sel[2]), .Z(N267) );
  GTECH_AND2 C512 ( .A(readC_sel[1]), .B(readC_sel[0]), .Z(N268) );
  GTECH_AND2 C513 ( .A(N267), .B(N268), .Z(N269) );
  GTECH_AND2 C619 ( .A(N303), .B(N304), .Z(N307) );
  GTECH_AND2 C620 ( .A(N305), .B(N306), .Z(N308) );
  GTECH_AND2 C621 ( .A(N307), .B(N308), .Z(N309) );
  GTECH_OR2 C623 ( .A(readD_sel[3]), .B(readD_sel[2]), .Z(N310) );
  GTECH_OR2 C624 ( .A(readD_sel[1]), .B(N306), .Z(N311) );
  GTECH_OR2 C625 ( .A(N310), .B(N311), .Z(N312) );
  GTECH_OR2 C629 ( .A(N305), .B(readD_sel[0]), .Z(N314) );
  GTECH_OR2 C630 ( .A(N310), .B(N314), .Z(N315) );
  GTECH_OR2 C635 ( .A(N305), .B(N306), .Z(N317) );
  GTECH_OR2 C636 ( .A(N310), .B(N317), .Z(N318) );
  GTECH_OR2 C639 ( .A(readD_sel[3]), .B(N304), .Z(N320) );
  GTECH_OR2 C640 ( .A(readD_sel[1]), .B(readD_sel[0]), .Z(N321) );
  GTECH_OR2 C641 ( .A(N320), .B(N321), .Z(N322) );
  GTECH_OR2 C647 ( .A(N320), .B(N311), .Z(N324) );
  GTECH_OR2 C653 ( .A(N320), .B(N314), .Z(N326) );
  GTECH_OR2 C660 ( .A(N320), .B(N317), .Z(N328) );
  GTECH_OR2 C663 ( .A(N303), .B(readD_sel[2]), .Z(N330) );
  GTECH_OR2 C665 ( .A(N330), .B(N321), .Z(N331) );
  GTECH_OR2 C671 ( .A(N330), .B(N311), .Z(N333) );
  GTECH_OR2 C677 ( .A(N330), .B(N314), .Z(N335) );
  GTECH_OR2 C684 ( .A(N330), .B(N317), .Z(N337) );
  GTECH_OR2 C688 ( .A(N303), .B(N304), .Z(N339) );
  GTECH_OR2 C690 ( .A(N339), .B(N321), .Z(N340) );
  GTECH_OR2 C697 ( .A(N339), .B(N311), .Z(N342) );
  GTECH_OR2 C704 ( .A(N339), .B(N314), .Z(N344) );
  GTECH_AND2 C706 ( .A(readD_sel[3]), .B(readD_sel[2]), .Z(N346) );
  GTECH_AND2 C707 ( .A(readD_sel[1]), .B(readD_sel[0]), .Z(N347) );
  GTECH_AND2 C708 ( .A(N346), .B(N347), .Z(N348) );
  \**SEQGEN**  r0_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[31]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[30]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[29]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[28]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[27]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[26]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[25]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[24]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[23]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[22]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[21]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[20]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[19]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[18]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[17]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[16]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[15]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[14]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[13]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[12]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[11]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[10]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r0_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(r0in[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r0[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N383) );
  \**SEQGEN**  r1_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[31]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[30]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[29]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[28]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[27]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[26]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[25]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[24]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[23]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[22]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[21]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[20]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[19]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[18]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[17]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[16]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[15]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[14]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[13]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[12]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[11]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[10]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r1_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(r1in[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r1[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N388) );
  \**SEQGEN**  r2_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[31]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[30]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[29]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[28]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[27]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[26]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[25]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[24]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[23]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[22]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[21]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[20]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[19]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[18]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[17]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[16]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[15]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[14]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[13]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[12]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[11]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[10]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r2_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(r2in[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r2[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N393) );
  \**SEQGEN**  r3_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[31]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[30]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[29]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[28]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[27]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[26]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[25]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[24]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[23]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[22]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[21]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[20]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[19]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[18]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[17]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[16]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[15]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[14]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[13]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[12]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[11]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[10]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r3_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(r3in[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r3[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N397) );
  \**SEQGEN**  r4_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[31]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[30]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[29]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[28]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[27]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[26]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[25]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[24]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[23]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[22]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[21]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[20]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[19]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[18]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[17]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[16]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[15]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[14]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[13]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[12]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[11]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[10]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r4_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(r4in[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r4[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N402) );
  \**SEQGEN**  r5_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[31]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[30]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[29]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[28]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[27]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[26]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[25]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[24]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[23]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[22]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[21]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[20]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[19]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[18]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[17]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[16]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[15]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[14]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[13]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[12]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[11]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[10]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r5_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(r5in[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r5[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N407) );
  \**SEQGEN**  r6_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[31]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[30]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[29]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[28]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[27]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[26]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[25]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[24]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[23]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[22]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[21]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[20]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[19]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[18]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[17]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[16]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[15]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[14]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[13]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[12]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[11]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[10]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r6_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(r6in[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r6[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N412) );
  \**SEQGEN**  r7_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[31]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[30]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[29]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[28]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[27]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[26]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[25]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[24]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[23]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[22]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[21]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[20]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[19]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[18]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[17]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[16]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[15]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[14]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[13]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[12]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[11]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[10]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r7_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(r7in[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r7[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  r8_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[31]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[30]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[29]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[28]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[27]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[26]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[25]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[24]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[23]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[22]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[21]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[20]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[19]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[18]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[17]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[16]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[15]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[14]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[13]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[12]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[11]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[10]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r8_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(r8in[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r8[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N423) );
  \**SEQGEN**  r9_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[31]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[30]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[29]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[28]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[27]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[26]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[25]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[24]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[23]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[22]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[21]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[20]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[19]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[18]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[17]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[16]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[15]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[14]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[13]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[12]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[11]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[10]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r9_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(r9in[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r9[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N428) );
  \**SEQGEN**  r10_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r10in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r10[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(r10in[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r10[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(r10in[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r10[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(r10in[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r10[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(r10in[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r10[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(r10in[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r10[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(r10in[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r10[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(r10in[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r10[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(r10in[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r10[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(r10in[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r10[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r10_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(r10in[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r10[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N433) );
  \**SEQGEN**  r11_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r11in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r11[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(r11in[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r11[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(r11in[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r11[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(r11in[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r11[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(r11in[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r11[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(r11in[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r11[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(r11in[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r11[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(r11in[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r11[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(r11in[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r11[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(r11in[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r11[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r11_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(r11in[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r11[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N438) );
  \**SEQGEN**  r12_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        r12in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        r12[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(r12in[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r12[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(r12in[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r12[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(r12in[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r12[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(r12in[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r12[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(r12in[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r12[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(r12in[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r12[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(r12in[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r12[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(r12in[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r12[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(r12in[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r12[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  r12_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(r12in[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(r12[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N443) );
  \**SEQGEN**  lr_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[31]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[30]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[29]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[28]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[27]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[26]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[25]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[24]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[23]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[22]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[21]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[20]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[19]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[18]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[17]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[16]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[15]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[14]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[13]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[12]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[11]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[10]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  lr_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(lrin[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(lr[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N454) );
  \**SEQGEN**  sp_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[31]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[30]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[29]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[28]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[27]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[26]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[25]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[24]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[23]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[22]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[21]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[20]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[19]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[18]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[17]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[16]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[15]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[14]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[13]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[12]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[11]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[10]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  sp_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(spin[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(sp_out[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  pc_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[31]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[30]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[29]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[28]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[27]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[26]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[25]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[24]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[23]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[22]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[21]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[20]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[19]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[18]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[17]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[16]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[15]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[14]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[13]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[12]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[11]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[10]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  pc_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(pcin[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(pc_out[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N468) );
  \**SEQGEN**  cpsr_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        next_cpsr_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        cpsr_out[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  cpsr_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        next_cpsr_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        cpsr_out[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  cpsr_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        next_cpsr_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        cpsr_out[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  cpsr_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        next_cpsr_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        cpsr_out[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  tmp1_reg_31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N464) );
  \**SEQGEN**  tmp1_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        tmp1in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        tmp1[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N464) );
  GTECH_OR2 C2169 ( .A(write2_sel[3]), .B(write2_sel[4]), .Z(N469) );
  GTECH_OR2 C2170 ( .A(write2_sel[2]), .B(N469), .Z(N470) );
  GTECH_OR2 C2171 ( .A(write2_sel[1]), .B(N470), .Z(N471) );
  GTECH_OR2 C2172 ( .A(write2_sel[0]), .B(N471), .Z(N472) );
  GTECH_NOT I_0 ( .A(N472), .Z(N473) );
  GTECH_OR2 C2174 ( .A(write1_sel[3]), .B(write1_sel[4]), .Z(N474) );
  GTECH_OR2 C2175 ( .A(write1_sel[2]), .B(N474), .Z(N475) );
  GTECH_OR2 C2176 ( .A(write1_sel[1]), .B(N475), .Z(N476) );
  GTECH_OR2 C2177 ( .A(write1_sel[0]), .B(N476), .Z(N477) );
  GTECH_NOT I_1 ( .A(N477), .Z(N478) );
  GTECH_NOT I_2 ( .A(write2_sel[0]), .Z(N479) );
  GTECH_OR2 C2183 ( .A(N479), .B(N471), .Z(N480) );
  GTECH_NOT I_3 ( .A(N480), .Z(N481) );
  GTECH_NOT I_4 ( .A(write1_sel[0]), .Z(N482) );
  GTECH_OR2 C2189 ( .A(N482), .B(N476), .Z(N483) );
  GTECH_NOT I_5 ( .A(N483), .Z(N484) );
  GTECH_NOT I_6 ( .A(write2_sel[1]), .Z(N485) );
  GTECH_OR2 C2194 ( .A(N485), .B(N470), .Z(N486) );
  GTECH_OR2 C2195 ( .A(write2_sel[0]), .B(N486), .Z(N487) );
  GTECH_NOT I_7 ( .A(N487), .Z(N488) );
  GTECH_NOT I_8 ( .A(write1_sel[1]), .Z(N489) );
  GTECH_OR2 C2200 ( .A(N489), .B(N475), .Z(N490) );
  GTECH_OR2 C2201 ( .A(write1_sel[0]), .B(N490), .Z(N491) );
  GTECH_NOT I_9 ( .A(N491), .Z(N492) );
  GTECH_OR2 C2214 ( .A(N482), .B(N490), .Z(N493) );
  GTECH_NOT I_10 ( .A(N493), .Z(N494) );
  GTECH_NOT I_11 ( .A(write2_sel[2]), .Z(N495) );
  GTECH_OR2 C2218 ( .A(N495), .B(N469), .Z(N496) );
  GTECH_OR2 C2219 ( .A(write2_sel[1]), .B(N496), .Z(N497) );
  GTECH_OR2 C2220 ( .A(write2_sel[0]), .B(N497), .Z(N498) );
  GTECH_NOT I_12 ( .A(N498), .Z(N499) );
  GTECH_NOT I_13 ( .A(write1_sel[2]), .Z(N500) );
  GTECH_OR2 C2224 ( .A(N500), .B(N474), .Z(N501) );
  GTECH_OR2 C2225 ( .A(write1_sel[1]), .B(N501), .Z(N502) );
  GTECH_OR2 C2226 ( .A(write1_sel[0]), .B(N502), .Z(N503) );
  GTECH_NOT I_14 ( .A(N503), .Z(N504) );
  GTECH_OR2 C2233 ( .A(N479), .B(N497), .Z(N505) );
  GTECH_NOT I_15 ( .A(N505), .Z(N506) );
  GTECH_OR2 C2240 ( .A(N482), .B(N502), .Z(N507) );
  GTECH_NOT I_16 ( .A(N507), .Z(N508) );
  GTECH_OR2 C2246 ( .A(N485), .B(N496), .Z(N509) );
  GTECH_OR2 C2247 ( .A(write2_sel[0]), .B(N509), .Z(N510) );
  GTECH_NOT I_17 ( .A(N510), .Z(N511) );
  GTECH_OR2 C2253 ( .A(N489), .B(N501), .Z(N512) );
  GTECH_OR2 C2254 ( .A(write1_sel[0]), .B(N512), .Z(N513) );
  GTECH_NOT I_18 ( .A(N513), .Z(N514) );
  GTECH_OR2 C2262 ( .A(N479), .B(N509), .Z(N515) );
  GTECH_NOT I_19 ( .A(N515), .Z(N516) );
  GTECH_OR2 C2270 ( .A(N482), .B(N512), .Z(N517) );
  GTECH_NOT I_20 ( .A(N517), .Z(N518) );
  GTECH_NOT I_21 ( .A(write2_sel[3]), .Z(N519) );
  GTECH_OR2 C2273 ( .A(N519), .B(write2_sel[4]), .Z(N520) );
  GTECH_OR2 C2274 ( .A(write2_sel[2]), .B(N520), .Z(N521) );
  GTECH_OR2 C2275 ( .A(write2_sel[1]), .B(N521), .Z(N522) );
  GTECH_OR2 C2276 ( .A(write2_sel[0]), .B(N522), .Z(N523) );
  GTECH_NOT I_22 ( .A(N523), .Z(N524) );
  GTECH_NOT I_23 ( .A(write1_sel[3]), .Z(N525) );
  GTECH_OR2 C2279 ( .A(N525), .B(write1_sel[4]), .Z(N526) );
  GTECH_OR2 C2280 ( .A(write1_sel[2]), .B(N526), .Z(N527) );
  GTECH_OR2 C2281 ( .A(write1_sel[1]), .B(N527), .Z(N528) );
  GTECH_OR2 C2282 ( .A(write1_sel[0]), .B(N528), .Z(N529) );
  GTECH_NOT I_24 ( .A(N529), .Z(N530) );
  GTECH_OR2 C2289 ( .A(N479), .B(N522), .Z(N531) );
  GTECH_NOT I_25 ( .A(N531), .Z(N532) );
  GTECH_OR2 C2296 ( .A(N482), .B(N528), .Z(N533) );
  GTECH_NOT I_26 ( .A(N533), .Z(N534) );
  GTECH_OR2 C2302 ( .A(N485), .B(N521), .Z(N535) );
  GTECH_OR2 C2303 ( .A(write2_sel[0]), .B(N535), .Z(N536) );
  GTECH_NOT I_27 ( .A(N536), .Z(N537) );
  GTECH_OR2 C2309 ( .A(N489), .B(N527), .Z(N538) );
  GTECH_OR2 C2310 ( .A(write1_sel[0]), .B(N538), .Z(N539) );
  GTECH_NOT I_28 ( .A(N539), .Z(N540) );
  GTECH_OR2 C2318 ( .A(N479), .B(N535), .Z(N541) );
  GTECH_NOT I_29 ( .A(N541), .Z(N542) );
  GTECH_OR2 C2326 ( .A(N482), .B(N538), .Z(N543) );
  GTECH_NOT I_30 ( .A(N543), .Z(N544) );
  GTECH_OR2 C2331 ( .A(N495), .B(N520), .Z(N545) );
  GTECH_OR2 C2332 ( .A(write2_sel[1]), .B(N545), .Z(N546) );
  GTECH_OR2 C2333 ( .A(write2_sel[0]), .B(N546), .Z(N547) );
  GTECH_NOT I_31 ( .A(N547), .Z(N548) );
  GTECH_OR2 C2338 ( .A(N500), .B(N526), .Z(N549) );
  GTECH_OR2 C2339 ( .A(write1_sel[1]), .B(N549), .Z(N550) );
  GTECH_OR2 C2340 ( .A(write1_sel[0]), .B(N550), .Z(N551) );
  GTECH_NOT I_32 ( .A(N551), .Z(N552) );
  GTECH_OR2 C2347 ( .A(N485), .B(N545), .Z(N553) );
  GTECH_OR2 C2348 ( .A(write2_sel[0]), .B(N553), .Z(N554) );
  GTECH_NOT I_33 ( .A(N554), .Z(N555) );
  GTECH_OR2 C2355 ( .A(N489), .B(N549), .Z(N556) );
  GTECH_OR2 C2356 ( .A(write1_sel[0]), .B(N556), .Z(N557) );
  GTECH_NOT I_34 ( .A(N557), .Z(N558) );
  GTECH_OR2 C2364 ( .A(N479), .B(N546), .Z(N559) );
  GTECH_NOT I_35 ( .A(N559), .Z(N560) );
  GTECH_OR2 C2372 ( .A(N482), .B(N550), .Z(N561) );
  GTECH_NOT I_36 ( .A(N561), .Z(N562) );
  GTECH_OR2 C2381 ( .A(N482), .B(N556), .Z(N563) );
  GTECH_NOT I_37 ( .A(N563), .Z(N564) );
  GTECH_OR2 C2390 ( .A(N479), .B(N553), .Z(N565) );
  GTECH_NOT I_38 ( .A(N565), .Z(N566) );
  GTECH_NOT I_39 ( .A(write2_sel[4]), .Z(N567) );
  GTECH_OR2 C2405 ( .A(N519), .B(N567), .Z(N568) );
  GTECH_OR2 C2406 ( .A(N495), .B(N568), .Z(N569) );
  GTECH_OR2 C2407 ( .A(N485), .B(N569), .Z(N570) );
  GTECH_OR2 C2408 ( .A(write2_sel[0]), .B(N570), .Z(N571) );
  GTECH_NOT I_40 ( .A(N571), .Z(N572) );
  GTECH_NOT I_41 ( .A(write1_sel[4]), .Z(N573) );
  GTECH_OR2 C2414 ( .A(N525), .B(N573), .Z(N574) );
  GTECH_OR2 C2415 ( .A(N500), .B(N574), .Z(N575) );
  GTECH_OR2 C2416 ( .A(N489), .B(N575), .Z(N576) );
  GTECH_OR2 C2417 ( .A(write1_sel[0]), .B(N576), .Z(N577) );
  GTECH_NOT I_42 ( .A(N577), .Z(N578) );
  SELECT_OP C2867 ( .DATA1(r0), .DATA2(r1), .DATA3(r2), .DATA4(r3), .DATA5(r4), 
        .DATA6(r5), .DATA7(r6), .DATA8(r7), .DATA9(r8), .DATA10(r9), .DATA11(
        r10), .DATA12(r11), .DATA13(r12), .DATA14(sp_out), .DATA15(lr), 
        .DATA16(pc_out), .DATA17(tmp1), .DATA18(immediate1_in), .DATA19({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CONTROL1(N0), .CONTROL2(
        N1), .CONTROL3(N2), .CONTROL4(N3), .CONTROL5(N4), .CONTROL6(N5), 
        .CONTROL7(N6), .CONTROL8(N7), .CONTROL9(N8), .CONTROL10(N9), 
        .CONTROL11(N10), .CONTROL12(N11), .CONTROL13(N12), .CONTROL14(N13), 
        .CONTROL15(N14), .CONTROL16(N15), .CONTROL17(N16), .CONTROL18(N17), 
        .CONTROL19(N18), .Z(regA_out) );
  GTECH_BUF B_0 ( .A(N98), .Z(N0) );
  GTECH_BUF B_1 ( .A(N103), .Z(N1) );
  GTECH_BUF B_2 ( .A(N107), .Z(N2) );
  GTECH_BUF B_3 ( .A(N109), .Z(N3) );
  GTECH_BUF B_4 ( .A(N113), .Z(N4) );
  GTECH_BUF B_5 ( .A(N115), .Z(N5) );
  GTECH_BUF B_6 ( .A(N119), .Z(N6) );
  GTECH_BUF B_7 ( .A(N121), .Z(N7) );
  GTECH_BUF B_8 ( .A(N125), .Z(N8) );
  GTECH_BUF B_9 ( .A(N127), .Z(N9) );
  GTECH_BUF B_10 ( .A(N130), .Z(N10) );
  GTECH_BUF B_11 ( .A(N132), .Z(N11) );
  GTECH_BUF B_12 ( .A(N135), .Z(N12) );
  GTECH_BUF B_13 ( .A(N137), .Z(N13) );
  GTECH_BUF B_14 ( .A(N140), .Z(N14) );
  GTECH_BUF B_15 ( .A(N142), .Z(N15) );
  GTECH_BUF B_16 ( .A(N146), .Z(N16) );
  GTECH_BUF B_17 ( .A(N150), .Z(N17) );
  GTECH_BUF B_18 ( .A(N157), .Z(N18) );
  SELECT_OP C2868 ( .DATA1(r0), .DATA2(r1), .DATA3(r2), .DATA4(r3), .DATA5(r4), 
        .DATA6(r5), .DATA7(r6), .DATA8(r7), .DATA9(r8), .DATA10(r9), .DATA11(
        r10), .DATA12(r11), .DATA13(r12), .DATA14(sp_out), .DATA15(lr), 
        .DATA16(pc_out), .DATA17(tmp1), .DATA18(immediate2_in), .DATA19({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CONTROL1(N19), .CONTROL2(
        N20), .CONTROL3(N21), .CONTROL4(N22), .CONTROL5(N23), .CONTROL6(N24), 
        .CONTROL7(N25), .CONTROL8(N26), .CONTROL9(N27), .CONTROL10(N28), 
        .CONTROL11(N29), .CONTROL12(N30), .CONTROL13(N31), .CONTROL14(N32), 
        .CONTROL15(N33), .CONTROL16(N34), .CONTROL17(N35), .CONTROL18(N36), 
        .CONTROL19(N37), .Z(regB_out) );
  GTECH_BUF B_19 ( .A(N163), .Z(N19) );
  GTECH_BUF B_20 ( .A(N168), .Z(N20) );
  GTECH_BUF B_21 ( .A(N172), .Z(N21) );
  GTECH_BUF B_22 ( .A(N174), .Z(N22) );
  GTECH_BUF B_23 ( .A(N178), .Z(N23) );
  GTECH_BUF B_24 ( .A(N180), .Z(N24) );
  GTECH_BUF B_25 ( .A(N184), .Z(N25) );
  GTECH_BUF B_26 ( .A(N186), .Z(N26) );
  GTECH_BUF B_27 ( .A(N190), .Z(N27) );
  GTECH_BUF B_28 ( .A(N192), .Z(N28) );
  GTECH_BUF B_29 ( .A(N195), .Z(N29) );
  GTECH_BUF B_30 ( .A(N197), .Z(N30) );
  GTECH_BUF B_31 ( .A(N200), .Z(N31) );
  GTECH_BUF B_32 ( .A(N202), .Z(N32) );
  GTECH_BUF B_33 ( .A(N205), .Z(N33) );
  GTECH_BUF B_34 ( .A(N207), .Z(N34) );
  GTECH_BUF B_35 ( .A(N211), .Z(N35) );
  GTECH_BUF B_36 ( .A(N215), .Z(N36) );
  GTECH_BUF B_37 ( .A(N222), .Z(N37) );
  SELECT_OP C2869 ( .DATA1(r0), .DATA2(r1), .DATA3(r2), .DATA4(r3), .DATA5(r4), 
        .DATA6(r5), .DATA7(r6), .DATA8(r7), .DATA9(r8), .DATA10(r9), .DATA11(
        r10), .DATA12(r11), .DATA13(r12), .DATA14(sp_out), .DATA15(lr), 
        .DATA16(pc_out), .CONTROL1(N38), .CONTROL2(N39), .CONTROL3(N40), 
        .CONTROL4(N41), .CONTROL5(N42), .CONTROL6(N43), .CONTROL7(N44), 
        .CONTROL8(N45), .CONTROL9(N46), .CONTROL10(N47), .CONTROL11(N48), 
        .CONTROL12(N49), .CONTROL13(N50), .CONTROL14(N51), .CONTROL15(N52), 
        .CONTROL16(N53), .Z({N301, N300, N299, N298, N297, N296, N295, N294, 
        N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, 
        N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270}) );
  GTECH_BUF B_38 ( .A(N230), .Z(N38) );
  GTECH_BUF B_39 ( .A(N234), .Z(N39) );
  GTECH_BUF B_40 ( .A(N237), .Z(N40) );
  GTECH_BUF B_41 ( .A(N240), .Z(N41) );
  GTECH_BUF B_42 ( .A(N244), .Z(N42) );
  GTECH_BUF B_43 ( .A(N246), .Z(N43) );
  GTECH_BUF B_44 ( .A(N248), .Z(N44) );
  GTECH_BUF B_45 ( .A(N250), .Z(N45) );
  GTECH_BUF B_46 ( .A(N253), .Z(N46) );
  GTECH_BUF B_47 ( .A(N255), .Z(N47) );
  GTECH_BUF B_48 ( .A(N257), .Z(N48) );
  GTECH_BUF B_49 ( .A(N259), .Z(N49) );
  GTECH_BUF B_50 ( .A(N262), .Z(N50) );
  GTECH_BUF B_51 ( .A(N264), .Z(N51) );
  GTECH_BUF B_52 ( .A(N266), .Z(N52) );
  GTECH_BUF B_53 ( .A(N269), .Z(N53) );
  SELECT_OP C2870 ( .DATA1({N301, N300, N299, N298, N297, N296, N295, N294, 
        N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, 
        N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270}), .DATA2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CONTROL1(N54), 
        .CONTROL2(N55), .Z(regC_out) );
  GTECH_BUF B_54 ( .A(N223), .Z(N54) );
  GTECH_BUF B_55 ( .A(readC_sel[4]), .Z(N55) );
  SELECT_OP C2871 ( .DATA1(r0), .DATA2(r1), .DATA3(r2), .DATA4(r3), .DATA5(r4), 
        .DATA6(r5), .DATA7(r6), .DATA8(r7), .DATA9(r8), .DATA10(r9), .DATA11(
        r10), .DATA12(r11), .DATA13(r12), .DATA14(sp_out), .DATA15(lr), 
        .DATA16(pc_out), .CONTROL1(N56), .CONTROL2(N57), .CONTROL3(N58), 
        .CONTROL4(N59), .CONTROL5(N60), .CONTROL6(N61), .CONTROL7(N62), 
        .CONTROL8(N63), .CONTROL9(N64), .CONTROL10(N65), .CONTROL11(N66), 
        .CONTROL12(N67), .CONTROL13(N68), .CONTROL14(N69), .CONTROL15(N70), 
        .CONTROL16(N71), .Z({N380, N379, N378, N377, N376, N375, N374, N373, 
        N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, 
        N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349}) );
  GTECH_BUF B_56 ( .A(N309), .Z(N56) );
  GTECH_BUF B_57 ( .A(N313), .Z(N57) );
  GTECH_BUF B_58 ( .A(N316), .Z(N58) );
  GTECH_BUF B_59 ( .A(N319), .Z(N59) );
  GTECH_BUF B_60 ( .A(N323), .Z(N60) );
  GTECH_BUF B_61 ( .A(N325), .Z(N61) );
  GTECH_BUF B_62 ( .A(N327), .Z(N62) );
  GTECH_BUF B_63 ( .A(N329), .Z(N63) );
  GTECH_BUF B_64 ( .A(N332), .Z(N64) );
  GTECH_BUF B_65 ( .A(N334), .Z(N65) );
  GTECH_BUF B_66 ( .A(N336), .Z(N66) );
  GTECH_BUF B_67 ( .A(N338), .Z(N67) );
  GTECH_BUF B_68 ( .A(N341), .Z(N68) );
  GTECH_BUF B_69 ( .A(N343), .Z(N69) );
  GTECH_BUF B_70 ( .A(N345), .Z(N70) );
  GTECH_BUF B_71 ( .A(N348), .Z(N71) );
  SELECT_OP C2872 ( .DATA1({N380, N379, N378, N377, N376, N375, N374, N373, 
        N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, 
        N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349}), .DATA2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CONTROL1(N72), 
        .CONTROL2(N73), .Z(regD_out) );
  GTECH_BUF B_72 ( .A(N302), .Z(N72) );
  GTECH_BUF B_73 ( .A(readD_sel[4]), .Z(N73) );
  SELECT_OP C2873 ( .DATA1(write1_in), .DATA2(write2_in), .CONTROL1(N74), 
        .CONTROL2(N385), .Z(r0in) );
  GTECH_BUF B_74 ( .A(N381), .Z(N74) );
  SELECT_OP C2874 ( .DATA1(write1_in), .DATA2(write2_in), .CONTROL1(N75), 
        .CONTROL2(N390), .Z(r1in) );
  GTECH_BUF B_75 ( .A(N386), .Z(N75) );
  SELECT_OP C2875 ( .DATA1(write1_in), .DATA2(write2_in), .CONTROL1(N76), 
        .CONTROL2(N395), .Z(r2in) );
  GTECH_BUF B_76 ( .A(N391), .Z(N76) );
  SELECT_OP C2876 ( .DATA1(write1_in), .DATA2(write2_in), .CONTROL1(N77), 
        .CONTROL2(N399), .Z(r3in) );
  GTECH_BUF B_77 ( .A(N396), .Z(N77) );
  SELECT_OP C2877 ( .DATA1(write1_in), .DATA2(write2_in), .CONTROL1(N78), 
        .CONTROL2(N404), .Z(r4in) );
  GTECH_BUF B_78 ( .A(N400), .Z(N78) );
  SELECT_OP C2878 ( .DATA1(write1_in), .DATA2(write2_in), .CONTROL1(N79), 
        .CONTROL2(N409), .Z(r5in) );
  GTECH_BUF B_79 ( .A(N405), .Z(N79) );
  SELECT_OP C2879 ( .DATA1(write1_in), .DATA2(write2_in), .CONTROL1(N80), 
        .CONTROL2(N414), .Z(r6in) );
  GTECH_BUF B_80 ( .A(N410), .Z(N80) );
  SELECT_OP C2880 ( .DATA1(write1_in), .DATA2(write2_in), .DATA3(r4), 
        .CONTROL1(N81), .CONTROL2(N420), .CONTROL3(N418), .Z(r7in) );
  GTECH_BUF B_81 ( .A(N415), .Z(N81) );
  SELECT_OP C2881 ( .DATA1(write1_in), .DATA2(write2_in), .CONTROL1(N82), 
        .CONTROL2(N425), .Z(r8in) );
  GTECH_BUF B_82 ( .A(N421), .Z(N82) );
  SELECT_OP C2882 ( .DATA1(write1_in), .DATA2(write2_in), .CONTROL1(N83), 
        .CONTROL2(N430), .Z(r9in) );
  GTECH_BUF B_83 ( .A(N426), .Z(N83) );
  SELECT_OP C2883 ( .DATA1(write1_in), .DATA2(write2_in), .CONTROL1(N84), 
        .CONTROL2(N435), .Z(r10in) );
  GTECH_BUF B_84 ( .A(N431), .Z(N84) );
  SELECT_OP C2884 ( .DATA1(write1_in), .DATA2(write2_in), .CONTROL1(N85), 
        .CONTROL2(N440), .Z(r11in) );
  GTECH_BUF B_85 ( .A(N436), .Z(N85) );
  SELECT_OP C2885 ( .DATA1(write1_in), .DATA2(write2_in), .CONTROL1(N86), 
        .CONTROL2(N445), .Z(r12in) );
  GTECH_BUF B_86 ( .A(N441), .Z(N86) );
  SELECT_OP C2886 ( .DATA1(write1_in), .DATA2(write2_in), .DATA3(next_sp_in), 
        .CONTROL1(N87), .CONTROL2(N451), .CONTROL3(N449), .Z(spin) );
  GTECH_BUF B_87 ( .A(N446), .Z(N87) );
  SELECT_OP C2887 ( .DATA1(write1_in), .DATA2(write2_in), .CONTROL1(N88), 
        .CONTROL2(N456), .Z(lrin) );
  GTECH_BUF B_88 ( .A(N452), .Z(N88) );
  SELECT_OP C2888 ( .DATA1(write1_in), .DATA2(write2_in), .CONTROL1(N89), 
        .CONTROL2(N460), .Z(pc_write_in) );
  GTECH_BUF B_89 ( .A(N459), .Z(N89) );
  SELECT_OP C2889 ( .DATA1(pc_write_in), .DATA2(next_pc_in), .CONTROL1(N90), 
        .CONTROL2(N91), .Z(pcin) );
  GTECH_BUF B_90 ( .A(pc_write_select), .Z(N90) );
  GTECH_BUF B_91 ( .A(N461), .Z(N91) );
  SELECT_OP C2890 ( .DATA1(write1_in), .DATA2(write2_in), .CONTROL1(N92), 
        .CONTROL2(N466), .Z(tmp1in) );
  GTECH_BUF B_92 ( .A(N462), .Z(N92) );
  GTECH_NOT I_43 ( .A(readA_sel[4]), .Z(N93) );
  GTECH_NOT I_44 ( .A(readA_sel[0]), .Z(N94) );
  GTECH_NOT I_45 ( .A(N102), .Z(N103) );
  GTECH_NOT I_46 ( .A(N106), .Z(N107) );
  GTECH_NOT I_47 ( .A(N108), .Z(N109) );
  GTECH_NOT I_48 ( .A(N112), .Z(N113) );
  GTECH_NOT I_49 ( .A(N114), .Z(N115) );
  GTECH_NOT I_50 ( .A(N118), .Z(N119) );
  GTECH_NOT I_51 ( .A(N120), .Z(N121) );
  GTECH_NOT I_52 ( .A(N124), .Z(N125) );
  GTECH_NOT I_53 ( .A(N126), .Z(N127) );
  GTECH_NOT I_54 ( .A(N129), .Z(N130) );
  GTECH_NOT I_55 ( .A(N131), .Z(N132) );
  GTECH_NOT I_56 ( .A(N134), .Z(N135) );
  GTECH_NOT I_57 ( .A(N136), .Z(N137) );
  GTECH_NOT I_58 ( .A(N139), .Z(N140) );
  GTECH_NOT I_59 ( .A(N141), .Z(N142) );
  GTECH_NOT I_60 ( .A(N145), .Z(N146) );
  GTECH_NOT I_61 ( .A(readA_sel[3]), .Z(N151) );
  GTECH_NOT I_62 ( .A(readA_sel[2]), .Z(N153) );
  GTECH_NOT I_63 ( .A(readA_sel[1]), .Z(N155) );
  GTECH_OR2 C2914 ( .A(N152), .B(N579), .Z(N157) );
  GTECH_OR2 C2915 ( .A(N154), .B(N156), .Z(N579) );
  GTECH_NOT I_64 ( .A(readB_sel[4]), .Z(N158) );
  GTECH_NOT I_65 ( .A(readB_sel[0]), .Z(N159) );
  GTECH_NOT I_66 ( .A(N167), .Z(N168) );
  GTECH_NOT I_67 ( .A(N171), .Z(N172) );
  GTECH_NOT I_68 ( .A(N173), .Z(N174) );
  GTECH_NOT I_69 ( .A(N177), .Z(N178) );
  GTECH_NOT I_70 ( .A(N179), .Z(N180) );
  GTECH_NOT I_71 ( .A(N183), .Z(N184) );
  GTECH_NOT I_72 ( .A(N185), .Z(N186) );
  GTECH_NOT I_73 ( .A(N189), .Z(N190) );
  GTECH_NOT I_74 ( .A(N191), .Z(N192) );
  GTECH_NOT I_75 ( .A(N194), .Z(N195) );
  GTECH_NOT I_76 ( .A(N196), .Z(N197) );
  GTECH_NOT I_77 ( .A(N199), .Z(N200) );
  GTECH_NOT I_78 ( .A(N201), .Z(N202) );
  GTECH_NOT I_79 ( .A(N204), .Z(N205) );
  GTECH_NOT I_80 ( .A(N206), .Z(N207) );
  GTECH_NOT I_81 ( .A(N210), .Z(N211) );
  GTECH_NOT I_82 ( .A(readB_sel[3]), .Z(N216) );
  GTECH_NOT I_83 ( .A(readB_sel[2]), .Z(N218) );
  GTECH_NOT I_84 ( .A(readB_sel[1]), .Z(N220) );
  GTECH_OR2 C2956 ( .A(N217), .B(N580), .Z(N222) );
  GTECH_OR2 C2957 ( .A(N219), .B(N221), .Z(N580) );
  GTECH_NOT I_85 ( .A(readC_sel[4]), .Z(N223) );
  GTECH_NOT I_86 ( .A(readC_sel[3]), .Z(N224) );
  GTECH_NOT I_87 ( .A(readC_sel[2]), .Z(N225) );
  GTECH_NOT I_88 ( .A(readC_sel[1]), .Z(N226) );
  GTECH_NOT I_89 ( .A(readC_sel[0]), .Z(N227) );
  GTECH_NOT I_90 ( .A(N233), .Z(N234) );
  GTECH_NOT I_91 ( .A(N236), .Z(N237) );
  GTECH_NOT I_92 ( .A(N239), .Z(N240) );
  GTECH_NOT I_93 ( .A(N243), .Z(N244) );
  GTECH_NOT I_94 ( .A(N245), .Z(N246) );
  GTECH_NOT I_95 ( .A(N247), .Z(N248) );
  GTECH_NOT I_96 ( .A(N249), .Z(N250) );
  GTECH_NOT I_97 ( .A(N252), .Z(N253) );
  GTECH_NOT I_98 ( .A(N254), .Z(N255) );
  GTECH_NOT I_99 ( .A(N256), .Z(N257) );
  GTECH_NOT I_100 ( .A(N258), .Z(N259) );
  GTECH_NOT I_101 ( .A(N261), .Z(N262) );
  GTECH_NOT I_102 ( .A(N263), .Z(N264) );
  GTECH_NOT I_103 ( .A(N265), .Z(N266) );
  GTECH_NOT I_104 ( .A(readD_sel[4]), .Z(N302) );
  GTECH_NOT I_105 ( .A(readD_sel[3]), .Z(N303) );
  GTECH_NOT I_106 ( .A(readD_sel[2]), .Z(N304) );
  GTECH_NOT I_107 ( .A(readD_sel[1]), .Z(N305) );
  GTECH_NOT I_108 ( .A(readD_sel[0]), .Z(N306) );
  GTECH_NOT I_109 ( .A(N312), .Z(N313) );
  GTECH_NOT I_110 ( .A(N315), .Z(N316) );
  GTECH_NOT I_111 ( .A(N318), .Z(N319) );
  GTECH_NOT I_112 ( .A(N322), .Z(N323) );
  GTECH_NOT I_113 ( .A(N324), .Z(N325) );
  GTECH_NOT I_114 ( .A(N326), .Z(N327) );
  GTECH_NOT I_115 ( .A(N328), .Z(N329) );
  GTECH_NOT I_116 ( .A(N331), .Z(N332) );
  GTECH_NOT I_117 ( .A(N333), .Z(N334) );
  GTECH_NOT I_118 ( .A(N335), .Z(N336) );
  GTECH_NOT I_119 ( .A(N337), .Z(N338) );
  GTECH_NOT I_120 ( .A(N340), .Z(N341) );
  GTECH_NOT I_121 ( .A(N342), .Z(N343) );
  GTECH_NOT I_122 ( .A(N344), .Z(N345) );
  GTECH_AND2 C3051 ( .A(N478), .B(write1_en), .Z(N381) );
  GTECH_AND2 C3052 ( .A(N473), .B(write2_en), .Z(N382) );
  GTECH_OR2 C3055 ( .A(N382), .B(N381), .Z(N383) );
  GTECH_NOT I_123 ( .A(N381), .Z(N384) );
  GTECH_AND2 C3058 ( .A(N382), .B(N384), .Z(N385) );
  GTECH_AND2 C3059 ( .A(N484), .B(write1_en), .Z(N386) );
  GTECH_AND2 C3060 ( .A(N481), .B(write2_en), .Z(N387) );
  GTECH_OR2 C3063 ( .A(N387), .B(N386), .Z(N388) );
  GTECH_NOT I_124 ( .A(N386), .Z(N389) );
  GTECH_AND2 C3066 ( .A(N387), .B(N389), .Z(N390) );
  GTECH_AND2 C3067 ( .A(N492), .B(write1_en), .Z(N391) );
  GTECH_AND2 C3068 ( .A(N488), .B(write2_en), .Z(N392) );
  GTECH_OR2 C3071 ( .A(N392), .B(N391), .Z(N393) );
  GTECH_NOT I_125 ( .A(N391), .Z(N394) );
  GTECH_AND2 C3074 ( .A(N392), .B(N394), .Z(N395) );
  GTECH_AND2 C3075 ( .A(N494), .B(write1_en), .Z(N396) );
  GTECH_OR2 C3077 ( .A(N392), .B(N396), .Z(N397) );
  GTECH_NOT I_126 ( .A(N396), .Z(N398) );
  GTECH_AND2 C3080 ( .A(N392), .B(N398), .Z(N399) );
  GTECH_AND2 C3081 ( .A(N504), .B(write1_en), .Z(N400) );
  GTECH_AND2 C3082 ( .A(N499), .B(write2_en), .Z(N401) );
  GTECH_OR2 C3085 ( .A(N401), .B(N400), .Z(N402) );
  GTECH_NOT I_127 ( .A(N400), .Z(N403) );
  GTECH_AND2 C3088 ( .A(N401), .B(N403), .Z(N404) );
  GTECH_AND2 C3089 ( .A(N508), .B(write1_en), .Z(N405) );
  GTECH_AND2 C3090 ( .A(N506), .B(write2_en), .Z(N406) );
  GTECH_OR2 C3093 ( .A(N406), .B(N405), .Z(N407) );
  GTECH_NOT I_128 ( .A(N405), .Z(N408) );
  GTECH_AND2 C3096 ( .A(N406), .B(N408), .Z(N409) );
  GTECH_AND2 C3097 ( .A(N514), .B(write1_en), .Z(N410) );
  GTECH_AND2 C3098 ( .A(N511), .B(write2_en), .Z(N411) );
  GTECH_OR2 C3101 ( .A(N411), .B(N410), .Z(N412) );
  GTECH_NOT I_129 ( .A(N410), .Z(N413) );
  GTECH_AND2 C3104 ( .A(N411), .B(N413), .Z(N414) );
  GTECH_AND2 C3105 ( .A(N518), .B(write1_en), .Z(N415) );
  GTECH_AND2 C3106 ( .A(N516), .B(write2_en), .Z(N416) );
  GTECH_OR2 C3109 ( .A(N416), .B(N415), .Z(N417) );
  GTECH_NOT I_130 ( .A(N417), .Z(N418) );
  GTECH_NOT I_131 ( .A(N415), .Z(N419) );
  GTECH_AND2 C3112 ( .A(N416), .B(N419), .Z(N420) );
  GTECH_AND2 C3113 ( .A(N530), .B(write1_en), .Z(N421) );
  GTECH_AND2 C3114 ( .A(N524), .B(write2_en), .Z(N422) );
  GTECH_OR2 C3117 ( .A(N422), .B(N421), .Z(N423) );
  GTECH_NOT I_132 ( .A(N421), .Z(N424) );
  GTECH_AND2 C3120 ( .A(N422), .B(N424), .Z(N425) );
  GTECH_AND2 C3121 ( .A(N534), .B(write1_en), .Z(N426) );
  GTECH_AND2 C3122 ( .A(N532), .B(write2_en), .Z(N427) );
  GTECH_OR2 C3125 ( .A(N427), .B(N426), .Z(N428) );
  GTECH_NOT I_133 ( .A(N426), .Z(N429) );
  GTECH_AND2 C3128 ( .A(N427), .B(N429), .Z(N430) );
  GTECH_AND2 C3129 ( .A(N540), .B(write1_en), .Z(N431) );
  GTECH_AND2 C3130 ( .A(N537), .B(write2_en), .Z(N432) );
  GTECH_OR2 C3133 ( .A(N432), .B(N431), .Z(N433) );
  GTECH_NOT I_134 ( .A(N431), .Z(N434) );
  GTECH_AND2 C3136 ( .A(N432), .B(N434), .Z(N435) );
  GTECH_AND2 C3137 ( .A(N544), .B(write1_en), .Z(N436) );
  GTECH_AND2 C3138 ( .A(N542), .B(write2_en), .Z(N437) );
  GTECH_OR2 C3141 ( .A(N437), .B(N436), .Z(N438) );
  GTECH_NOT I_135 ( .A(N436), .Z(N439) );
  GTECH_AND2 C3144 ( .A(N437), .B(N439), .Z(N440) );
  GTECH_AND2 C3145 ( .A(N552), .B(write1_en), .Z(N441) );
  GTECH_AND2 C3146 ( .A(N548), .B(write2_en), .Z(N442) );
  GTECH_OR2 C3149 ( .A(N442), .B(N441), .Z(N443) );
  GTECH_NOT I_136 ( .A(N441), .Z(N444) );
  GTECH_AND2 C3152 ( .A(N442), .B(N444), .Z(N445) );
  GTECH_AND2 C3153 ( .A(N562), .B(write1_en), .Z(N446) );
  GTECH_AND2 C3154 ( .A(N560), .B(write2_en), .Z(N447) );
  GTECH_OR2 C3157 ( .A(N447), .B(N446), .Z(N448) );
  GTECH_NOT I_137 ( .A(N448), .Z(N449) );
  GTECH_NOT I_138 ( .A(N446), .Z(N450) );
  GTECH_AND2 C3160 ( .A(N447), .B(N450), .Z(N451) );
  GTECH_AND2 C3161 ( .A(N558), .B(write1_en), .Z(N452) );
  GTECH_AND2 C3162 ( .A(N555), .B(write2_en), .Z(N453) );
  GTECH_OR2 C3165 ( .A(N453), .B(N452), .Z(N454) );
  GTECH_NOT I_139 ( .A(N452), .Z(N455) );
  GTECH_AND2 C3168 ( .A(N453), .B(N455), .Z(N456) );
  GTECH_OR2 C3169 ( .A(N581), .B(N582), .Z(pc_write_select) );
  GTECH_AND2 C3170 ( .A(write1_en), .B(N564), .Z(N581) );
  GTECH_AND2 C3171 ( .A(write2_en), .B(N566), .Z(N582) );
  GTECH_OR2 C3172 ( .A(N612), .B(next_pc_en[0]), .Z(N457) );
  GTECH_OR2 C3173 ( .A(N611), .B(next_pc_en[1]), .Z(N612) );
  GTECH_OR2 C3174 ( .A(N610), .B(next_pc_en[2]), .Z(N611) );
  GTECH_OR2 C3175 ( .A(N609), .B(next_pc_en[3]), .Z(N610) );
  GTECH_OR2 C3176 ( .A(N608), .B(next_pc_en[4]), .Z(N609) );
  GTECH_OR2 C3177 ( .A(N607), .B(next_pc_en[5]), .Z(N608) );
  GTECH_OR2 C3178 ( .A(N606), .B(next_pc_en[6]), .Z(N607) );
  GTECH_OR2 C3179 ( .A(N605), .B(next_pc_en[7]), .Z(N606) );
  GTECH_OR2 C3180 ( .A(N604), .B(next_pc_en[8]), .Z(N605) );
  GTECH_OR2 C3181 ( .A(N603), .B(next_pc_en[9]), .Z(N604) );
  GTECH_OR2 C3182 ( .A(N602), .B(next_pc_en[10]), .Z(N603) );
  GTECH_OR2 C3183 ( .A(N601), .B(next_pc_en[11]), .Z(N602) );
  GTECH_OR2 C3184 ( .A(N600), .B(next_pc_en[12]), .Z(N601) );
  GTECH_OR2 C3185 ( .A(N599), .B(next_pc_en[13]), .Z(N600) );
  GTECH_OR2 C3186 ( .A(N598), .B(next_pc_en[14]), .Z(N599) );
  GTECH_OR2 C3187 ( .A(N597), .B(next_pc_en[15]), .Z(N598) );
  GTECH_OR2 C3188 ( .A(N596), .B(next_pc_en[16]), .Z(N597) );
  GTECH_OR2 C3189 ( .A(N595), .B(next_pc_en[17]), .Z(N596) );
  GTECH_OR2 C3190 ( .A(N594), .B(next_pc_en[18]), .Z(N595) );
  GTECH_OR2 C3191 ( .A(N593), .B(next_pc_en[19]), .Z(N594) );
  GTECH_OR2 C3192 ( .A(N592), .B(next_pc_en[20]), .Z(N593) );
  GTECH_OR2 C3193 ( .A(N591), .B(next_pc_en[21]), .Z(N592) );
  GTECH_OR2 C3194 ( .A(N590), .B(next_pc_en[22]), .Z(N591) );
  GTECH_OR2 C3195 ( .A(N589), .B(next_pc_en[23]), .Z(N590) );
  GTECH_OR2 C3196 ( .A(N588), .B(next_pc_en[24]), .Z(N589) );
  GTECH_OR2 C3197 ( .A(N587), .B(next_pc_en[25]), .Z(N588) );
  GTECH_OR2 C3198 ( .A(N586), .B(next_pc_en[26]), .Z(N587) );
  GTECH_OR2 C3199 ( .A(N585), .B(next_pc_en[27]), .Z(N586) );
  GTECH_OR2 C3200 ( .A(N584), .B(next_pc_en[28]), .Z(N585) );
  GTECH_OR2 C3201 ( .A(N583), .B(next_pc_en[29]), .Z(N584) );
  GTECH_OR2 C3202 ( .A(next_pc_en[31]), .B(next_pc_en[30]), .Z(N583) );
  GTECH_NOT I_140 ( .A(N457), .Z(N458) );
  GTECH_AND2 C3205 ( .A(write1_en), .B(N564), .Z(N459) );
  GTECH_NOT I_141 ( .A(N459), .Z(N460) );
  GTECH_NOT I_142 ( .A(pc_write_select), .Z(N461) );
  GTECH_AND2 C3211 ( .A(N578), .B(write1_en), .Z(N462) );
  GTECH_AND2 C3212 ( .A(N572), .B(write2_en), .Z(N463) );
  GTECH_OR2 C3215 ( .A(N463), .B(N462), .Z(N464) );
  GTECH_NOT I_143 ( .A(N462), .Z(N465) );
  GTECH_AND2 C3218 ( .A(N463), .B(N465), .Z(N466) );
  GTECH_AND2 C3232 ( .A(N458), .B(N461), .Z(N467) );
  GTECH_NOT I_144 ( .A(N467), .Z(N468) );
endmodule

