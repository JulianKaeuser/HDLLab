
module ALU_VARIABLE ( a, b, op, c_in, result, c_out, z, n, v );
  input [31:0] a;
  input [31:0] b;
  input [3:0] op;
  output [31:0] result;
  input c_in;
  output c_out, z, n, v;
  wire   mult_x_18_n1010, mult_x_18_n1006, mult_x_18_n1002, mult_x_18_n998,
         mult_x_18_n994, mult_x_18_n990, mult_x_18_n986, mult_x_18_n979,
         mult_x_18_n978, mult_x_18_n975, mult_x_18_n974, mult_x_18_n971,
         mult_x_18_n970, mult_x_18_n969, mult_x_18_n967, mult_x_18_n966,
         mult_x_18_n963, mult_x_18_n962, mult_x_18_n959, mult_x_18_n958,
         mult_x_18_n957, mult_x_18_n955, mult_x_18_n954, mult_x_18_n950,
         mult_x_18_n948, mult_x_18_n946, mult_x_18_n945, mult_x_18_n944,
         mult_x_18_n942, mult_x_18_n941, mult_x_18_n940, mult_x_18_n939,
         mult_x_18_n938, mult_x_18_n937, mult_x_18_n936, mult_x_18_n935,
         mult_x_18_n934, mult_x_18_n933, mult_x_18_n932, mult_x_18_n931,
         mult_x_18_n930, mult_x_18_n929, mult_x_18_n928, mult_x_18_n927,
         mult_x_18_n926, mult_x_18_n925, mult_x_18_n923, mult_x_18_n922,
         mult_x_18_n921, mult_x_18_n920, mult_x_18_n919, mult_x_18_n918,
         mult_x_18_n917, mult_x_18_n916, mult_x_18_n915, mult_x_18_n914,
         mult_x_18_n912, mult_x_18_n911, mult_x_18_n910, mult_x_18_n909,
         mult_x_18_n908, mult_x_18_n907, mult_x_18_n906, mult_x_18_n905,
         mult_x_18_n904, mult_x_18_n903, mult_x_18_n902, mult_x_18_n901,
         mult_x_18_n900, mult_x_18_n899, mult_x_18_n898, mult_x_18_n894,
         mult_x_18_n893, mult_x_18_n892, mult_x_18_n891, mult_x_18_n890,
         mult_x_18_n889, mult_x_18_n888, mult_x_18_n887, mult_x_18_n886,
         mult_x_18_n885, mult_x_18_n884, mult_x_18_n883, mult_x_18_n882,
         mult_x_18_n881, mult_x_18_n880, mult_x_18_n879, mult_x_18_n878,
         mult_x_18_n877, mult_x_18_n875, mult_x_18_n874, mult_x_18_n873,
         mult_x_18_n871, mult_x_18_n870, mult_x_18_n869, mult_x_18_n867,
         mult_x_18_n865, mult_x_18_n863, mult_x_18_n862, mult_x_18_n861,
         mult_x_18_n859, mult_x_18_n858, mult_x_18_n857, mult_x_18_n855,
         mult_x_18_n854, mult_x_18_n853, mult_x_18_n852, mult_x_18_n851,
         mult_x_18_n850, mult_x_18_n847, mult_x_18_n846, mult_x_18_n845,
         mult_x_18_n844, mult_x_18_n843, mult_x_18_n842, mult_x_18_n841,
         mult_x_18_n840, mult_x_18_n839, mult_x_18_n838, mult_x_18_n837,
         mult_x_18_n836, mult_x_18_n835, mult_x_18_n834, mult_x_18_n833,
         mult_x_18_n832, mult_x_18_n831, mult_x_18_n830, mult_x_18_n829,
         mult_x_18_n827, mult_x_18_n826, mult_x_18_n825, mult_x_18_n824,
         mult_x_18_n823, mult_x_18_n822, mult_x_18_n821, mult_x_18_n820,
         mult_x_18_n819, mult_x_18_n818, mult_x_18_n817, mult_x_18_n816,
         mult_x_18_n815, mult_x_18_n814, mult_x_18_n813, mult_x_18_n812,
         mult_x_18_n811, mult_x_18_n810, mult_x_18_n806, mult_x_18_n804,
         mult_x_18_n802, mult_x_18_n800, mult_x_18_n798, mult_x_18_n796,
         mult_x_18_n795, mult_x_18_n794, mult_x_18_n793, mult_x_18_n791,
         mult_x_18_n790, mult_x_18_n789, mult_x_18_n788, mult_x_18_n787,
         mult_x_18_n786, mult_x_18_n785, mult_x_18_n784, mult_x_18_n783,
         mult_x_18_n782, mult_x_18_n781, mult_x_18_n780, mult_x_18_n779,
         mult_x_18_n778, mult_x_18_n775, mult_x_18_n774, mult_x_18_n773,
         mult_x_18_n772, mult_x_18_n771, mult_x_18_n770, mult_x_18_n769,
         mult_x_18_n768, mult_x_18_n767, mult_x_18_n766, mult_x_18_n765,
         mult_x_18_n763, mult_x_18_n762, mult_x_18_n761, mult_x_18_n759,
         mult_x_18_n758, mult_x_18_n757, mult_x_18_n755, mult_x_18_n754,
         mult_x_18_n751, mult_x_18_n750, mult_x_18_n749, mult_x_18_n748,
         mult_x_18_n747, mult_x_18_n746, mult_x_18_n745, mult_x_18_n743,
         mult_x_18_n742, mult_x_18_n741, mult_x_18_n740, mult_x_18_n739,
         mult_x_18_n738, mult_x_18_n734, mult_x_18_n733, mult_x_18_n731,
         mult_x_18_n730, mult_x_18_n725, mult_x_18_n721, mult_x_18_n719,
         mult_x_18_n717, mult_x_18_n716, mult_x_18_n715, mult_x_18_n707,
         mult_x_18_n704, mult_x_18_n703, mult_x_18_n702, mult_x_18_n701,
         mult_x_18_n700, mult_x_18_n699, mult_x_18_n698, mult_x_18_n697,
         mult_x_18_n696, mult_x_18_n695, mult_x_18_n694, mult_x_18_n693,
         mult_x_18_n692, mult_x_18_n691, mult_x_18_n690, mult_x_18_n689,
         mult_x_18_n688, mult_x_18_n687, mult_x_18_n686, mult_x_18_n685,
         mult_x_18_n684, mult_x_18_n683, mult_x_18_n682, mult_x_18_n681,
         mult_x_18_n680, mult_x_18_n679, mult_x_18_n678, mult_x_18_n677,
         mult_x_18_n676, mult_x_18_n675, mult_x_18_n674, mult_x_18_n673,
         mult_x_18_n672, mult_x_18_n671, mult_x_18_n670, mult_x_18_n669,
         mult_x_18_n668, mult_x_18_n667, mult_x_18_n666, mult_x_18_n665,
         mult_x_18_n664, mult_x_18_n663, mult_x_18_n662, mult_x_18_n661,
         mult_x_18_n660, mult_x_18_n659, mult_x_18_n658, mult_x_18_n657,
         mult_x_18_n656, mult_x_18_n655, mult_x_18_n654, mult_x_18_n653,
         mult_x_18_n652, mult_x_18_n651, mult_x_18_n650, mult_x_18_n649,
         mult_x_18_n648, mult_x_18_n647, mult_x_18_n646, mult_x_18_n645,
         mult_x_18_n644, mult_x_18_n643, mult_x_18_n642, mult_x_18_n641,
         mult_x_18_n640, mult_x_18_n639, mult_x_18_n638, mult_x_18_n637,
         mult_x_18_n636, mult_x_18_n635, mult_x_18_n634, mult_x_18_n633,
         mult_x_18_n632, mult_x_18_n631, mult_x_18_n630, mult_x_18_n629,
         mult_x_18_n628, mult_x_18_n627, mult_x_18_n626, mult_x_18_n625,
         mult_x_18_n624, mult_x_18_n623, mult_x_18_n622, mult_x_18_n621,
         mult_x_18_n620, mult_x_18_n619, mult_x_18_n618, mult_x_18_n617,
         mult_x_18_n616, mult_x_18_n615, mult_x_18_n614, mult_x_18_n613,
         mult_x_18_n612, mult_x_18_n611, mult_x_18_n610, mult_x_18_n609,
         mult_x_18_n608, mult_x_18_n607, mult_x_18_n606, mult_x_18_n605,
         mult_x_18_n604, mult_x_18_n603, mult_x_18_n602, mult_x_18_n601,
         mult_x_18_n600, mult_x_18_n599, mult_x_18_n598, mult_x_18_n597,
         mult_x_18_n596, mult_x_18_n595, mult_x_18_n594, mult_x_18_n593,
         mult_x_18_n592, mult_x_18_n591, mult_x_18_n590, mult_x_18_n589,
         mult_x_18_n588, mult_x_18_n587, mult_x_18_n586, mult_x_18_n585,
         mult_x_18_n584, mult_x_18_n583, mult_x_18_n582, mult_x_18_n581,
         mult_x_18_n580, mult_x_18_n579, mult_x_18_n578, mult_x_18_n577,
         mult_x_18_n576, mult_x_18_n575, mult_x_18_n574, mult_x_18_n573,
         mult_x_18_n572, mult_x_18_n571, mult_x_18_n570, mult_x_18_n569,
         mult_x_18_n568, mult_x_18_n567, mult_x_18_n566, mult_x_18_n565,
         mult_x_18_n564, mult_x_18_n563, mult_x_18_n562, mult_x_18_n561,
         mult_x_18_n560, mult_x_18_n559, mult_x_18_n558, mult_x_18_n557,
         mult_x_18_n556, mult_x_18_n555, mult_x_18_n554, mult_x_18_n553,
         mult_x_18_n552, mult_x_18_n551, mult_x_18_n550, mult_x_18_n549,
         mult_x_18_n548, mult_x_18_n547, mult_x_18_n546, mult_x_18_n545,
         mult_x_18_n544, mult_x_18_n543, mult_x_18_n542, mult_x_18_n541,
         mult_x_18_n540, mult_x_18_n539, mult_x_18_n538, mult_x_18_n537,
         mult_x_18_n536, mult_x_18_n535, mult_x_18_n534, mult_x_18_n533,
         mult_x_18_n532, mult_x_18_n531, mult_x_18_n530, mult_x_18_n529,
         mult_x_18_n528, mult_x_18_n527, mult_x_18_n526, mult_x_18_n525,
         mult_x_18_n524, mult_x_18_n523, mult_x_18_n522, mult_x_18_n521,
         mult_x_18_n520, mult_x_18_n519, mult_x_18_n518, mult_x_18_n517,
         mult_x_18_n516, mult_x_18_n515, mult_x_18_n514, mult_x_18_n513,
         mult_x_18_n512, mult_x_18_n511, mult_x_18_n510, mult_x_18_n509,
         mult_x_18_n508, mult_x_18_n507, mult_x_18_n506, mult_x_18_n505,
         mult_x_18_n504, mult_x_18_n503, mult_x_18_n502, mult_x_18_n501,
         mult_x_18_n500, mult_x_18_n499, mult_x_18_n498, mult_x_18_n497,
         mult_x_18_n496, mult_x_18_n495, mult_x_18_n494, mult_x_18_n493,
         mult_x_18_n492, mult_x_18_n491, mult_x_18_n490, mult_x_18_n489,
         mult_x_18_n488, mult_x_18_n487, mult_x_18_n486, mult_x_18_n485,
         mult_x_18_n484, mult_x_18_n483, mult_x_18_n482, mult_x_18_n481,
         mult_x_18_n480, mult_x_18_n479, mult_x_18_n478, mult_x_18_n477,
         mult_x_18_n476, mult_x_18_n475, mult_x_18_n474, mult_x_18_n473,
         mult_x_18_n472, mult_x_18_n471, mult_x_18_n470, mult_x_18_n469,
         mult_x_18_n468, mult_x_18_n467, mult_x_18_n466, mult_x_18_n465,
         mult_x_18_n464, mult_x_18_n463, mult_x_18_n462, mult_x_18_n461,
         mult_x_18_n460, mult_x_18_n459, mult_x_18_n458, mult_x_18_n457,
         mult_x_18_n456, mult_x_18_n455, mult_x_18_n454, mult_x_18_n453,
         mult_x_18_n452, mult_x_18_n451, mult_x_18_n450, mult_x_18_n449,
         mult_x_18_n448, mult_x_18_n447, mult_x_18_n446, mult_x_18_n445,
         mult_x_18_n444, mult_x_18_n443, mult_x_18_n442, mult_x_18_n441,
         mult_x_18_n440, mult_x_18_n439, mult_x_18_n438, mult_x_18_n437,
         mult_x_18_n436, mult_x_18_n435, mult_x_18_n434, mult_x_18_n433,
         mult_x_18_n432, mult_x_18_n431, mult_x_18_n430, mult_x_18_n429,
         mult_x_18_n428, mult_x_18_n427, mult_x_18_n426, mult_x_18_n425,
         mult_x_18_n424, mult_x_18_n423, mult_x_18_n422, mult_x_18_n421,
         mult_x_18_n420, mult_x_18_n419, mult_x_18_n418, mult_x_18_n417,
         mult_x_18_n416, mult_x_18_n415, mult_x_18_n414, mult_x_18_n413,
         mult_x_18_n412, mult_x_18_n411, mult_x_18_n410, mult_x_18_n409,
         mult_x_18_n408, mult_x_18_n407, mult_x_18_n406, mult_x_18_n405,
         mult_x_18_n404, mult_x_18_n403, mult_x_18_n402, mult_x_18_n401,
         mult_x_18_n400, mult_x_18_n399, mult_x_18_n398, mult_x_18_n397,
         mult_x_18_n396, mult_x_18_n395, mult_x_18_n394, mult_x_18_n393,
         mult_x_18_n392, mult_x_18_n391, mult_x_18_n390, mult_x_18_n389,
         mult_x_18_n388, mult_x_18_n387, mult_x_18_n386, mult_x_18_n385,
         mult_x_18_n384, mult_x_18_n383, mult_x_18_n381, mult_x_18_n380,
         mult_x_18_n379, mult_x_18_n378, mult_x_18_n377, mult_x_18_n376,
         mult_x_18_n375, mult_x_18_n374, mult_x_18_n373, mult_x_18_n372,
         mult_x_18_n371, mult_x_18_n370, mult_x_18_n369, mult_x_18_n368,
         mult_x_18_n367, mult_x_18_n366, mult_x_18_n365, mult_x_18_n364,
         mult_x_18_n363, mult_x_18_n362, mult_x_18_n361, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978;
  tri   [3:0] op;

  CMPE42D1BWP12T mult_x_18_U486 ( .A(mult_x_18_n725), .B(mult_x_18_n922), .C(
        mult_x_18_n978), .CIX(mult_x_18_n702), .D(mult_x_18_n701), .CO(
        mult_x_18_n698), .COX(mult_x_18_n697), .S(mult_x_18_n699) );
  CMPE42D1BWP12T mult_x_18_U460 ( .A(mult_x_18_n888), .B(mult_x_18_n865), .C(
        mult_x_18_n969), .CIX(mult_x_18_n636), .D(mult_x_18_n642), .CO(
        mult_x_18_n629), .COX(mult_x_18_n628), .S(mult_x_18_n630) );
  CMPE42D1BWP12T mult_x_18_U455 ( .A(mult_x_18_n887), .B(mult_x_18_n939), .C(
        mult_x_18_n912), .CIX(mult_x_18_n625), .D(mult_x_18_n621), .CO(
        mult_x_18_n616), .COX(mult_x_18_n615), .S(mult_x_18_n617) );
  CMPE42D1BWP12T mult_x_18_U473 ( .A(mult_x_18_n670), .B(mult_x_18_n944), .C(
        mult_x_18_n671), .CIX(mult_x_18_n675), .D(mult_x_18_n668), .CO(
        mult_x_18_n664), .COX(mult_x_18_n663), .S(mult_x_18_n665) );
  CMPE42D1BWP12T mult_x_18_U449 ( .A(mult_x_18_n616), .B(mult_x_18_n605), .C(
        mult_x_18_n613), .CIX(mult_x_18_n609), .D(mult_x_18_n602), .CO(
        mult_x_18_n598), .COX(mult_x_18_n597), .S(mult_x_18_n599) );
  CMPE42D1BWP12T mult_x_18_U410 ( .A(mult_x_18_n514), .B(mult_x_18_n496), .C(
        mult_x_18_n511), .CIX(mult_x_18_n507), .D(mult_x_18_n493), .CO(
        mult_x_18_n489), .COX(mult_x_18_n488), .S(mult_x_18_n490) );
  CMPE42D1BWP12T mult_x_18_U469 ( .A(mult_x_18_n660), .B(mult_x_18_n662), .C(
        mult_x_18_n663), .CIX(mult_x_18_n658), .D(mult_x_18_n667), .CO(
        mult_x_18_n654), .COX(mult_x_18_n653), .S(mult_x_18_n655) );
  INVD1BWP12T U3 ( .I(a[27]), .ZN(n1816) );
  ND2D1BWP12T U4 ( .A1(n2671), .A2(n2977), .ZN(n2699) );
  INVD1BWP12T U5 ( .I(n1717), .ZN(n852) );
  MAOI22D0BWP12T U6 ( .A1(n2932), .A2(n2720), .B1(n2719), .B2(n2718), .ZN(
        n2727) );
  MOAI22D0BWP12T U7 ( .A1(n2725), .A2(n2806), .B1(n2722), .B2(b[21]), .ZN(
        n2723) );
  HA1D0BWP12T U8 ( .A(n1347), .B(n1346), .CO(mult_x_18_n595), .S(
        mult_x_18_n596) );
  HA1D0BWP12T U9 ( .A(n1307), .B(n1306), .CO(mult_x_18_n620), .S(
        mult_x_18_n621) );
  HA1D0BWP12T U10 ( .A(n1341), .B(n1340), .CO(mult_x_18_n642), .S(
        mult_x_18_n643) );
  HA1D0BWP12T U11 ( .A(n1313), .B(n1312), .CO(mult_x_18_n677), .S(
        mult_x_18_n678) );
  XNR2D1BWP12T U12 ( .A1(a[25]), .A2(n2477), .ZN(n1215) );
  HA1D0BWP12T U13 ( .A(n1335), .B(n1334), .CO(mult_x_18_n690), .S(
        mult_x_18_n691) );
  HA1D0BWP12T U14 ( .A(n1295), .B(n1294), .CO(mult_x_18_n700), .S(
        mult_x_18_n701) );
  INVD1BWP12T U15 ( .I(n2477), .ZN(n557) );
  XNR2D1BWP12T U16 ( .A1(a[25]), .A2(b[6]), .ZN(n1043) );
  CMPE42D1BWP12T U17 ( .A(mult_x_18_n517), .B(mult_x_18_n499), .C(
        mult_x_18_n490), .CIX(mult_x_18_n504), .D(mult_x_18_n508), .CO(
        mult_x_18_n486), .COX(mult_x_18_n485), .S(mult_x_18_n487) );
  CMPE42D1BWP12T U18 ( .A(mult_x_18_n629), .B(mult_x_18_n617), .C(
        mult_x_18_n626), .CIX(mult_x_18_n622), .D(mult_x_18_n614), .CO(
        mult_x_18_n610), .COX(mult_x_18_n609), .S(mult_x_18_n611) );
  CMPE42D1BWP12T U19 ( .A(mult_x_18_n604), .B(mult_x_18_n591), .C(
        mult_x_18_n601), .CIX(mult_x_18_n597), .D(mult_x_18_n588), .CO(
        mult_x_18_n584), .COX(mult_x_18_n583), .S(mult_x_18_n585) );
  OAI21D1BWP12T U20 ( .A1(n1397), .A2(n1396), .B(n1417), .ZN(n2343) );
  ND2D1BWP12T U21 ( .A1(n1870), .A2(n1869), .ZN(n1398) );
  CKBD1BWP12T U22 ( .I(n2527), .Z(n528) );
  INVD1BWP12T U23 ( .I(n2528), .ZN(n569) );
  CKBD1BWP12T U24 ( .I(n2527), .Z(n570) );
  NR2D1BWP12T U25 ( .A1(n1891), .A2(n472), .ZN(n1400) );
  NR2D1BWP12T U26 ( .A1(n803), .A2(n1398), .ZN(n2001) );
  INVD1BWP12T U27 ( .I(b[6]), .ZN(n564) );
  INVD2BWP12T U28 ( .I(n750), .ZN(n1872) );
  INVD1BWP12T U29 ( .I(b[4]), .ZN(n466) );
  INVD1BWP12T U30 ( .I(b[3]), .ZN(n539) );
  NR2D1BWP12T U31 ( .A1(n2528), .A2(b[6]), .ZN(n505) );
  OAI21D1BWP12T U32 ( .A1(n946), .A2(n945), .B(n953), .ZN(n1010) );
  NR2D1BWP12T U33 ( .A1(n2620), .A2(n563), .ZN(n1625) );
  INVD1BWP12T U34 ( .I(n2231), .ZN(n1558) );
  INVD1BWP12T U35 ( .I(b[14]), .ZN(n2275) );
  INVD1BWP12T U36 ( .I(b[13]), .ZN(n2278) );
  INVD1BWP12T U37 ( .I(b[15]), .ZN(n2276) );
  INVD1BWP12T U38 ( .I(a[17]), .ZN(n2683) );
  XNR2XD4BWP12T U39 ( .A1(n2594), .A2(n2308), .ZN(n2644) );
  ND2D1BWP12T U40 ( .A1(n2397), .A2(n2967), .ZN(n1379) );
  INVD1BWP12T U41 ( .I(n1804), .ZN(n1536) );
  AOI21D1BWP12T U42 ( .A1(n693), .A2(n611), .B(n610), .ZN(n1665) );
  OR2XD1BWP12T U43 ( .A1(mult_x_18_n540), .A2(mult_x_18_n554), .Z(n1669) );
  OR2XD1BWP12T U44 ( .A1(mult_x_18_n571), .A2(mult_x_18_n584), .Z(n1723) );
  OAI21D1BWP12T U45 ( .A1(n1794), .A2(n1793), .B(n2337), .ZN(n783) );
  INVD2BWP12T U46 ( .I(n2234), .ZN(n2609) );
  INVD1BWP12T U47 ( .I(a[18]), .ZN(n2705) );
  INVD1BWP12T U48 ( .I(b[18]), .ZN(n2703) );
  INVD1BWP12T U49 ( .I(n2598), .ZN(n2277) );
  OAI21D1BWP12T U50 ( .A1(n2369), .A2(n637), .B(n636), .ZN(n2350) );
  INVD1BWP12T U51 ( .I(n2897), .ZN(n2899) );
  OR2XD1BWP12T U52 ( .A1(mult_x_18_n687), .A2(mult_x_18_n693), .Z(n589) );
  ND2D1BWP12T U53 ( .A1(n476), .A2(n2080), .ZN(n1997) );
  INVD1BWP12T U54 ( .I(b[9]), .ZN(n2283) );
  INVD1BWP12T U55 ( .I(n2605), .ZN(n571) );
  INVD1BWP12T U56 ( .I(n616), .ZN(n2450) );
  INR2D1BWP12T U57 ( .A1(n471), .B1(n1870), .ZN(n1891) );
  OR2XD1BWP12T U58 ( .A1(n2639), .A2(n2831), .Z(n2052) );
  IND2D1BWP12T U59 ( .A1(n2831), .B1(n2639), .ZN(n1926) );
  CKBD1BWP12T U60 ( .I(n466), .Z(n2870) );
  CKBD1BWP12T U61 ( .I(n539), .Z(n2827) );
  INVD1BWP12T U62 ( .I(n2949), .ZN(n2825) );
  NR2D1BWP12T U63 ( .A1(n2115), .A2(n2310), .ZN(n2058) );
  AOI21D1BWP12T U64 ( .A1(n1424), .A2(n1423), .B(n1422), .ZN(n1428) );
  XNR2D1BWP12T U65 ( .A1(n1683), .A2(n1682), .ZN(n2671) );
  INVD1BWP12T U66 ( .I(n2115), .ZN(n2174) );
  FA1D0BWP12T U67 ( .A(n2725), .B(b[21]), .CI(n2335), .CO(n767), .S(n2716) );
  OAI211D1BWP12T U68 ( .A1(n2822), .A2(n852), .B(n851), .C(n850), .ZN(
        result[14]) );
  FA1D0BWP12T U69 ( .A(n2310), .B(n674), .CI(n2916), .CO(n2917), .S(n2398) );
  TPNR3D1BWP12T U70 ( .A1(op[2]), .A2(n535), .A3(n534), .ZN(n2967) );
  FA1D0BWP12T U71 ( .A(a[31]), .B(b[31]), .CI(n2918), .CO(n2919), .S(n632) );
  INVD1BWP12T U72 ( .I(n2878), .ZN(n2940) );
  FA1D0BWP12T U73 ( .A(n2310), .B(b[31]), .CI(n2658), .CO(n2659), .S(n2471) );
  FA1D0BWP12T U74 ( .A(a[29]), .B(n2292), .CI(n1497), .CO(n1349), .S(n2461) );
  FA1D0BWP12T U75 ( .A(n2310), .B(b[31]), .CI(n2660), .CO(n2661), .S(n2463) );
  FA1D0BWP12T U76 ( .A(a[30]), .B(b[30]), .CI(n1350), .CO(n2918), .S(n1805) );
  FA1D0BWP12T U77 ( .A(a[28]), .B(b[28]), .CI(n1456), .CO(n1498), .S(n1803) );
  FA1D0BWP12T U78 ( .A(a[29]), .B(b[29]), .CI(n1498), .CO(n1350), .S(n1804) );
  INVD1BWP12T U79 ( .I(n632), .ZN(n2466) );
  FA1D0BWP12T U80 ( .A(a[25]), .B(n2269), .CI(n732), .CO(n1591), .S(n1656) );
  FA1D0BWP12T U81 ( .A(mult_x_18_n385), .B(mult_x_18_n363), .CI(n2593), .CO(
        n2655), .S(n2656) );
  MAOI22D0BWP12T U82 ( .A1(n2173), .A2(n985), .B1(n2119), .B2(n994), .ZN(n1)
         );
  CKND2D0BWP12T U83 ( .A1(n2170), .A2(n999), .ZN(n2) );
  OAI211D0BWP12T U84 ( .A1(n2116), .A2(n986), .B(n1), .C(n2), .ZN(n2139) );
  CKND2D0BWP12T U85 ( .A1(n2142), .A2(n1999), .ZN(n3) );
  AOI222D0BWP12T U86 ( .A1(n2002), .A2(n2140), .B1(n2000), .B2(n2143), .C1(
        n2001), .C2(n2141), .ZN(n4) );
  AOI21D0BWP12T U87 ( .A1(n3), .A2(n4), .B(n2025), .ZN(n5) );
  AOI211D0BWP12T U88 ( .A1(n1966), .A2(n2033), .B(n2006), .C(n5), .ZN(n6) );
  OAI21D0BWP12T U89 ( .A1(n1997), .A2(n2510), .B(n6), .ZN(n2802) );
  CKND2D0BWP12T U90 ( .A1(n953), .A2(n954), .ZN(n7) );
  MAOI22D0BWP12T U91 ( .A1(n955), .A2(n7), .B1(n955), .B2(n7), .ZN(n2380) );
  NR2D0BWP12T U92 ( .A1(n1934), .A2(n1926), .ZN(n8) );
  AOI211D0BWP12T U93 ( .A1(n1929), .A2(n1920), .B(n8), .C(n2868), .ZN(n9) );
  OA21D0BWP12T U94 ( .A1(n1919), .A2(n2827), .B(n9), .Z(n2896) );
  CKND2D0BWP12T U95 ( .A1(n1434), .A2(n1430), .ZN(n10) );
  MAOI22D0BWP12T U96 ( .A1(n1435), .A2(n10), .B1(n1435), .B2(n10), .ZN(n2454)
         );
  CKND0BWP12T U97 ( .I(n1749), .ZN(n11) );
  INR3D0BWP12T U98 ( .A1(n635), .B1(n1772), .B2(n1748), .ZN(n12) );
  AOI211D0BWP12T U99 ( .A1(n635), .A2(n11), .B(n12), .C(n1751), .ZN(n13) );
  CKND2D0BWP12T U100 ( .A1(n2346), .A2(n2347), .ZN(n14) );
  MAOI22D0BWP12T U101 ( .A1(n13), .A2(n14), .B1(n13), .B2(n14), .ZN(n2888) );
  IAO21D0BWP12T U102 ( .A1(n1707), .A2(n1708), .B(n1709), .ZN(n2473) );
  CKND2D0BWP12T U103 ( .A1(n1595), .A2(n1594), .ZN(n15) );
  MOAI22D0BWP12T U104 ( .A1(n1596), .A2(n15), .B1(n1596), .B2(n15), .ZN(n2695)
         );
  CKND0BWP12T U105 ( .I(n2814), .ZN(n16) );
  AOI22D0BWP12T U106 ( .A1(n2967), .A2(n2702), .B1(n2701), .B2(n16), .ZN(n17)
         );
  OAI21D0BWP12T U107 ( .A1(a[18]), .A2(n2944), .B(n2949), .ZN(n18) );
  AOI22D0BWP12T U108 ( .A1(b[18]), .A2(n18), .B1(n2704), .B2(n2786), .ZN(n19)
         );
  MOAI22D0BWP12T U109 ( .A1(n2703), .A2(n2951), .B1(n2703), .B2(n2948), .ZN(
        n20) );
  CKND0BWP12T U110 ( .I(n2705), .ZN(n21) );
  OAI32D0BWP12T U111 ( .A1(n2705), .A2(n2825), .A3(n20), .B1(n2947), .B2(n21), 
        .ZN(n22) );
  AOI22D0BWP12T U112 ( .A1(n2706), .A2(n2775), .B1(n2940), .B2(n2709), .ZN(n23) );
  AOI22D0BWP12T U113 ( .A1(n2707), .A2(n2905), .B1(n2866), .B2(n2710), .ZN(n24) );
  AN4D0BWP12T U114 ( .A1(n19), .A2(n22), .A3(n23), .A4(n24), .Z(n25) );
  OA211D0BWP12T U115 ( .A1(n2708), .A2(n2964), .B(n17), .C(n25), .Z(n2713) );
  OA22D0BWP12T U116 ( .A1(n2603), .A2(n1320), .B1(n2604), .B2(n1321), .Z(n26)
         );
  OA22D0BWP12T U117 ( .A1(n2647), .A2(n1322), .B1(n2649), .B2(n1323), .Z(n27)
         );
  NR2D0BWP12T U118 ( .A1(n26), .A2(n27), .ZN(mult_x_18_n536) );
  MAOI22D0BWP12T U119 ( .A1(n26), .A2(n27), .B1(n26), .B2(n27), .ZN(
        mult_x_18_n537) );
  OA22D0BWP12T U120 ( .A1(n2052), .A2(n1862), .B1(n1861), .B2(n1926), .Z(n2055) );
  CKND0BWP12T U121 ( .I(n2165), .ZN(n28) );
  AOI22D0BWP12T U122 ( .A1(n2173), .A2(n2172), .B1(n2170), .B2(n2171), .ZN(n29) );
  AOI22D0BWP12T U123 ( .A1(n2169), .A2(n2168), .B1(n2166), .B2(n2167), .ZN(n30) );
  AO21D0BWP12T U124 ( .A1(n29), .A2(n30), .B(n2202), .Z(n31) );
  OAI31D0BWP12T U125 ( .A1(n2200), .A2(n2175), .A3(n28), .B(n31), .ZN(n32) );
  AOI211D0BWP12T U126 ( .A1(n2868), .A2(n2902), .B(n2174), .C(n32), .ZN(n2787)
         );
  CKND2D0BWP12T U127 ( .A1(n2342), .A2(n2341), .ZN(n33) );
  MOAI22D0BWP12T U128 ( .A1(n2343), .A2(n33), .B1(n2343), .B2(n33), .ZN(n2693)
         );
  AOI222D0BWP12T U129 ( .A1(n1999), .A2(n987), .B1(n2001), .B2(n986), .C1(
        n2000), .C2(n1000), .ZN(n34) );
  IOA21D0BWP12T U130 ( .A1(n2002), .A2(n994), .B(n34), .ZN(n2526) );
  CKND2D0BWP12T U131 ( .A1(n848), .A2(n847), .ZN(n35) );
  MOAI22D0BWP12T U132 ( .A1(n849), .A2(n35), .B1(n849), .B2(n35), .ZN(n2455)
         );
  CKND2D0BWP12T U133 ( .A1(n2349), .A2(n2348), .ZN(n36) );
  MOAI22D0BWP12T U134 ( .A1(n1747), .A2(n36), .B1(n1747), .B2(n36), .ZN(n2515)
         );
  CKND2D0BWP12T U135 ( .A1(n869), .A2(n868), .ZN(n37) );
  MOAI22D0BWP12T U136 ( .A1(n1709), .A2(n37), .B1(n1709), .B2(n37), .ZN(n1710)
         );
  CKND2D0BWP12T U137 ( .A1(n1561), .A2(n1557), .ZN(n38) );
  MOAI22D0BWP12T U138 ( .A1(n1558), .A2(n38), .B1(n1558), .B2(n38), .ZN(n1607)
         );
  IAO21D0BWP12T U139 ( .A1(n1933), .A2(n1851), .B(n1574), .ZN(n1859) );
  CKND0BWP12T U140 ( .I(n2025), .ZN(n39) );
  CKND0BWP12T U141 ( .I(n2017), .ZN(n40) );
  AOI22D0BWP12T U142 ( .A1(n1966), .A2(n39), .B1(n1948), .B2(n40), .ZN(n41) );
  OA211D0BWP12T U143 ( .A1(n1997), .A2(n2829), .B(n2014), .C(n41), .Z(n1989)
         );
  CKND2D0BWP12T U144 ( .A1(n1417), .A2(n1418), .ZN(n42) );
  MAOI22D0BWP12T U145 ( .A1(n1397), .A2(n42), .B1(n1397), .B2(n42), .ZN(n2383)
         );
  CKND0BWP12T U146 ( .I(n2639), .ZN(n43) );
  OAI222D0BWP12T U147 ( .A1(n43), .A2(n901), .B1(n2126), .B2(n2118), .C1(n763), 
        .C2(n2116), .ZN(n44) );
  IAO21D0BWP12T U148 ( .A1(n2128), .A2(n2117), .B(n44), .ZN(n2581) );
  CKND2D0BWP12T U149 ( .A1(n2415), .A2(n1595), .ZN(n45) );
  MAOI22D0BWP12T U150 ( .A1(n2416), .A2(n45), .B1(n2416), .B2(n45), .ZN(n2692)
         );
  CKND2D0BWP12T U151 ( .A1(n1012), .A2(n1011), .ZN(n46) );
  MOAI22D0BWP12T U152 ( .A1(n1010), .A2(n46), .B1(n1010), .B2(n46), .ZN(n1792)
         );
  CKND2D0BWP12T U153 ( .A1(n1685), .A2(n1684), .ZN(n47) );
  MOAI22D0BWP12T U154 ( .A1(n1686), .A2(n47), .B1(n1686), .B2(n47), .ZN(n2504)
         );
  CKND2D0BWP12T U155 ( .A1(n924), .A2(n921), .ZN(n48) );
  MAOI22D0BWP12T U156 ( .A1(n925), .A2(n48), .B1(n925), .B2(n48), .ZN(n1600)
         );
  MUX2ND0BWP12T U157 ( .I0(n2948), .I1(n2478), .S(n2231), .ZN(n49) );
  AOI31D0BWP12T U158 ( .A1(n2949), .A2(n49), .A3(n2878), .B(n2603), .ZN(n50)
         );
  OAI22D0BWP12T U159 ( .A1(n2302), .A2(n2806), .B1(n2285), .B2(n2949), .ZN(n51) );
  AOI211D0BWP12T U160 ( .A1(n2258), .A2(n2480), .B(n50), .C(n51), .ZN(n52) );
  CKND0BWP12T U161 ( .I(n2822), .ZN(n53) );
  AOI22D0BWP12T U162 ( .A1(n2358), .A2(n2967), .B1(n1711), .B2(n53), .ZN(n54)
         );
  OAI211D0BWP12T U163 ( .A1(n2964), .A2(n1975), .B(n52), .C(n54), .ZN(n55) );
  AOI22D0BWP12T U164 ( .A1(n1562), .A2(n2893), .B1(n2858), .B2(n1758), .ZN(n56) );
  CKND2D0BWP12T U165 ( .A1(n1607), .A2(n2855), .ZN(n57) );
  OAI211D0BWP12T U166 ( .A1(n2901), .A2(n2194), .B(n56), .C(n57), .ZN(n58) );
  AOI211D0BWP12T U167 ( .A1(n2425), .A2(n2866), .B(n55), .C(n58), .ZN(n59) );
  OAI21D0BWP12T U168 ( .A1(n2058), .A2(n1922), .B(n2905), .ZN(n60) );
  OAI211D0BWP12T U169 ( .A1(n2061), .A2(n2495), .B(n59), .C(n60), .ZN(
        result[0]) );
  OAI22D0BWP12T U170 ( .A1(n1881), .A2(n1933), .B1(n1882), .B2(n1930), .ZN(n61) );
  IAO21D0BWP12T U171 ( .A1(n1927), .A2(n2052), .B(n61), .ZN(n62) );
  OA211D0BWP12T U172 ( .A1(n1883), .A2(n1926), .B(n2870), .C(n62), .Z(n2053)
         );
  CKND2D0BWP12T U173 ( .A1(n1441), .A2(n1442), .ZN(n63) );
  MAOI22D0BWP12T U174 ( .A1(n2626), .A2(n63), .B1(n2626), .B2(n63), .ZN(n1826)
         );
  AOI222D0BWP12T U175 ( .A1(n2002), .A2(n2172), .B1(n2000), .B2(n2168), .C1(
        n2001), .C2(n2171), .ZN(n64) );
  CKND2D0BWP12T U176 ( .A1(n2167), .A2(n1999), .ZN(n65) );
  AOI21D0BWP12T U177 ( .A1(n65), .A2(n64), .B(n2025), .ZN(n66) );
  AOI211D0BWP12T U178 ( .A1(n1991), .A2(n2033), .B(n2006), .C(n66), .ZN(n67)
         );
  OAI21D0BWP12T U179 ( .A1(n1997), .A2(n2904), .B(n67), .ZN(n2772) );
  AOI21D0BWP12T U180 ( .A1(n2370), .A2(n2374), .B(n2371), .ZN(n68) );
  CKND2D0BWP12T U181 ( .A1(n2372), .A2(n2351), .ZN(n69) );
  MAOI22D0BWP12T U182 ( .A1(n68), .A2(n69), .B1(n68), .B2(n69), .ZN(n2587) );
  CKND2D0BWP12T U183 ( .A1(n1394), .A2(n1393), .ZN(n70) );
  MOAI22D0BWP12T U184 ( .A1(n1395), .A2(n70), .B1(n1395), .B2(n70), .ZN(n2453)
         );
  CKND2D0BWP12T U185 ( .A1(n1438), .A2(n1437), .ZN(n71) );
  MOAI22D0BWP12T U186 ( .A1(n1436), .A2(n71), .B1(n1436), .B2(n71), .ZN(n1790)
         );
  CKND2D0BWP12T U187 ( .A1(n1661), .A2(n1663), .ZN(n72) );
  MOAI22D0BWP12T U188 ( .A1(n1662), .A2(n72), .B1(n1662), .B2(n72), .ZN(n2767)
         );
  CKND2D0BWP12T U189 ( .A1(n809), .A2(n808), .ZN(n73) );
  MOAI22D0BWP12T U190 ( .A1(n810), .A2(n73), .B1(n810), .B2(n73), .ZN(n1651)
         );
  IOA21D0BWP12T U191 ( .A1(n1891), .A2(n2079), .B(n2046), .ZN(n2746) );
  OA22D0BWP12T U192 ( .A1(n2603), .A2(n1086), .B1(n2604), .B2(n1183), .Z(n74)
         );
  OA22D0BWP12T U193 ( .A1(n2647), .A2(n1251), .B1(n2649), .B2(n1180), .Z(n75)
         );
  NR2D0BWP12T U194 ( .A1(n74), .A2(n75), .ZN(mult_x_18_n465) );
  MAOI22D0BWP12T U195 ( .A1(n74), .A2(n75), .B1(n74), .B2(n75), .ZN(
        mult_x_18_n466) );
  IND2D0BWP12T U196 ( .A1(n2482), .B1(n2603), .ZN(n906) );
  IAO21D0BWP12T U197 ( .A1(n2870), .A2(n950), .B(n951), .ZN(n1902) );
  CKND2D0BWP12T U198 ( .A1(n2412), .A2(n2411), .ZN(n76) );
  MOAI22D0BWP12T U199 ( .A1(n2413), .A2(n76), .B1(n2413), .B2(n76), .ZN(n2710)
         );
  CKND2D0BWP12T U200 ( .A1(n818), .A2(n819), .ZN(n77) );
  MAOI22D0BWP12T U201 ( .A1(n817), .A2(n77), .B1(n817), .B2(n77), .ZN(n1791)
         );
  OAI21D0BWP12T U202 ( .A1(n1664), .A2(n1665), .B(n1663), .ZN(n78) );
  CKND2D0BWP12T U203 ( .A1(n1666), .A2(n1667), .ZN(n79) );
  MOAI22D0BWP12T U204 ( .A1(n78), .A2(n79), .B1(n78), .B2(n79), .ZN(n2799) );
  CKND0BWP12T U205 ( .I(n1799), .ZN(n80) );
  MOAI22D0BWP12T U206 ( .A1(n2065), .A2(n2718), .B1(n2786), .B2(n2196), .ZN(
        n81) );
  AOI21D0BWP12T U207 ( .A1(n737), .A2(n2948), .B(n2825), .ZN(n82) );
  OAI32D0BWP12T U208 ( .A1(n2232), .A2(n737), .A3(n2951), .B1(n82), .B2(n2232), 
        .ZN(n83) );
  AOI211D0BWP12T U209 ( .A1(n2569), .A2(n2932), .B(n2807), .C(n83), .ZN(n84)
         );
  OAI21D0BWP12T U210 ( .A1(n2944), .A2(a[22]), .B(n2949), .ZN(n85) );
  AOI22D0BWP12T U211 ( .A1(b[22]), .A2(n85), .B1(n2232), .B2(n2947), .ZN(n86)
         );
  OAI211D0BWP12T U212 ( .A1(n2038), .A2(n2964), .B(n84), .C(n86), .ZN(n87) );
  AOI211D0BWP12T U213 ( .A1(n1839), .A2(n2940), .B(n81), .C(n87), .ZN(n88) );
  CKND2D0BWP12T U214 ( .A1(n2967), .A2(n2389), .ZN(n89) );
  OAI211D0BWP12T U215 ( .A1(n2814), .A2(n80), .B(n88), .C(n89), .ZN(n768) );
  OAI21D0BWP12T U216 ( .A1(n1639), .A2(n1635), .B(n1636), .ZN(n90) );
  AOI21D0BWP12T U217 ( .A1(n424), .A2(n90), .B(n1638), .ZN(n91) );
  CKND2D0BWP12T U218 ( .A1(n1641), .A2(n2449), .ZN(n92) );
  MAOI22D0BWP12T U219 ( .A1(n91), .A2(n92), .B1(n91), .B2(n92), .ZN(n2913) );
  CKND2D0BWP12T U220 ( .A1(n2376), .A2(n1774), .ZN(n93) );
  AOI21D0BWP12T U221 ( .A1(n2370), .A2(n2374), .B(n2371), .ZN(n94) );
  OAI21D0BWP12T U222 ( .A1(n2373), .A2(n94), .B(n2372), .ZN(n95) );
  MOAI22D0BWP12T U223 ( .A1(n93), .A2(n95), .B1(n93), .B2(n95), .ZN(n2536) );
  OA22D0BWP12T U224 ( .A1(n2603), .A2(n1316), .B1(n2604), .B2(n1317), .Z(n96)
         );
  OA22D0BWP12T U225 ( .A1(n2647), .A2(n1318), .B1(n2649), .B2(n1319), .Z(n97)
         );
  NR2D0BWP12T U226 ( .A1(n96), .A2(n97), .ZN(mult_x_18_n502) );
  MAOI22D0BWP12T U227 ( .A1(n96), .A2(n97), .B1(n96), .B2(n97), .ZN(
        mult_x_18_n503) );
  CMPE42D1BWP12T U228 ( .A(mult_x_18_n932), .B(mult_x_18_n761), .C(
        mult_x_18_n817), .CIX(mult_x_18_n530), .D(mult_x_18_n880), .CO(
        mult_x_18_n514), .COX(mult_x_18_n513), .S(mult_x_18_n515) );
  INR3D0BWP12T U229 ( .A1(n1832), .B1(n2830), .B2(n906), .ZN(n1573) );
  MAOI22D0BWP12T U230 ( .A1(n1885), .A2(n1443), .B1(n1994), .B2(n2964), .ZN(
        n98) );
  OAI21D0BWP12T U231 ( .A1(n2944), .A2(a[14]), .B(n2949), .ZN(n99) );
  AOI22D0BWP12T U232 ( .A1(b[14]), .A2(n99), .B1(n1441), .B2(n2947), .ZN(n100)
         );
  CKND2D0BWP12T U233 ( .A1(n2275), .A2(n2948), .ZN(n101) );
  OAI211D0BWP12T U234 ( .A1(n2951), .A2(n2275), .B(n2949), .C(n101), .ZN(n102)
         );
  AOI22D0BWP12T U235 ( .A1(a[14]), .A2(n102), .B1(n1837), .B2(n2940), .ZN(n103) );
  OA211D0BWP12T U236 ( .A1(n2942), .A2(n2208), .B(n100), .C(n103), .Z(n104) );
  OAI211D0BWP12T U237 ( .A1(n2071), .A2(n2957), .B(n98), .C(n104), .ZN(n841)
         );
  OA222D0BWP12T U238 ( .A1(n1890), .A2(n1926), .B1(n1861), .B2(n1930), .C1(
        n1862), .C2(n1933), .Z(n105) );
  OA211D0BWP12T U239 ( .A1(n1889), .A2(n2052), .B(n105), .C(n2870), .Z(n537)
         );
  CKND2D0BWP12T U240 ( .A1(n2342), .A2(n2341), .ZN(n106) );
  MOAI22D0BWP12T U241 ( .A1(n1746), .A2(n106), .B1(n1746), .B2(n106), .ZN(
        n2694) );
  CKND2D0BWP12T U242 ( .A1(n970), .A2(n969), .ZN(n107) );
  MOAI22D0BWP12T U243 ( .A1(n971), .A2(n107), .B1(n971), .B2(n107), .ZN(n1716)
         );
  OAI211D1BWP12T U244 ( .A1(n2466), .A2(n2814), .B(n683), .C(n682), .ZN(n108)
         );
  AOI21D0BWP12T U245 ( .A1(n2463), .A2(n2866), .B(n108), .ZN(n109) );
  CKND2D0BWP12T U246 ( .A1(n2855), .A2(n2471), .ZN(n110) );
  OAI211D1BWP12T U247 ( .A1(n2822), .A2(n1742), .B(n109), .C(n110), .ZN(
        result[31]) );
  NR4D0BWP12T U248 ( .A1(n2867), .A2(n2559), .A3(n2444), .A4(n2523), .ZN(n111)
         );
  OR4D0BWP12T U249 ( .A1(n2424), .A2(n2973), .A3(n2491), .A4(n2425), .Z(n112)
         );
  NR4D0BWP12T U250 ( .A1(n2432), .A2(n2592), .A3(n2843), .A4(n112), .ZN(n113)
         );
  NR4D0BWP12T U251 ( .A1(n2884), .A2(n2516), .A3(n2418), .A4(n2417), .ZN(n114)
         );
  NR3D0BWP12T U252 ( .A1(n2453), .A2(n2455), .A3(n2454), .ZN(n115) );
  ND4D0BWP12T U253 ( .A1(n111), .A2(n113), .A3(n114), .A4(n115), .ZN(n116) );
  OR4D0BWP12T U254 ( .A1(n2710), .A2(n2456), .A3(n2692), .A4(n116), .Z(n117)
         );
  OR4D0BWP12T U255 ( .A1(n2736), .A2(n2457), .A3(n2926), .A4(n117), .Z(n118)
         );
  OR4D0BWP12T U256 ( .A1(n2458), .A2(n2939), .A3(n2762), .A4(n118), .Z(n119)
         );
  OR4D0BWP12T U257 ( .A1(n2459), .A2(n2796), .A3(n2817), .A4(n119), .Z(n2460)
         );
  CKND0BWP12T U258 ( .I(n2705), .ZN(n120) );
  NR2D0BWP12T U259 ( .A1(a[16]), .A2(n2679), .ZN(n121) );
  CKND2D0BWP12T U260 ( .A1(n121), .A2(n1405), .ZN(n122) );
  NR2D0BWP12T U261 ( .A1(n120), .A2(n122), .ZN(n788) );
  MAOI22D0BWP12T U262 ( .A1(n120), .A2(n122), .B1(n120), .B2(n122), .ZN(n2709)
         );
  IND2D0BWP12T U263 ( .A1(n2174), .B1(n2961), .ZN(n123) );
  AO21D0BWP12T U264 ( .A1(n2135), .A2(n123), .B(n2048), .Z(n2047) );
  IAO21D0BWP12T U265 ( .A1(n2871), .A2(n562), .B(n1589), .ZN(n2437) );
  IAO21D0BWP12T U266 ( .A1(n2482), .A2(n2231), .B(n2258), .ZN(n1000) );
  CKND2D0BWP12T U267 ( .A1(n1675), .A2(n1674), .ZN(n124) );
  MOAI22D0BWP12T U268 ( .A1(n1721), .A2(n124), .B1(n1721), .B2(n124), .ZN(
        n2700) );
  CKND2D0BWP12T U269 ( .A1(n921), .A2(n920), .ZN(n125) );
  MOAI22D0BWP12T U270 ( .A1(n922), .A2(n125), .B1(n922), .B2(n125), .ZN(n2417)
         );
  NR3D0BWP12T U271 ( .A1(n2935), .A2(n1797), .A3(n2715), .ZN(n126) );
  NR4D0BWP12T U272 ( .A1(n1759), .A2(n2490), .A3(n1758), .A4(n2814), .ZN(n127)
         );
  NR4D0BWP12T U273 ( .A1(n2859), .A2(n1767), .A3(n2888), .A4(n1753), .ZN(n128)
         );
  NR4D0BWP12T U274 ( .A1(n2846), .A2(n2541), .A3(n2561), .A4(n2588), .ZN(n129)
         );
  IND4D0BWP12T U275 ( .A1(n1789), .B1(n127), .B2(n128), .B3(n129), .ZN(n130)
         );
  NR4D0BWP12T U276 ( .A1(n2515), .A2(n1792), .A3(n1791), .A4(n130), .ZN(n131)
         );
  NR4D0BWP12T U277 ( .A1(n2701), .A2(n1795), .A3(n2694), .A4(n1790), .ZN(n132)
         );
  NR3D0BWP12T U278 ( .A1(n2969), .A2(n2741), .A3(n1799), .ZN(n133) );
  ND4D0BWP12T U279 ( .A1(n126), .A2(n131), .A3(n132), .A4(n133), .ZN(n134) );
  OR4D0BWP12T U280 ( .A1(n2768), .A2(n2800), .A3(n1801), .A4(n134), .Z(n1802)
         );
  CMPE42D1BWP12T U281 ( .A(mult_x_18_n842), .B(mult_x_18_n806), .C(
        mult_x_18_n886), .CIX(mult_x_18_n615), .D(mult_x_18_n911), .CO(
        mult_x_18_n604), .COX(mult_x_18_n603), .S(mult_x_18_n605) );
  CKND2D0BWP12T U282 ( .A1(n2242), .A2(n976), .ZN(n135) );
  MAOI22D0BWP12T U283 ( .A1(n2643), .A2(n135), .B1(n2643), .B2(n135), .ZN(
        n1836) );
  NR2D0BWP12T U284 ( .A1(n1884), .A2(n1886), .ZN(n136) );
  OAI22D0BWP12T U285 ( .A1(n2842), .A2(n136), .B1(n1949), .B2(n2964), .ZN(n137) );
  OAI21D0BWP12T U286 ( .A1(n2944), .A2(n2626), .B(n2949), .ZN(n138) );
  AOI22D0BWP12T U287 ( .A1(b[15]), .A2(n138), .B1(n2240), .B2(n2947), .ZN(n139) );
  OAI21D0BWP12T U288 ( .A1(n2276), .A2(n2951), .B(n2949), .ZN(n140) );
  AOI32D0BWP12T U289 ( .A1(n2948), .A2(n2626), .A3(n2276), .B1(n140), .B2(
        n2626), .ZN(n141) );
  OAI211D0BWP12T U290 ( .A1(n2942), .A2(n2206), .B(n139), .C(n141), .ZN(n142)
         );
  AOI211D0BWP12T U291 ( .A1(n2940), .A2(n1826), .B(n137), .C(n142), .ZN(n143)
         );
  OA21D0BWP12T U292 ( .A1(n2070), .A2(n2957), .B(n143), .Z(n1449) );
  OA222D0BWP12T U293 ( .A1(n1903), .A2(n1930), .B1(n1904), .B2(n2052), .C1(
        n1914), .C2(n1926), .Z(n144) );
  OA211D0BWP12T U294 ( .A1(n1912), .A2(n1933), .B(n144), .C(n2870), .Z(n2048)
         );
  CKND2D0BWP12T U295 ( .A1(n1423), .A2(n815), .ZN(n145) );
  MOAI22D0BWP12T U296 ( .A1(n1424), .A2(n145), .B1(n1424), .B2(n145), .ZN(
        n1717) );
  CKND2D0BWP12T U297 ( .A1(n1647), .A2(n2412), .ZN(n146) );
  MAOI22D0BWP12T U298 ( .A1(n1648), .A2(n146), .B1(n1648), .B2(n146), .ZN(
        n2711) );
  CKND2D0BWP12T U299 ( .A1(n2443), .A2(n1618), .ZN(n147) );
  AOI21D0BWP12T U300 ( .A1(n2437), .A2(n2441), .B(n2438), .ZN(n148) );
  OAI21D0BWP12T U301 ( .A1(n2440), .A2(n148), .B(n2439), .ZN(n149) );
  MOAI22D0BWP12T U302 ( .A1(n147), .A2(n149), .B1(n147), .B2(n149), .ZN(n2523)
         );
  CKND2D0BWP12T U303 ( .A1(n1577), .A2(n1585), .ZN(n150) );
  IOA21D0BWP12T U304 ( .A1(n2374), .A2(n1764), .B(n2366), .ZN(n151) );
  MOAI22D0BWP12T U305 ( .A1(n150), .A2(n151), .B1(n150), .B2(n151), .ZN(n2365)
         );
  CMPE42D1BWP12T U306 ( .A(mult_x_18_n998), .B(mult_x_18_n791), .C(
        mult_x_18_n967), .CIX(mult_x_18_n618), .D(mult_x_18_n620), .CO(
        mult_x_18_n607), .COX(mult_x_18_n606), .S(mult_x_18_n608) );
  INR2D0BWP12T U307 ( .A1(n833), .B1(n834), .ZN(n976) );
  NR2D0BWP12T U308 ( .A1(a[16]), .A2(n1830), .ZN(n152) );
  MOAI22D0BWP12T U309 ( .A1(n2679), .A2(n152), .B1(n2679), .B2(n152), .ZN(
        n2672) );
  CKND0BWP12T U310 ( .I(n2868), .ZN(n153) );
  OAI21D0BWP12T U311 ( .A1(a[31]), .A2(n153), .B(n2115), .ZN(n2068) );
  MOAI22D0BWP12T U312 ( .A1(n2639), .A2(n870), .B1(n2639), .B2(n876), .ZN(
        n2770) );
  OAI21D0BWP12T U313 ( .A1(n2345), .A2(n2369), .B(n2344), .ZN(n154) );
  CKND2D0BWP12T U314 ( .A1(n2346), .A2(n2347), .ZN(n155) );
  MOAI22D0BWP12T U315 ( .A1(n154), .A2(n155), .B1(n154), .B2(n155), .ZN(n2892)
         );
  CKND2D0BWP12T U316 ( .A1(n1561), .A2(n1560), .ZN(n156) );
  MOAI22D0BWP12T U317 ( .A1(n2231), .A2(n156), .B1(n2231), .B2(n156), .ZN(
        n1758) );
  OAI21D0BWP12T U318 ( .A1(n2944), .A2(a[20]), .B(n2949), .ZN(n157) );
  AOI22D0BWP12T U319 ( .A1(b[20]), .A2(n157), .B1(n2929), .B2(n2947), .ZN(n158) );
  OAI21D0BWP12T U320 ( .A1(n2410), .A2(n2951), .B(n2949), .ZN(n159) );
  AOI32D0BWP12T U321 ( .A1(n2948), .A2(a[20]), .A3(n2410), .B1(n159), .B2(
        a[20]), .ZN(n160) );
  OAI211D0BWP12T U322 ( .A1(n2942), .A2(n2930), .B(n158), .C(n160), .ZN(n161)
         );
  MAOI22D0BWP12T U323 ( .A1(n2940), .A2(n2927), .B1(n2957), .B2(n2933), .ZN(
        n162) );
  CKND2D0BWP12T U324 ( .A1(n2931), .A2(n2932), .ZN(n163) );
  OAI211D0BWP12T U325 ( .A1(n2928), .A2(n2964), .B(n162), .C(n163), .ZN(n164)
         );
  AOI211D0BWP12T U326 ( .A1(n2967), .A2(n2934), .B(n161), .C(n164), .ZN(n2936)
         );
  CKND2D0BWP12T U327 ( .A1(n1598), .A2(n1597), .ZN(n165) );
  MOAI22D0BWP12T U328 ( .A1(n1599), .A2(n165), .B1(n1599), .B2(n165), .ZN(
        n2517) );
  OA222D0BWP12T U329 ( .A1(n1889), .A2(n1926), .B1(n1862), .B2(n1930), .C1(
        n1890), .C2(n1933), .Z(n166) );
  OA211D0BWP12T U330 ( .A1(n1897), .A2(n2052), .B(n166), .C(n2870), .Z(n1977)
         );
  OR4D0BWP12T U331 ( .A1(n2822), .A2(n1710), .A3(n2473), .A4(n1711), .Z(n167)
         );
  OR4D0BWP12T U332 ( .A1(n1712), .A2(n2883), .A3(n2854), .A4(n167), .Z(n168)
         );
  OR4D0BWP12T U333 ( .A1(n2568), .A2(n1713), .A3(n2542), .A4(n168), .Z(n169)
         );
  NR4D0BWP12T U334 ( .A1(n2567), .A2(n1714), .A3(n2915), .A4(n169), .ZN(n170)
         );
  NR3D0BWP12T U335 ( .A1(n1715), .A2(n1716), .A3(n2504), .ZN(n171) );
  NR3D0BWP12T U336 ( .A1(n1718), .A2(n1717), .A3(n2671), .ZN(n172) );
  ND4D0BWP12T U337 ( .A1(n427), .A2(n170), .A3(n171), .A4(n172), .ZN(n173) );
  OR4D0BWP12T U338 ( .A1(n2700), .A2(n2938), .A3(n1726), .A4(n173), .Z(n174)
         );
  OR4D0BWP12T U339 ( .A1(n2978), .A2(n1735), .A3(n2740), .A4(n174), .Z(n175)
         );
  OR4D0BWP12T U340 ( .A1(n2767), .A2(n1736), .A3(n2799), .A4(n175), .Z(n1737)
         );
  NR2D0BWP12T U341 ( .A1(n2636), .A2(n2231), .ZN(n176) );
  MAOI22D0BWP12T U342 ( .A1(a[29]), .A2(n176), .B1(n2248), .B2(n2638), .ZN(
        n275) );
  CMPE42D1BWP12T U343 ( .A(mult_x_18_n931), .B(mult_x_18_n716), .C(
        mult_x_18_n816), .CIX(mult_x_18_n513), .D(mult_x_18_n835), .CO(
        mult_x_18_n495), .COX(mult_x_18_n494), .S(mult_x_18_n496) );
  OAI22D0BWP12T U344 ( .A1(n471), .A2(n2098), .B1(n2639), .B2(n2097), .ZN(n177) );
  OAI21D0BWP12T U345 ( .A1(n2831), .A2(n177), .B(n2099), .ZN(n2782) );
  AOI21D0BWP12T U346 ( .A1(n2368), .A2(n633), .B(n634), .ZN(n178) );
  IOA21D0BWP12T U347 ( .A1(n533), .A2(b[9]), .B(n635), .ZN(n179) );
  MAOI22D0BWP12T U348 ( .A1(n178), .A2(n179), .B1(n178), .B2(n179), .ZN(n2377)
         );
  IND2D0BWP12T U349 ( .A1(n2620), .B1(n2869), .ZN(n1820) );
  CKND2D0BWP12T U350 ( .A1(n1832), .A2(n1833), .ZN(n180) );
  MAOI22D0BWP12T U351 ( .A1(n2830), .A2(n180), .B1(n2830), .B2(n180), .ZN(
        n2845) );
  CKND2D0BWP12T U352 ( .A1(n1417), .A2(n1418), .ZN(n181) );
  MAOI22D0BWP12T U353 ( .A1(n1419), .A2(n181), .B1(n1419), .B2(n181), .ZN(
        n1795) );
  CKND2D0BWP12T U354 ( .A1(n1669), .A2(n734), .ZN(n182) );
  MOAI22D0BWP12T U355 ( .A1(n1670), .A2(n182), .B1(n1670), .B2(n182), .ZN(
        n1735) );
  CKND2D0BWP12T U356 ( .A1(n782), .A2(n2948), .ZN(n183) );
  OAI211D0BWP12T U357 ( .A1(n2951), .A2(n782), .B(n2949), .C(n183), .ZN(n184)
         );
  AOI22D0BWP12T U358 ( .A1(n1866), .A2(n2932), .B1(n2091), .B2(n1373), .ZN(
        n185) );
  OAI21D0BWP12T U359 ( .A1(n2944), .A2(n2609), .B(n2949), .ZN(n186) );
  MAOI22D0BWP12T U360 ( .A1(b[19]), .A2(n186), .B1(n2609), .B2(n2806), .ZN(
        n187) );
  OAI211D0BWP12T U361 ( .A1(n2942), .A2(n2190), .B(n185), .C(n187), .ZN(n188)
         );
  AOI211D0BWP12T U362 ( .A1(n2609), .A2(n184), .B(n2807), .C(n188), .ZN(n189)
         );
  CKND0BWP12T U363 ( .I(n2964), .ZN(n190) );
  AOI22D0BWP12T U364 ( .A1(n1827), .A2(n2940), .B1(n1989), .B2(n190), .ZN(n191) );
  CKND0BWP12T U365 ( .I(n2814), .ZN(n192) );
  AOI22D0BWP12T U366 ( .A1(n2967), .A2(n2387), .B1(n1797), .B2(n192), .ZN(n193) );
  ND3D0BWP12T U367 ( .A1(n189), .A2(n191), .A3(n193), .ZN(n807) );
  NR4D0BWP12T U368 ( .A1(n1600), .A2(n2517), .A3(n1642), .A4(n2913), .ZN(n194)
         );
  NR4D0BWP12T U369 ( .A1(n1606), .A2(n2476), .A3(n1607), .A4(n2657), .ZN(n195)
         );
  NR2D0BWP12T U370 ( .A1(n2856), .A2(n2539), .ZN(n196) );
  NR4D0BWP12T U371 ( .A1(n1634), .A2(n2570), .A3(n2824), .A4(n2558), .ZN(n197)
         );
  ND4D0BWP12T U372 ( .A1(n194), .A2(n195), .A3(n196), .A4(n197), .ZN(n198) );
  OR4D0BWP12T U373 ( .A1(n1644), .A2(n1643), .A3(n1645), .A4(n198), .Z(n199)
         );
  OR4D0BWP12T U374 ( .A1(n1649), .A2(n2711), .A3(n2695), .A4(n199), .Z(n200)
         );
  OR4D0BWP12T U375 ( .A1(n2737), .A2(n1651), .A3(n2937), .A4(n200), .Z(n201)
         );
  OR4D0BWP12T U376 ( .A1(n2975), .A2(n2763), .A3(n1653), .A4(n201), .Z(n1655)
         );
  MAOI22D0BWP12T U377 ( .A1(n711), .A2(n2001), .B1(n1959), .B2(n792), .ZN(
        n2027) );
  CKND0BWP12T U378 ( .I(n2639), .ZN(n202) );
  CKND0BWP12T U379 ( .I(n471), .ZN(n203) );
  AOI22D0BWP12T U380 ( .A1(n1882), .A2(n202), .B1(n2051), .B2(n203), .ZN(n1852) );
  MUX2ND0BWP12T U381 ( .I0(n2184), .I1(n2189), .S(n2827), .ZN(n204) );
  NR2D0BWP12T U382 ( .A1(n2135), .A2(n204), .ZN(n2210) );
  CKND2D0BWP12T U383 ( .A1(n2367), .A2(n2368), .ZN(n205) );
  MAOI22D0BWP12T U384 ( .A1(n2369), .A2(n205), .B1(n2369), .B2(n205), .ZN(
        n2553) );
  MOAI22D0BWP12T U385 ( .A1(a[29]), .A2(n2868), .B1(a[29]), .B2(n2868), .ZN(
        n206) );
  OAI22D0BWP12T U386 ( .A1(n2638), .A2(n2637), .B1(n2636), .B2(n206), .ZN(n207) );
  MOAI22D0BWP12T U387 ( .A1(a[31]), .A2(n2639), .B1(a[31]), .B2(n2639), .ZN(
        n208) );
  OAI22D0BWP12T U388 ( .A1(n2642), .A2(n2641), .B1(n2640), .B2(n208), .ZN(n209) );
  MAOI22D0BWP12T U389 ( .A1(n207), .A2(n209), .B1(n207), .B2(n209), .ZN(n210)
         );
  MAOI22D0BWP12T U390 ( .A1(mult_x_18_n370), .A2(n210), .B1(mult_x_18_n370), 
        .B2(n210), .ZN(n211) );
  MOAI22D0BWP12T U391 ( .A1(n2643), .A2(b[20]), .B1(n2643), .B2(b[20]), .ZN(
        n212) );
  OAI22D0BWP12T U392 ( .A1(n2646), .A2(n2645), .B1(n2644), .B2(n212), .ZN(n213) );
  MOAI22D0BWP12T U393 ( .A1(n2679), .A2(b[16]), .B1(n2679), .B2(b[16]), .ZN(
        n214) );
  OAI22D0BWP12T U394 ( .A1(n2649), .A2(n2648), .B1(n2647), .B2(n214), .ZN(n215) );
  MOAI22D0BWP12T U395 ( .A1(n213), .A2(n215), .B1(n213), .B2(n215), .ZN(n216)
         );
  MOAI22D0BWP12T U396 ( .A1(n2830), .A2(b[30]), .B1(n2830), .B2(b[30]), .ZN(
        n217) );
  OAI22D0BWP12T U397 ( .A1(n2652), .A2(n2651), .B1(n2650), .B2(n217), .ZN(n218) );
  MAOI22D0BWP12T U398 ( .A1(n216), .A2(n218), .B1(n216), .B2(n218), .ZN(n219)
         );
  MAOI22D0BWP12T U399 ( .A1(n211), .A2(n219), .B1(n211), .B2(n219), .ZN(n220)
         );
  MAOI22D0BWP12T U400 ( .A1(mult_x_18_n380), .A2(n220), .B1(mult_x_18_n380), 
        .B2(n220), .ZN(n221) );
  MAOI22D0BWP12T U401 ( .A1(mult_x_18_n371), .A2(n221), .B1(mult_x_18_n371), 
        .B2(n221), .ZN(n2653) );
  OAI21D0BWP12T U402 ( .A1(n2944), .A2(a[27]), .B(n2949), .ZN(n222) );
  MAOI22D0BWP12T U403 ( .A1(b[27]), .A2(n222), .B1(a[27]), .B2(n2806), .ZN(
        n223) );
  CKND2D0BWP12T U404 ( .A1(n2805), .A2(n2948), .ZN(n224) );
  OAI211D0BWP12T U405 ( .A1(n2951), .A2(n2805), .B(n2949), .C(n224), .ZN(n225)
         );
  MOAI22D0BWP12T U406 ( .A1(n2957), .A2(n2803), .B1(n2804), .B2(n2932), .ZN(
        n226) );
  AOI211D0BWP12T U407 ( .A1(a[27]), .A2(n225), .B(n2807), .C(n226), .ZN(n227)
         );
  OAI211D0BWP12T U408 ( .A1(n2942), .A2(n2808), .B(n223), .C(n227), .ZN(n2809)
         );
  CKND0BWP12T U409 ( .I(n2449), .ZN(n228) );
  OA21D0BWP12T U410 ( .A1(n2447), .A2(n228), .B(n2448), .Z(n229) );
  OAI31D0BWP12T U411 ( .A1(n2450), .A2(n2446), .A3(n228), .B(n229), .ZN(n230)
         );
  CKND2D0BWP12T U412 ( .A1(n2452), .A2(n1598), .ZN(n231) );
  MOAI22D0BWP12T U413 ( .A1(n230), .A2(n231), .B1(n230), .B2(n231), .ZN(n2516)
         );
  CKND2D0BWP12T U414 ( .A1(n1688), .A2(n1687), .ZN(n232) );
  MOAI22D0BWP12T U415 ( .A1(n1689), .A2(n232), .B1(n1689), .B2(n232), .ZN(
        n2915) );
  INR3D0BWP12T U416 ( .A1(n2578), .B1(n1820), .B2(n1835), .ZN(n233) );
  MOAI22D0BWP12T U417 ( .A1(n2527), .A2(n233), .B1(n2527), .B2(n233), .ZN(
        n2522) );
  AOI21D0BWP12T U418 ( .A1(n1778), .A2(n1786), .B(n1780), .ZN(n234) );
  CKND2D0BWP12T U419 ( .A1(n1781), .A2(n1585), .ZN(n235) );
  MAOI22D0BWP12T U420 ( .A1(n234), .A2(n235), .B1(n234), .B2(n235), .ZN(n1767)
         );
  AOI21D0BWP12T U421 ( .A1(n2866), .A2(n2796), .B(n2795), .ZN(n236) );
  CKND2D0BWP12T U422 ( .A1(n2855), .A2(n2797), .ZN(n237) );
  OAI211D1BWP12T U423 ( .A1(n2822), .A2(n2798), .B(n236), .C(n237), .ZN(
        result[26]) );
  CMPE42D1BWP12T U424 ( .A(mult_x_18_n938), .B(mult_x_18_n863), .C(
        mult_x_18_n823), .CIX(mult_x_18_n608), .D(mult_x_18_n612), .CO(
        mult_x_18_n601), .COX(mult_x_18_n600), .S(mult_x_18_n602) );
  OA21D1BWP12T U425 ( .A1(n2097), .A2(n1933), .B(n1993), .Z(n875) );
  CKND0BWP12T U426 ( .I(a[31]), .ZN(n238) );
  MAOI22D0BWP12T U427 ( .A1(n2639), .A2(n238), .B1(n2639), .B2(n2098), .ZN(
        n822) );
  AOI22D0BWP12T U428 ( .A1(n2017), .A2(n1505), .B1(n1998), .B2(n2012), .ZN(
        n239) );
  AOI21D0BWP12T U429 ( .A1(n239), .A2(n1997), .B(n1901), .ZN(n1995) );
  OAI22D0BWP12T U430 ( .A1(n2603), .A2(n2602), .B1(n2604), .B2(n1037), .ZN(
        n240) );
  IND2D0BWP12T U431 ( .A1(n2231), .B1(a[31]), .ZN(n241) );
  OAI22D0BWP12T U432 ( .A1(n2310), .A2(n2642), .B1(n2640), .B2(n241), .ZN(n242) );
  MAOI22D0BWP12T U433 ( .A1(n240), .A2(n242), .B1(n240), .B2(n242), .ZN(
        mult_x_18_n383) );
  AN2D0BWP12T U434 ( .A1(n240), .A2(n242), .Z(n2625) );
  CKND2D0BWP12T U435 ( .A1(a[28]), .A2(a[29]), .ZN(n243) );
  OAI211D0BWP12T U436 ( .A1(a[28]), .A2(a[29]), .B(n2636), .C(n243), .ZN(n2638) );
  OAI22D0BWP12T U437 ( .A1(n2831), .A2(n2180), .B1(n2875), .B2(n2827), .ZN(
        n244) );
  NR2D0BWP12T U438 ( .A1(n2135), .A2(n244), .ZN(n2209) );
  MAOI22D0BWP12T U439 ( .A1(n2827), .A2(n2139), .B1(n2827), .B2(n2844), .ZN(
        n2514) );
  CKND2D0BWP12T U440 ( .A1(n1764), .A2(n2366), .ZN(n245) );
  MOAI22D0BWP12T U441 ( .A1(n2374), .A2(n245), .B1(n2374), .B2(n245), .ZN(
        n2857) );
  CKND2D0BWP12T U442 ( .A1(n953), .A2(n954), .ZN(n246) );
  MAOI22D0BWP12T U443 ( .A1(n946), .A2(n246), .B1(n946), .B2(n246), .ZN(n1789)
         );
  CKND0BWP12T U444 ( .I(n2973), .ZN(n247) );
  AOI222D0BWP12T U445 ( .A1(n1416), .A2(n2035), .B1(n2011), .B2(n2031), .C1(
        n2033), .C2(n2018), .ZN(n248) );
  MAOI22D0BWP12T U446 ( .A1(n2940), .A2(n1831), .B1(n2964), .B2(n248), .ZN(
        n249) );
  AOI22D0BWP12T U447 ( .A1(n1542), .A2(n2960), .B1(n2383), .B2(n2967), .ZN(
        n250) );
  OAI211D0BWP12T U448 ( .A1(n2207), .A2(n2942), .B(n249), .C(n250), .ZN(n251)
         );
  NR2D0BWP12T U449 ( .A1(n2951), .A2(n2270), .ZN(n252) );
  AOI211D0BWP12T U450 ( .A1(n2270), .A2(n2948), .B(n2825), .C(n252), .ZN(n253)
         );
  OAI21D0BWP12T U451 ( .A1(a[16]), .A2(n2944), .B(n2949), .ZN(n254) );
  AOI22D0BWP12T U452 ( .A1(b[16]), .A2(n254), .B1(n2947), .B2(n2235), .ZN(n255) );
  OAI211D0BWP12T U453 ( .A1(n2235), .A2(n253), .B(n2682), .C(n255), .ZN(n256)
         );
  AOI211D0BWP12T U454 ( .A1(n2453), .A2(n247), .B(n251), .C(n256), .ZN(n257)
         );
  IOA21D0BWP12T U455 ( .A1(n1795), .A2(n2858), .B(n257), .ZN(n1420) );
  CKND2D0BWP12T U456 ( .A1(n2899), .A2(n2948), .ZN(n258) );
  OAI211D0BWP12T U457 ( .A1(n2951), .A2(n2899), .B(n2949), .C(n258), .ZN(n259)
         );
  OAI21D0BWP12T U458 ( .A1(n2944), .A2(n2900), .B(n2949), .ZN(n260) );
  AOI22D0BWP12T U459 ( .A1(n2897), .A2(n260), .B1(n2898), .B2(n2947), .ZN(n261) );
  AOI21D0BWP12T U460 ( .A1(n2895), .A2(n2894), .B(n2893), .ZN(n262) );
  MAOI22D0BWP12T U461 ( .A1(n2904), .A2(n2903), .B1(n2896), .B2(n262), .ZN(
        n263) );
  OAI211D0BWP12T U462 ( .A1(n2902), .A2(n2901), .B(n261), .C(n263), .ZN(n264)
         );
  AOI21D0BWP12T U463 ( .A1(n2900), .A2(n259), .B(n264), .ZN(n2908) );
  OAI21D0BWP12T U464 ( .A1(n1635), .A2(n1639), .B(n1636), .ZN(n265) );
  CKND2D0BWP12T U465 ( .A1(n1637), .A2(n424), .ZN(n266) );
  MOAI22D0BWP12T U466 ( .A1(n265), .A2(n266), .B1(n265), .B2(n266), .ZN(n1642)
         );
  CKND2D0BWP12T U467 ( .A1(n1691), .A2(n1690), .ZN(n267) );
  MOAI22D0BWP12T U468 ( .A1(n1692), .A2(n267), .B1(n1692), .B2(n267), .ZN(
        n2567) );
  OA22D0BWP12T U469 ( .A1(n1925), .A2(n2052), .B1(n1924), .B2(n2827), .Z(n268)
         );
  OA211D0BWP12T U470 ( .A1(n1927), .A2(n1926), .B(n2870), .C(n268), .Z(n2540)
         );
  NR2D0BWP12T U471 ( .A1(n1820), .A2(n1835), .ZN(n269) );
  MOAI22D0BWP12T U472 ( .A1(n2574), .A2(n269), .B1(n2574), .B2(n269), .ZN(
        n2586) );
  CKND2D0BWP12T U473 ( .A1(n1590), .A2(n1587), .ZN(n270) );
  IOA21D0BWP12T U474 ( .A1(n2441), .A2(n1612), .B(n2433), .ZN(n271) );
  MOAI22D0BWP12T U475 ( .A1(n270), .A2(n271), .B1(n270), .B2(n271), .ZN(n2432)
         );
  AOI21D0BWP12T U476 ( .A1(n2866), .A2(n2458), .B(n731), .ZN(n272) );
  CKND2D0BWP12T U477 ( .A1(n2855), .A2(n1656), .ZN(n273) );
  OAI211D1BWP12T U478 ( .A1(n2822), .A2(n733), .B(n272), .C(n273), .ZN(
        result[25]) );
  OA22D0BWP12T U479 ( .A1(n2603), .A2(n1030), .B1(n2604), .B2(n1085), .Z(n274)
         );
  NR2D0BWP12T U480 ( .A1(n274), .A2(n275), .ZN(mult_x_18_n425) );
  MAOI22D0BWP12T U481 ( .A1(n274), .A2(n275), .B1(n274), .B2(n275), .ZN(
        mult_x_18_n426) );
  CMPE42D1BWP12T U482 ( .A(mult_x_18_n919), .B(mult_x_18_n946), .C(
        mult_x_18_n975), .CIX(mult_x_18_n684), .D(mult_x_18_n685), .CO(
        mult_x_18_n680), .COX(mult_x_18_n679), .S(mult_x_18_n681) );
  OAI21D0BWP12T U483 ( .A1(n2639), .A2(n1881), .B(n2827), .ZN(n276) );
  IAO21D0BWP12T U484 ( .A1(n471), .A2(n1882), .B(n276), .ZN(n806) );
  CKND0BWP12T U485 ( .I(n2830), .ZN(n277) );
  OAI32D0BWP12T U486 ( .A1(n277), .A2(n2650), .A3(n2231), .B1(n2652), .B2(n277), .ZN(n443) );
  CKND2D0BWP12T U487 ( .A1(a[31]), .A2(a[30]), .ZN(n278) );
  OAI211D0BWP12T U488 ( .A1(a[31]), .A2(a[30]), .B(n2640), .C(n278), .ZN(n2642) );
  CKND2D0BWP12T U489 ( .A1(n1012), .A2(n1011), .ZN(n279) );
  MOAI22D0BWP12T U490 ( .A1(n1013), .A2(n279), .B1(n1013), .B2(n279), .ZN(
        n2381) );
  CKND0BWP12T U491 ( .I(n2831), .ZN(n280) );
  MAOI22D0BWP12T U492 ( .A1(n2163), .A2(n280), .B1(n2164), .B2(n2827), .ZN(
        n2902) );
  IOA21D0BWP12T U493 ( .A1(n876), .A2(n863), .B(n766), .ZN(n2569) );
  CKND2D0BWP12T U494 ( .A1(n2337), .A2(n2338), .ZN(n281) );
  MAOI22D0BWP12T U495 ( .A1(n1794), .A2(n281), .B1(n1794), .B2(n281), .ZN(
        n2701) );
  OR4D0BWP12T U496 ( .A1(n1834), .A2(n2845), .A3(n2487), .A4(n2878), .Z(n282)
         );
  NR4D0BWP12T U497 ( .A1(n1831), .A2(n1836), .A3(n2709), .A4(n282), .ZN(n283)
         );
  NR3D0BWP12T U498 ( .A1(n2927), .A2(n1837), .A3(n2672), .ZN(n284) );
  NR4D0BWP12T U499 ( .A1(n1825), .A2(n2887), .A3(n2505), .A4(n1824), .ZN(n285)
         );
  NR4D0BWP12T U500 ( .A1(n2543), .A2(n1821), .A3(n2586), .A4(n2522), .ZN(n286)
         );
  IND3D0BWP12T U501 ( .A1(n1826), .B1(n285), .B2(n286), .ZN(n287) );
  NR4D0BWP12T U502 ( .A1(n1839), .A2(n1827), .A3(n2731), .A4(n287), .ZN(n288)
         );
  ND4D0BWP12T U503 ( .A1(n426), .A2(n283), .A3(n284), .A4(n288), .ZN(n289) );
  OR4D0BWP12T U504 ( .A1(n1840), .A2(n2941), .A3(n2756), .A4(n289), .Z(n290)
         );
  OR4D0BWP12T U505 ( .A1(n1841), .A2(n2811), .A3(n2790), .A4(n290), .Z(n1842)
         );
  NR2D0BWP12T U506 ( .A1(n2951), .A2(n2511), .ZN(n291) );
  AOI211D0BWP12T U507 ( .A1(n2511), .A2(n2948), .B(n2825), .C(n291), .ZN(n292)
         );
  OAI21D0BWP12T U508 ( .A1(n2944), .A2(n2594), .B(n2949), .ZN(n293) );
  AOI22D0BWP12T U509 ( .A1(n2512), .A2(n2947), .B1(b[11]), .B2(n293), .ZN(n294) );
  AOI22D0BWP12T U510 ( .A1(n2509), .A2(n2905), .B1(n2903), .B2(n2510), .ZN(
        n295) );
  OAI211D0BWP12T U511 ( .A1(n2512), .A2(n292), .B(n294), .C(n295), .ZN(n296)
         );
  CKND0BWP12T U512 ( .I(n2507), .ZN(n297) );
  MOAI22D0BWP12T U513 ( .A1(n2842), .A2(n297), .B1(n2513), .B2(n2514), .ZN(
        n298) );
  AOI211D0BWP12T U514 ( .A1(n2515), .A2(n2858), .B(n296), .C(n298), .ZN(n2519)
         );
  OAI21D0BWP12T U515 ( .A1(n2446), .A2(n2450), .B(n2447), .ZN(n299) );
  CKND2D0BWP12T U516 ( .A1(n2448), .A2(n2449), .ZN(n300) );
  MOAI22D0BWP12T U517 ( .A1(n299), .A2(n300), .B1(n299), .B2(n300), .ZN(n2884)
         );
  CKND2D0BWP12T U518 ( .A1(n1694), .A2(n1693), .ZN(n301) );
  MOAI22D0BWP12T U519 ( .A1(n1695), .A2(n301), .B1(n1695), .B2(n301), .ZN(
        n2542) );
  AOI21D0BWP12T U520 ( .A1(n1621), .A2(n1629), .B(n1623), .ZN(n302) );
  CKND2D0BWP12T U521 ( .A1(n1624), .A2(n1587), .ZN(n303) );
  MAOI22D0BWP12T U522 ( .A1(n302), .A2(n303), .B1(n302), .B2(n303), .ZN(n1634)
         );
  OAI21D0BWP12T U523 ( .A1(n2944), .A2(n2871), .B(n2949), .ZN(n304) );
  AOI22D0BWP12T U524 ( .A1(n2869), .A2(n2947), .B1(n2868), .B2(n304), .ZN(n305) );
  OAI21D0BWP12T U525 ( .A1(n2870), .A2(n2951), .B(n2949), .ZN(n306) );
  AOI32D0BWP12T U526 ( .A1(n2948), .A2(n2871), .A3(n2870), .B1(n306), .B2(
        n2871), .ZN(n307) );
  OAI211D0BWP12T U527 ( .A1(n2873), .A2(n2872), .B(n305), .C(n307), .ZN(n308)
         );
  AOI21D0BWP12T U528 ( .A1(n2874), .A2(n2875), .B(n308), .ZN(n2876) );
  CKND0BWP12T U529 ( .I(n2926), .ZN(n309) );
  CKND2D0BWP12T U530 ( .A1(n2858), .A2(n2935), .ZN(n310) );
  OAI211D0BWP12T U531 ( .A1(n2973), .A2(n309), .B(n2936), .C(n310), .ZN(n311)
         );
  AOI21D1BWP12T U532 ( .A1(n2937), .A2(n2855), .B(n311), .ZN(n312) );
  IOA21D0BWP12T U533 ( .A1(n2977), .A2(n2938), .B(n312), .ZN(result[20]) );
  INR3D0BWP12T U534 ( .A1(n1311), .B1(n2900), .B2(n1822), .ZN(n833) );
  CKND0BWP12T U535 ( .I(n1870), .ZN(n313) );
  MAOI22D0BWP12T U536 ( .A1(a[29]), .A2(n313), .B1(n1871), .B2(n2251), .ZN(
        n1004) );
  CKND0BWP12T U537 ( .I(n2639), .ZN(n314) );
  MAOI22D0BWP12T U538 ( .A1(n1903), .A2(n314), .B1(n471), .B2(n934), .ZN(n1858) );
  CMPE42D1BWP12T U539 ( .A(mult_x_18_n691), .B(mult_x_18_n920), .C(
        mult_x_18_n695), .CIX(mult_x_18_n692), .D(mult_x_18_n689), .CO(
        mult_x_18_n686), .COX(mult_x_18_n685), .S(mult_x_18_n687) );
  OAI22D0BWP12T U540 ( .A1(n2603), .A2(n435), .B1(n2604), .B2(n437), .ZN(n315)
         );
  MOAI22D0BWP12T U541 ( .A1(n2830), .A2(n2231), .B1(n2830), .B2(n2231), .ZN(
        n316) );
  OAI22D0BWP12T U542 ( .A1(n2652), .A2(n316), .B1(n2650), .B2(n436), .ZN(n317)
         );
  MAOI22D0BWP12T U543 ( .A1(n315), .A2(n317), .B1(n315), .B2(n317), .ZN(n444)
         );
  AN2D0BWP12T U544 ( .A1(n315), .A2(n317), .Z(n445) );
  CKND0BWP12T U545 ( .I(n2482), .ZN(n318) );
  OAI21D0BWP12T U546 ( .A1(n2231), .A2(n318), .B(n2604), .ZN(n1707) );
  AOI21D0BWP12T U547 ( .A1(n2868), .A2(n2066), .B(n837), .ZN(n319) );
  AOI21D0BWP12T U548 ( .A1(n2115), .A2(n319), .B(n2058), .ZN(n2071) );
  CKND0BWP12T U549 ( .I(n2770), .ZN(n320) );
  OAI21D0BWP12T U550 ( .A1(n2868), .A2(n320), .B(n2202), .ZN(n321) );
  CKND0BWP12T U551 ( .I(n1998), .ZN(n322) );
  AOI22D0BWP12T U552 ( .A1(n1992), .A2(n2508), .B1(n2031), .B2(n1991), .ZN(
        n323) );
  OA211D0BWP12T U553 ( .A1(n1990), .A2(n322), .B(n2014), .C(n323), .Z(n324) );
  AOI21D0BWP12T U554 ( .A1(n1993), .A2(n321), .B(n324), .ZN(n2708) );
  IAO21D0BWP12T U555 ( .A1(n2830), .A2(n561), .B(n1610), .ZN(n1621) );
  CKND0BWP12T U556 ( .I(n1413), .ZN(n325) );
  OA222D0BWP12T U557 ( .A1(n325), .A2(n2128), .B1(n2126), .B2(n2117), .C1(n471), .C2(n1547), .Z(n2875) );
  OAI21D0BWP12T U558 ( .A1(n2360), .A2(n2361), .B(n2359), .ZN(n326) );
  CKND2D0BWP12T U559 ( .A1(n2363), .A2(n1769), .ZN(n327) );
  MOAI22D0BWP12T U560 ( .A1(n326), .A2(n327), .B1(n326), .B2(n327), .ZN(n2838)
         );
  CKND2D0BWP12T U561 ( .A1(n785), .A2(n784), .ZN(n328) );
  MOAI22D0BWP12T U562 ( .A1(n783), .A2(n328), .B1(n783), .B2(n328), .ZN(n1797)
         );
  MOAI22D0BWP12T U563 ( .A1(n2594), .A2(b[22]), .B1(n2594), .B2(b[22]), .ZN(
        n329) );
  OAI22D0BWP12T U564 ( .A1(n2597), .A2(n2596), .B1(n2595), .B2(n329), .ZN(n330) );
  AOI21D0BWP12T U565 ( .A1(n2604), .A2(n2603), .B(n2602), .ZN(n331) );
  MOAI22D0BWP12T U566 ( .A1(n2725), .A2(n2598), .B1(n2725), .B2(n2598), .ZN(
        n332) );
  OAI22D0BWP12T U567 ( .A1(n2601), .A2(n2600), .B1(n2599), .B2(n332), .ZN(n333) );
  MOAI22D0BWP12T U568 ( .A1(n331), .A2(n333), .B1(n331), .B2(n333), .ZN(n334)
         );
  MOAI22D0BWP12T U569 ( .A1(a[25]), .A2(n2605), .B1(a[25]), .B2(n2605), .ZN(
        n335) );
  OAI22D0BWP12T U570 ( .A1(n2608), .A2(n2607), .B1(n2606), .B2(n335), .ZN(n336) );
  MAOI22D0BWP12T U571 ( .A1(n334), .A2(n336), .B1(n334), .B2(n336), .ZN(n337)
         );
  MAOI22D0BWP12T U572 ( .A1(n330), .A2(n337), .B1(n330), .B2(n337), .ZN(n338)
         );
  MAOI22D0BWP12T U573 ( .A1(mult_x_18_n379), .A2(n338), .B1(mult_x_18_n379), 
        .B2(n338), .ZN(n339) );
  MAOI22D0BWP12T U574 ( .A1(mult_x_18_n374), .A2(mult_x_18_n377), .B1(
        mult_x_18_n374), .B2(mult_x_18_n377), .ZN(n340) );
  MOAI22D0BWP12T U575 ( .A1(n2609), .A2(b[14]), .B1(n2609), .B2(b[14]), .ZN(
        n341) );
  OAI22D0BWP12T U576 ( .A1(n2612), .A2(n2611), .B1(n2610), .B2(n341), .ZN(n342) );
  MOAI22D0BWP12T U577 ( .A1(n2613), .A2(b[24]), .B1(n2613), .B2(b[24]), .ZN(
        n343) );
  OAI22D0BWP12T U578 ( .A1(n2616), .A2(n2615), .B1(n2614), .B2(n343), .ZN(n344) );
  MOAI22D0BWP12T U579 ( .A1(a[27]), .A2(b[6]), .B1(a[27]), .B2(b[6]), .ZN(n345) );
  OAI22D0BWP12T U580 ( .A1(n2619), .A2(n2618), .B1(n2617), .B2(n345), .ZN(n346) );
  MAOI22D0BWP12T U581 ( .A1(n344), .A2(n346), .B1(n344), .B2(n346), .ZN(n347)
         );
  MOAI22D0BWP12T U582 ( .A1(n2620), .A2(b[28]), .B1(n2620), .B2(b[28]), .ZN(
        n348) );
  OAI22D0BWP12T U583 ( .A1(n2623), .A2(n2622), .B1(n2621), .B2(n348), .ZN(n349) );
  MAOI22D0BWP12T U584 ( .A1(n347), .A2(n349), .B1(n347), .B2(n349), .ZN(n350)
         );
  MAOI22D0BWP12T U585 ( .A1(n342), .A2(n350), .B1(n342), .B2(n350), .ZN(n351)
         );
  MAOI22D0BWP12T U586 ( .A1(mult_x_18_n376), .A2(n351), .B1(mult_x_18_n376), 
        .B2(n351), .ZN(n352) );
  MAOI22D0BWP12T U587 ( .A1(n340), .A2(n352), .B1(n340), .B2(n352), .ZN(n353)
         );
  MAOI22D0BWP12T U588 ( .A1(n339), .A2(n353), .B1(n339), .B2(n353), .ZN(n354)
         );
  MAOI22D0BWP12T U589 ( .A1(mult_x_18_n367), .A2(n354), .B1(mult_x_18_n367), 
        .B2(n354), .ZN(n2624) );
  CKND2D0BWP12T U590 ( .A1(n1727), .A2(n1728), .ZN(n355) );
  MAOI22D0BWP12T U591 ( .A1(n1729), .A2(n355), .B1(n1729), .B2(n355), .ZN(n427) );
  CKND2D0BWP12T U592 ( .A1(n1391), .A2(n1394), .ZN(n356) );
  MAOI22D0BWP12T U593 ( .A1(n1392), .A2(n356), .B1(n1392), .B2(n356), .ZN(
        n1649) );
  CKND2D0BWP12T U594 ( .A1(n2435), .A2(n2436), .ZN(n357) );
  MAOI22D0BWP12T U595 ( .A1(n2450), .A2(n357), .B1(n2450), .B2(n357), .ZN(
        n2559) );
  OAI22D0BWP12T U596 ( .A1(n1934), .A2(n1933), .B1(n1932), .B2(n2052), .ZN(
        n358) );
  AOI211D0BWP12T U597 ( .A1(n1929), .A2(n2049), .B(n2868), .C(n358), .ZN(n359)
         );
  OA21D0BWP12T U598 ( .A1(n1931), .A2(n1930), .B(n359), .Z(n2585) );
  NR2D0BWP12T U599 ( .A1(n2871), .A2(n1835), .ZN(n360) );
  MOAI22D0BWP12T U600 ( .A1(n2620), .A2(n360), .B1(n2620), .B2(n360), .ZN(
        n1825) );
  OAI211D0BWP12T U601 ( .A1(n2532), .A2(n2533), .B(n2531), .C(n2530), .ZN(n361) );
  AOI21D0BWP12T U602 ( .A1(n2967), .A2(n2536), .B(n361), .ZN(n362) );
  AOI21D0BWP12T U603 ( .A1(n2746), .A2(n2894), .B(n2893), .ZN(n363) );
  AOI22D0BWP12T U604 ( .A1(n2538), .A2(n2886), .B1(n2855), .B2(n2539), .ZN(
        n364) );
  CKND0BWP12T U605 ( .I(n2957), .ZN(n365) );
  AOI22D0BWP12T U606 ( .A1(n2858), .A2(n2541), .B1(n2537), .B2(n365), .ZN(n366) );
  OAI211D0BWP12T U607 ( .A1(n2540), .A2(n363), .B(n364), .C(n366), .ZN(n367)
         );
  CKND0BWP12T U608 ( .I(n2522), .ZN(n368) );
  MOAI22D0BWP12T U609 ( .A1(n2878), .A2(n368), .B1(n2866), .B2(n2523), .ZN(
        n369) );
  AOI211D0BWP12T U610 ( .A1(n2977), .A2(n2542), .B(n367), .C(n369), .ZN(n370)
         );
  OAI211D0BWP12T U611 ( .A1(n2535), .A2(n2534), .B(n362), .C(n370), .ZN(
        result[7]) );
  IOA21D0BWP12T U612 ( .A1(n1870), .A2(a[31]), .B(n1849), .ZN(n2098) );
  IOA21D0BWP12T U613 ( .A1(n750), .A2(a[31]), .B(n1004), .ZN(n1863) );
  CMPE42D1BWP12T U614 ( .A(mult_x_18_n921), .B(mult_x_18_n948), .C(
        mult_x_18_n700), .CIX(mult_x_18_n697), .D(mult_x_18_n696), .CO(
        mult_x_18_n693), .COX(mult_x_18_n692), .S(mult_x_18_n694) );
  OA22D1BWP12T U615 ( .A1(n471), .A2(n854), .B1(n853), .B2(n2639), .Z(n871) );
  IOA21D0BWP12T U616 ( .A1(n2057), .A2(n2827), .B(n2956), .ZN(n2101) );
  IAO21D0BWP12T U617 ( .A1(n2827), .A2(n1854), .B(n806), .ZN(n1866) );
  IND2D0BWP12T U618 ( .A1(n1822), .B1(n1823), .ZN(n371) );
  MAOI22D0BWP12T U619 ( .A1(n2900), .A2(n371), .B1(n2900), .B2(n371), .ZN(
        n2887) );
  IND2D0BWP12T U620 ( .A1(n548), .B1(n671), .ZN(n2949) );
  IND4D0BWP12T U621 ( .A1(n2514), .B1(n2195), .B2(n2902), .B3(n2194), .ZN(n372) );
  AOI211D0BWP12T U622 ( .A1(n2198), .A2(n372), .B(n2197), .C(n2196), .ZN(n2325) );
  MOAI22D0BWP12T U623 ( .A1(n2626), .A2(b[18]), .B1(n2626), .B2(b[18]), .ZN(
        n373) );
  OAI22D0BWP12T U624 ( .A1(n2629), .A2(n2628), .B1(n2627), .B2(n373), .ZN(n374) );
  MOAI22D0BWP12T U625 ( .A1(n2747), .A2(n2897), .B1(n2747), .B2(n2897), .ZN(
        n375) );
  OAI22D0BWP12T U626 ( .A1(n2632), .A2(n2631), .B1(n2630), .B2(n375), .ZN(n376) );
  MAOI22D0BWP12T U627 ( .A1(n374), .A2(n376), .B1(n374), .B2(n376), .ZN(n377)
         );
  MOAI22D0BWP12T U628 ( .A1(n2633), .A2(b[26]), .B1(n2633), .B2(b[26]), .ZN(
        n378) );
  OAI22D0BWP12T U629 ( .A1(n2635), .A2(n2634), .B1(n1025), .B2(n378), .ZN(n379) );
  MAOI22D0BWP12T U630 ( .A1(n377), .A2(n379), .B1(n377), .B2(n379), .ZN(n380)
         );
  MAOI22D0BWP12T U631 ( .A1(n2625), .A2(n380), .B1(n2625), .B2(n380), .ZN(n381) );
  MAOI22D0BWP12T U632 ( .A1(mult_x_18_n373), .A2(n381), .B1(mult_x_18_n373), 
        .B2(n381), .ZN(n382) );
  MAOI22D0BWP12T U633 ( .A1(mult_x_18_n364), .A2(n382), .B1(mult_x_18_n364), 
        .B2(n382), .ZN(n2654) );
  CKND2D0BWP12T U634 ( .A1(n2349), .A2(n2348), .ZN(n383) );
  MOAI22D0BWP12T U635 ( .A1(n2350), .A2(n383), .B1(n2350), .B2(n383), .ZN(
        n2506) );
  OAI21D0BWP12T U636 ( .A1(n1748), .A2(n1772), .B(n1749), .ZN(n384) );
  CKND2D0BWP12T U637 ( .A1(n1750), .A2(n635), .ZN(n385) );
  MOAI22D0BWP12T U638 ( .A1(n384), .A2(n385), .B1(n384), .B2(n385), .ZN(n1753)
         );
  CKND2D0BWP12T U639 ( .A1(n1608), .A2(n1618), .ZN(n386) );
  MAOI22D0BWP12T U640 ( .A1(n1639), .A2(n386), .B1(n1639), .B2(n386), .ZN(
        n2539) );
  AO222D0BWP12T U641 ( .A1(n2173), .A2(n986), .B1(n2170), .B2(n987), .C1(n1000), .C2(n2166), .Z(n2184) );
  CKND2D0BWP12T U642 ( .A1(n1702), .A2(n1701), .ZN(n387) );
  MOAI22D0BWP12T U643 ( .A1(n1703), .A2(n387), .B1(n1703), .B2(n387), .ZN(
        n2883) );
  OAI21D0BWP12T U644 ( .A1(n2427), .A2(n2428), .B(n2426), .ZN(n388) );
  CKND2D0BWP12T U645 ( .A1(n2430), .A2(n2431), .ZN(n389) );
  MOAI22D0BWP12T U646 ( .A1(n388), .A2(n389), .B1(n388), .B2(n389), .ZN(n2843)
         );
  CKND0BWP12T U647 ( .I(n2855), .ZN(n390) );
  CKND0BWP12T U648 ( .I(n2866), .ZN(n391) );
  OAI22D0BWP12T U649 ( .A1(n2659), .A2(n390), .B1(n2661), .B2(n391), .ZN(n2922) );
  OAI211D0BWP12T U650 ( .A1(n2585), .A2(n2584), .B(n2583), .C(n2582), .ZN(n392) );
  INVD1BWP12T U651 ( .I(n2568), .ZN(n393) );
  OAI22D1BWP12T U652 ( .A1(n2822), .A2(n393), .B1(n2591), .B2(n2957), .ZN(n394) );
  AOI211D1BWP12T U653 ( .A1(n2586), .A2(n2940), .B(n392), .C(n394), .ZN(n395)
         );
  CKND2D0BWP12T U654 ( .A1(n2590), .A2(n2886), .ZN(n396) );
  CKND2D0BWP12T U655 ( .A1(n2866), .A2(n2592), .ZN(n397) );
  ND4D1BWP12T U656 ( .A1(n2589), .A2(n395), .A3(n396), .A4(n397), .ZN(
        result[6]) );
  CMPE42D1BWP12T U657 ( .A(mult_x_18_n652), .B(mult_x_18_n942), .C(
        mult_x_18_n649), .CIX(mult_x_18_n653), .D(mult_x_18_n657), .CO(
        mult_x_18_n645), .COX(mult_x_18_n644), .S(mult_x_18_n646) );
  AOI222D0BWP12T U658 ( .A1(n1999), .A2(n1512), .B1(n2001), .B2(n1513), .C1(
        n2000), .C2(n792), .ZN(n398) );
  IOA21D0BWP12T U659 ( .A1(n2002), .A2(n1511), .B(n398), .ZN(n1966) );
  CKND0BWP12T U660 ( .I(n1640), .ZN(n399) );
  OAI21D0BWP12T U661 ( .A1(n2301), .A2(n2283), .B(n399), .ZN(n685) );
  CMPE42D1BWP12T U662 ( .A(mult_x_18_n1010), .B(mult_x_18_n923), .C(
        mult_x_18_n950), .CIX(mult_x_18_n707), .D(mult_x_18_n979), .CO(
        mult_x_18_n703), .COX(mult_x_18_n702), .S(mult_x_18_n704) );
  INR2D0BWP12T U663 ( .A1(n2385), .B1(n2909), .ZN(n842) );
  AOI21D0BWP12T U664 ( .A1(n1998), .A2(n1970), .B(n2508), .ZN(n400) );
  OAI32D0BWP12T U665 ( .A1(n1902), .A2(n2034), .A3(n1998), .B1(n400), .B2(
        n1902), .ZN(n1982) );
  MAOI22D0BWP12T U666 ( .A1(n2827), .A2(n2201), .B1(n2827), .B2(n2474), .ZN(
        n2195) );
  IAO21D0BWP12T U667 ( .A1(n2871), .A2(n2868), .B(n1576), .ZN(n2370) );
  IOA21D0BWP12T U668 ( .A1(n2831), .A2(n822), .B(n766), .ZN(n2076) );
  OA21D0BWP12T U669 ( .A1(n2231), .A2(n2302), .B(n2355), .Z(n2358) );
  IND2D0BWP12T U670 ( .A1(n2264), .B1(n2944), .ZN(n2948) );
  NR3D0BWP12T U671 ( .A1(n1855), .A2(n2804), .A3(n1981), .ZN(n401) );
  ND4D0BWP12T U672 ( .A1(n1918), .A2(n2063), .A3(n401), .A4(n1961), .ZN(n402)
         );
  NR3D0BWP12T U673 ( .A1(n2706), .A2(n1964), .A3(n402), .ZN(n1888) );
  INR3D0BWP12T U674 ( .A1(n1823), .B1(n2900), .B2(n1822), .ZN(n403) );
  MOAI22D0BWP12T U675 ( .A1(n2594), .A2(n403), .B1(n2594), .B2(n403), .ZN(
        n2505) );
  AOI21D0BWP12T U676 ( .A1(n1618), .A2(n1619), .B(n1617), .ZN(n404) );
  IOA21D0BWP12T U677 ( .A1(n571), .A2(a[8]), .B(n1620), .ZN(n405) );
  MAOI22D0BWP12T U678 ( .A1(n404), .A2(n405), .B1(n404), .B2(n405), .ZN(n2558)
         );
  CKND2D0BWP12T U679 ( .A1(n1771), .A2(n1774), .ZN(n406) );
  MAOI22D0BWP12T U680 ( .A1(n1772), .A2(n406), .B1(n1772), .B2(n406), .ZN(
        n2541) );
  AOI21D0BWP12T U681 ( .A1(n2437), .A2(n2441), .B(n2438), .ZN(n407) );
  CKND2D0BWP12T U682 ( .A1(n2439), .A2(n2419), .ZN(n408) );
  MAOI22D0BWP12T U683 ( .A1(n407), .A2(n408), .B1(n407), .B2(n408), .ZN(n2592)
         );
  IND2D0BWP12T U684 ( .A1(n1704), .B1(n1705), .ZN(n409) );
  MAOI22D0BWP12T U685 ( .A1(n1706), .A2(n409), .B1(n1706), .B2(n409), .ZN(
        n2854) );
  MAOI22D0BWP12T U686 ( .A1(mult_x_18_n365), .A2(mult_x_18_n368), .B1(
        mult_x_18_n365), .B2(mult_x_18_n368), .ZN(n410) );
  MAOI22D0BWP12T U687 ( .A1(n2654), .A2(n2653), .B1(n2654), .B2(n2653), .ZN(
        n411) );
  MAOI22D0BWP12T U688 ( .A1(n410), .A2(n411), .B1(n410), .B2(n411), .ZN(n412)
         );
  MAOI22D0BWP12T U689 ( .A1(n2624), .A2(n412), .B1(n2624), .B2(n412), .ZN(n413) );
  MAOI22D0BWP12T U690 ( .A1(mult_x_18_n361), .A2(n413), .B1(mult_x_18_n361), 
        .B2(n413), .ZN(n414) );
  MAOI22D0BWP12T U691 ( .A1(n414), .A2(mult_x_18_n362), .B1(n414), .B2(
        mult_x_18_n362), .ZN(n415) );
  MAOI22D0BWP12T U692 ( .A1(n2655), .A2(n415), .B1(n2655), .B2(n415), .ZN(
        n2925) );
  NR2D0BWP12T U693 ( .A1(n1978), .A2(n2495), .ZN(n416) );
  AOI22D0BWP12T U694 ( .A1(n1906), .A2(n416), .B1(n2858), .B2(n1767), .ZN(n417) );
  MOAI22D0BWP12T U695 ( .A1(n1977), .A2(n1578), .B1(n2365), .B2(n2967), .ZN(
        n418) );
  OAI211D0BWP12T U696 ( .A1(n2257), .A2(n1583), .B(n1582), .C(n1581), .ZN(n419) );
  AOI211D0BWP12T U697 ( .A1(n2874), .A2(n2184), .B(n418), .C(n419), .ZN(n420)
         );
  AOI22D0BWP12T U698 ( .A1(n2866), .A2(n2432), .B1(n2855), .B2(n1634), .ZN(
        n421) );
  AOI22D0BWP12T U699 ( .A1(n2940), .A2(n1825), .B1(n2977), .B2(n1712), .ZN(
        n422) );
  AN4D0BWP12T U700 ( .A1(n417), .A2(n420), .A3(n421), .A4(n422), .Z(n423) );
  OAI21D0BWP12T U701 ( .A1(n2103), .A2(n2957), .B(n423), .ZN(result[5]) );
  FA1D2BWP12T U702 ( .A(a[25]), .B(b[25]), .CI(n700), .CO(n1743), .S(n1801) );
  FA1D2BWP12T U703 ( .A(a[22]), .B(b[22]), .CI(n738), .CO(n1744), .S(n1799) );
  TPOAI22D1BWP12T U704 ( .A1(n2616), .A2(n1153), .B1(n2614), .B2(n1122), .ZN(
        mult_x_18_n892) );
  TPOAI22D1BWP12T U705 ( .A1(n2616), .A2(n1050), .B1(n2614), .B2(n1099), .ZN(
        n1052) );
  TPNR2D1BWP12T U706 ( .A1(b[11]), .A2(n2897), .ZN(n501) );
  INVD1BWP12T U707 ( .I(b[11]), .ZN(n2511) );
  INVD2BWP12T U708 ( .I(b[5]), .ZN(n2284) );
  INVD4BWP12T U709 ( .I(a[25]), .ZN(n2253) );
  OR2XD1BWP12T U710 ( .A1(n521), .A2(n2283), .Z(n424) );
  INVD3BWP12T U711 ( .I(n2233), .ZN(n2725) );
  XNR2XD4BWP12T U712 ( .A1(n2620), .A2(n2574), .ZN(n1025) );
  INVD1BWP12T U713 ( .I(a[4]), .ZN(n2869) );
  OR2XD1BWP12T U714 ( .A1(mult_x_18_n539), .A2(mult_x_18_n523), .Z(n425) );
  OR2XD1BWP12T U715 ( .A1(n570), .A2(n569), .Z(n1618) );
  XNR2D1BWP12T U716 ( .A1(n1835), .A2(n2871), .ZN(n426) );
  NR2D1BWP12T U717 ( .A1(n516), .A2(n563), .ZN(n1589) );
  BUFFD2BWP12T U718 ( .I(a[2]), .Z(n2303) );
  INVD2BWP12T U719 ( .I(a[1]), .ZN(n2481) );
  INVD8BWP12T U720 ( .I(n2481), .ZN(n2482) );
  XNR2XD4BWP12T U721 ( .A1(n2303), .A2(n2482), .ZN(n2650) );
  INVD3BWP12T U722 ( .I(a[3]), .ZN(n2835) );
  INVD9BWP12T U723 ( .I(n2835), .ZN(n2830) );
  XOR2D1BWP12T U724 ( .A1(n2303), .A2(n2830), .Z(n428) );
  ND2D8BWP12T U725 ( .A1(n2650), .A2(n428), .ZN(n2652) );
  INVD1P75BWP12T U726 ( .I(b[2]), .ZN(n471) );
  INVD8BWP12T U727 ( .I(n471), .ZN(n2639) );
  XNR2D1BWP12T U728 ( .A1(n2830), .A2(n2639), .ZN(n434) );
  INVD4BWP12T U729 ( .I(n539), .ZN(n2831) );
  XNR2D1BWP12T U730 ( .A1(n2830), .A2(n2831), .ZN(n1147) );
  OAI22D1BWP12T U731 ( .A1(n2652), .A2(n434), .B1(n2650), .B2(n1147), .ZN(n450) );
  CKND3BWP12T U732 ( .I(a[5]), .ZN(n2257) );
  INVD8BWP12T U733 ( .I(n2257), .ZN(n2620) );
  INVD2BWP12T U734 ( .I(n2869), .ZN(n2871) );
  XOR2D1BWP12T U735 ( .A1(n2620), .A2(n2871), .Z(n429) );
  XNR2XD4BWP12T U736 ( .A1(n2871), .A2(n2830), .ZN(n2621) );
  ND2XD8BWP12T U737 ( .A1(n429), .A2(n2621), .ZN(n2623) );
  CKND2BWP12T U738 ( .I(b[0]), .ZN(n2285) );
  INVD9BWP12T U739 ( .I(n2285), .ZN(n2231) );
  XNR2D1BWP12T U740 ( .A1(n2620), .A2(n2231), .ZN(n430) );
  INVD1BWP12T U741 ( .I(b[1]), .ZN(n2483) );
  INVD4BWP12T U742 ( .I(n2483), .ZN(n2477) );
  XNR2D1BWP12T U743 ( .A1(n2620), .A2(n2477), .ZN(n1112) );
  OAI22D1BWP12T U744 ( .A1(n2623), .A2(n430), .B1(n1112), .B2(n2621), .ZN(n449) );
  BUFFD2BWP12T U745 ( .I(a[0]), .Z(n2302) );
  INVD4BWP12T U746 ( .I(n2302), .ZN(n2603) );
  TPND2D3BWP12T U747 ( .A1(n2482), .A2(n2603), .ZN(n2604) );
  INVD6BWP12T U748 ( .I(n466), .ZN(n2868) );
  XNR2D1BWP12T U749 ( .A1(n2482), .A2(n2868), .ZN(n433) );
  XNR2D1BWP12T U750 ( .A1(n2482), .A2(b[5]), .ZN(n1125) );
  OAI22D1BWP12T U751 ( .A1(n2604), .A2(n433), .B1(n1125), .B2(n2603), .ZN(
        n1315) );
  CKND0BWP12T U752 ( .I(n2620), .ZN(n432) );
  IND2D1BWP12T U753 ( .A1(n2231), .B1(n2620), .ZN(n431) );
  OAI22D1BWP12T U754 ( .A1(n2623), .A2(n432), .B1(n2621), .B2(n431), .ZN(n1314) );
  NR2D1BWP12T U755 ( .A1(mult_x_18_n704), .A2(n456), .ZN(n1696) );
  XNR2D1BWP12T U756 ( .A1(n2482), .A2(n2831), .ZN(n435) );
  OAI22D1BWP12T U757 ( .A1(n2604), .A2(n435), .B1(n433), .B2(n2603), .ZN(n453)
         );
  INR2D1BWP12T U758 ( .A1(n2231), .B1(n2621), .ZN(n452) );
  XNR2D1BWP12T U759 ( .A1(n2830), .A2(n2477), .ZN(n436) );
  OAI22D1BWP12T U760 ( .A1(n2652), .A2(n436), .B1(n2650), .B2(n434), .ZN(n451)
         );
  XNR2D1BWP12T U761 ( .A1(n2482), .A2(n2639), .ZN(n437) );
  OR2XD1BWP12T U762 ( .A1(n446), .A2(n445), .Z(n1702) );
  NR2D1BWP12T U763 ( .A1(n444), .A2(n443), .ZN(n1704) );
  XNR2D1BWP12T U764 ( .A1(n2482), .A2(n2477), .ZN(n438) );
  OAI22D1BWP12T U765 ( .A1(n2604), .A2(n438), .B1(n437), .B2(n2603), .ZN(n441)
         );
  INR2D1BWP12T U766 ( .A1(n2231), .B1(n2650), .ZN(n440) );
  OR2XD1BWP12T U767 ( .A1(n441), .A2(n440), .Z(n869) );
  OAI22D1BWP12T U768 ( .A1(n2604), .A2(n2231), .B1(n438), .B2(n2603), .ZN(
        n1708) );
  INVD1BWP12T U769 ( .I(n1708), .ZN(n439) );
  INR2D1BWP12T U770 ( .A1(n1707), .B1(n439), .ZN(n1709) );
  ND2D1BWP12T U771 ( .A1(n441), .A2(n440), .ZN(n868) );
  INVD1BWP12T U772 ( .I(n868), .ZN(n442) );
  AOI21D1BWP12T U773 ( .A1(n869), .A2(n1709), .B(n442), .ZN(n1706) );
  ND2D1BWP12T U774 ( .A1(n444), .A2(n443), .ZN(n1705) );
  OAI21D1BWP12T U775 ( .A1(n1704), .A2(n1706), .B(n1705), .ZN(n1703) );
  ND2D1BWP12T U776 ( .A1(n446), .A2(n445), .ZN(n1701) );
  INVD1BWP12T U777 ( .I(n1701), .ZN(n447) );
  AOI21D1BWP12T U778 ( .A1(n1702), .A2(n1703), .B(n447), .ZN(n1566) );
  FA1D0BWP12T U779 ( .A(n450), .B(n449), .CI(n448), .CO(n456), .S(n455) );
  FA1D0BWP12T U780 ( .A(n453), .B(n452), .CI(n451), .CO(n454), .S(n446) );
  NR2D1BWP12T U781 ( .A1(n455), .A2(n454), .ZN(n1563) );
  ND2D1BWP12T U782 ( .A1(n455), .A2(n454), .ZN(n1564) );
  OA21D1BWP12T U783 ( .A1(n1566), .A2(n1563), .B(n1564), .Z(n1699) );
  ND2D1BWP12T U784 ( .A1(mult_x_18_n704), .A2(n456), .ZN(n1697) );
  OAI21D1BWP12T U785 ( .A1(n1696), .A2(n1699), .B(n1697), .ZN(n1695) );
  OR2D1BWP12T U786 ( .A1(mult_x_18_n699), .A2(mult_x_18_n703), .Z(n1694) );
  ND2D1BWP12T U787 ( .A1(mult_x_18_n699), .A2(mult_x_18_n703), .ZN(n1693) );
  INVD1BWP12T U788 ( .I(n1693), .ZN(n457) );
  AOI21D1BWP12T U789 ( .A1(n1695), .A2(n1694), .B(n457), .ZN(n591) );
  INVD1BWP12T U790 ( .I(n591), .ZN(n1692) );
  OR2XD1BWP12T U791 ( .A1(mult_x_18_n698), .A2(mult_x_18_n694), .Z(n1691) );
  ND2D1BWP12T U792 ( .A1(mult_x_18_n698), .A2(mult_x_18_n694), .ZN(n1690) );
  INVD1BWP12T U793 ( .I(n1690), .ZN(n588) );
  AOI21D1BWP12T U794 ( .A1(n1692), .A2(n1691), .B(n588), .ZN(n459) );
  ND2D1BWP12T U795 ( .A1(mult_x_18_n687), .A2(mult_x_18_n693), .ZN(n586) );
  ND2D1BWP12T U796 ( .A1(n589), .A2(n586), .ZN(n458) );
  XOR2XD1BWP12T U797 ( .A1(n459), .A2(n458), .Z(n1713) );
  INVD1BWP12T U798 ( .I(op[2]), .ZN(n670) );
  ND2D1BWP12T U799 ( .A1(op[3]), .A2(op[0]), .ZN(n535) );
  NR3D1BWP12T U800 ( .A1(op[1]), .A2(n670), .A3(n535), .ZN(n2977) );
  CKND2D1BWP12T U801 ( .A1(n1713), .A2(n2977), .ZN(n577) );
  OR2XD4BWP12T U802 ( .A1(n2231), .A2(n2477), .Z(n1870) );
  INVD2BWP12T U803 ( .I(a[21]), .ZN(n2233) );
  CKND2D4BWP12T U804 ( .A1(n2477), .A2(n2231), .ZN(n1869) );
  CKND1BWP12T U805 ( .I(a[24]), .ZN(n2946) );
  OAI22D0BWP12T U806 ( .A1(n1870), .A2(n2233), .B1(n1869), .B2(n2946), .ZN(
        n461) );
  INVD2BWP12T U807 ( .I(a[23]), .ZN(n2751) );
  IND2D1BWP12T U808 ( .A1(n2231), .B1(n2477), .ZN(n826) );
  INVD2P3BWP12T U809 ( .I(n826), .ZN(n750) );
  IND2D1BWP12T U810 ( .A1(n2477), .B1(n2231), .ZN(n825) );
  INVD1BWP12T U811 ( .I(n825), .ZN(n751) );
  INVD2BWP12T U812 ( .I(n751), .ZN(n1871) );
  CKND1BWP12T U813 ( .I(a[22]), .ZN(n2232) );
  OAI22D1BWP12T U814 ( .A1(n2751), .A2(n1872), .B1(n1871), .B2(n2232), .ZN(
        n460) );
  NR2D1BWP12T U815 ( .A1(n461), .A2(n460), .ZN(n1861) );
  ND2D1BWP12T U816 ( .A1(n2639), .A2(n2831), .ZN(n1930) );
  INVD2BWP12T U817 ( .I(a[13]), .ZN(n2241) );
  CKND1BWP12T U818 ( .I(a[16]), .ZN(n2235) );
  OAI22D0BWP12T U819 ( .A1(n1870), .A2(n2241), .B1(n1869), .B2(n2235), .ZN(
        n463) );
  INVD2BWP12T U820 ( .I(a[15]), .ZN(n2240) );
  OAI22D1BWP12T U821 ( .A1(n1872), .A2(n2240), .B1(n1871), .B2(n1441), .ZN(
        n462) );
  NR2D1BWP12T U822 ( .A1(n463), .A2(n462), .ZN(n1890) );
  OAI22D1BWP12T U823 ( .A1(n1870), .A2(n2683), .B1(n1871), .B2(n2705), .ZN(
        n465) );
  INVD2BWP12T U824 ( .I(a[19]), .ZN(n2234) );
  CKND1BWP12T U825 ( .I(a[20]), .ZN(n2929) );
  TPOAI22D0BWP12T U826 ( .A1(n1872), .A2(n2234), .B1(n1869), .B2(n2929), .ZN(
        n464) );
  NR2D1BWP12T U827 ( .A1(n465), .A2(n464), .ZN(n1862) );
  IND2D1BWP12T U828 ( .A1(n2639), .B1(n2831), .ZN(n1933) );
  INVD2BWP12T U829 ( .I(a[9]), .ZN(n2243) );
  BUFFD2BWP12T U830 ( .I(a[12]), .Z(n2308) );
  INVD1BWP12T U831 ( .I(n2308), .ZN(n2242) );
  OAI22D1BWP12T U832 ( .A1(n1870), .A2(n2243), .B1(n1869), .B2(n2242), .ZN(
        n468) );
  INVD2BWP12T U833 ( .I(a[11]), .ZN(n2512) );
  INVD1BWP12T U834 ( .I(a[10]), .ZN(n2898) );
  TPOAI22D0BWP12T U835 ( .A1(n1872), .A2(n2512), .B1(n1871), .B2(n2898), .ZN(
        n467) );
  NR2D1BWP12T U836 ( .A1(n468), .A2(n467), .ZN(n1889) );
  INVD1BWP12T U837 ( .I(a[29]), .ZN(n2248) );
  INVD1BWP12T U838 ( .I(a[30]), .ZN(n2251) );
  INVD1BWP12T U839 ( .I(a[31]), .ZN(n2310) );
  INVD1BWP12T U840 ( .I(n1863), .ZN(n1851) );
  CKND1BWP12T U841 ( .I(a[26]), .ZN(n2779) );
  TPOAI22D0BWP12T U842 ( .A1(n1870), .A2(n2253), .B1(n1871), .B2(n2779), .ZN(
        n470) );
  INVD1BWP12T U843 ( .I(a[27]), .ZN(n2252) );
  CKND1BWP12T U844 ( .I(a[28]), .ZN(n2249) );
  OAI22D0BWP12T U845 ( .A1(n1872), .A2(n2252), .B1(n1869), .B2(n2249), .ZN(
        n469) );
  NR2D1BWP12T U846 ( .A1(n470), .A2(n469), .ZN(n1570) );
  OAI22D1BWP12T U847 ( .A1(n1851), .A2(n1926), .B1(n1570), .B2(n2052), .ZN(
        n1855) );
  NR2D0BWP12T U848 ( .A1(n1855), .A2(n2870), .ZN(n477) );
  ND2D1BWP12T U849 ( .A1(n1870), .A2(n2639), .ZN(n803) );
  INVD1BWP12T U850 ( .I(n803), .ZN(n472) );
  ND2D1BWP12T U851 ( .A1(n1400), .A2(n1398), .ZN(n1959) );
  INVD1BWP12T U852 ( .I(n1959), .ZN(n1999) );
  CKMUX2D1BWP12T U853 ( .I0(n2620), .I1(n2871), .S(n2231), .Z(n986) );
  INVD1BWP12T U854 ( .I(n986), .ZN(n1001) );
  NR2D1BWP12T U855 ( .A1(n1398), .A2(n472), .ZN(n2000) );
  MUX2D1BWP12T U856 ( .I0(n2830), .I1(n2303), .S(n2231), .Z(n987) );
  INVD1BWP12T U857 ( .I(n987), .ZN(n1003) );
  AOI22D0BWP12T U858 ( .A1(n1999), .A2(n1001), .B1(n2000), .B2(n1003), .ZN(
        n475) );
  INVD1BWP12T U859 ( .I(n1398), .ZN(n473) );
  OR2D2BWP12T U860 ( .A1(n1400), .A2(n473), .Z(n1940) );
  INVD2BWP12T U861 ( .I(n1940), .ZN(n2002) );
  INVD4BWP12T U862 ( .I(n2243), .ZN(n2301) );
  MUX2NXD0BWP12T U863 ( .I0(n2301), .I1(a[8]), .S(n2231), .ZN(n999) );
  NR2D1BWP12T U864 ( .A1(n1400), .A2(n1398), .ZN(n1945) );
  CKND3BWP12T U865 ( .I(a[7]), .ZN(n2532) );
  INVD4BWP12T U866 ( .I(n2532), .ZN(n2527) );
  BUFFD2BWP12T U867 ( .I(a[6]), .Z(n2574) );
  CKMUX2D1BWP12T U868 ( .I0(n2527), .I1(n2574), .S(n2231), .Z(n994) );
  INVD1BWP12T U869 ( .I(n994), .ZN(n789) );
  AOI22D0BWP12T U870 ( .A1(n2002), .A2(n999), .B1(n1945), .B2(n789), .ZN(n474)
         );
  ND2D1BWP12T U871 ( .A1(n475), .A2(n474), .ZN(n2024) );
  TPNR2D0BWP12T U872 ( .A1(n2285), .A2(n2302), .ZN(n2258) );
  ND2D1BWP12T U873 ( .A1(n2002), .A2(n1000), .ZN(n2021) );
  INVD1BWP12T U874 ( .I(n1891), .ZN(n648) );
  XNR2D2BWP12T U875 ( .A1(n648), .A2(n2831), .ZN(n2017) );
  INVD1BWP12T U876 ( .I(n2017), .ZN(n1998) );
  MUX2NXD0BWP12T U877 ( .I0(n2024), .I1(n2021), .S(n1998), .ZN(n714) );
  ND2D1BWP12T U878 ( .A1(n648), .A2(n2868), .ZN(n476) );
  ND2D1BWP12T U879 ( .A1(n2831), .A2(n2868), .ZN(n2080) );
  MOAI22D0BWP12T U880 ( .A1(n537), .A2(n477), .B1(n714), .B2(n1997), .ZN(n1972) );
  CKND1BWP12T U881 ( .I(op[3]), .ZN(n544) );
  ND2D1BWP12T U882 ( .A1(op[2]), .A2(n544), .ZN(n573) );
  CKND0BWP12T U883 ( .I(n573), .ZN(n478) );
  INVD1BWP12T U884 ( .I(op[0]), .ZN(n547) );
  INVD1BWP12T U885 ( .I(op[1]), .ZN(n534) );
  NR2D1BWP12T U886 ( .A1(n547), .A2(n534), .ZN(n536) );
  ND2D1BWP12T U887 ( .A1(n478), .A2(n536), .ZN(n2964) );
  INVD1BWP12T U888 ( .I(n2964), .ZN(n2894) );
  NR3D1BWP12T U889 ( .A1(op[1]), .A2(n547), .A3(n573), .ZN(n2858) );
  INVD1BWP12T U890 ( .I(n2858), .ZN(n2814) );
  NR2D1BWP12T U891 ( .A1(n2482), .A2(n2477), .ZN(n1754) );
  NR2XD0BWP12T U892 ( .A1(n2639), .A2(n2303), .ZN(n887) );
  NR2D1BWP12T U893 ( .A1(n1754), .A2(n887), .ZN(n480) );
  NR2XD0BWP12T U894 ( .A1(n2302), .A2(c_in), .ZN(n1559) );
  CKND2D1BWP12T U895 ( .A1(n2302), .A2(c_in), .ZN(n1560) );
  OAI21D1BWP12T U896 ( .A1(n1558), .A2(n1559), .B(n1560), .ZN(n886) );
  CKND2D1BWP12T U897 ( .A1(n2482), .A2(n2477), .ZN(n1755) );
  CKND2D1BWP12T U898 ( .A1(n2639), .A2(n2303), .ZN(n888) );
  OAI21D1BWP12T U899 ( .A1(n1755), .A2(n887), .B(n888), .ZN(n479) );
  AOI21D1BWP12T U900 ( .A1(n480), .A2(n886), .B(n479), .ZN(n1584) );
  CKBD1BWP12T U901 ( .I(n2830), .Z(n481) );
  NR2D1BWP12T U902 ( .A1(n481), .A2(n2831), .ZN(n1760) );
  NR2D1BWP12T U903 ( .A1(n2868), .A2(n2871), .ZN(n1762) );
  NR2D1BWP12T U904 ( .A1(n1760), .A2(n1762), .ZN(n1778) );
  CKBD1BWP12T U905 ( .I(n2620), .Z(n482) );
  NR2D1BWP12T U906 ( .A1(n482), .A2(b[5]), .ZN(n1782) );
  INVD1BWP12T U907 ( .I(b[6]), .ZN(n2572) );
  NR2D1BWP12T U908 ( .A1(b[6]), .A2(n2574), .ZN(n2373) );
  NR2D1BWP12T U909 ( .A1(n1782), .A2(n2373), .ZN(n484) );
  ND2D1BWP12T U910 ( .A1(n1778), .A2(n484), .ZN(n486) );
  CKND2D1BWP12T U911 ( .A1(n481), .A2(n2831), .ZN(n1768) );
  CKND2D1BWP12T U912 ( .A1(n2868), .A2(n2871), .ZN(n1763) );
  OAI21D1BWP12T U913 ( .A1(n1768), .A2(n1762), .B(n1763), .ZN(n1780) );
  ND2D1BWP12T U914 ( .A1(n482), .A2(b[5]), .ZN(n1781) );
  ND2D1BWP12T U915 ( .A1(b[6]), .A2(n2574), .ZN(n2372) );
  OAI21D1BWP12T U916 ( .A1(n1781), .A2(n2373), .B(n2372), .ZN(n483) );
  TPAOI21D1BWP12T U917 ( .A1(n484), .A2(n1780), .B(n483), .ZN(n485) );
  TPOAI21D1BWP12T U918 ( .A1(n1584), .A2(n486), .B(n485), .ZN(n1775) );
  CKND3BWP12T U919 ( .I(n1775), .ZN(n1772) );
  INVD1BWP12T U920 ( .I(b[7]), .ZN(n2525) );
  INVD2BWP12T U921 ( .I(n2525), .ZN(n2528) );
  OR2XD1BWP12T U922 ( .A1(n528), .A2(n2528), .Z(n1774) );
  INVD1BWP12T U923 ( .I(b[8]), .ZN(n2545) );
  INVD2BWP12T U924 ( .I(n2545), .ZN(n2605) );
  OR2XD1BWP12T U925 ( .A1(n2605), .A2(a[8]), .Z(n2368) );
  ND2D1BWP12T U926 ( .A1(n1774), .A2(n2368), .ZN(n1748) );
  CKND2D1BWP12T U927 ( .A1(n528), .A2(n2528), .ZN(n1771) );
  INVD1BWP12T U928 ( .I(n1771), .ZN(n1773) );
  CKND2D1BWP12T U929 ( .A1(n2605), .A2(a[8]), .ZN(n2367) );
  INVD1BWP12T U930 ( .I(n2367), .ZN(n634) );
  AOI21D1BWP12T U931 ( .A1(n1773), .A2(n2368), .B(n634), .ZN(n1749) );
  CKBD1BWP12T U932 ( .I(n2301), .Z(n487) );
  NR2D1BWP12T U933 ( .A1(n487), .A2(b[9]), .ZN(n627) );
  ND2D1BWP12T U934 ( .A1(n487), .A2(b[9]), .ZN(n1750) );
  AOI22D1BWP12T U935 ( .A1(n1972), .A2(n2894), .B1(n2858), .B2(n1753), .ZN(
        n576) );
  CKND0BWP12T U936 ( .I(n535), .ZN(n543) );
  NR2D1BWP12T U937 ( .A1(op[2]), .A2(op[1]), .ZN(n545) );
  ND2D1BWP12T U938 ( .A1(n543), .A2(n545), .ZN(n2878) );
  INVD8BWP12T U939 ( .I(n2527), .ZN(n1119) );
  INVD1BWP12T U940 ( .I(n2574), .ZN(n2578) );
  ND2D1BWP12T U941 ( .A1(n1119), .A2(n2578), .ZN(n488) );
  NR2D1BWP12T U942 ( .A1(n1820), .A2(n488), .ZN(n489) );
  INVD1BWP12T U943 ( .I(n2303), .ZN(n1832) );
  ND2D1BWP12T U944 ( .A1(n489), .A2(n1573), .ZN(n834) );
  INVD1BWP12T U945 ( .I(n834), .ZN(n1823) );
  INVD1BWP12T U946 ( .I(a[8]), .ZN(n2550) );
  CKND2D0BWP12T U947 ( .A1(n1823), .A2(n2550), .ZN(n490) );
  CKXOR2D0BWP12T U948 ( .A1(n490), .A2(n2301), .Z(n1824) );
  CKND0BWP12T U949 ( .I(n1004), .ZN(n492) );
  ND2D1BWP12T U950 ( .A1(n2639), .A2(n2477), .ZN(n2116) );
  NR2D0BWP12T U951 ( .A1(n2116), .A2(n2310), .ZN(n491) );
  AOI21D0BWP12T U952 ( .A1(n492), .A2(n2639), .B(n491), .ZN(n493) );
  OAI21D1BWP12T U953 ( .A1(n2639), .A2(n1570), .B(n493), .ZN(n2057) );
  TPNR2D0BWP12T U954 ( .A1(b[31]), .A2(b[30]), .ZN(n496) );
  TPNR2D0BWP12T U955 ( .A1(b[29]), .A2(b[28]), .ZN(n495) );
  TPNR2D0BWP12T U956 ( .A1(b[27]), .A2(b[26]), .ZN(n494) );
  ND4D1BWP12T U957 ( .A1(n496), .A2(n495), .A3(n494), .A4(n2284), .ZN(n510) );
  TPNR2D0BWP12T U958 ( .A1(b[25]), .A2(b[24]), .ZN(n500) );
  TPNR2D0BWP12T U959 ( .A1(b[23]), .A2(b[22]), .ZN(n499) );
  TPNR2D0BWP12T U960 ( .A1(b[21]), .A2(b[20]), .ZN(n498) );
  NR2XD0BWP12T U961 ( .A1(b[19]), .A2(b[18]), .ZN(n497) );
  ND4D1BWP12T U962 ( .A1(n500), .A2(n499), .A3(n498), .A4(n497), .ZN(n509) );
  TPNR2D0BWP12T U963 ( .A1(b[17]), .A2(b[16]), .ZN(n504) );
  TPNR2D0BWP12T U964 ( .A1(b[15]), .A2(b[14]), .ZN(n503) );
  BUFFD2BWP12T U965 ( .I(b[12]), .Z(n2598) );
  NR2D1BWP12T U966 ( .A1(b[13]), .A2(n2598), .ZN(n502) );
  BUFFD2BWP12T U967 ( .I(b[10]), .Z(n2897) );
  ND4D1BWP12T U968 ( .A1(n504), .A2(n503), .A3(n502), .A4(n501), .ZN(n508) );
  NR2D1BWP12T U969 ( .A1(b[9]), .A2(n2605), .ZN(n506) );
  CKND2D1BWP12T U970 ( .A1(n506), .A2(n505), .ZN(n507) );
  NR4D2BWP12T U971 ( .A1(n510), .A2(n509), .A3(n508), .A4(n507), .ZN(n2115) );
  CKND0BWP12T U972 ( .I(n2080), .ZN(n2154) );
  NR2D1BWP12T U973 ( .A1(n2174), .A2(n2154), .ZN(n2187) );
  OAI21D0BWP12T U974 ( .A1(n2870), .A2(n2057), .B(n2187), .ZN(n511) );
  ND2D1BWP12T U975 ( .A1(n2831), .A2(a[31]), .ZN(n2099) );
  AOI21D0BWP12T U976 ( .A1(n511), .A2(n2099), .B(n537), .ZN(n512) );
  NR2D0BWP12T U977 ( .A1(n512), .A2(n2058), .ZN(n2072) );
  NR2D1BWP12T U978 ( .A1(op[0]), .A2(op[1]), .ZN(n671) );
  INVD1BWP12T U979 ( .I(n671), .ZN(n513) );
  NR2D1BWP12T U980 ( .A1(n573), .A2(n513), .ZN(n2905) );
  INVD1BWP12T U981 ( .I(n2905), .ZN(n2957) );
  NR2D1BWP12T U982 ( .A1(n1558), .A2(n2302), .ZN(n2422) );
  NR2D1BWP12T U983 ( .A1(n2482), .A2(n557), .ZN(n2420) );
  CKND2D1BWP12T U984 ( .A1(n2482), .A2(n557), .ZN(n2421) );
  OAI21D1BWP12T U985 ( .A1(n2422), .A2(n2420), .B(n2421), .ZN(n904) );
  INVD1P75BWP12T U986 ( .I(n2831), .ZN(n561) );
  NR2D1BWP12T U987 ( .A1(n2830), .A2(n561), .ZN(n2429) );
  INVD1P75BWP12T U988 ( .I(n2639), .ZN(n558) );
  NR2D1BWP12T U989 ( .A1(n558), .A2(n2303), .ZN(n2427) );
  NR2D1BWP12T U990 ( .A1(n2429), .A2(n2427), .ZN(n515) );
  CKND2D1BWP12T U991 ( .A1(n558), .A2(n2303), .ZN(n2426) );
  ND2D1BWP12T U992 ( .A1(n2830), .A2(n561), .ZN(n2430) );
  OAI21D1BWP12T U993 ( .A1(n2429), .A2(n2426), .B(n2430), .ZN(n514) );
  AOI21D1BWP12T U994 ( .A1(n904), .A2(n515), .B(n514), .ZN(n1588) );
  CKBD1BWP12T U995 ( .I(n2620), .Z(n516) );
  INVD2P3BWP12T U996 ( .I(b[5]), .ZN(n563) );
  INVD1P75BWP12T U997 ( .I(n2868), .ZN(n562) );
  NR2D1BWP12T U998 ( .A1(n570), .A2(n569), .ZN(n2442) );
  NR2D1BWP12T U999 ( .A1(n564), .A2(n2574), .ZN(n2440) );
  NR2D1BWP12T U1000 ( .A1(n2442), .A2(n2440), .ZN(n518) );
  CKND2D1BWP12T U1001 ( .A1(n2437), .A2(n518), .ZN(n520) );
  ND2D1BWP12T U1002 ( .A1(n562), .A2(n2871), .ZN(n2433) );
  ND2D1BWP12T U1003 ( .A1(n516), .A2(n563), .ZN(n1590) );
  OAI21D1BWP12T U1004 ( .A1(n1589), .A2(n2433), .B(n1590), .ZN(n2438) );
  ND2D1BWP12T U1005 ( .A1(n564), .A2(n2574), .ZN(n2439) );
  ND2D1BWP12T U1006 ( .A1(n570), .A2(n569), .ZN(n2443) );
  OAI21D1BWP12T U1007 ( .A1(n2442), .A2(n2439), .B(n2443), .ZN(n517) );
  AOI21D1BWP12T U1008 ( .A1(n2438), .A2(n518), .B(n517), .ZN(n519) );
  OAI21D1BWP12T U1009 ( .A1(n1588), .A2(n520), .B(n519), .ZN(n616) );
  OR2XD1BWP12T U1010 ( .A1(n571), .A2(a[8]), .Z(n2436) );
  CKND2D1BWP12T U1011 ( .A1(n571), .A2(a[8]), .ZN(n2435) );
  INVD1BWP12T U1012 ( .I(n2435), .ZN(n618) );
  TPAOI21D0BWP12T U1013 ( .A1(n616), .A2(n2436), .B(n618), .ZN(n523) );
  CKBD1BWP12T U1014 ( .I(n2301), .Z(n521) );
  CKND2D1BWP12T U1015 ( .A1(n521), .A2(n2283), .ZN(n617) );
  CKND2D1BWP12T U1016 ( .A1(n424), .A2(n617), .ZN(n522) );
  XOR2XD1BWP12T U1017 ( .A1(n523), .A2(n522), .Z(n2444) );
  ND3D1BWP12T U1018 ( .A1(op[1]), .A2(n547), .A3(n670), .ZN(n542) );
  NR2D1BWP12T U1019 ( .A1(n544), .A2(n542), .ZN(n2866) );
  MOAI22D0BWP12T U1020 ( .A1(n2072), .A2(n2957), .B1(n2444), .B2(n2866), .ZN(
        n556) );
  CKND2D1BWP12T U1021 ( .A1(n2231), .A2(n2302), .ZN(n2355) );
  NR2D1BWP12T U1022 ( .A1(n2482), .A2(n2477), .ZN(n2352) );
  CKND2D1BWP12T U1023 ( .A1(n2482), .A2(n2477), .ZN(n2353) );
  OAI21D1BWP12T U1024 ( .A1(n2355), .A2(n2352), .B(n2353), .ZN(n892) );
  CKBD1BWP12T U1025 ( .I(n2830), .Z(n524) );
  NR2D1BWP12T U1026 ( .A1(n524), .A2(n2831), .ZN(n2362) );
  NR2XD0BWP12T U1027 ( .A1(n2639), .A2(n2303), .ZN(n2360) );
  NR2D1BWP12T U1028 ( .A1(n2362), .A2(n2360), .ZN(n526) );
  CKND2D1BWP12T U1029 ( .A1(n2639), .A2(n2303), .ZN(n2359) );
  CKND2D1BWP12T U1030 ( .A1(n524), .A2(n2831), .ZN(n2363) );
  OAI21D1BWP12T U1031 ( .A1(n2362), .A2(n2359), .B(n2363), .ZN(n525) );
  AOI21D1BWP12T U1032 ( .A1(n892), .A2(n526), .B(n525), .ZN(n1575) );
  CKBD1BWP12T U1033 ( .I(n2620), .Z(n527) );
  NR2D1BWP12T U1034 ( .A1(n527), .A2(b[5]), .ZN(n1576) );
  NR2D1BWP12T U1035 ( .A1(n528), .A2(n2528), .ZN(n2375) );
  NR2D1BWP12T U1036 ( .A1(n2375), .A2(n2373), .ZN(n530) );
  ND2D1BWP12T U1037 ( .A1(n2370), .A2(n530), .ZN(n532) );
  CKND2D1BWP12T U1038 ( .A1(n2868), .A2(n2871), .ZN(n2366) );
  CKND2D1BWP12T U1039 ( .A1(n527), .A2(b[5]), .ZN(n1577) );
  OAI21D1BWP12T U1040 ( .A1(n1576), .A2(n2366), .B(n1577), .ZN(n2371) );
  CKND2D1BWP12T U1041 ( .A1(n528), .A2(n2528), .ZN(n2376) );
  OAI21D1BWP12T U1042 ( .A1(n2375), .A2(n2372), .B(n2376), .ZN(n529) );
  AOI21D1BWP12T U1043 ( .A1(n2371), .A2(n530), .B(n529), .ZN(n531) );
  OAI21D1BWP12T U1044 ( .A1(n1575), .A2(n532), .B(n531), .ZN(n633) );
  CKBD1BWP12T U1045 ( .I(n2301), .Z(n533) );
  OR2XD1BWP12T U1046 ( .A1(n533), .A2(b[9]), .Z(n635) );
  ND3D1BWP12T U1047 ( .A1(n536), .A2(n544), .A3(n670), .ZN(n2495) );
  INVD1BWP12T U1048 ( .I(n2495), .ZN(n2886) );
  CKND2D0BWP12T U1049 ( .A1(n1855), .A2(n2115), .ZN(n538) );
  CKND2D2BWP12T U1050 ( .A1(n2115), .A2(n2870), .ZN(n2135) );
  AOI21D0BWP12T U1051 ( .A1(n538), .A2(n2135), .B(n537), .ZN(n1936) );
  INVD0BWP12T U1052 ( .I(n999), .ZN(n982) );
  OR2D2BWP12T U1053 ( .A1(n2639), .A2(n2477), .Z(n2126) );
  IND2D1BWP12T U1054 ( .A1(n2639), .B1(n2477), .ZN(n2128) );
  OAI22D0BWP12T U1055 ( .A1(n982), .A2(n2126), .B1(n994), .B2(n2128), .ZN(n541) );
  NR2D1BWP12T U1056 ( .A1(n471), .A2(n2477), .ZN(n2166) );
  INVD1BWP12T U1057 ( .I(n2166), .ZN(n2119) );
  OAI22D0BWP12T U1058 ( .A1(n2119), .A2(n986), .B1(n987), .B2(n2116), .ZN(n540) );
  NR2D1BWP12T U1059 ( .A1(n541), .A2(n540), .ZN(n2201) );
  INVD1BWP12T U1060 ( .I(n2126), .ZN(n2173) );
  ND2D1BWP12T U1061 ( .A1(n1000), .A2(n2173), .ZN(n2474) );
  NR2D1BWP12T U1062 ( .A1(op[3]), .A2(n542), .ZN(n2786) );
  INVD1BWP12T U1063 ( .I(n2786), .ZN(n2942) );
  NR2D1BWP12T U1064 ( .A1(n2135), .A2(n2942), .ZN(n2513) );
  INVD1BWP12T U1065 ( .I(n2513), .ZN(n2901) );
  ND3D1BWP12T U1066 ( .A1(n543), .A2(op[2]), .A3(op[1]), .ZN(n2806) );
  INVD1BWP12T U1067 ( .I(n2806), .ZN(n2947) );
  AN3D1BWP12T U1068 ( .A1(op[0]), .A2(n545), .A3(n544), .Z(n2480) );
  INVD1BWP12T U1069 ( .I(n2480), .ZN(n2944) );
  CKND2D1BWP12T U1070 ( .A1(op[3]), .A2(op[2]), .ZN(n548) );
  OAI21D0BWP12T U1071 ( .A1(n2301), .A2(n2944), .B(n2949), .ZN(n546) );
  AOI22D0BWP12T U1072 ( .A1(n2947), .A2(n2243), .B1(n546), .B2(b[9]), .ZN(n552) );
  ND2D1BWP12T U1073 ( .A1(n671), .A2(n670), .ZN(n2951) );
  ND2D1BWP12T U1074 ( .A1(op[1]), .A2(n547), .ZN(n572) );
  NR2D0BWP12T U1075 ( .A1(n572), .A2(n548), .ZN(n2264) );
  TPND2D0BWP12T U1076 ( .A1(n2283), .A2(n2948), .ZN(n549) );
  OAI211D0BWP12T U1077 ( .A1(n2283), .A2(n2951), .B(n549), .C(n2949), .ZN(n550) );
  CKND2D0BWP12T U1078 ( .A1(n550), .A2(n2301), .ZN(n551) );
  OAI211D1BWP12T U1079 ( .A1(n2195), .A2(n2901), .B(n552), .C(n551), .ZN(n553)
         );
  AOI21D1BWP12T U1080 ( .A1(n2886), .A2(n1936), .B(n553), .ZN(n554) );
  IOA21D1BWP12T U1081 ( .A1(n2377), .A2(n2967), .B(n554), .ZN(n555) );
  AOI211D1BWP12T U1082 ( .A1(n2940), .A2(n1824), .B(n556), .C(n555), .ZN(n575)
         );
  NR2D1BWP12T U1083 ( .A1(n2482), .A2(n557), .ZN(n1601) );
  NR2D1BWP12T U1084 ( .A1(n558), .A2(n2303), .ZN(n881) );
  NR2D1BWP12T U1085 ( .A1(n1601), .A2(n881), .ZN(n560) );
  NR2XD0BWP12T U1086 ( .A1(n2302), .A2(c_in), .ZN(n1556) );
  CKND2D1BWP12T U1087 ( .A1(n2302), .A2(c_in), .ZN(n1557) );
  OAI21D1BWP12T U1088 ( .A1(n2231), .A2(n1556), .B(n1557), .ZN(n880) );
  CKND2D1BWP12T U1089 ( .A1(n2482), .A2(n557), .ZN(n1602) );
  CKND2D1BWP12T U1090 ( .A1(n558), .A2(n2303), .ZN(n882) );
  OAI21D1BWP12T U1091 ( .A1(n881), .A2(n1602), .B(n882), .ZN(n559) );
  AOI21D1BWP12T U1092 ( .A1(n560), .A2(n880), .B(n559), .ZN(n1586) );
  NR2D1BWP12T U1093 ( .A1(n562), .A2(n2871), .ZN(n1610) );
  NR2D1BWP12T U1094 ( .A1(n564), .A2(n2574), .ZN(n1630) );
  NR2D1BWP12T U1095 ( .A1(n1625), .A2(n1630), .ZN(n566) );
  CKND2D1BWP12T U1096 ( .A1(n1621), .A2(n566), .ZN(n568) );
  ND2D1BWP12T U1097 ( .A1(n2830), .A2(n561), .ZN(n1615) );
  CKND2D1BWP12T U1098 ( .A1(n562), .A2(n2871), .ZN(n1611) );
  OAI21D1BWP12T U1099 ( .A1(n1610), .A2(n1615), .B(n1611), .ZN(n1623) );
  ND2D1BWP12T U1100 ( .A1(n2620), .A2(n563), .ZN(n1624) );
  ND2D1BWP12T U1101 ( .A1(n564), .A2(n2574), .ZN(n1631) );
  OAI21D1BWP12T U1102 ( .A1(n1624), .A2(n1630), .B(n1631), .ZN(n565) );
  AOI21D1BWP12T U1103 ( .A1(n566), .A2(n1623), .B(n565), .ZN(n567) );
  OAI21D1BWP12T U1104 ( .A1(n1586), .A2(n568), .B(n567), .ZN(n1619) );
  INVD1BWP12T U1105 ( .I(n1619), .ZN(n1639) );
  OR2XD1BWP12T U1106 ( .A1(n571), .A2(a[8]), .Z(n1620) );
  ND2D1BWP12T U1107 ( .A1(n1618), .A2(n1620), .ZN(n1635) );
  ND2D1BWP12T U1108 ( .A1(n570), .A2(n569), .ZN(n1608) );
  INVD1BWP12T U1109 ( .I(n1608), .ZN(n1617) );
  AOI21D1BWP12T U1110 ( .A1(n1617), .A2(n1620), .B(n618), .ZN(n1636) );
  ND2D1BWP12T U1111 ( .A1(n2301), .A2(n2283), .ZN(n1637) );
  NR2D1BWP12T U1112 ( .A1(n573), .A2(n572), .ZN(n2855) );
  CKND2D1BWP12T U1113 ( .A1(n1642), .A2(n2855), .ZN(n574) );
  ND4D1BWP12T U1114 ( .A1(n577), .A2(n576), .A3(n575), .A4(n574), .ZN(
        result[9]) );
  INVD6BWP12T U1115 ( .I(n2512), .ZN(n2594) );
  INVD6BWP12T U1116 ( .I(n2241), .ZN(n2643) );
  XOR2D1BWP12T U1117 ( .A1(n2308), .A2(n2643), .Z(n578) );
  CKND2D2BWP12T U1118 ( .A1(n2644), .A2(n578), .ZN(n2646) );
  XNR2D0BWP12T U1119 ( .A1(n2643), .A2(b[17]), .ZN(n1271) );
  XNR2XD0BWP12T U1120 ( .A1(n2643), .A2(b[18]), .ZN(n583) );
  TPOAI22D0BWP12T U1121 ( .A1(n2646), .A2(n1271), .B1(n2644), .B2(n583), .ZN(
        mult_x_18_n830) );
  INVD6BWP12T U1122 ( .I(n2683), .ZN(n2679) );
  XNR2XD4BWP12T U1123 ( .A1(n2679), .A2(a[18]), .ZN(n2610) );
  CKXOR2D1BWP12T U1124 ( .A1(a[18]), .A2(n2609), .Z(n579) );
  ND2D1BWP12T U1125 ( .A1(n2610), .A2(n579), .ZN(n2612) );
  XNR2XD1BWP12T U1126 ( .A1(n2609), .A2(n2897), .ZN(n1282) );
  XNR2XD1BWP12T U1127 ( .A1(n2609), .A2(b[11]), .ZN(n580) );
  TPOAI22D0BWP12T U1128 ( .A1(n2612), .A2(n1282), .B1(n2610), .B2(n580), .ZN(
        mult_x_18_n780) );
  XNR2XD0BWP12T U1129 ( .A1(n2609), .A2(n2598), .ZN(n1035) );
  TPOAI22D0BWP12T U1130 ( .A1(n2612), .A2(n580), .B1(n2610), .B2(n1035), .ZN(
        mult_x_18_n779) );
  XNR2D0BWP12T U1131 ( .A1(n2482), .A2(b[29]), .ZN(n1030) );
  XNR2D0BWP12T U1132 ( .A1(n2482), .A2(b[30]), .ZN(n1037) );
  OAI22D0BWP12T U1133 ( .A1(n2604), .A2(n1030), .B1(n1037), .B2(n2603), .ZN(
        mult_x_18_n986) );
  XNR2D2BWP12T U1134 ( .A1(a[22]), .A2(n2725), .ZN(n2630) );
  INVD3BWP12T U1135 ( .I(n2751), .ZN(n2747) );
  XOR2XD1BWP12T U1136 ( .A1(n2747), .A2(a[22]), .Z(n581) );
  CKND2D2BWP12T U1137 ( .A1(n2630), .A2(n581), .ZN(n2632) );
  XNR2XD1BWP12T U1138 ( .A1(n2747), .A2(n2528), .ZN(n1090) );
  XNR2XD1BWP12T U1139 ( .A1(n2747), .A2(n2605), .ZN(n1042) );
  OAI22D1BWP12T U1140 ( .A1(n2632), .A2(n1090), .B1(n1042), .B2(n2630), .ZN(
        mult_x_18_n755) );
  INVD6BWP12T U1141 ( .I(n2240), .ZN(n2626) );
  XNR2D2BWP12T U1142 ( .A1(n2626), .A2(a[16]), .ZN(n2647) );
  XOR2XD1BWP12T U1143 ( .A1(n2679), .A2(a[16]), .Z(n582) );
  ND2D4BWP12T U1144 ( .A1(n2647), .A2(n582), .ZN(n2649) );
  XNR2XD0BWP12T U1145 ( .A1(n2679), .A2(b[14]), .ZN(n1286) );
  XNR2XD0BWP12T U1146 ( .A1(n2679), .A2(b[15]), .ZN(n2648) );
  OAI22D0BWP12T U1147 ( .A1(n2649), .A2(n1286), .B1(n2648), .B2(n2647), .ZN(
        mult_x_18_n793) );
  XNR2XD0BWP12T U1148 ( .A1(n2643), .A2(b[19]), .ZN(n2645) );
  OAI22D0BWP12T U1149 ( .A1(n2646), .A2(n583), .B1(n2644), .B2(n2645), .ZN(
        mult_x_18_n829) );
  XNR2XD4BWP12T U1150 ( .A1(a[14]), .A2(n2643), .ZN(n2627) );
  CKXOR2D1BWP12T U1151 ( .A1(a[14]), .A2(n2626), .Z(n584) );
  CKND2D3BWP12T U1152 ( .A1(n2627), .A2(n584), .ZN(n2629) );
  XNR2XD0BWP12T U1153 ( .A1(n2626), .A2(b[14]), .ZN(n1031) );
  XNR2XD0BWP12T U1154 ( .A1(n2626), .A2(b[15]), .ZN(n1032) );
  TPOAI22D0BWP12T U1155 ( .A1(n2629), .A2(n1031), .B1(n2627), .B2(n1032), .ZN(
        mult_x_18_n812) );
  INVD1BWP12T U1156 ( .I(n2977), .ZN(n2822) );
  CKND2D1BWP12T U1157 ( .A1(n425), .A2(n1669), .ZN(n609) );
  NR2D1BWP12T U1158 ( .A1(mult_x_18_n585), .A2(mult_x_18_n598), .ZN(n776) );
  NR2D1BWP12T U1159 ( .A1(mult_x_18_n599), .A2(mult_x_18_n610), .ZN(n774) );
  NR2D1BWP12T U1160 ( .A1(n776), .A2(n774), .ZN(n1720) );
  CKND2D1BWP12T U1161 ( .A1(n1723), .A2(n1720), .ZN(n605) );
  OR2D2BWP12T U1162 ( .A1(mult_x_18_n635), .A2(mult_x_18_n645), .Z(n1426) );
  OR2D2BWP12T U1163 ( .A1(mult_x_18_n654), .A2(mult_x_18_n646), .Z(n1423) );
  CKND2D1BWP12T U1164 ( .A1(n1426), .A2(n1423), .ZN(n600) );
  NR2D1BWP12T U1165 ( .A1(mult_x_18_n665), .A2(mult_x_18_n672), .ZN(n585) );
  INVD1BWP12T U1166 ( .I(n585), .ZN(n917) );
  OR2XD1BWP12T U1167 ( .A1(mult_x_18_n673), .A2(mult_x_18_n680), .Z(n1685) );
  ND2D1BWP12T U1168 ( .A1(n917), .A2(n1685), .ZN(n596) );
  CKND2D1BWP12T U1169 ( .A1(n589), .A2(n1691), .ZN(n592) );
  INVD1BWP12T U1170 ( .I(n586), .ZN(n587) );
  AOI21D1BWP12T U1171 ( .A1(n589), .A2(n588), .B(n587), .ZN(n590) );
  TPOAI21D1BWP12T U1172 ( .A1(n592), .A2(n591), .B(n590), .ZN(n1689) );
  OR2D1BWP12T U1173 ( .A1(mult_x_18_n681), .A2(mult_x_18_n686), .Z(n1688) );
  ND2D1BWP12T U1174 ( .A1(mult_x_18_n681), .A2(mult_x_18_n686), .ZN(n1687) );
  INVD1BWP12T U1175 ( .I(n1687), .ZN(n593) );
  AOI21D1BWP12T U1176 ( .A1(n1689), .A2(n1688), .B(n593), .ZN(n914) );
  ND2D1BWP12T U1177 ( .A1(mult_x_18_n673), .A2(mult_x_18_n680), .ZN(n1684) );
  INVD1BWP12T U1178 ( .I(n1684), .ZN(n915) );
  ND2D1BWP12T U1179 ( .A1(mult_x_18_n665), .A2(mult_x_18_n672), .ZN(n916) );
  INVD1BWP12T U1180 ( .I(n916), .ZN(n594) );
  TPAOI21D1BWP12T U1181 ( .A1(n917), .A2(n915), .B(n594), .ZN(n595) );
  TPOAI21D1BWP12T U1182 ( .A1(n596), .A2(n914), .B(n595), .ZN(n971) );
  OR2XD1BWP12T U1183 ( .A1(mult_x_18_n655), .A2(mult_x_18_n664), .Z(n970) );
  ND2D1BWP12T U1184 ( .A1(mult_x_18_n655), .A2(mult_x_18_n664), .ZN(n969) );
  INVD1BWP12T U1185 ( .I(n969), .ZN(n597) );
  TPAOI21D1BWP12T U1186 ( .A1(n971), .A2(n970), .B(n597), .ZN(n814) );
  ND2D1BWP12T U1187 ( .A1(mult_x_18_n654), .A2(mult_x_18_n646), .ZN(n815) );
  INVD1BWP12T U1188 ( .I(n815), .ZN(n1422) );
  ND2D1BWP12T U1189 ( .A1(mult_x_18_n635), .A2(mult_x_18_n645), .ZN(n1425) );
  INVD1BWP12T U1190 ( .I(n1425), .ZN(n598) );
  TPAOI21D1BWP12T U1191 ( .A1(n1426), .A2(n1422), .B(n598), .ZN(n599) );
  TPOAI21D1BWP12T U1192 ( .A1(n600), .A2(n814), .B(n599), .ZN(n1387) );
  NR2D1BWP12T U1193 ( .A1(mult_x_18_n623), .A2(mult_x_18_n611), .ZN(n1679) );
  NR2D1BWP12T U1194 ( .A1(mult_x_18_n624), .A2(mult_x_18_n634), .ZN(n1677) );
  NR2D1BWP12T U1195 ( .A1(n1679), .A2(n1677), .ZN(n602) );
  ND2D1BWP12T U1196 ( .A1(mult_x_18_n624), .A2(mult_x_18_n634), .ZN(n1676) );
  ND2D1BWP12T U1197 ( .A1(mult_x_18_n623), .A2(mult_x_18_n611), .ZN(n1680) );
  OAI21D1BWP12T U1198 ( .A1(n1679), .A2(n1676), .B(n1680), .ZN(n601) );
  TPAOI21D1BWP12T U1199 ( .A1(n1387), .A2(n602), .B(n601), .ZN(n773) );
  ND2D1BWP12T U1200 ( .A1(mult_x_18_n599), .A2(mult_x_18_n610), .ZN(n1674) );
  ND2D1BWP12T U1201 ( .A1(mult_x_18_n585), .A2(mult_x_18_n598), .ZN(n777) );
  OAI21D1BWP12T U1202 ( .A1(n776), .A2(n1674), .B(n777), .ZN(n1719) );
  ND2D1BWP12T U1203 ( .A1(mult_x_18_n571), .A2(mult_x_18_n584), .ZN(n1722) );
  INVD1BWP12T U1204 ( .I(n1722), .ZN(n603) );
  AOI21D1BWP12T U1205 ( .A1(n1723), .A2(n1719), .B(n603), .ZN(n604) );
  OAI21D1BWP12T U1206 ( .A1(n605), .A2(n773), .B(n604), .ZN(n1729) );
  OR2D1BWP12T U1207 ( .A1(mult_x_18_n555), .A2(mult_x_18_n570), .Z(n1728) );
  ND2D1BWP12T U1208 ( .A1(mult_x_18_n555), .A2(mult_x_18_n570), .ZN(n1727) );
  INVD1BWP12T U1209 ( .I(n1727), .ZN(n606) );
  AOI21D1BWP12T U1210 ( .A1(n1729), .A2(n1728), .B(n606), .ZN(n735) );
  ND2D1BWP12T U1211 ( .A1(mult_x_18_n540), .A2(mult_x_18_n554), .ZN(n734) );
  INVD1BWP12T U1212 ( .I(n734), .ZN(n1668) );
  ND2D1BWP12T U1213 ( .A1(mult_x_18_n539), .A2(mult_x_18_n523), .ZN(n1671) );
  INVD1BWP12T U1214 ( .I(n1671), .ZN(n607) );
  AOI21D1BWP12T U1215 ( .A1(n425), .A2(n1668), .B(n607), .ZN(n608) );
  TPOAI21D1BWP12T U1216 ( .A1(n609), .A2(n735), .B(n608), .ZN(n693) );
  NR2XD0BWP12T U1217 ( .A1(mult_x_18_n487), .A2(mult_x_18_n505), .ZN(n694) );
  NR2D1BWP12T U1218 ( .A1(mult_x_18_n506), .A2(mult_x_18_n522), .ZN(n1730) );
  NR2D1BWP12T U1219 ( .A1(n694), .A2(n1730), .ZN(n611) );
  ND2D1BWP12T U1220 ( .A1(mult_x_18_n506), .A2(mult_x_18_n522), .ZN(n1731) );
  ND2D1BWP12T U1221 ( .A1(mult_x_18_n487), .A2(mult_x_18_n505), .ZN(n695) );
  OAI21D1BWP12T U1222 ( .A1(n694), .A2(n1731), .B(n695), .ZN(n610) );
  INVD1BWP12T U1223 ( .I(n1665), .ZN(n1662) );
  NR2D1BWP12T U1224 ( .A1(mult_x_18_n486), .A2(mult_x_18_n469), .ZN(n1664) );
  INVD1BWP12T U1225 ( .I(n1664), .ZN(n1661) );
  OR2XD1BWP12T U1226 ( .A1(mult_x_18_n468), .A2(mult_x_18_n449), .Z(n1667) );
  AN2XD1BWP12T U1227 ( .A1(n1661), .A2(n1667), .Z(n615) );
  ND2D1BWP12T U1228 ( .A1(mult_x_18_n486), .A2(mult_x_18_n469), .ZN(n1663) );
  CKND0BWP12T U1229 ( .I(n1663), .ZN(n613) );
  ND2D1BWP12T U1230 ( .A1(mult_x_18_n468), .A2(mult_x_18_n449), .ZN(n1666) );
  INVD1BWP12T U1231 ( .I(n1666), .ZN(n612) );
  AO21D1BWP12T U1232 ( .A1(n1667), .A2(n613), .B(n612), .Z(n614) );
  AO21D1BWP12T U1233 ( .A1(n1662), .A2(n615), .B(n614), .Z(n1454) );
  INVD1BWP12T U1234 ( .I(n2656), .ZN(n1742) );
  INVD1BWP12T U1235 ( .I(b[23]), .ZN(n2406) );
  INVD1BWP12T U1236 ( .I(b[22]), .ZN(n737) );
  INVD1BWP12T U1237 ( .I(b[21]), .ZN(n2408) );
  INVD1BWP12T U1238 ( .I(b[20]), .ZN(n2410) );
  INVD1BWP12T U1239 ( .I(b[19]), .ZN(n782) );
  NR2D1BWP12T U1240 ( .A1(n2594), .A2(n2511), .ZN(n2451) );
  INVD2BWP12T U1241 ( .I(n2898), .ZN(n2900) );
  NR2D1BWP12T U1242 ( .A1(n2899), .A2(n2900), .ZN(n2445) );
  OR2XD1BWP12T U1243 ( .A1(n2451), .A2(n2445), .Z(n620) );
  ND2D1BWP12T U1244 ( .A1(n424), .A2(n2436), .ZN(n2446) );
  OR2XD1BWP12T U1245 ( .A1(n620), .A2(n2446), .Z(n622) );
  AOI21D1BWP12T U1246 ( .A1(n424), .A2(n618), .B(n1638), .ZN(n2447) );
  CKND2D1BWP12T U1247 ( .A1(n2899), .A2(n2900), .ZN(n2448) );
  CKND2D1BWP12T U1248 ( .A1(n2594), .A2(n2511), .ZN(n2452) );
  OA21D1BWP12T U1249 ( .A1(n2451), .A2(n2448), .B(n2452), .Z(n619) );
  OA21D1BWP12T U1250 ( .A1(n2447), .A2(n620), .B(n619), .Z(n621) );
  RCOAI21D1BWP12T U1251 ( .A1(n2450), .A2(n622), .B(n621), .ZN(n922) );
  OR2XD1BWP12T U1252 ( .A1(n2277), .A2(n2308), .Z(n921) );
  CKND2D1BWP12T U1253 ( .A1(n2277), .A2(n2308), .ZN(n920) );
  INVD1BWP12T U1254 ( .I(n920), .ZN(n623) );
  TPAOI21D1BWP12T U1255 ( .A1(n922), .A2(n921), .B(n623), .ZN(n975) );
  NR2XD0BWP12T U1256 ( .A1(n2643), .A2(n2278), .ZN(n972) );
  ND2D1BWP12T U1257 ( .A1(n2643), .A2(n2278), .ZN(n973) );
  TPOAI21D1BWP12T U1258 ( .A1(n975), .A2(n972), .B(n973), .ZN(n849) );
  OR2XD1BWP12T U1259 ( .A1(n2275), .A2(a[14]), .Z(n848) );
  CKND2D1BWP12T U1260 ( .A1(n2275), .A2(a[14]), .ZN(n847) );
  INVD1BWP12T U1261 ( .I(n847), .ZN(n624) );
  TPAOI21D1BWP12T U1262 ( .A1(n849), .A2(n848), .B(n624), .ZN(n1435) );
  NR2D1BWP12T U1263 ( .A1(n2626), .A2(n2276), .ZN(n1433) );
  ND2D1BWP12T U1264 ( .A1(n2626), .A2(n2276), .ZN(n1434) );
  TPOAI21D1BWP12T U1265 ( .A1(n1435), .A2(n1433), .B(n1434), .ZN(n1395) );
  INVD1BWP12T U1266 ( .I(b[16]), .ZN(n2270) );
  OR2XD1BWP12T U1267 ( .A1(n2270), .A2(a[16]), .Z(n1394) );
  CKND2D1BWP12T U1268 ( .A1(n2270), .A2(a[16]), .ZN(n1393) );
  INVD1BWP12T U1269 ( .I(n1393), .ZN(n625) );
  AOI21D1BWP12T U1270 ( .A1(n1395), .A2(n1394), .B(n625), .ZN(n2416) );
  INVD1BWP12T U1271 ( .I(b[17]), .ZN(n2678) );
  NR2D0BWP12T U1272 ( .A1(n2679), .A2(n2678), .ZN(n2414) );
  CKND2D1BWP12T U1273 ( .A1(n2679), .A2(n2678), .ZN(n2415) );
  OAI21D1BWP12T U1274 ( .A1(n2416), .A2(n2414), .B(n2415), .ZN(n2413) );
  OR2XD1BWP12T U1275 ( .A1(n2703), .A2(a[18]), .Z(n2412) );
  CKND2D1BWP12T U1276 ( .A1(n2703), .A2(a[18]), .ZN(n2411) );
  INVD1BWP12T U1277 ( .I(n2411), .ZN(n626) );
  AO21D1BWP12T U1278 ( .A1(n2413), .A2(n2412), .B(n626), .Z(n781) );
  NR2D1BWP12T U1279 ( .A1(n2897), .A2(n2900), .ZN(n1752) );
  OR2XD1BWP12T U1280 ( .A1(n627), .A2(n1752), .Z(n629) );
  OR2XD1BWP12T U1281 ( .A1(n629), .A2(n1748), .Z(n631) );
  ND2D1BWP12T U1282 ( .A1(n2897), .A2(n2900), .ZN(n2346) );
  OA21D1BWP12T U1283 ( .A1(n1750), .A2(n1752), .B(n2346), .Z(n628) );
  OA21D1BWP12T U1284 ( .A1(n629), .A2(n1749), .B(n628), .Z(n630) );
  TPOAI21D2BWP12T U1285 ( .A1(n1772), .A2(n631), .B(n630), .ZN(n1747) );
  OR2XD1BWP12T U1286 ( .A1(n2594), .A2(b[11]), .Z(n2349) );
  ND2D1BWP12T U1287 ( .A1(n2594), .A2(b[11]), .ZN(n2348) );
  INVD1BWP12T U1288 ( .I(n2348), .ZN(n638) );
  AOI21D1BWP12T U1289 ( .A1(n1747), .A2(n2349), .B(n638), .ZN(n946) );
  NR2D1BWP12T U1290 ( .A1(n2598), .A2(n2308), .ZN(n945) );
  ND2D1BWP12T U1291 ( .A1(n2598), .A2(n2308), .ZN(n953) );
  OR2XD1BWP12T U1292 ( .A1(n2643), .A2(b[13]), .Z(n1012) );
  ND2D1BWP12T U1293 ( .A1(n2643), .A2(b[13]), .ZN(n1011) );
  INVD1BWP12T U1294 ( .I(n1011), .ZN(n639) );
  TPAOI21D2BWP12T U1295 ( .A1(n1010), .A2(n1012), .B(n639), .ZN(n817) );
  NR2D1BWP12T U1296 ( .A1(a[14]), .A2(b[14]), .ZN(n816) );
  ND2D1BWP12T U1297 ( .A1(a[14]), .A2(b[14]), .ZN(n818) );
  TPOAI21D2BWP12T U1298 ( .A1(n817), .A2(n816), .B(n818), .ZN(n1436) );
  OR2XD1BWP12T U1299 ( .A1(n2626), .A2(b[15]), .Z(n1438) );
  ND2D1BWP12T U1300 ( .A1(n2626), .A2(b[15]), .ZN(n1437) );
  INVD1BWP12T U1301 ( .I(n1437), .ZN(n640) );
  TPAOI21D2BWP12T U1302 ( .A1(n1436), .A2(n1438), .B(n640), .ZN(n1419) );
  NR2D1BWP12T U1303 ( .A1(a[16]), .A2(b[16]), .ZN(n1396) );
  ND2D1BWP12T U1304 ( .A1(a[16]), .A2(b[16]), .ZN(n1417) );
  OAI21D1BWP12T U1305 ( .A1(n1419), .A2(n1396), .B(n1417), .ZN(n1746) );
  OR2XD1BWP12T U1306 ( .A1(n2679), .A2(b[17]), .Z(n2342) );
  ND2D1BWP12T U1307 ( .A1(n2679), .A2(b[17]), .ZN(n2341) );
  INVD1BWP12T U1308 ( .I(n2341), .ZN(n641) );
  TPAOI21D2BWP12T U1309 ( .A1(n1746), .A2(n2342), .B(n641), .ZN(n1794) );
  NR2D1BWP12T U1310 ( .A1(a[18]), .A2(b[18]), .ZN(n1793) );
  ND2D1BWP12T U1311 ( .A1(a[18]), .A2(b[18]), .ZN(n2337) );
  OR2XD1BWP12T U1312 ( .A1(n2609), .A2(b[19]), .Z(n785) );
  ND2D1BWP12T U1313 ( .A1(n2609), .A2(b[19]), .ZN(n784) );
  INVD1BWP12T U1314 ( .I(n784), .ZN(n642) );
  AO21D1BWP12T U1315 ( .A1(n783), .A2(n785), .B(n642), .Z(n1745) );
  INVD1BWP12T U1316 ( .I(n633), .ZN(n2369) );
  ND2D1BWP12T U1317 ( .A1(n635), .A2(n2368), .ZN(n2345) );
  OR2XD1BWP12T U1318 ( .A1(n2345), .A2(n1752), .Z(n637) );
  AOI21D1BWP12T U1319 ( .A1(n635), .A2(n634), .B(n1751), .ZN(n2344) );
  OA21D1BWP12T U1320 ( .A1(n2344), .A2(n1752), .B(n2346), .Z(n636) );
  TPAOI21D2BWP12T U1321 ( .A1(n2350), .A2(n2349), .B(n638), .ZN(n955) );
  TPOAI21D2BWP12T U1322 ( .A1(n955), .A2(n945), .B(n953), .ZN(n1013) );
  TPAOI21D2BWP12T U1323 ( .A1(n1013), .A2(n1012), .B(n639), .ZN(n821) );
  TPOAI21D2BWP12T U1324 ( .A1(n821), .A2(n816), .B(n818), .ZN(n1440) );
  TPAOI21D2BWP12T U1325 ( .A1(n1440), .A2(n1438), .B(n640), .ZN(n1397) );
  TPAOI21D1BWP12T U1326 ( .A1(n2343), .A2(n2342), .B(n641), .ZN(n2340) );
  TPOAI21D1BWP12T U1327 ( .A1(n2340), .A2(n1793), .B(n2337), .ZN(n787) );
  AO21D1BWP12T U1328 ( .A1(n787), .A2(n785), .B(n642), .Z(n2336) );
  ND2D1BWP12T U1329 ( .A1(n2398), .A2(n2967), .ZN(n683) );
  INVD1BWP12T U1330 ( .I(a[25]), .ZN(n1108) );
  INVD1BWP12T U1331 ( .I(a[20]), .ZN(n1829) );
  INVD1BWP12T U1332 ( .I(n2609), .ZN(n1223) );
  INVD8BWP12T U1333 ( .I(n2301), .ZN(n1049) );
  ND2D1BWP12T U1334 ( .A1(n1049), .A2(n2550), .ZN(n1822) );
  INVD1BWP12T U1335 ( .I(n2594), .ZN(n1311) );
  INVD1BWP12T U1336 ( .I(n2643), .ZN(n1061) );
  CKND2D1BWP12T U1337 ( .A1(n1061), .A2(n2242), .ZN(n835) );
  INVD1BWP12T U1338 ( .I(n2626), .ZN(n1219) );
  CKND0BWP12T U1339 ( .I(a[14]), .ZN(n1441) );
  TPND2D0BWP12T U1340 ( .A1(n1219), .A2(n1441), .ZN(n643) );
  NR2XD0BWP12T U1341 ( .A1(n835), .A2(n643), .ZN(n644) );
  CKND2D1BWP12T U1342 ( .A1(n833), .A2(n644), .ZN(n645) );
  NR2D1BWP12T U1343 ( .A1(n645), .A2(n834), .ZN(n1405) );
  XNR2D1BWP12T U1344 ( .A1(n2665), .A2(a[31]), .ZN(n2666) );
  NR2D1BWP12T U1345 ( .A1(n2017), .A2(n1997), .ZN(n2008) );
  ND2D1BWP12T U1346 ( .A1(n1998), .A2(n1997), .ZN(n2023) );
  MUX2XD0BWP12T U1347 ( .I0(n2609), .I1(a[18]), .S(n2231), .Z(n657) );
  MUX2NXD0BWP12T U1348 ( .I0(n2725), .I1(a[20]), .S(n2231), .ZN(n2143) );
  MUX2NXD0BWP12T U1349 ( .I0(n2679), .I1(a[16]), .S(n2231), .ZN(n1513) );
  AOI22D0BWP12T U1350 ( .A1(n2001), .A2(n2143), .B1(n2000), .B2(n1513), .ZN(
        n647) );
  MUX2NXD0BWP12T U1351 ( .I0(n2747), .I1(a[22]), .S(n2231), .ZN(n2142) );
  TPND2D0BWP12T U1352 ( .A1(n2002), .A2(n2142), .ZN(n646) );
  OAI211D0BWP12T U1353 ( .A1(n657), .A2(n1959), .B(n647), .C(n646), .ZN(n1987)
         );
  OR2XD1BWP12T U1354 ( .A1(n2831), .A2(n2868), .Z(n2202) );
  NR2D1BWP12T U1355 ( .A1(n648), .A2(n2202), .ZN(n2006) );
  NR2D0BWP12T U1356 ( .A1(n1997), .A2(n2006), .ZN(n649) );
  ND2D1BWP12T U1357 ( .A1(n649), .A2(n2017), .ZN(n2022) );
  MUX2NXD0BWP12T U1358 ( .I0(n2626), .I1(a[14]), .S(n2231), .ZN(n1512) );
  TPNR2D0BWP12T U1359 ( .A1(n1940), .A2(n1512), .ZN(n652) );
  MUX2NXD0BWP12T U1360 ( .I0(n2594), .I1(n2900), .S(n2231), .ZN(n985) );
  NR2D0BWP12T U1361 ( .A1(n1959), .A2(n985), .ZN(n651) );
  INVD1BWP12T U1362 ( .I(n2000), .ZN(n1941) );
  INVD1BWP12T U1363 ( .I(n2001), .ZN(n1501) );
  MUX2NXD0BWP12T U1364 ( .I0(n2643), .I1(n2308), .S(n2231), .ZN(n792) );
  OAI22D0BWP12T U1365 ( .A1(n1941), .A2(n999), .B1(n1501), .B2(n792), .ZN(n650) );
  NR3D1BWP12T U1366 ( .A1(n652), .A2(n651), .A3(n650), .ZN(n1986) );
  CKND2D3BWP12T U1367 ( .A1(n2017), .A2(n1997), .ZN(n2025) );
  MUX2NXD0BWP12T U1368 ( .I0(a[27]), .I1(a[26]), .S(n2231), .ZN(n2140) );
  TPNR2D0BWP12T U1369 ( .A1(n1959), .A2(n2140), .ZN(n654) );
  MUX2NXD0BWP12T U1370 ( .I0(a[25]), .I1(a[24]), .S(n2231), .ZN(n2141) );
  MUX2NXD0BWP12T U1371 ( .I0(a[29]), .I1(a[28]), .S(n2231), .ZN(n664) );
  TPOAI22D0BWP12T U1372 ( .A1(n1941), .A2(n2141), .B1(n1501), .B2(n664), .ZN(
        n653) );
  AOI211D0BWP12T U1373 ( .A1(n2002), .A2(a[30]), .B(n654), .C(n653), .ZN(n655)
         );
  OAI222D1BWP12T U1374 ( .A1(n2023), .A2(n1987), .B1(n2022), .B2(n1986), .C1(
        n2025), .C2(n655), .ZN(n1952) );
  AOI21D1BWP12T U1375 ( .A1(n2008), .A2(n2526), .B(n1952), .ZN(n656) );
  NR2D1BWP12T U1376 ( .A1(n656), .A2(n2964), .ZN(n681) );
  NR2D1BWP12T U1377 ( .A1(n2135), .A2(n2495), .ZN(n2775) );
  NR2D1BWP12T U1378 ( .A1(n2868), .A2(n2964), .ZN(n2893) );
  NR2D1BWP12T U1379 ( .A1(n2775), .A2(n2893), .ZN(n2675) );
  ND3D0BWP12T U1380 ( .A1(n1891), .A2(a[31]), .A3(n2827), .ZN(n1850) );
  NR2D1BWP12T U1381 ( .A1(n2827), .A2(n2868), .ZN(n2155) );
  INVD1BWP12T U1382 ( .I(n2128), .ZN(n2170) );
  AOI22D0BWP12T U1383 ( .A1(n2170), .A2(n2143), .B1(n2142), .B2(n2173), .ZN(
        n659) );
  INVD1BWP12T U1384 ( .I(n2116), .ZN(n2169) );
  INVD1BWP12T U1385 ( .I(n657), .ZN(n1511) );
  AOI22D0BWP12T U1386 ( .A1(n2169), .A2(n1513), .B1(n1511), .B2(n2166), .ZN(
        n658) );
  ND2D1BWP12T U1387 ( .A1(n659), .A2(n658), .ZN(n2177) );
  INVD1BWP12T U1388 ( .I(n792), .ZN(n996) );
  INVD0BWP12T U1389 ( .I(n1512), .ZN(n711) );
  OAI22D0BWP12T U1390 ( .A1(n996), .A2(n2128), .B1(n711), .B2(n2126), .ZN(n661) );
  NR2D0BWP12T U1391 ( .A1(n982), .A2(n2116), .ZN(n660) );
  RCAOI211D0BWP12T U1392 ( .A1(n2166), .A2(n985), .B(n661), .C(n660), .ZN(
        n2176) );
  IND2XD1BWP12T U1393 ( .A1(n2831), .B1(n2868), .ZN(n2159) );
  OAI22D0BWP12T U1394 ( .A1(n1000), .A2(n2116), .B1(n986), .B2(n2128), .ZN(
        n663) );
  NR2XD0BWP12T U1395 ( .A1(n994), .A2(n2126), .ZN(n662) );
  AOI211D1BWP12T U1396 ( .A1(n2166), .A2(n1003), .B(n663), .C(n662), .ZN(n2179) );
  OAI22D0BWP12T U1397 ( .A1(n2176), .A2(n2159), .B1(n2179), .B2(n2080), .ZN(
        n669) );
  CKND0BWP12T U1398 ( .I(n2006), .ZN(n1360) );
  CKND0BWP12T U1399 ( .I(n2140), .ZN(n1516) );
  CKND2D1BWP12T U1400 ( .A1(n2173), .A2(n2231), .ZN(n1548) );
  OAI22D0BWP12T U1401 ( .A1(n1516), .A2(n2119), .B1(a[30]), .B2(n1548), .ZN(
        n666) );
  INVD0BWP12T U1402 ( .I(n2141), .ZN(n1518) );
  INVD0BWP12T U1403 ( .I(n664), .ZN(n1517) );
  OAI22D0BWP12T U1404 ( .A1(n1518), .A2(n2116), .B1(n1517), .B2(n2128), .ZN(
        n665) );
  INVD1BWP12T U1405 ( .I(n2202), .ZN(n2769) );
  OAI21D0BWP12T U1406 ( .A1(n666), .A2(n665), .B(n2769), .ZN(n667) );
  OAI211D0BWP12T U1407 ( .A1(a[31]), .A2(n1360), .B(n667), .C(n2115), .ZN(n668) );
  AOI211D1BWP12T U1408 ( .A1(n2155), .A2(n2177), .B(n669), .C(n668), .ZN(n2197) );
  ND2D1BWP12T U1409 ( .A1(n2197), .A2(n2786), .ZN(n679) );
  XNR2XD1BWP12T U1410 ( .A1(a[31]), .A2(b[31]), .ZN(n2663) );
  INVD1BWP12T U1411 ( .I(n2663), .ZN(n677) );
  CKND0BWP12T U1412 ( .I(b[31]), .ZN(n674) );
  TPND2D0BWP12T U1413 ( .A1(n674), .A2(n670), .ZN(n672) );
  AOI22D0BWP12T U1414 ( .A1(n672), .A2(n671), .B1(n2264), .B2(n674), .ZN(n673)
         );
  NR2D0BWP12T U1415 ( .A1(n673), .A2(n2310), .ZN(n676) );
  TPOAI22D0BWP12T U1416 ( .A1(n674), .A2(n2949), .B1(a[31]), .B2(n2806), .ZN(
        n675) );
  AOI211D1BWP12T U1417 ( .A1(n677), .A2(n2480), .B(n676), .C(n675), .ZN(n678)
         );
  OAI211D1BWP12T U1418 ( .A1(n2675), .A2(n1850), .B(n679), .C(n678), .ZN(n680)
         );
  AOI211D1BWP12T U1419 ( .A1(n2666), .A2(n2940), .B(n681), .C(n680), .ZN(n682)
         );
  NR2D1BWP12T U1420 ( .A1(n2899), .A2(n2900), .ZN(n1640) );
  OR2D0BWP12T U1421 ( .A1(n685), .A2(n1635), .Z(n687) );
  CKND2D1BWP12T U1422 ( .A1(n2899), .A2(n2900), .ZN(n1641) );
  OA21D1BWP12T U1423 ( .A1(n1637), .A2(n1640), .B(n1641), .Z(n684) );
  OA21D1BWP12T U1424 ( .A1(n685), .A2(n1636), .B(n684), .Z(n686) );
  OAI21D1BWP12T U1425 ( .A1(n1639), .A2(n687), .B(n686), .ZN(n1599) );
  OR2XD1BWP12T U1426 ( .A1(n2594), .A2(n2511), .Z(n1598) );
  ND2D1BWP12T U1427 ( .A1(n2594), .A2(n2511), .ZN(n1597) );
  INVD1BWP12T U1428 ( .I(n1597), .ZN(n688) );
  AOI21D1BWP12T U1429 ( .A1(n1599), .A2(n1598), .B(n688), .ZN(n925) );
  NR2XD0BWP12T U1430 ( .A1(n2277), .A2(n2308), .ZN(n923) );
  ND2D1BWP12T U1431 ( .A1(n2277), .A2(n2308), .ZN(n924) );
  OAI21D1BWP12T U1432 ( .A1(n925), .A2(n923), .B(n924), .ZN(n1017) );
  OR2XD1BWP12T U1433 ( .A1(n2643), .A2(n2278), .Z(n1015) );
  ND2D1BWP12T U1434 ( .A1(n2643), .A2(n2278), .ZN(n1014) );
  INVD1BWP12T U1435 ( .I(n1014), .ZN(n689) );
  AOI21D1BWP12T U1436 ( .A1(n1017), .A2(n1015), .B(n689), .ZN(n846) );
  NR2D1BWP12T U1437 ( .A1(n2275), .A2(a[14]), .ZN(n843) );
  ND2D1BWP12T U1438 ( .A1(n2275), .A2(a[14]), .ZN(n844) );
  TPOAI21D1BWP12T U1439 ( .A1(n846), .A2(n843), .B(n844), .ZN(n1432) );
  OR2XD1BWP12T U1440 ( .A1(n2626), .A2(n2276), .Z(n1430) );
  ND2D1BWP12T U1441 ( .A1(n2626), .A2(n2276), .ZN(n1429) );
  INVD1BWP12T U1442 ( .I(n1429), .ZN(n690) );
  AOI21D1BWP12T U1443 ( .A1(n1432), .A2(n1430), .B(n690), .ZN(n1392) );
  NR2D1BWP12T U1444 ( .A1(n2270), .A2(a[16]), .ZN(n1390) );
  ND2D1BWP12T U1445 ( .A1(n2270), .A2(a[16]), .ZN(n1391) );
  RCOAI21D1BWP12T U1446 ( .A1(n1392), .A2(n1390), .B(n1391), .ZN(n1596) );
  OR2XD1BWP12T U1447 ( .A1(n2679), .A2(n2678), .Z(n1595) );
  ND2D1BWP12T U1448 ( .A1(n2679), .A2(n2678), .ZN(n1594) );
  INVD1BWP12T U1449 ( .I(n1594), .ZN(n691) );
  AOI21D1BWP12T U1450 ( .A1(n1596), .A2(n1595), .B(n691), .ZN(n1648) );
  NR2D1BWP12T U1451 ( .A1(n2703), .A2(a[18]), .ZN(n1646) );
  ND2D1BWP12T U1452 ( .A1(n2703), .A2(a[18]), .ZN(n1647) );
  OAI21D1BWP12T U1453 ( .A1(n1648), .A2(n1646), .B(n1647), .ZN(n810) );
  OR2XD1BWP12T U1454 ( .A1(n2609), .A2(n782), .Z(n809) );
  ND2D1BWP12T U1455 ( .A1(n2609), .A2(n782), .ZN(n808) );
  INVD1BWP12T U1456 ( .I(n808), .ZN(n692) );
  AO21D1BWP12T U1457 ( .A1(n810), .A2(n809), .B(n692), .Z(n1593) );
  CKBD0BWP12T U1458 ( .I(result[31]), .Z(n) );
  INVD1BWP12T U1459 ( .I(n693), .ZN(n1734) );
  OAI21D1BWP12T U1460 ( .A1(n1734), .A2(n1730), .B(n1731), .ZN(n698) );
  INVD1BWP12T U1461 ( .I(n694), .ZN(n696) );
  ND2D1BWP12T U1462 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNR2XD1BWP12T U1463 ( .A1(n698), .A2(n697), .ZN(n1736) );
  INVD1BWP12T U1464 ( .I(n1736), .ZN(n733) );
  FA1D0BWP12T U1465 ( .A(a[25]), .B(n2269), .CI(n699), .CO(n2403), .S(n2458)
         );
  INVD1BWP12T U1466 ( .I(n1801), .ZN(n730) );
  HA1D1BWP12T U1467 ( .A(n1108), .B(n701), .CO(n1817), .S(n1840) );
  AOI22D0BWP12T U1468 ( .A1(n2173), .A2(n1513), .B1(n1512), .B2(n2170), .ZN(
        n703) );
  AOI22D0BWP12T U1469 ( .A1(n2166), .A2(n792), .B1(n985), .B2(n2169), .ZN(n702) );
  ND2D1BWP12T U1470 ( .A1(n703), .A2(n702), .ZN(n2199) );
  AOI22D0BWP12T U1471 ( .A1(n1511), .A2(n2169), .B1(n2166), .B2(n2143), .ZN(
        n705) );
  AOI22D0BWP12T U1472 ( .A1(n2173), .A2(n2141), .B1(n2142), .B2(n2170), .ZN(
        n704) );
  AOI21D0BWP12T U1473 ( .A1(n705), .A2(n704), .B(n2202), .ZN(n706) );
  AO211D0BWP12T U1474 ( .A1(n2155), .A2(n2199), .B(n706), .C(n2174), .Z(n707)
         );
  AOI21D1BWP12T U1475 ( .A1(n2868), .A2(n2195), .B(n707), .ZN(n2192) );
  INVD1BWP12T U1476 ( .I(n2192), .ZN(n725) );
  CKND2D0BWP12T U1477 ( .A1(n1999), .A2(n2143), .ZN(n709) );
  AOI22D0BWP12T U1478 ( .A1(n2000), .A2(n1511), .B1(n2001), .B2(n2142), .ZN(
        n708) );
  OAI211D0BWP12T U1479 ( .A1(n1518), .A2(n1940), .B(n709), .C(n708), .ZN(n710)
         );
  INVD1BWP12T U1480 ( .I(n2025), .ZN(n2031) );
  AOI21D0BWP12T U1481 ( .A1(n710), .A2(n2031), .B(n2006), .ZN(n713) );
  INVD1BWP12T U1482 ( .I(n2023), .ZN(n2033) );
  INVD0BWP12T U1483 ( .I(n1513), .ZN(n1508) );
  INVD0BWP12T U1484 ( .I(n985), .ZN(n995) );
  AOI22D0BWP12T U1485 ( .A1(n2002), .A2(n1508), .B1(n995), .B2(n2000), .ZN(
        n2026) );
  TPND3D0BWP12T U1486 ( .A1(n2027), .A2(n2033), .A3(n2026), .ZN(n712) );
  OAI211D0BWP12T U1487 ( .A1(n1997), .A2(n714), .B(n713), .C(n712), .ZN(n716)
         );
  ND2XD0BWP12T U1488 ( .A1(n1570), .A2(n471), .ZN(n1860) );
  OAI211D0BWP12T U1489 ( .A1(n471), .A2(n1863), .B(n1860), .C(n2769), .ZN(n715) );
  CKND2D1BWP12T U1490 ( .A1(n716), .A2(n715), .ZN(n1953) );
  ND2D1BWP12T U1491 ( .A1(n1953), .A2(n2894), .ZN(n724) );
  ND2D1BWP12T U1492 ( .A1(n2135), .A2(a[31]), .ZN(n2094) );
  INVD1BWP12T U1493 ( .I(n2094), .ZN(n2783) );
  INVD1BWP12T U1494 ( .I(n2099), .ZN(n2079) );
  NR2D1BWP12T U1495 ( .A1(n2783), .A2(n2079), .ZN(n2956) );
  INVD1BWP12T U1496 ( .I(n2068), .ZN(n2084) );
  NR2D1BWP12T U1497 ( .A1(n2084), .A2(n2058), .ZN(n2095) );
  NR2D1BWP12T U1498 ( .A1(n2095), .A2(n2957), .ZN(n2781) );
  CKND0BWP12T U1499 ( .I(b[25]), .ZN(n2269) );
  TPNR2D0BWP12T U1500 ( .A1(n2269), .A2(n2951), .ZN(n717) );
  RCAOI211D0BWP12T U1501 ( .A1(n2269), .A2(n2948), .B(n717), .C(n2825), .ZN(
        n721) );
  CKND2D0BWP12T U1502 ( .A1(n2775), .A2(n1855), .ZN(n720) );
  OAI21D0BWP12T U1503 ( .A1(a[25]), .A2(n2944), .B(n2949), .ZN(n718) );
  AOI22D0BWP12T U1504 ( .A1(n2947), .A2(n2253), .B1(n718), .B2(b[25]), .ZN(
        n719) );
  OAI211D0BWP12T U1505 ( .A1(n721), .A2(n2253), .B(n720), .C(n719), .ZN(n722)
         );
  AOI21D1BWP12T U1506 ( .A1(n2101), .A2(n2781), .B(n722), .ZN(n723) );
  OAI211D1BWP12T U1507 ( .A1(n725), .A2(n2942), .B(n724), .C(n723), .ZN(n726)
         );
  AOI21D1BWP12T U1508 ( .A1(n1840), .A2(n2940), .B(n726), .ZN(n729) );
  FA1D2BWP12T U1509 ( .A(a[25]), .B(b[25]), .CI(n727), .CO(n2332), .S(n2391)
         );
  ND2D1BWP12T U1510 ( .A1(n2391), .A2(n2967), .ZN(n728) );
  OAI211D1BWP12T U1511 ( .A1(n2814), .A2(n730), .B(n729), .C(n728), .ZN(n731)
         );
  INVD1BWP12T U1512 ( .I(n2855), .ZN(n2657) );
  INVD1BWP12T U1513 ( .I(n735), .ZN(n1670) );
  INVD1BWP12T U1514 ( .I(n1735), .ZN(n772) );
  FA1D1BWP12T U1515 ( .A(n737), .B(a[22]), .CI(n736), .CO(n2405), .S(n2457) );
  HA1D0BWP12T U1516 ( .A(n2232), .B(n739), .CO(n1819), .S(n1839) );
  MUX2NXD0BWP12T U1517 ( .I0(n2303), .I1(n2482), .S(n2231), .ZN(n1413) );
  MUX2D1BWP12T U1518 ( .I0(n2871), .I1(n2830), .S(n2231), .Z(n2117) );
  CKND2D1BWP12T U1519 ( .A1(n750), .A2(n2302), .ZN(n899) );
  INVD1BWP12T U1520 ( .I(n899), .ZN(n763) );
  AOI22D0BWP12T U1521 ( .A1(n2001), .A2(n2117), .B1(n1400), .B2(n763), .ZN(
        n741) );
  MUX2D1BWP12T U1522 ( .I0(n2574), .I1(n2620), .S(n2231), .Z(n2118) );
  ND2D1BWP12T U1523 ( .A1(n2002), .A2(n2118), .ZN(n740) );
  OAI211D1BWP12T U1524 ( .A1(n1413), .A2(n1959), .B(n741), .C(n740), .ZN(n2573) );
  INVD1BWP12T U1525 ( .I(n2022), .ZN(n2035) );
  CKMUX2D1BWP12T U1526 ( .I0(n2308), .I1(n2594), .S(n2231), .Z(n2125) );
  MUX2NXD0BWP12T U1527 ( .I0(a[8]), .I1(n2527), .S(n2231), .ZN(n1944) );
  INVD1BWP12T U1528 ( .I(n1944), .ZN(n2120) );
  AOI22D0BWP12T U1529 ( .A1(n2001), .A2(n2125), .B1(n2000), .B2(n2120), .ZN(
        n743) );
  MUX2NXD0BWP12T U1530 ( .I0(a[14]), .I1(n2643), .S(n2231), .ZN(n1466) );
  INVD1BWP12T U1531 ( .I(n1466), .ZN(n2124) );
  TPND2D0BWP12T U1532 ( .A1(n2002), .A2(n2124), .ZN(n742) );
  CKND2D1BWP12T U1533 ( .A1(n743), .A2(n742), .ZN(n745) );
  CKMUX2D1BWP12T U1534 ( .I0(n2900), .I1(n2301), .S(n2231), .Z(n2121) );
  INVD1BWP12T U1535 ( .I(n2121), .ZN(n1408) );
  TPNR2D0BWP12T U1536 ( .A1(n1959), .A2(n1408), .ZN(n744) );
  NR2D1BWP12T U1537 ( .A1(n745), .A2(n744), .ZN(n1356) );
  INVD0BWP12T U1538 ( .I(n1356), .ZN(n749) );
  MUX2XD0BWP12T U1539 ( .I0(a[22]), .I1(n2725), .S(n2231), .Z(n1471) );
  MUX2D0BWP12T U1540 ( .I0(a[16]), .I1(n2626), .S(n2231), .Z(n1460) );
  INVD1BWP12T U1541 ( .I(n1460), .ZN(n2127) );
  MUX2NXD0BWP12T U1542 ( .I0(a[20]), .I1(n2609), .S(n2231), .ZN(n2168) );
  OAI22D1BWP12T U1543 ( .A1(n1941), .A2(n2127), .B1(n1501), .B2(n2168), .ZN(
        n747) );
  MUX2NXD0BWP12T U1544 ( .I0(a[18]), .I1(n2679), .S(n2231), .ZN(n2149) );
  TPNR2D0BWP12T U1545 ( .A1(n1959), .A2(n2149), .ZN(n746) );
  AOI211D1BWP12T U1546 ( .A1(n1471), .A2(n2002), .B(n747), .C(n746), .ZN(n1355) );
  INVD1BWP12T U1547 ( .I(n1355), .ZN(n748) );
  AOI222D1BWP12T U1548 ( .A1(n2573), .A2(n2035), .B1(n749), .B2(n2033), .C1(
        n748), .C2(n2031), .ZN(n2038) );
  OAI22D1BWP12T U1549 ( .A1(n1870), .A2(n2251), .B1(n1871), .B2(n2310), .ZN(
        n876) );
  INVD1BWP12T U1550 ( .I(n876), .ZN(n1849) );
  AOI22D1BWP12T U1551 ( .A1(n2747), .A2(n751), .B1(n750), .B2(a[24]), .ZN(n755) );
  INR2XD0BWP12T U1552 ( .A1(a[22]), .B1(n1870), .ZN(n753) );
  NR2XD0BWP12T U1553 ( .A1(n1869), .A2(n2253), .ZN(n752) );
  NR2D1BWP12T U1554 ( .A1(n753), .A2(n752), .ZN(n754) );
  ND2D1BWP12T U1555 ( .A1(n755), .A2(n754), .ZN(n854) );
  INVD1BWP12T U1556 ( .I(n2052), .ZN(n1920) );
  MUX2D1BWP12T U1557 ( .I0(a[26]), .I1(a[27]), .S(n2231), .Z(n933) );
  NR2D1BWP12T U1558 ( .A1(n1872), .A2(a[28]), .ZN(n757) );
  NR2D0BWP12T U1559 ( .A1(n1869), .A2(a[29]), .ZN(n756) );
  NR2D1BWP12T U1560 ( .A1(n757), .A2(n756), .ZN(n758) );
  TPOAI21D0BWP12T U1561 ( .A1(n2477), .A2(n933), .B(n758), .ZN(n870) );
  INVD1BWP12T U1562 ( .I(n870), .ZN(n2097) );
  INVD1BWP12T U1563 ( .I(n1926), .ZN(n2049) );
  AOI22D1BWP12T U1564 ( .A1(n854), .A2(n1920), .B1(n2097), .B2(n2049), .ZN(
        n766) );
  INVD1BWP12T U1565 ( .I(n2076), .ZN(n2065) );
  NR2D1BWP12T U1566 ( .A1(n2068), .A2(n2957), .ZN(n1373) );
  INVD1BWP12T U1567 ( .I(n1373), .ZN(n2718) );
  AOI22D0BWP12T U1568 ( .A1(n2173), .A2(n1466), .B1(n1408), .B2(n2166), .ZN(
        n760) );
  INVD1BWP12T U1569 ( .I(n2125), .ZN(n1956) );
  AOI22D0BWP12T U1570 ( .A1(n2170), .A2(n1956), .B1(n1944), .B2(n2169), .ZN(
        n759) );
  ND2D1BWP12T U1571 ( .A1(n760), .A2(n759), .ZN(n1363) );
  AOI22D0BWP12T U1572 ( .A1(n2170), .A2(n2168), .B1(n2149), .B2(n2166), .ZN(
        n762) );
  INVD1BWP12T U1573 ( .I(n1471), .ZN(n2167) );
  AOI22D0BWP12T U1574 ( .A1(n2173), .A2(n2167), .B1(n2127), .B2(n2169), .ZN(
        n761) );
  CKND2D1BWP12T U1575 ( .A1(n762), .A2(n761), .ZN(n1362) );
  INVD0BWP12T U1576 ( .I(n1362), .ZN(n764) );
  CKND2D1BWP12T U1577 ( .A1(n899), .A2(n1413), .ZN(n901) );
  OAI22D0BWP12T U1578 ( .A1(n764), .A2(n2202), .B1(n2581), .B2(n2870), .ZN(
        n765) );
  INVD1BWP12T U1579 ( .I(n2187), .ZN(n2204) );
  RCAOI211D0BWP12T U1580 ( .A1(n2831), .A2(n1363), .B(n765), .C(n2204), .ZN(
        n2196) );
  INVD1BWP12T U1581 ( .I(n2675), .ZN(n2932) );
  INVD1BWP12T U1582 ( .I(n1933), .ZN(n863) );
  NR2D1BWP12T U1583 ( .A1(n2094), .A2(n2957), .ZN(n2807) );
  FA1D2BWP12T U1584 ( .A(a[22]), .B(b[22]), .CI(n767), .CO(n2334), .S(n2389)
         );
  AOI21D1BWP12T U1585 ( .A1(n2866), .A2(n2457), .B(n768), .ZN(n771) );
  FA1D1BWP12T U1586 ( .A(n737), .B(a[22]), .CI(n769), .CO(n1592), .S(n1653) );
  ND2D1BWP12T U1587 ( .A1(n1653), .A2(n2855), .ZN(n770) );
  OAI211D2BWP12T U1588 ( .A1(n2822), .A2(n772), .B(n771), .C(n770), .ZN(
        result[22]) );
  INVD1P75BWP12T U1589 ( .I(n773), .ZN(n1721) );
  INVD1BWP12T U1590 ( .I(n774), .ZN(n1675) );
  INVD1BWP12T U1591 ( .I(n1674), .ZN(n775) );
  AOI21D1BWP12T U1592 ( .A1(n1721), .A2(n1675), .B(n775), .ZN(n780) );
  INVD0BWP12T U1593 ( .I(n776), .ZN(n778) );
  CKND2D1BWP12T U1594 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2XD1BWP12T U1595 ( .A1(n780), .A2(n779), .Z(n1726) );
  INVD1P75BWP12T U1596 ( .I(n1726), .ZN(n813) );
  FA1D0BWP12T U1597 ( .A(n2609), .B(n782), .CI(n781), .CO(n2409), .S(n2456) );
  CKND2D0BWP12T U1598 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNR2XD1BWP12T U1599 ( .A1(n787), .A2(n786), .ZN(n2387) );
  HA1D1BWP12T U1600 ( .A(n1223), .B(n788), .CO(n1828), .S(n1827) );
  AOI22D1BWP12T U1601 ( .A1(n1999), .A2(n789), .B1(n1945), .B2(n999), .ZN(n791) );
  TPAOI22D0BWP12T U1602 ( .A1(n2002), .A2(n985), .B1(n2000), .B2(n1001), .ZN(
        n790) );
  ND2D1BWP12T U1603 ( .A1(n791), .A2(n790), .ZN(n1948) );
  AOI22D1BWP12T U1604 ( .A1(n2002), .A2(n987), .B1(n1945), .B2(n1000), .ZN(
        n1973) );
  INVD1BWP12T U1605 ( .I(n1973), .ZN(n2829) );
  NR2D1BWP12T U1606 ( .A1(n2008), .A2(n2006), .ZN(n2014) );
  AOI22D1BWP12T U1607 ( .A1(n987), .A2(n2173), .B1(n1000), .B2(n2170), .ZN(
        n2138) );
  OAI31D0BWP12T U1608 ( .A1(n2831), .A2(n2138), .A3(n2174), .B(n2135), .ZN(
        n796) );
  AOI22D0BWP12T U1609 ( .A1(n1511), .A2(n2173), .B1(n2170), .B2(n1513), .ZN(
        n794) );
  AOI22D0BWP12T U1610 ( .A1(n2169), .A2(n792), .B1(n1512), .B2(n2166), .ZN(
        n793) );
  ND2D1BWP12T U1611 ( .A1(n794), .A2(n793), .ZN(n2147) );
  AOI22D0BWP12T U1612 ( .A1(n2155), .A2(n2139), .B1(n2147), .B2(n2769), .ZN(
        n795) );
  ND2D1BWP12T U1613 ( .A1(n796), .A2(n795), .ZN(n2190) );
  OAI22D0BWP12T U1614 ( .A1(n1870), .A2(n2234), .B1(n1869), .B2(n2232), .ZN(
        n798) );
  TPOAI22D0BWP12T U1615 ( .A1(n1872), .A2(n2233), .B1(n1871), .B2(n2929), .ZN(
        n797) );
  NR2D1BWP12T U1616 ( .A1(n798), .A2(n797), .ZN(n1881) );
  OAI22D0BWP12T U1617 ( .A1(n1870), .A2(n2751), .B1(n1869), .B2(n2779), .ZN(
        n800) );
  TPOAI22D0BWP12T U1618 ( .A1(n1872), .A2(n2253), .B1(n1871), .B2(n2946), .ZN(
        n799) );
  NR2D1BWP12T U1619 ( .A1(n800), .A2(n799), .ZN(n1882) );
  OAI22D0BWP12T U1620 ( .A1(n1870), .A2(n2252), .B1(n1869), .B2(n2251), .ZN(
        n802) );
  TPOAI22D0BWP12T U1621 ( .A1(n1872), .A2(n2248), .B1(n1871), .B2(n2249), .ZN(
        n801) );
  NR2D1BWP12T U1622 ( .A1(n802), .A2(n801), .ZN(n2051) );
  IOA21D0BWP12T U1623 ( .A1(n2639), .A2(n2310), .B(n803), .ZN(n804) );
  TPAOI21D0BWP12T U1624 ( .A1(n2051), .A2(n471), .B(n804), .ZN(n1854) );
  NR2D0BWP12T U1625 ( .A1(n1930), .A2(a[31]), .ZN(n805) );
  AOI211D1BWP12T U1626 ( .A1(n863), .A2(n2051), .B(n806), .C(n805), .ZN(n2091)
         );
  AOI21D1BWP12T U1627 ( .A1(n2866), .A2(n2456), .B(n807), .ZN(n812) );
  ND2D1BWP12T U1628 ( .A1(n1651), .A2(n2855), .ZN(n811) );
  OAI211D2BWP12T U1629 ( .A1(n2822), .A2(n813), .B(n812), .C(n811), .ZN(
        result[19]) );
  INVD1BWP12T U1630 ( .I(n814), .ZN(n1424) );
  INVD1BWP12T U1631 ( .I(n816), .ZN(n819) );
  TPND2D0BWP12T U1632 ( .A1(n819), .A2(n818), .ZN(n820) );
  XOR2XD1BWP12T U1633 ( .A1(n821), .A2(n820), .Z(n2385) );
  CKND0BWP12T U1634 ( .I(n2967), .ZN(n2909) );
  TPAOI21D0BWP12T U1635 ( .A1(n822), .A2(n2827), .B(n2079), .ZN(n2066) );
  CKND2D0BWP12T U1636 ( .A1(n854), .A2(n471), .ZN(n824) );
  CKND2D0BWP12T U1637 ( .A1(n2097), .A2(n2639), .ZN(n823) );
  AOI31D0BWP12T U1638 ( .A1(n824), .A2(n2870), .A3(n823), .B(n2769), .ZN(n832)
         );
  OAI22D1BWP12T U1639 ( .A1(n1870), .A2(n2705), .B1(n1869), .B2(n2233), .ZN(
        n828) );
  TPOAI22D0BWP12T U1640 ( .A1(n826), .A2(n2929), .B1(n825), .B2(n2234), .ZN(
        n827) );
  NR2D1BWP12T U1641 ( .A1(n828), .A2(n827), .ZN(n1931) );
  OAI22D0BWP12T U1642 ( .A1(n1870), .A2(n1441), .B1(n1869), .B2(n2683), .ZN(
        n830) );
  OAI22D0BWP12T U1643 ( .A1(n1872), .A2(n2235), .B1(n1871), .B2(n2240), .ZN(
        n829) );
  NR2D1BWP12T U1644 ( .A1(n830), .A2(n829), .ZN(n1934) );
  OAI22D0BWP12T U1645 ( .A1(n1931), .A2(n1926), .B1(n1934), .B2(n2052), .ZN(
        n831) );
  NR2D1BWP12T U1646 ( .A1(n832), .A2(n831), .ZN(n837) );
  INVD1BWP12T U1647 ( .I(n976), .ZN(n926) );
  NR2D1BWP12T U1648 ( .A1(n926), .A2(n835), .ZN(n1442) );
  XNR2XD1BWP12T U1649 ( .A1(n1442), .A2(a[14]), .ZN(n1837) );
  AOI21D0BWP12T U1650 ( .A1(n876), .A2(n1920), .B(n2870), .ZN(n836) );
  NR2D1BWP12T U1651 ( .A1(n837), .A2(n836), .ZN(n1885) );
  CKAN2D1BWP12T U1652 ( .A1(n2115), .A2(n2886), .Z(n1443) );
  NR2D0BWP12T U1653 ( .A1(n2573), .A2(n2017), .ZN(n838) );
  INVD1BWP12T U1654 ( .I(n1997), .ZN(n2508) );
  AOI211D0BWP12T U1655 ( .A1(n2017), .A2(n1356), .B(n838), .C(n2508), .ZN(n839) );
  NR2D1BWP12T U1656 ( .A1(n839), .A2(n1885), .ZN(n1994) );
  CKND2D0BWP12T U1657 ( .A1(n1363), .A2(n2827), .ZN(n840) );
  INVD1BWP12T U1658 ( .I(n2135), .ZN(n2198) );
  OAI211D0BWP12T U1659 ( .A1(n2581), .A2(n2827), .B(n840), .C(n2198), .ZN(
        n2208) );
  AOI211D1BWP12T U1660 ( .A1(n1791), .A2(n2858), .B(n842), .C(n841), .ZN(n851)
         );
  TPND2D0BWP12T U1661 ( .A1(n848), .A2(n844), .ZN(n845) );
  CKXOR2D1BWP12T U1662 ( .A1(n846), .A2(n845), .Z(n1644) );
  AOI22D1BWP12T U1663 ( .A1(n1644), .A2(n2855), .B1(n2866), .B2(n2455), .ZN(
        n850) );
  INVD1BWP12T U1664 ( .I(n1931), .ZN(n853) );
  INVD1BWP12T U1665 ( .I(n871), .ZN(n1919) );
  CKND2D1BWP12T U1666 ( .A1(n1919), .A2(n2827), .ZN(n1993) );
  TPOAI21D0BWP12T U1667 ( .A1(n1930), .A2(n2098), .B(n875), .ZN(n2069) );
  OAI21D0BWP12T U1668 ( .A1(n2069), .A2(n2174), .B(n2135), .ZN(n867) );
  OAI22D1BWP12T U1669 ( .A1(n1870), .A2(n2578), .B1(n1869), .B2(n2243), .ZN(
        n856) );
  OAI22D1BWP12T U1670 ( .A1(n1872), .A2(n2550), .B1(n1871), .B2(n2532), .ZN(
        n855) );
  NR2D1BWP12T U1671 ( .A1(n856), .A2(n855), .ZN(n1932) );
  NR2D1BWP12T U1672 ( .A1(n2128), .A2(n2231), .ZN(n1894) );
  AOI21D0BWP12T U1673 ( .A1(n1891), .A2(n1832), .B(n2831), .ZN(n857) );
  IOA21D0BWP12T U1674 ( .A1(n1894), .A2(n2869), .B(n857), .ZN(n860) );
  INR2D1BWP12T U1675 ( .A1(n2231), .B1(n2128), .ZN(n1893) );
  INVD1BWP12T U1676 ( .I(n1893), .ZN(n858) );
  OAI22D1BWP12T U1677 ( .A1(n858), .A2(n2620), .B1(n2830), .B2(n1548), .ZN(
        n859) );
  AOI211D1BWP12T U1678 ( .A1(n2639), .A2(n1932), .B(n860), .C(n859), .ZN(n866)
         );
  OAI22D0BWP12T U1679 ( .A1(n1870), .A2(n2900), .B1(n2643), .B2(n1869), .ZN(
        n862) );
  OAI22D0BWP12T U1680 ( .A1(n2308), .A2(n1872), .B1(n1871), .B2(n2594), .ZN(
        n861) );
  NR2D1BWP12T U1681 ( .A1(n862), .A2(n861), .ZN(n1929) );
  AOI21D1BWP12T U1682 ( .A1(n1929), .A2(n863), .B(n2868), .ZN(n864) );
  OAI21D1BWP12T U1683 ( .A1(n1934), .A2(n1930), .B(n864), .ZN(n865) );
  NR2D1BWP12T U1684 ( .A1(n866), .A2(n865), .ZN(n874) );
  INVD1BWP12T U1685 ( .I(n874), .ZN(n878) );
  AOI21D0BWP12T U1686 ( .A1(n867), .A2(n878), .B(n2058), .ZN(n2090) );
  CKND2D1BWP12T U1687 ( .A1(n1710), .A2(n2977), .ZN(n913) );
  OAI22D0BWP12T U1688 ( .A1(n871), .A2(n2159), .B1(n2080), .B2(n2770), .ZN(
        n873) );
  NR2D0BWP12T U1689 ( .A1(n1400), .A2(n899), .ZN(n872) );
  OA21D1BWP12T U1690 ( .A1(n2002), .A2(n872), .B(n901), .Z(n1946) );
  INVD1BWP12T U1691 ( .I(n1946), .ZN(n1992) );
  OAI22D1BWP12T U1692 ( .A1(n874), .A2(n873), .B1(n1992), .B2(n2025), .ZN(
        n1971) );
  OA21D1BWP12T U1693 ( .A1(n876), .A2(n1930), .B(n875), .Z(n2706) );
  INVD1BWP12T U1694 ( .I(n2706), .ZN(n877) );
  RCOAI21D0BWP12T U1695 ( .A1(n877), .A2(n2174), .B(n2135), .ZN(n879) );
  ND2D1BWP12T U1696 ( .A1(n879), .A2(n878), .ZN(n1937) );
  NR2D1BWP12T U1697 ( .A1(n1937), .A2(n2495), .ZN(n911) );
  INVD1BWP12T U1698 ( .I(n880), .ZN(n1604) );
  OAI21D0BWP12T U1699 ( .A1(n1604), .A2(n1601), .B(n1602), .ZN(n885) );
  CKND0BWP12T U1700 ( .I(n881), .ZN(n883) );
  ND2XD0BWP12T U1701 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNR2XD1BWP12T U1702 ( .A1(n885), .A2(n884), .ZN(n1606) );
  INVD1BWP12T U1703 ( .I(n1606), .ZN(n909) );
  INVD1BWP12T U1704 ( .I(n886), .ZN(n1756) );
  OAI21D0BWP12T U1705 ( .A1(n1756), .A2(n1754), .B(n1755), .ZN(n890) );
  CKND2D0BWP12T U1706 ( .A1(n893), .A2(n888), .ZN(n889) );
  XNR2XD1BWP12T U1707 ( .A1(n890), .A2(n889), .ZN(n1759) );
  NR2D0BWP12T U1708 ( .A1(n471), .A2(n2951), .ZN(n891) );
  AOI211D0BWP12T U1709 ( .A1(n471), .A2(n2948), .B(n891), .C(n2825), .ZN(n898)
         );
  INVD1BWP12T U1710 ( .I(n892), .ZN(n2361) );
  INVD0BWP12T U1711 ( .I(n2360), .ZN(n893) );
  CKND2D1BWP12T U1712 ( .A1(n893), .A2(n2359), .ZN(n894) );
  XOR2XD1BWP12T U1713 ( .A1(n2361), .A2(n894), .Z(n2357) );
  CKND2D0BWP12T U1714 ( .A1(n2357), .A2(n2967), .ZN(n897) );
  OAI21D0BWP12T U1715 ( .A1(n2303), .A2(n2944), .B(n2949), .ZN(n895) );
  AOI22D0BWP12T U1716 ( .A1(n2947), .A2(n1832), .B1(n895), .B2(n2639), .ZN(
        n896) );
  OAI211D1BWP12T U1717 ( .A1(n898), .A2(n1832), .B(n897), .C(n896), .ZN(n903)
         );
  ND2D1BWP12T U1718 ( .A1(n2513), .A2(n2827), .ZN(n2535) );
  OAI21D0BWP12T U1719 ( .A1(n899), .A2(n2639), .B(n2126), .ZN(n900) );
  CKND2D1BWP12T U1720 ( .A1(n901), .A2(n900), .ZN(n2164) );
  NR2XD0BWP12T U1721 ( .A1(n2535), .A2(n2164), .ZN(n902) );
  AOI211D1BWP12T U1722 ( .A1(n1759), .A2(n2858), .B(n903), .C(n902), .ZN(n908)
         );
  INVD1BWP12T U1723 ( .I(n904), .ZN(n2428) );
  CKND2D1BWP12T U1724 ( .A1(n883), .A2(n2426), .ZN(n905) );
  XOR2D1BWP12T U1725 ( .A1(n2428), .A2(n905), .Z(n2424) );
  INVD0BWP12T U1726 ( .I(n906), .ZN(n1833) );
  XNR2XD0BWP12T U1727 ( .A1(n1833), .A2(n2303), .ZN(n1834) );
  AOI22D0BWP12T U1728 ( .A1(n2424), .A2(n2866), .B1(n1834), .B2(n2940), .ZN(
        n907) );
  OAI211D1BWP12T U1729 ( .A1(n2657), .A2(n909), .B(n908), .C(n907), .ZN(n910)
         );
  AOI211D1BWP12T U1730 ( .A1(n2894), .A2(n1971), .B(n911), .C(n910), .ZN(n912)
         );
  OAI211D1BWP12T U1731 ( .A1(n2090), .A2(n2957), .B(n913), .C(n912), .ZN(
        result[2]) );
  INVD1BWP12T U1732 ( .I(n914), .ZN(n1686) );
  AOI21D1BWP12T U1733 ( .A1(n1686), .A2(n1685), .B(n915), .ZN(n919) );
  ND2D1BWP12T U1734 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2XD1BWP12T U1735 ( .A1(n919), .A2(n918), .Z(n1714) );
  INVD1BWP12T U1736 ( .I(n1600), .ZN(n949) );
  XOR2XD1BWP12T U1737 ( .A1(n926), .A2(n2308), .Z(n1821) );
  CKND0BWP12T U1738 ( .I(n2117), .ZN(n928) );
  INR2D1BWP12T U1739 ( .A1(n2302), .B1(n1870), .ZN(n1547) );
  CKND0BWP12T U1740 ( .I(n1547), .ZN(n927) );
  OAI222D1BWP12T U1741 ( .A1(n928), .A2(n1940), .B1(n927), .B2(n1891), .C1(
        n1413), .C2(n1501), .ZN(n2036) );
  INVD1BWP12T U1742 ( .I(n2036), .ZN(n1970) );
  TPND2D0BWP12T U1743 ( .A1(n1999), .A2(n2120), .ZN(n931) );
  AOI22D0BWP12T U1744 ( .A1(n2001), .A2(n2121), .B1(n2000), .B2(n2118), .ZN(
        n930) );
  TPND2D0BWP12T U1745 ( .A1(n2002), .A2(n2125), .ZN(n929) );
  ND3D1BWP12T U1746 ( .A1(n931), .A2(n930), .A3(n929), .ZN(n2034) );
  TPOAI22D0BWP12T U1747 ( .A1(n1870), .A2(n2946), .B1(n1871), .B2(n2253), .ZN(
        n932) );
  AOI21D1BWP12T U1748 ( .A1(n2477), .A2(n933), .B(n932), .ZN(n1848) );
  INVD0BWP12T U1749 ( .I(n1848), .ZN(n934) );
  TPOAI22D0BWP12T U1750 ( .A1(n1870), .A2(n2929), .B1(n1872), .B2(n2232), .ZN(
        n936) );
  TPOAI22D0BWP12T U1751 ( .A1(n1871), .A2(n2233), .B1(n1869), .B2(n2751), .ZN(
        n935) );
  NR2D1BWP12T U1752 ( .A1(n936), .A2(n935), .ZN(n1903) );
  OAI22D0BWP12T U1753 ( .A1(n1870), .A2(n2235), .B1(n1871), .B2(n2683), .ZN(
        n938) );
  OAI22D0BWP12T U1754 ( .A1(n1872), .A2(n2705), .B1(n1869), .B2(n2234), .ZN(
        n937) );
  NR2D1BWP12T U1755 ( .A1(n938), .A2(n937), .ZN(n1912) );
  TPNR2D0BWP12T U1756 ( .A1(n1912), .A2(n1926), .ZN(n942) );
  OAI22D0BWP12T U1757 ( .A1(n1870), .A2(n2242), .B1(n1869), .B2(n2240), .ZN(
        n940) );
  OAI22D0BWP12T U1758 ( .A1(n1872), .A2(n1441), .B1(n1871), .B2(n2241), .ZN(
        n939) );
  NR2D1BWP12T U1759 ( .A1(n940), .A2(n939), .ZN(n1914) );
  OAI21D0BWP12T U1760 ( .A1(n1914), .A2(n2052), .B(n2870), .ZN(n941) );
  AOI211D1BWP12T U1761 ( .A1(n1858), .A2(n2831), .B(n942), .C(n941), .ZN(n951)
         );
  OAI22D0BWP12T U1762 ( .A1(n1870), .A2(n2249), .B1(n1869), .B2(n2310), .ZN(
        n944) );
  TPOAI22D0BWP12T U1763 ( .A1(n2251), .A2(n1872), .B1(n1871), .B2(n2248), .ZN(
        n943) );
  NR2D1BWP12T U1764 ( .A1(n944), .A2(n943), .ZN(n1856) );
  NR2D1BWP12T U1765 ( .A1(n1856), .A2(n2052), .ZN(n950) );
  MAOI22D0BWP12T U1766 ( .A1(n1821), .A2(n2940), .B1(n1982), .B2(n2964), .ZN(
        n948) );
  INVD1BWP12T U1767 ( .I(n945), .ZN(n954) );
  ND2D1BWP12T U1768 ( .A1(n1789), .A2(n2858), .ZN(n947) );
  OAI211D1BWP12T U1769 ( .A1(n2657), .A2(n949), .B(n948), .C(n947), .ZN(n967)
         );
  AOI21D0BWP12T U1770 ( .A1(a[31]), .A2(n2052), .B(n950), .ZN(n1479) );
  AOI211D1BWP12T U1771 ( .A1(n2868), .A2(n1479), .B(n951), .C(n2174), .ZN(n952) );
  NR2D0BWP12T U1772 ( .A1(n952), .A2(n2058), .ZN(n2060) );
  CKND2D1BWP12T U1773 ( .A1(n2380), .A2(n2967), .ZN(n965) );
  TPNR2D0BWP12T U1774 ( .A1(n2277), .A2(n2951), .ZN(n956) );
  RCAOI211D0BWP12T U1775 ( .A1(n2277), .A2(n2948), .B(n956), .C(n2825), .ZN(
        n962) );
  OAI22D0BWP12T U1776 ( .A1(n2118), .A2(n2116), .B1(n2125), .B2(n2126), .ZN(
        n958) );
  OAI22D0BWP12T U1777 ( .A1(n2119), .A2(n2120), .B1(n2121), .B2(n2128), .ZN(
        n957) );
  NR2D1BWP12T U1778 ( .A1(n958), .A2(n957), .ZN(n2180) );
  ND2D1BWP12T U1779 ( .A1(n2209), .A2(n2786), .ZN(n961) );
  OAI21D0BWP12T U1780 ( .A1(n2308), .A2(n2944), .B(n2949), .ZN(n959) );
  AOI22D0BWP12T U1781 ( .A1(n2947), .A2(n2242), .B1(n959), .B2(n2598), .ZN(
        n960) );
  OAI211D1BWP12T U1782 ( .A1(n962), .A2(n2242), .B(n961), .C(n960), .ZN(n963)
         );
  AOI21D1BWP12T U1783 ( .A1(n1902), .A2(n1443), .B(n963), .ZN(n964) );
  OAI211D1BWP12T U1784 ( .A1(n2060), .A2(n2957), .B(n965), .C(n964), .ZN(n966)
         );
  AOI211D1BWP12T U1785 ( .A1(n2866), .A2(n2417), .B(n967), .C(n966), .ZN(n968)
         );
  IOA21D1BWP12T U1786 ( .A1(n1714), .A2(n2977), .B(n968), .ZN(result[12]) );
  CKND2D1BWP12T U1787 ( .A1(n1716), .A2(n2977), .ZN(n1021) );
  CKND2D0BWP12T U1788 ( .A1(n1015), .A2(n973), .ZN(n974) );
  XOR2XD1BWP12T U1789 ( .A1(n975), .A2(n974), .Z(n2418) );
  CKND2D0BWP12T U1790 ( .A1(n1863), .A2(n1920), .ZN(n980) );
  OAI22D0BWP12T U1791 ( .A1(n1570), .A2(n1930), .B1(n1862), .B2(n1926), .ZN(
        n979) );
  OAI21D0BWP12T U1792 ( .A1(n1861), .A2(n1933), .B(n2870), .ZN(n978) );
  NR2D0BWP12T U1793 ( .A1(n1890), .A2(n2052), .ZN(n977) );
  NR3D1BWP12T U1794 ( .A1(n979), .A2(n978), .A3(n977), .ZN(n1006) );
  AOI21D1BWP12T U1795 ( .A1(n2868), .A2(n980), .B(n1006), .ZN(n1901) );
  NR2D0BWP12T U1796 ( .A1(n2278), .A2(n2951), .ZN(n981) );
  AOI211D0BWP12T U1797 ( .A1(n2278), .A2(n2948), .B(n981), .C(n2825), .ZN(n991) );
  OAI22D0BWP12T U1798 ( .A1(n982), .A2(n2119), .B1(n994), .B2(n2116), .ZN(n984) );
  NR2D0BWP12T U1799 ( .A1(n996), .A2(n2126), .ZN(n983) );
  AOI211D1BWP12T U1800 ( .A1(n2170), .A2(n985), .B(n984), .C(n983), .ZN(n2189)
         );
  CKND2D1BWP12T U1801 ( .A1(n2210), .A2(n2786), .ZN(n990) );
  OAI21D0BWP12T U1802 ( .A1(n2643), .A2(n2944), .B(n2949), .ZN(n988) );
  AOI22D0BWP12T U1803 ( .A1(n2947), .A2(n2241), .B1(n988), .B2(b[13]), .ZN(
        n989) );
  OAI211D0BWP12T U1804 ( .A1(n991), .A2(n2241), .B(n990), .C(n989), .ZN(n992)
         );
  RCAOI21D0BWP12T U1805 ( .A1(n1901), .A2(n1443), .B(n992), .ZN(n993) );
  IOA21D1BWP12T U1806 ( .A1(n2940), .A2(n1836), .B(n993), .ZN(n1009) );
  AOI22D0BWP12T U1807 ( .A1(n995), .A2(n2001), .B1(n2000), .B2(n994), .ZN(n998) );
  TPND2D0BWP12T U1808 ( .A1(n2002), .A2(n996), .ZN(n997) );
  OAI211D0BWP12T U1809 ( .A1(n999), .A2(n1959), .B(n998), .C(n997), .ZN(n2016)
         );
  INVD1BWP12T U1810 ( .I(n2016), .ZN(n1505) );
  CKND0BWP12T U1811 ( .I(n1000), .ZN(n1002) );
  OAI222D1BWP12T U1812 ( .A1(n1003), .A2(n1501), .B1(n1002), .B2(n1959), .C1(
        n1001), .C2(n1940), .ZN(n1947) );
  INVD1BWP12T U1813 ( .I(n1947), .ZN(n2012) );
  OAI22D0BWP12T U1814 ( .A1(n1004), .A2(n2639), .B1(n2173), .B2(n2310), .ZN(
        n1571) );
  CKND2D0BWP12T U1815 ( .A1(n1571), .A2(n2827), .ZN(n1524) );
  AOI21D0BWP12T U1816 ( .A1(n1524), .A2(n2099), .B(n2174), .ZN(n1005) );
  NR2D0BWP12T U1817 ( .A1(n1005), .A2(n2198), .ZN(n1007) );
  INVD1BWP12T U1818 ( .I(n2058), .ZN(n2105) );
  TPOAI21D0BWP12T U1819 ( .A1(n1007), .A2(n1006), .B(n2105), .ZN(n2104) );
  MOAI22D0BWP12T U1820 ( .A1(n1995), .A2(n2964), .B1(n2905), .B2(n2104), .ZN(
        n1008) );
  RCAOI211D0BWP12T U1821 ( .A1(n2418), .A2(n2866), .B(n1009), .C(n1008), .ZN(
        n1020) );
  AOI22D1BWP12T U1822 ( .A1(n2858), .A2(n1792), .B1(n2381), .B2(n2967), .ZN(
        n1019) );
  CKND2D1BWP12T U1823 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNR2D1BWP12T U1824 ( .A1(n1017), .A2(n1016), .ZN(n1645) );
  CKND2D1BWP12T U1825 ( .A1(n1645), .A2(n2855), .ZN(n1018) );
  ND4D1BWP12T U1826 ( .A1(n1021), .A2(n1020), .A3(n1019), .A4(n1018), .ZN(
        result[13]) );
  INVD15BWP12T U1827 ( .I(n1119), .ZN(n2633) );
  XNR2XD8BWP12T U1828 ( .A1(a[8]), .A2(n2633), .ZN(n1022) );
  BUFFXD12BWP12T U1829 ( .I(n1022), .Z(n2614) );
  INVD15BWP12T U1830 ( .I(n1049), .ZN(n2613) );
  XOR2D2BWP12T U1831 ( .A1(a[8]), .A2(n2613), .Z(n1023) );
  ND2D4BWP12T U1832 ( .A1(n2614), .A2(n1023), .ZN(n2616) );
  XNR2D0BWP12T U1833 ( .A1(n2613), .A2(b[22]), .ZN(n1024) );
  XNR2D0BWP12T U1834 ( .A1(n2613), .A2(b[23]), .ZN(n2615) );
  OAI22D0BWP12T U1835 ( .A1(n2616), .A2(n1024), .B1(n2614), .B2(n2615), .ZN(
        mult_x_18_n873) );
  XNR2D0BWP12T U1836 ( .A1(n2613), .A2(b[21]), .ZN(n1280) );
  TPOAI22D0BWP12T U1837 ( .A1(n2616), .A2(n1280), .B1(n2614), .B2(n1024), .ZN(
        mult_x_18_n874) );
  XOR2D1BWP12T U1838 ( .A1(n2633), .A2(n2574), .Z(n1026) );
  TPND2D8BWP12T U1839 ( .A1(n1025), .A2(n1026), .ZN(n2635) );
  XNR2D1BWP12T U1840 ( .A1(n2633), .A2(b[5]), .ZN(n1139) );
  XNR2D1BWP12T U1841 ( .A1(n2633), .A2(b[6]), .ZN(n1203) );
  OAI22D1BWP12T U1842 ( .A1(n2635), .A2(n1139), .B1(n1025), .B2(n1203), .ZN(
        mult_x_18_n917) );
  XOR2D1BWP12T U1843 ( .A1(n2594), .A2(n2900), .Z(n1027) );
  XNR2XD4BWP12T U1844 ( .A1(n2613), .A2(n2900), .ZN(n2595) );
  TPND2D8BWP12T U1845 ( .A1(n1027), .A2(n2595), .ZN(n2597) );
  XNR2D0BWP12T U1846 ( .A1(n2594), .A2(b[19]), .ZN(n1253) );
  XNR2D0BWP12T U1847 ( .A1(n2594), .A2(b[20]), .ZN(n1029) );
  OAI22D0BWP12T U1848 ( .A1(n2597), .A2(n1253), .B1(n1029), .B2(n2595), .ZN(
        mult_x_18_n851) );
  XNR2D1BWP12T U1849 ( .A1(n2594), .A2(n2477), .ZN(n1160) );
  XNR2D1BWP12T U1850 ( .A1(n2594), .A2(n2639), .ZN(n1327) );
  OAI22D1BWP12T U1851 ( .A1(n2597), .A2(n1160), .B1(n1327), .B2(n2595), .ZN(
        mult_x_18_n869) );
  XNR2D0BWP12T U1852 ( .A1(n2633), .A2(b[23]), .ZN(n1268) );
  XNR2D0BWP12T U1853 ( .A1(n2633), .A2(b[24]), .ZN(n1028) );
  TPOAI22D0BWP12T U1854 ( .A1(n2635), .A2(n1268), .B1(n1025), .B2(n1028), .ZN(
        mult_x_18_n899) );
  XNR2D0BWP12T U1855 ( .A1(n2633), .A2(b[25]), .ZN(n2634) );
  OAI22D0BWP12T U1856 ( .A1(n2635), .A2(n1028), .B1(n1025), .B2(n2634), .ZN(
        mult_x_18_n898) );
  XNR2D0BWP12T U1857 ( .A1(n2594), .A2(b[21]), .ZN(n2596) );
  OAI22D0BWP12T U1858 ( .A1(n2597), .A2(n1029), .B1(n2596), .B2(n2595), .ZN(
        mult_x_18_n850) );
  XNR2D0BWP12T U1859 ( .A1(n2482), .A2(b[26]), .ZN(n1183) );
  XNR2D0BWP12T U1860 ( .A1(n2482), .A2(b[27]), .ZN(n1086) );
  XNR2D1BWP12T U1861 ( .A1(n2679), .A2(n2897), .ZN(n1180) );
  XNR2XD1BWP12T U1862 ( .A1(n2679), .A2(b[11]), .ZN(n1251) );
  XNR2D0BWP12T U1863 ( .A1(n2482), .A2(b[28]), .ZN(n1085) );
  XNR2XD1BWP12T U1864 ( .A1(a[28]), .A2(a[27]), .ZN(n2636) );
  XNR2XD0BWP12T U1865 ( .A1(n2626), .A2(b[13]), .ZN(n1275) );
  TPOAI22D0BWP12T U1866 ( .A1(n2629), .A2(n1275), .B1(n2627), .B2(n1031), .ZN(
        mult_x_18_n813) );
  XNR2XD0BWP12T U1867 ( .A1(n2626), .A2(b[16]), .ZN(n1033) );
  TPOAI22D0BWP12T U1868 ( .A1(n2629), .A2(n1032), .B1(n2627), .B2(n1033), .ZN(
        mult_x_18_n811) );
  XNR2XD1BWP12T U1869 ( .A1(n2620), .A2(b[25]), .ZN(n1269) );
  XNR2D0BWP12T U1870 ( .A1(n2620), .A2(b[26]), .ZN(n1034) );
  OAI22D0BWP12T U1871 ( .A1(n2623), .A2(n1269), .B1(n1034), .B2(n2621), .ZN(
        mult_x_18_n926) );
  XNR2D0BWP12T U1872 ( .A1(n2830), .A2(b[27]), .ZN(n1092) );
  XNR2D0BWP12T U1873 ( .A1(n2830), .A2(b[28]), .ZN(n1036) );
  TPOAI22D0BWP12T U1874 ( .A1(n2652), .A2(n1092), .B1(n2650), .B2(n1036), .ZN(
        mult_x_18_n955) );
  XNR2XD0BWP12T U1875 ( .A1(n2626), .A2(b[17]), .ZN(n2628) );
  OAI22D0BWP12T U1876 ( .A1(n2629), .A2(n1033), .B1(n2627), .B2(n2628), .ZN(
        mult_x_18_n810) );
  XNR2D0BWP12T U1877 ( .A1(n2620), .A2(b[27]), .ZN(n2622) );
  OAI22D0BWP12T U1878 ( .A1(n2623), .A2(n1034), .B1(n2622), .B2(n2621), .ZN(
        mult_x_18_n925) );
  XNR2XD0BWP12T U1879 ( .A1(n2609), .A2(b[13]), .ZN(n2611) );
  OAI22D0BWP12T U1880 ( .A1(n2612), .A2(n1035), .B1(n2610), .B2(n2611), .ZN(
        mult_x_18_n778) );
  XNR2D1BWP12T U1881 ( .A1(n2620), .A2(n2897), .ZN(n1244) );
  XNR2D1BWP12T U1882 ( .A1(n2620), .A2(b[11]), .ZN(n1114) );
  TPOAI22D1BWP12T U1883 ( .A1(n2623), .A2(n1244), .B1(n1114), .B2(n2621), .ZN(
        mult_x_18_n941) );
  XNR2D0BWP12T U1884 ( .A1(n2830), .A2(b[29]), .ZN(n2651) );
  OAI22D0BWP12T U1885 ( .A1(n2652), .A2(n1036), .B1(n2650), .B2(n2651), .ZN(
        mult_x_18_n954) );
  XNR2XD0BWP12T U1886 ( .A1(n2482), .A2(b[31]), .ZN(n2602) );
  XNR2D0BWP12T U1887 ( .A1(a[29]), .A2(a[30]), .ZN(n2640) );
  XNR2XD1BWP12T U1888 ( .A1(n2830), .A2(b[25]), .ZN(n1235) );
  XNR2XD1BWP12T U1889 ( .A1(n2830), .A2(b[26]), .ZN(n1093) );
  TPOAI22D0BWP12T U1890 ( .A1(n2652), .A2(n1235), .B1(n2650), .B2(n1093), .ZN(
        mult_x_18_n957) );
  XNR2D2BWP12T U1891 ( .A1(a[20]), .A2(n2609), .ZN(n2599) );
  CKXOR2D1BWP12T U1892 ( .A1(a[20]), .A2(n2725), .Z(n1038) );
  CKND2D3BWP12T U1893 ( .A1(n2599), .A2(n1038), .ZN(n2601) );
  XNR2XD1BWP12T U1894 ( .A1(n2725), .A2(n2897), .ZN(n1039) );
  XNR2XD0BWP12T U1895 ( .A1(n2725), .A2(b[11]), .ZN(n2600) );
  OAI22D0BWP12T U1896 ( .A1(n2601), .A2(n1039), .B1(n2599), .B2(n2600), .ZN(
        mult_x_18_n765) );
  XNR2XD1BWP12T U1897 ( .A1(n2725), .A2(b[9]), .ZN(n1256) );
  TPOAI22D0BWP12T U1898 ( .A1(n2601), .A2(n1256), .B1(n2599), .B2(n1039), .ZN(
        mult_x_18_n766) );
  XNR2XD1BWP12T U1899 ( .A1(a[29]), .A2(n2639), .ZN(n1233) );
  XNR2D0BWP12T U1900 ( .A1(a[29]), .A2(n2831), .ZN(n2637) );
  OAI22D0BWP12T U1901 ( .A1(n2638), .A2(n1233), .B1(n2637), .B2(n2636), .ZN(
        mult_x_18_n733) );
  XNR2D2BWP12T U1902 ( .A1(n2747), .A2(a[24]), .ZN(n2606) );
  XOR2XD1BWP12T U1903 ( .A1(a[25]), .A2(a[24]), .Z(n1040) );
  ND2D1BWP12T U1904 ( .A1(n2606), .A2(n1040), .ZN(n2608) );
  XNR2D0BWP12T U1905 ( .A1(a[25]), .A2(n2528), .ZN(n2607) );
  OAI22D0BWP12T U1906 ( .A1(n2608), .A2(n1043), .B1(n2606), .B2(n2607), .ZN(
        mult_x_18_n745) );
  XNR2D1BWP12T U1907 ( .A1(a[26]), .A2(a[25]), .ZN(n2617) );
  CKXOR2D1BWP12T U1908 ( .A1(a[26]), .A2(a[27]), .Z(n1041) );
  ND2D1BWP12T U1909 ( .A1(n2617), .A2(n1041), .ZN(n2619) );
  XNR2XD0BWP12T U1910 ( .A1(a[27]), .A2(n2868), .ZN(n1288) );
  XNR2XD1BWP12T U1911 ( .A1(a[27]), .A2(b[5]), .ZN(n2618) );
  OAI22D0BWP12T U1912 ( .A1(n2619), .A2(n1288), .B1(n2617), .B2(n2618), .ZN(
        mult_x_18_n738) );
  XNR2XD0BWP12T U1913 ( .A1(n2747), .A2(b[9]), .ZN(n2631) );
  OAI22D0BWP12T U1914 ( .A1(n2632), .A2(n1042), .B1(n2631), .B2(n2630), .ZN(
        mult_x_18_n754) );
  XNR2XD1BWP12T U1915 ( .A1(a[25]), .A2(b[5]), .ZN(n1246) );
  TPOAI22D0BWP12T U1916 ( .A1(n2608), .A2(n1246), .B1(n2606), .B2(n1043), .ZN(
        mult_x_18_n746) );
  IND2D0BWP12T U1917 ( .A1(n2231), .B1(n2725), .ZN(n1044) );
  OAI22D1BWP12T U1918 ( .A1(n2601), .A2(n2233), .B1(n2599), .B2(n1044), .ZN(
        n1047) );
  XNR2D1BWP12T U1919 ( .A1(n2594), .A2(n2897), .ZN(n1193) );
  XNR2D1BWP12T U1920 ( .A1(n2594), .A2(b[11]), .ZN(n1131) );
  OAI22D1BWP12T U1921 ( .A1(n2597), .A2(n1193), .B1(n1131), .B2(n2595), .ZN(
        n1046) );
  XNR2XD1BWP12T U1922 ( .A1(n2830), .A2(b[18]), .ZN(n1077) );
  XNR2D1BWP12T U1923 ( .A1(n2830), .A2(b[19]), .ZN(n1105) );
  OAI22D1BWP12T U1924 ( .A1(n2652), .A2(n1077), .B1(n2650), .B2(n1105), .ZN(
        n1045) );
  FA1D0BWP12T U1925 ( .A(n1047), .B(n1046), .CI(n1045), .CO(mult_x_18_n565), 
        .S(mult_x_18_n566) );
  INR2D1BWP12T U1926 ( .A1(n2231), .B1(n2630), .ZN(mult_x_18_n763) );
  IND2XD1BWP12T U1927 ( .A1(n2231), .B1(n2613), .ZN(n1048) );
  OAI22D1BWP12T U1928 ( .A1(n2616), .A2(n1049), .B1(n2614), .B2(n1048), .ZN(
        n1053) );
  XNR2D1BWP12T U1929 ( .A1(n2613), .A2(n2231), .ZN(n1050) );
  XNR2D1BWP12T U1930 ( .A1(n2613), .A2(n2477), .ZN(n1099) );
  XNR2D1BWP12T U1931 ( .A1(n2830), .A2(b[6]), .ZN(n1066) );
  XNR2D1BWP12T U1932 ( .A1(n2830), .A2(n2528), .ZN(n1190) );
  OAI22D1BWP12T U1933 ( .A1(n2652), .A2(n1066), .B1(n2650), .B2(n1190), .ZN(
        n1051) );
  FA1D0BWP12T U1934 ( .A(n1053), .B(n1052), .CI(n1051), .CO(mult_x_18_n688), 
        .S(mult_x_18_n689) );
  XNR2D1BWP12T U1935 ( .A1(n2482), .A2(b[15]), .ZN(n1336) );
  XNR2D1BWP12T U1936 ( .A1(n2482), .A2(b[16]), .ZN(n1303) );
  OAI22D1BWP12T U1937 ( .A1(n2604), .A2(n1336), .B1(n1303), .B2(n2603), .ZN(
        n1056) );
  INR2D1BWP12T U1938 ( .A1(n2231), .B1(n2647), .ZN(n1055) );
  XNR2D1BWP12T U1939 ( .A1(n2633), .A2(b[9]), .ZN(n1128) );
  XNR2XD1BWP12T U1940 ( .A1(n2633), .A2(n2897), .ZN(n1149) );
  OAI22D1BWP12T U1941 ( .A1(n2635), .A2(n1128), .B1(n1025), .B2(n1149), .ZN(
        n1054) );
  FA1D0BWP12T U1942 ( .A(n1056), .B(n1055), .CI(n1054), .CO(mult_x_18_n631), 
        .S(mult_x_18_n632) );
  XNR2D1BWP12T U1943 ( .A1(n2482), .A2(b[11]), .ZN(n1308) );
  XNR2D1BWP12T U1944 ( .A1(n2482), .A2(n2598), .ZN(n1325) );
  OAI22D1BWP12T U1945 ( .A1(n2604), .A2(n1308), .B1(n1325), .B2(n2603), .ZN(
        n1059) );
  INR2D1BWP12T U1946 ( .A1(n2231), .B1(n2644), .ZN(n1058) );
  XNR2D1BWP12T U1947 ( .A1(n2830), .A2(b[9]), .ZN(n1144) );
  XNR2D1BWP12T U1948 ( .A1(n2830), .A2(n2897), .ZN(n1062) );
  OAI22D1BWP12T U1949 ( .A1(n2652), .A2(n1144), .B1(n2650), .B2(n1062), .ZN(
        n1057) );
  FA1D0BWP12T U1950 ( .A(n1059), .B(n1058), .CI(n1057), .CO(mult_x_18_n669), 
        .S(mult_x_18_n670) );
  IND2D1BWP12T U1951 ( .A1(n2231), .B1(n2643), .ZN(n1060) );
  OAI22D1BWP12T U1952 ( .A1(n2646), .A2(n1061), .B1(n2644), .B2(n1060), .ZN(
        n1065) );
  XNR2D1BWP12T U1953 ( .A1(n2620), .A2(n2605), .ZN(n1191) );
  XNR2D1BWP12T U1954 ( .A1(n2620), .A2(b[9]), .ZN(n1245) );
  OAI22D1BWP12T U1955 ( .A1(n2623), .A2(n1191), .B1(n1245), .B2(n2621), .ZN(
        n1064) );
  XNR2D1BWP12T U1956 ( .A1(n2830), .A2(b[11]), .ZN(n1100) );
  OAI22D1BWP12T U1957 ( .A1(n2652), .A2(n1062), .B1(n2650), .B2(n1100), .ZN(
        n1063) );
  FA1D0BWP12T U1958 ( .A(n1065), .B(n1064), .CI(n1063), .CO(mult_x_18_n659), 
        .S(mult_x_18_n660) );
  XNR2D1BWP12T U1959 ( .A1(n2482), .A2(n2528), .ZN(n1290) );
  XNR2XD1BWP12T U1960 ( .A1(n2482), .A2(n2605), .ZN(n1331) );
  OAI22D1BWP12T U1961 ( .A1(n2604), .A2(n1290), .B1(n1331), .B2(n2603), .ZN(
        n1069) );
  INR2D1BWP12T U1962 ( .A1(n2231), .B1(n2614), .ZN(n1068) );
  XNR2D1BWP12T U1963 ( .A1(n2830), .A2(b[5]), .ZN(n1137) );
  OAI22D1BWP12T U1964 ( .A1(n2652), .A2(n1137), .B1(n2650), .B2(n1066), .ZN(
        n1067) );
  FA1D0BWP12T U1965 ( .A(n1069), .B(n1068), .CI(n1067), .CO(mult_x_18_n695), 
        .S(mult_x_18_n696) );
  XNR2D1BWP12T U1966 ( .A1(n2482), .A2(b[23]), .ZN(n1320) );
  XNR2D1BWP12T U1967 ( .A1(n2482), .A2(b[24]), .ZN(n1317) );
  OAI22D1BWP12T U1968 ( .A1(n2604), .A2(n1320), .B1(n1317), .B2(n2603), .ZN(
        n1072) );
  INR2D1BWP12T U1969 ( .A1(n2231), .B1(n2606), .ZN(n1071) );
  XNR2XD1BWP12T U1970 ( .A1(n2830), .A2(b[21]), .ZN(n1208) );
  XNR2XD1BWP12T U1971 ( .A1(n2830), .A2(b[22]), .ZN(n1081) );
  OAI22D1BWP12T U1972 ( .A1(n2652), .A2(n1208), .B1(n2650), .B2(n1081), .ZN(
        n1070) );
  FA1D0BWP12T U1973 ( .A(n1072), .B(n1071), .CI(n1070), .CO(mult_x_18_n519), 
        .S(mult_x_18_n520) );
  INR2D1BWP12T U1974 ( .A1(n2231), .B1(n2595), .ZN(mult_x_18_n871) );
  INR2D1BWP12T U1975 ( .A1(n2231), .B1(n1025), .ZN(mult_x_18_n923) );
  XNR2D1BWP12T U1976 ( .A1(n2594), .A2(b[6]), .ZN(n1145) );
  XNR2D1BWP12T U1977 ( .A1(n2594), .A2(n2528), .ZN(n1168) );
  OAI22D1BWP12T U1978 ( .A1(n2597), .A2(n1145), .B1(n1168), .B2(n2595), .ZN(
        n1076) );
  XNR2D1BWP12T U1979 ( .A1(n2679), .A2(n2231), .ZN(n1073) );
  XNR2D1BWP12T U1980 ( .A1(n2679), .A2(n2477), .ZN(n1126) );
  OAI22D1BWP12T U1981 ( .A1(n2649), .A2(n1073), .B1(n1126), .B2(n2647), .ZN(
        n1075) );
  XNR2D1BWP12T U1982 ( .A1(n2830), .A2(b[14]), .ZN(n1132) );
  XNR2D1BWP12T U1983 ( .A1(n2830), .A2(b[15]), .ZN(n1098) );
  OAI22D1BWP12T U1984 ( .A1(n2652), .A2(n1132), .B1(n2650), .B2(n1098), .ZN(
        n1074) );
  FA1D0BWP12T U1985 ( .A(n1076), .B(n1075), .CI(n1074), .CO(mult_x_18_n618), 
        .S(mult_x_18_n619) );
  INR2D1BWP12T U1986 ( .A1(n2231), .B1(n2610), .ZN(mult_x_18_n791) );
  XNR2XD1BWP12T U1987 ( .A1(n2482), .A2(b[19]), .ZN(n1342) );
  XNR2D1BWP12T U1988 ( .A1(n2482), .A2(b[20]), .ZN(n1297) );
  OAI22D1BWP12T U1989 ( .A1(n2604), .A2(n1342), .B1(n1297), .B2(n2603), .ZN(
        n1080) );
  INR2D1BWP12T U1990 ( .A1(n2231), .B1(n2599), .ZN(n1079) );
  XNR2XD1BWP12T U1991 ( .A1(n2830), .A2(b[17]), .ZN(n1120) );
  OAI22D1BWP12T U1992 ( .A1(n2652), .A2(n1120), .B1(n2650), .B2(n1077), .ZN(
        n1078) );
  FA1D0BWP12T U1993 ( .A(n1080), .B(n1079), .CI(n1078), .CO(mult_x_18_n581), 
        .S(mult_x_18_n582) );
  XNR2D0BWP12T U1994 ( .A1(n2594), .A2(b[14]), .ZN(n1158) );
  XNR2D0BWP12T U1995 ( .A1(n2594), .A2(b[15]), .ZN(n1221) );
  OAI22D1BWP12T U1996 ( .A1(n2597), .A2(n1158), .B1(n1221), .B2(n2595), .ZN(
        n1084) );
  XNR2D1BWP12T U1997 ( .A1(n2747), .A2(n2639), .ZN(n1116) );
  XNR2D1BWP12T U1998 ( .A1(n2747), .A2(n2831), .ZN(n1152) );
  OAI22D1BWP12T U1999 ( .A1(n2632), .A2(n1116), .B1(n1152), .B2(n2630), .ZN(
        n1083) );
  XNR2XD1BWP12T U2000 ( .A1(n2830), .A2(b[23]), .ZN(n1141) );
  OAI22D1BWP12T U2001 ( .A1(n2652), .A2(n1081), .B1(n2650), .B2(n1141), .ZN(
        n1082) );
  FA1D0BWP12T U2002 ( .A(n1084), .B(n1083), .CI(n1082), .CO(mult_x_18_n500), 
        .S(mult_x_18_n501) );
  INR2D1BWP12T U2003 ( .A1(n2231), .B1(n2627), .ZN(mult_x_18_n827) );
  INR2D1BWP12T U2004 ( .A1(n2231), .B1(n2617), .ZN(mult_x_18_n743) );
  OAI22D0BWP12T U2005 ( .A1(n2604), .A2(n1086), .B1(n1085), .B2(n2603), .ZN(
        n1089) );
  INR2D1BWP12T U2006 ( .A1(n2231), .B1(n2636), .ZN(n1088) );
  XNR2D0BWP12T U2007 ( .A1(n2613), .A2(b[19]), .ZN(n1258) );
  XNR2D0BWP12T U2008 ( .A1(n2613), .A2(b[20]), .ZN(n1281) );
  OAI22D1BWP12T U2009 ( .A1(n2616), .A2(n1258), .B1(n2614), .B2(n1281), .ZN(
        n1087) );
  FA1D0BWP12T U2010 ( .A(n1089), .B(n1088), .CI(n1087), .CO(mult_x_18_n445), 
        .S(mult_x_18_n446) );
  XNR2D1BWP12T U2011 ( .A1(n2747), .A2(b[6]), .ZN(n1261) );
  OAI22D1BWP12T U2012 ( .A1(n2632), .A2(n1261), .B1(n1090), .B2(n2630), .ZN(
        n1096) );
  XNR2XD1BWP12T U2013 ( .A1(a[29]), .A2(n2231), .ZN(n1091) );
  XNR2XD1BWP12T U2014 ( .A1(a[29]), .A2(n2477), .ZN(n1234) );
  OAI22D1BWP12T U2015 ( .A1(n2638), .A2(n1091), .B1(n1234), .B2(n2636), .ZN(
        n1095) );
  TPOAI22D0BWP12T U2016 ( .A1(n2652), .A2(n1093), .B1(n2650), .B2(n1092), .ZN(
        n1094) );
  FA1D0BWP12T U2017 ( .A(n1096), .B(n1095), .CI(n1094), .CO(mult_x_18_n423), 
        .S(mult_x_18_n424) );
  INR2D1BWP12T U2018 ( .A1(n2231), .B1(n2640), .ZN(mult_x_18_n731) );
  XNR2D1BWP12T U2019 ( .A1(n2747), .A2(n2231), .ZN(n1097) );
  XNR2D1BWP12T U2020 ( .A1(n2747), .A2(n2477), .ZN(n1117) );
  OAI22D1BWP12T U2021 ( .A1(n2632), .A2(n1097), .B1(n1117), .B2(n2630), .ZN(
        mult_x_18_n762) );
  XNR2XD1BWP12T U2022 ( .A1(n2613), .A2(b[14]), .ZN(n1181) );
  XNR2XD1BWP12T U2023 ( .A1(n2613), .A2(b[15]), .ZN(n1196) );
  OAI22D1BWP12T U2024 ( .A1(n2616), .A2(n1181), .B1(n2614), .B2(n1196), .ZN(
        mult_x_18_n881) );
  XNR2D1BWP12T U2025 ( .A1(n2482), .A2(b[21]), .ZN(n1296) );
  XNR2D1BWP12T U2026 ( .A1(n2482), .A2(b[22]), .ZN(n1321) );
  OAI22D1BWP12T U2027 ( .A1(n2604), .A2(n1296), .B1(n1321), .B2(n2603), .ZN(
        mult_x_18_n994) );
  XNR2D1BWP12T U2028 ( .A1(n2679), .A2(b[5]), .ZN(n1298) );
  XNR2D1BWP12T U2029 ( .A1(n2679), .A2(b[6]), .ZN(n1323) );
  OAI22D1BWP12T U2030 ( .A1(n2649), .A2(n1298), .B1(n1323), .B2(n2647), .ZN(
        mult_x_18_n802) );
  XNR2D1BWP12T U2031 ( .A1(n2620), .A2(b[16]), .ZN(n1172) );
  XNR2D1BWP12T U2032 ( .A1(n2620), .A2(b[17]), .ZN(n1134) );
  OAI22D1BWP12T U2033 ( .A1(n2623), .A2(n1172), .B1(n1134), .B2(n2621), .ZN(
        mult_x_18_n935) );
  XNR2XD1BWP12T U2034 ( .A1(n2725), .A2(n2639), .ZN(n1226) );
  XNR2D1BWP12T U2035 ( .A1(n2725), .A2(n2831), .ZN(n1127) );
  OAI22D1BWP12T U2036 ( .A1(n2601), .A2(n1226), .B1(n2599), .B2(n1127), .ZN(
        mult_x_18_n773) );
  XNR2D1BWP12T U2037 ( .A1(n2830), .A2(b[16]), .ZN(n1121) );
  OAI22D1BWP12T U2038 ( .A1(n2652), .A2(n1098), .B1(n2650), .B2(n1121), .ZN(
        mult_x_18_n967) );
  XNR2D1BWP12T U2039 ( .A1(n2626), .A2(n2605), .ZN(n1103) );
  XNR2D1BWP12T U2040 ( .A1(n2626), .A2(b[9]), .ZN(n1206) );
  OAI22D1BWP12T U2041 ( .A1(n2629), .A2(n1103), .B1(n2627), .B2(n1206), .ZN(
        mult_x_18_n818) );
  XNR2D1BWP12T U2042 ( .A1(n2609), .A2(n2639), .ZN(n1241) );
  XNR2D1BWP12T U2043 ( .A1(n2609), .A2(n2831), .ZN(n1104) );
  OAI22D1BWP12T U2044 ( .A1(n2612), .A2(n1241), .B1(n2610), .B2(n1104), .ZN(
        mult_x_18_n788) );
  XNR2XD1BWP12T U2045 ( .A1(n2633), .A2(b[15]), .ZN(n1186) );
  XNR2XD1BWP12T U2046 ( .A1(n2633), .A2(b[16]), .ZN(n1102) );
  OAI22D1BWP12T U2047 ( .A1(n2635), .A2(n1186), .B1(n1025), .B2(n1102), .ZN(
        mult_x_18_n907) );
  XNR2D1BWP12T U2048 ( .A1(n2643), .A2(b[9]), .ZN(n1266) );
  XNR2D1BWP12T U2049 ( .A1(n2643), .A2(n2897), .ZN(n1212) );
  OAI22D1BWP12T U2050 ( .A1(n2646), .A2(n1266), .B1(n2644), .B2(n1212), .ZN(
        mult_x_18_n838) );
  XNR2D1BWP12T U2051 ( .A1(n2594), .A2(n2598), .ZN(n1130) );
  XNR2D0BWP12T U2052 ( .A1(n2594), .A2(b[13]), .ZN(n1159) );
  OAI22D1BWP12T U2053 ( .A1(n2597), .A2(n1130), .B1(n1159), .B2(n2595), .ZN(
        mult_x_18_n858) );
  XNR2XD1BWP12T U2054 ( .A1(n2633), .A2(b[17]), .ZN(n1101) );
  XNR2XD1BWP12T U2055 ( .A1(n2633), .A2(b[18]), .ZN(n1205) );
  OAI22D1BWP12T U2056 ( .A1(n2635), .A2(n1101), .B1(n1025), .B2(n1205), .ZN(
        mult_x_18_n905) );
  XNR2D1BWP12T U2057 ( .A1(n2613), .A2(n2639), .ZN(n1154) );
  OAI22D1BWP12T U2058 ( .A1(n2616), .A2(n1099), .B1(n2614), .B2(n1154), .ZN(
        mult_x_18_n894) );
  XNR2D1BWP12T U2059 ( .A1(n2620), .A2(n2598), .ZN(n1113) );
  XNR2D1BWP12T U2060 ( .A1(n2620), .A2(b[13]), .ZN(n1148) );
  OAI22D1BWP12T U2061 ( .A1(n2623), .A2(n1113), .B1(n1148), .B2(n2621), .ZN(
        mult_x_18_n939) );
  XNR2D1BWP12T U2062 ( .A1(n2613), .A2(n2605), .ZN(n1106) );
  XNR2D1BWP12T U2063 ( .A1(n2613), .A2(b[9]), .ZN(n1111) );
  OAI22D1BWP12T U2064 ( .A1(n2616), .A2(n1106), .B1(n2614), .B2(n1111), .ZN(
        mult_x_18_n887) );
  XNR2D1BWP12T U2065 ( .A1(n2830), .A2(n2598), .ZN(n1136) );
  OAI22D1BWP12T U2066 ( .A1(n2652), .A2(n1100), .B1(n2650), .B2(n1136), .ZN(
        mult_x_18_n971) );
  XNR2D1BWP12T U2067 ( .A1(n2594), .A2(n2831), .ZN(n1326) );
  XNR2D1BWP12T U2068 ( .A1(n2594), .A2(n2868), .ZN(n1339) );
  OAI22D1BWP12T U2069 ( .A1(n2597), .A2(n1326), .B1(n1339), .B2(n2595), .ZN(
        mult_x_18_n867) );
  XNR2D1BWP12T U2070 ( .A1(n2482), .A2(b[17]), .ZN(n1302) );
  XNR2D1BWP12T U2071 ( .A1(n2482), .A2(b[18]), .ZN(n1343) );
  OAI22D1BWP12T U2072 ( .A1(n2604), .A2(n1302), .B1(n1343), .B2(n2603), .ZN(
        mult_x_18_n998) );
  OAI22D1BWP12T U2073 ( .A1(n2635), .A2(n1102), .B1(n1025), .B2(n1101), .ZN(
        mult_x_18_n906) );
  XNR2D1BWP12T U2074 ( .A1(n2626), .A2(n2528), .ZN(n1156) );
  OAI22D1BWP12T U2075 ( .A1(n2629), .A2(n1156), .B1(n2627), .B2(n1103), .ZN(
        mult_x_18_n819) );
  XNR2D1BWP12T U2076 ( .A1(n2620), .A2(n2831), .ZN(n1292) );
  XNR2D1BWP12T U2077 ( .A1(n2620), .A2(n2868), .ZN(n1333) );
  OAI22D1BWP12T U2078 ( .A1(n2623), .A2(n1292), .B1(n1333), .B2(n2621), .ZN(
        mult_x_18_n948) );
  XNR2D1BWP12T U2079 ( .A1(n2609), .A2(n2868), .ZN(n1115) );
  OAI22D1BWP12T U2080 ( .A1(n2612), .A2(n1104), .B1(n2610), .B2(n1115), .ZN(
        mult_x_18_n787) );
  XNR2XD1BWP12T U2081 ( .A1(n2830), .A2(b[20]), .ZN(n1209) );
  OAI22D1BWP12T U2082 ( .A1(n2652), .A2(n1105), .B1(n2650), .B2(n1209), .ZN(
        mult_x_18_n963) );
  XNR2D1BWP12T U2083 ( .A1(n2613), .A2(n2528), .ZN(n1213) );
  OAI22D1BWP12T U2084 ( .A1(n2616), .A2(n1213), .B1(n2614), .B2(n1106), .ZN(
        mult_x_18_n888) );
  XNR2XD1BWP12T U2085 ( .A1(n2620), .A2(b[20]), .ZN(n1109) );
  XNR2XD1BWP12T U2086 ( .A1(n2620), .A2(b[21]), .ZN(n1199) );
  OAI22D1BWP12T U2087 ( .A1(n2623), .A2(n1109), .B1(n1199), .B2(n2621), .ZN(
        mult_x_18_n931) );
  IND2D0BWP12T U2088 ( .A1(n2231), .B1(a[25]), .ZN(n1107) );
  OAI22D1BWP12T U2089 ( .A1(n2608), .A2(n1108), .B1(n2606), .B2(n1107), .ZN(
        mult_x_18_n716) );
  XNR2XD1BWP12T U2090 ( .A1(n2643), .A2(b[11]), .ZN(n1211) );
  XNR2XD1BWP12T U2091 ( .A1(n2643), .A2(n2598), .ZN(n1230) );
  OAI22D1BWP12T U2092 ( .A1(n2646), .A2(n1211), .B1(n2644), .B2(n1230), .ZN(
        mult_x_18_n836) );
  XNR2XD1BWP12T U2093 ( .A1(n2620), .A2(b[19]), .ZN(n1197) );
  OAI22D1BWP12T U2094 ( .A1(n2623), .A2(n1197), .B1(n1109), .B2(n2621), .ZN(
        mult_x_18_n932) );
  XNR2D1BWP12T U2095 ( .A1(n2482), .A2(b[9]), .ZN(n1330) );
  XNR2D1BWP12T U2096 ( .A1(n2482), .A2(n2897), .ZN(n1309) );
  OAI22D1BWP12T U2097 ( .A1(n2604), .A2(n1330), .B1(n1309), .B2(n2603), .ZN(
        mult_x_18_n1006) );
  XNR2D1BWP12T U2098 ( .A1(n2613), .A2(n2831), .ZN(n1153) );
  XNR2D1BWP12T U2099 ( .A1(n2613), .A2(n2868), .ZN(n1122) );
  XNR2D1BWP12T U2100 ( .A1(n2679), .A2(n2528), .ZN(n1322) );
  XNR2D1BWP12T U2101 ( .A1(n2679), .A2(n2605), .ZN(n1319) );
  OAI22D1BWP12T U2102 ( .A1(n2649), .A2(n1322), .B1(n1319), .B2(n2647), .ZN(
        mult_x_18_n800) );
  XNR2D1BWP12T U2103 ( .A1(n2626), .A2(n2868), .ZN(n1169) );
  XNR2D1BWP12T U2104 ( .A1(n2626), .A2(b[5]), .ZN(n1238) );
  OAI22D1BWP12T U2105 ( .A1(n2629), .A2(n1169), .B1(n2627), .B2(n1238), .ZN(
        mult_x_18_n822) );
  XNR2D1BWP12T U2106 ( .A1(n2679), .A2(n2831), .ZN(n1344) );
  XNR2D1BWP12T U2107 ( .A1(n2679), .A2(n2868), .ZN(n1299) );
  OAI22D1BWP12T U2108 ( .A1(n2649), .A2(n1344), .B1(n1299), .B2(n2647), .ZN(
        mult_x_18_n804) );
  XNR2D1BWP12T U2109 ( .A1(n2633), .A2(n2231), .ZN(n1110) );
  XNR2D1BWP12T U2110 ( .A1(n2633), .A2(n2477), .ZN(n1129) );
  OAI22D1BWP12T U2111 ( .A1(n2635), .A2(n1110), .B1(n1025), .B2(n1129), .ZN(
        mult_x_18_n922) );
  XNR2XD1BWP12T U2112 ( .A1(n2613), .A2(n2897), .ZN(n1176) );
  OAI22D1BWP12T U2113 ( .A1(n2616), .A2(n1111), .B1(n2614), .B2(n1176), .ZN(
        mult_x_18_n886) );
  XNR2D1BWP12T U2114 ( .A1(n2620), .A2(n2639), .ZN(n1293) );
  OAI22D1BWP12T U2115 ( .A1(n2623), .A2(n1112), .B1(n1293), .B2(n2621), .ZN(
        mult_x_18_n950) );
  OAI22D1BWP12T U2116 ( .A1(n2623), .A2(n1114), .B1(n1113), .B2(n2621), .ZN(
        mult_x_18_n940) );
  XNR2D1BWP12T U2117 ( .A1(n2609), .A2(b[5]), .ZN(n1201) );
  OAI22D1BWP12T U2118 ( .A1(n2612), .A2(n1115), .B1(n2610), .B2(n1201), .ZN(
        mult_x_18_n786) );
  OAI22D1BWP12T U2119 ( .A1(n2632), .A2(n1117), .B1(n1116), .B2(n2630), .ZN(
        mult_x_18_n761) );
  XNR2D1BWP12T U2120 ( .A1(n2620), .A2(b[6]), .ZN(n1140) );
  XNR2D1BWP12T U2121 ( .A1(n2620), .A2(n2528), .ZN(n1192) );
  OAI22D1BWP12T U2122 ( .A1(n2623), .A2(n1140), .B1(n1192), .B2(n2621), .ZN(
        mult_x_18_n945) );
  IND2XD1BWP12T U2123 ( .A1(n2231), .B1(n2633), .ZN(n1118) );
  OAI22D1BWP12T U2124 ( .A1(n2635), .A2(n1119), .B1(n1025), .B2(n1118), .ZN(
        mult_x_18_n725) );
  OAI22D1BWP12T U2125 ( .A1(n2652), .A2(n1121), .B1(n2650), .B2(n1120), .ZN(
        mult_x_18_n966) );
  XNR2D1BWP12T U2126 ( .A1(n2613), .A2(b[5]), .ZN(n1123) );
  OAI22D1BWP12T U2127 ( .A1(n2616), .A2(n1122), .B1(n2614), .B2(n1123), .ZN(
        mult_x_18_n891) );
  XNR2D1BWP12T U2128 ( .A1(n2613), .A2(b[6]), .ZN(n1214) );
  OAI22D1BWP12T U2129 ( .A1(n2616), .A2(n1123), .B1(n2614), .B2(n1214), .ZN(
        mult_x_18_n890) );
  XNR2XD1BWP12T U2130 ( .A1(n2633), .A2(n2598), .ZN(n1184) );
  XNR2XD1BWP12T U2131 ( .A1(n2633), .A2(b[13]), .ZN(n1177) );
  OAI22D1BWP12T U2132 ( .A1(n2635), .A2(n1184), .B1(n1025), .B2(n1177), .ZN(
        mult_x_18_n910) );
  XNR2D1BWP12T U2133 ( .A1(n2725), .A2(n2231), .ZN(n1124) );
  XNR2D1BWP12T U2134 ( .A1(n2725), .A2(n2477), .ZN(n1227) );
  OAI22D1BWP12T U2135 ( .A1(n2601), .A2(n1124), .B1(n2599), .B2(n1227), .ZN(
        mult_x_18_n775) );
  XNR2D1BWP12T U2136 ( .A1(n2482), .A2(b[6]), .ZN(n1291) );
  OAI22D1BWP12T U2137 ( .A1(n2604), .A2(n1125), .B1(n1291), .B2(n2603), .ZN(
        mult_x_18_n1010) );
  XNR2D1BWP12T U2138 ( .A1(n2725), .A2(b[6]), .ZN(n1224) );
  XNR2D1BWP12T U2139 ( .A1(n2725), .A2(n2528), .ZN(n1243) );
  OAI22D1BWP12T U2140 ( .A1(n2601), .A2(n1224), .B1(n2599), .B2(n1243), .ZN(
        mult_x_18_n769) );
  XNR2D1BWP12T U2141 ( .A1(n2679), .A2(n2639), .ZN(n1345) );
  OAI22D1BWP12T U2142 ( .A1(n2649), .A2(n1126), .B1(n1345), .B2(n2647), .ZN(
        mult_x_18_n806) );
  XNR2D1BWP12T U2143 ( .A1(n2725), .A2(n2868), .ZN(n1171) );
  OAI22D1BWP12T U2144 ( .A1(n2601), .A2(n1127), .B1(n2599), .B2(n1171), .ZN(
        mult_x_18_n772) );
  XNR2XD1BWP12T U2145 ( .A1(n2613), .A2(n2598), .ZN(n1239) );
  XNR2XD1BWP12T U2146 ( .A1(n2613), .A2(b[13]), .ZN(n1182) );
  OAI22D1BWP12T U2147 ( .A1(n2616), .A2(n1239), .B1(n2614), .B2(n1182), .ZN(
        mult_x_18_n883) );
  XNR2D1BWP12T U2148 ( .A1(n2633), .A2(n2605), .ZN(n1200) );
  OAI22D1BWP12T U2149 ( .A1(n2635), .A2(n1200), .B1(n1025), .B2(n1128), .ZN(
        mult_x_18_n914) );
  XNR2D1BWP12T U2150 ( .A1(n2633), .A2(n2639), .ZN(n1163) );
  OAI22D1BWP12T U2151 ( .A1(n2635), .A2(n1129), .B1(n1025), .B2(n1163), .ZN(
        mult_x_18_n921) );
  OAI22D1BWP12T U2152 ( .A1(n2597), .A2(n1131), .B1(n1130), .B2(n2595), .ZN(
        mult_x_18_n859) );
  XNR2D1BWP12T U2153 ( .A1(n2830), .A2(b[13]), .ZN(n1135) );
  OAI22D1BWP12T U2154 ( .A1(n2652), .A2(n1135), .B1(n2650), .B2(n1132), .ZN(
        mult_x_18_n969) );
  XNR2D1BWP12T U2155 ( .A1(n2643), .A2(n2868), .ZN(n1178) );
  XNR2D1BWP12T U2156 ( .A1(n2643), .A2(b[5]), .ZN(n1143) );
  OAI22D1BWP12T U2157 ( .A1(n2646), .A2(n1178), .B1(n2644), .B2(n1143), .ZN(
        mult_x_18_n843) );
  XNR2D1BWP12T U2158 ( .A1(n2482), .A2(b[13]), .ZN(n1324) );
  XNR2D1BWP12T U2159 ( .A1(n2482), .A2(b[14]), .ZN(n1337) );
  OAI22D1BWP12T U2160 ( .A1(n2604), .A2(n1324), .B1(n1337), .B2(n2603), .ZN(
        mult_x_18_n1002) );
  XNR2D1BWP12T U2161 ( .A1(n2609), .A2(n2231), .ZN(n1133) );
  XNR2D1BWP12T U2162 ( .A1(n2609), .A2(n2477), .ZN(n1242) );
  OAI22D1BWP12T U2163 ( .A1(n2612), .A2(n1133), .B1(n2610), .B2(n1242), .ZN(
        mult_x_18_n790) );
  XNR2XD1BWP12T U2164 ( .A1(n2620), .A2(b[18]), .ZN(n1198) );
  OAI22D1BWP12T U2165 ( .A1(n2623), .A2(n1134), .B1(n1198), .B2(n2621), .ZN(
        mult_x_18_n934) );
  OAI22D1BWP12T U2166 ( .A1(n2652), .A2(n1136), .B1(n2650), .B2(n1135), .ZN(
        mult_x_18_n970) );
  XNR2D1BWP12T U2167 ( .A1(n2830), .A2(n2868), .ZN(n1146) );
  OAI22D1BWP12T U2168 ( .A1(n2652), .A2(n1146), .B1(n2650), .B2(n1137), .ZN(
        mult_x_18_n978) );
  XNR2XD1BWP12T U2169 ( .A1(a[25]), .A2(n2231), .ZN(n1138) );
  OAI22D1BWP12T U2170 ( .A1(n2608), .A2(n1138), .B1(n2606), .B2(n1215), .ZN(
        mult_x_18_n751) );
  XNR2D1BWP12T U2171 ( .A1(n2633), .A2(n2868), .ZN(n1151) );
  OAI22D1BWP12T U2172 ( .A1(n2635), .A2(n1151), .B1(n1025), .B2(n1139), .ZN(
        mult_x_18_n918) );
  XNR2D1BWP12T U2173 ( .A1(n2620), .A2(b[5]), .ZN(n1332) );
  OAI22D1BWP12T U2174 ( .A1(n2623), .A2(n1332), .B1(n1140), .B2(n2621), .ZN(
        mult_x_18_n946) );
  XNR2XD1BWP12T U2175 ( .A1(n2830), .A2(b[24]), .ZN(n1236) );
  OAI22D1BWP12T U2176 ( .A1(n2652), .A2(n1141), .B1(n2650), .B2(n1236), .ZN(
        mult_x_18_n959) );
  XNR2XD1BWP12T U2177 ( .A1(n2613), .A2(b[16]), .ZN(n1195) );
  XNR2XD1BWP12T U2178 ( .A1(n2613), .A2(b[17]), .ZN(n1142) );
  OAI22D1BWP12T U2179 ( .A1(n2616), .A2(n1195), .B1(n2614), .B2(n1142), .ZN(
        mult_x_18_n879) );
  XNR2XD1BWP12T U2180 ( .A1(n2613), .A2(b[18]), .ZN(n1259) );
  OAI22D1BWP12T U2181 ( .A1(n2616), .A2(n1142), .B1(n2614), .B2(n1259), .ZN(
        mult_x_18_n878) );
  XNR2D1BWP12T U2182 ( .A1(n2643), .A2(b[6]), .ZN(n1179) );
  OAI22D1BWP12T U2183 ( .A1(n2646), .A2(n1143), .B1(n2644), .B2(n1179), .ZN(
        mult_x_18_n842) );
  XNR2D1BWP12T U2184 ( .A1(n2830), .A2(n2605), .ZN(n1189) );
  OAI22D1BWP12T U2185 ( .A1(n2652), .A2(n1189), .B1(n2650), .B2(n1144), .ZN(
        mult_x_18_n974) );
  XNR2D1BWP12T U2186 ( .A1(n2594), .A2(b[5]), .ZN(n1338) );
  OAI22D1BWP12T U2187 ( .A1(n2597), .A2(n1338), .B1(n1145), .B2(n2595), .ZN(
        mult_x_18_n865) );
  OAI22D1BWP12T U2188 ( .A1(n2652), .A2(n1147), .B1(n2650), .B2(n1146), .ZN(
        mult_x_18_n979) );
  XNR2XD1BWP12T U2189 ( .A1(n2620), .A2(b[14]), .ZN(n1164) );
  OAI22D1BWP12T U2190 ( .A1(n2623), .A2(n1148), .B1(n1164), .B2(n2621), .ZN(
        mult_x_18_n938) );
  XNR2D1BWP12T U2191 ( .A1(n2594), .A2(n2605), .ZN(n1167) );
  XNR2D1BWP12T U2192 ( .A1(n2594), .A2(b[9]), .ZN(n1194) );
  OAI22D1BWP12T U2193 ( .A1(n2597), .A2(n1167), .B1(n1194), .B2(n2595), .ZN(
        mult_x_18_n862) );
  XNR2XD1BWP12T U2194 ( .A1(n2633), .A2(b[11]), .ZN(n1185) );
  OAI22D1BWP12T U2195 ( .A1(n2635), .A2(n1149), .B1(n1025), .B2(n1185), .ZN(
        mult_x_18_n912) );
  XNR2D1BWP12T U2196 ( .A1(n2643), .A2(n2231), .ZN(n1150) );
  XNR2D1BWP12T U2197 ( .A1(n2643), .A2(n2477), .ZN(n1155) );
  OAI22D1BWP12T U2198 ( .A1(n2646), .A2(n1150), .B1(n2644), .B2(n1155), .ZN(
        mult_x_18_n847) );
  XNR2D1BWP12T U2199 ( .A1(n2633), .A2(n2831), .ZN(n1162) );
  OAI22D1BWP12T U2200 ( .A1(n2635), .A2(n1162), .B1(n1025), .B2(n1151), .ZN(
        mult_x_18_n919) );
  XNR2XD1BWP12T U2201 ( .A1(n2747), .A2(n2868), .ZN(n1228) );
  OAI22D1BWP12T U2202 ( .A1(n2632), .A2(n1152), .B1(n1228), .B2(n2630), .ZN(
        mult_x_18_n759) );
  OAI22D1BWP12T U2203 ( .A1(n2616), .A2(n1154), .B1(n2614), .B2(n1153), .ZN(
        mult_x_18_n893) );
  XNR2D1BWP12T U2204 ( .A1(n2643), .A2(n2639), .ZN(n1217) );
  OAI22D1BWP12T U2205 ( .A1(n2646), .A2(n1155), .B1(n2644), .B2(n1217), .ZN(
        mult_x_18_n846) );
  XNR2D1BWP12T U2206 ( .A1(n2626), .A2(n2639), .ZN(n1174) );
  XNR2D1BWP12T U2207 ( .A1(n2626), .A2(n2831), .ZN(n1170) );
  OAI22D1BWP12T U2208 ( .A1(n2629), .A2(n1174), .B1(n2627), .B2(n1170), .ZN(
        mult_x_18_n824) );
  XNR2D1BWP12T U2209 ( .A1(n2626), .A2(b[6]), .ZN(n1237) );
  OAI22D1BWP12T U2210 ( .A1(n2629), .A2(n1237), .B1(n2627), .B2(n1156), .ZN(
        mult_x_18_n820) );
  IND2D0BWP12T U2211 ( .A1(n2231), .B1(a[27]), .ZN(n1157) );
  OAI22D1BWP12T U2212 ( .A1(n2619), .A2(n1816), .B1(n2617), .B2(n1157), .ZN(
        mult_x_18_n715) );
  OAI22D1BWP12T U2213 ( .A1(n2597), .A2(n1159), .B1(n1158), .B2(n2595), .ZN(
        mult_x_18_n857) );
  XNR2D1BWP12T U2214 ( .A1(n2594), .A2(n2231), .ZN(n1161) );
  OAI22D1BWP12T U2215 ( .A1(n2597), .A2(n1161), .B1(n1160), .B2(n2595), .ZN(
        mult_x_18_n870) );
  OAI22D1BWP12T U2216 ( .A1(n2635), .A2(n1163), .B1(n1025), .B2(n1162), .ZN(
        mult_x_18_n920) );
  XNR2XD1BWP12T U2217 ( .A1(n2620), .A2(b[15]), .ZN(n1173) );
  OAI22D1BWP12T U2218 ( .A1(n2623), .A2(n1164), .B1(n1173), .B2(n2621), .ZN(
        mult_x_18_n937) );
  XNR2D1BWP12T U2219 ( .A1(n2626), .A2(n2231), .ZN(n1165) );
  XNR2D1BWP12T U2220 ( .A1(n2626), .A2(n2477), .ZN(n1175) );
  OAI22D1BWP12T U2221 ( .A1(n2629), .A2(n1165), .B1(n2627), .B2(n1175), .ZN(
        mult_x_18_n826) );
  IND2XD0BWP12T U2222 ( .A1(n2231), .B1(n2747), .ZN(n1166) );
  OAI22D1BWP12T U2223 ( .A1(n2632), .A2(n2751), .B1(n2630), .B2(n1166), .ZN(
        mult_x_18_n717) );
  OAI22D1BWP12T U2224 ( .A1(n2597), .A2(n1168), .B1(n1167), .B2(n2595), .ZN(
        mult_x_18_n863) );
  OAI22D1BWP12T U2225 ( .A1(n2629), .A2(n1170), .B1(n2627), .B2(n1169), .ZN(
        mult_x_18_n823) );
  XNR2D1BWP12T U2226 ( .A1(n2725), .A2(b[5]), .ZN(n1225) );
  OAI22D1BWP12T U2227 ( .A1(n2601), .A2(n1171), .B1(n2599), .B2(n1225), .ZN(
        mult_x_18_n771) );
  OAI22D1BWP12T U2228 ( .A1(n2623), .A2(n1173), .B1(n1172), .B2(n2621), .ZN(
        mult_x_18_n936) );
  OAI22D1BWP12T U2229 ( .A1(n2629), .A2(n1175), .B1(n2627), .B2(n1174), .ZN(
        mult_x_18_n825) );
  XNR2XD1BWP12T U2230 ( .A1(n2613), .A2(b[11]), .ZN(n1240) );
  OAI22D1BWP12T U2231 ( .A1(n2616), .A2(n1176), .B1(n2614), .B2(n1240), .ZN(
        mult_x_18_n885) );
  XNR2XD1BWP12T U2232 ( .A1(n2633), .A2(b[14]), .ZN(n1187) );
  OAI22D1BWP12T U2233 ( .A1(n2635), .A2(n1177), .B1(n1025), .B2(n1187), .ZN(
        mult_x_18_n909) );
  XNR2D1BWP12T U2234 ( .A1(n2643), .A2(n2831), .ZN(n1216) );
  OAI22D1BWP12T U2235 ( .A1(n2646), .A2(n1216), .B1(n2644), .B2(n1178), .ZN(
        mult_x_18_n844) );
  XNR2D0BWP12T U2236 ( .A1(n2643), .A2(b[13]), .ZN(n1229) );
  XNR2D0BWP12T U2237 ( .A1(n2643), .A2(b[14]), .ZN(n1248) );
  OAI22D1BWP12T U2238 ( .A1(n2646), .A2(n1229), .B1(n2644), .B2(n1248), .ZN(
        mult_x_18_n834) );
  XNR2D1BWP12T U2239 ( .A1(n2643), .A2(n2528), .ZN(n1188) );
  OAI22D1BWP12T U2240 ( .A1(n2646), .A2(n1179), .B1(n2644), .B2(n1188), .ZN(
        mult_x_18_n841) );
  XNR2D1BWP12T U2241 ( .A1(n2679), .A2(b[9]), .ZN(n1318) );
  OAI22D1BWP12T U2242 ( .A1(n2649), .A2(n1318), .B1(n1180), .B2(n2647), .ZN(
        mult_x_18_n798) );
  OAI22D1BWP12T U2243 ( .A1(n2616), .A2(n1182), .B1(n2614), .B2(n1181), .ZN(
        mult_x_18_n882) );
  XNR2D0BWP12T U2244 ( .A1(n2482), .A2(b[25]), .ZN(n1316) );
  OAI22D1BWP12T U2245 ( .A1(n2604), .A2(n1316), .B1(n1183), .B2(n2603), .ZN(
        mult_x_18_n990) );
  OAI22D1BWP12T U2246 ( .A1(n2635), .A2(n1185), .B1(n1025), .B2(n1184), .ZN(
        mult_x_18_n911) );
  OAI22D1BWP12T U2247 ( .A1(n2635), .A2(n1187), .B1(n1025), .B2(n1186), .ZN(
        mult_x_18_n908) );
  XNR2D1BWP12T U2248 ( .A1(n2643), .A2(n2605), .ZN(n1267) );
  OAI22D1BWP12T U2249 ( .A1(n2646), .A2(n1188), .B1(n2644), .B2(n1267), .ZN(
        mult_x_18_n840) );
  OAI22D1BWP12T U2250 ( .A1(n2652), .A2(n1190), .B1(n2650), .B2(n1189), .ZN(
        mult_x_18_n975) );
  OAI22D1BWP12T U2251 ( .A1(n2623), .A2(n1192), .B1(n1191), .B2(n2621), .ZN(
        mult_x_18_n944) );
  OAI22D1BWP12T U2252 ( .A1(n2597), .A2(n1194), .B1(n1193), .B2(n2595), .ZN(
        mult_x_18_n861) );
  OAI22D1BWP12T U2253 ( .A1(n2616), .A2(n1196), .B1(n2614), .B2(n1195), .ZN(
        mult_x_18_n880) );
  OAI22D1BWP12T U2254 ( .A1(n2623), .A2(n1198), .B1(n1197), .B2(n2621), .ZN(
        mult_x_18_n933) );
  XNR2XD1BWP12T U2255 ( .A1(n2620), .A2(b[22]), .ZN(n1204) );
  OAI22D1BWP12T U2256 ( .A1(n2623), .A2(n1199), .B1(n1204), .B2(n2621), .ZN(
        mult_x_18_n930) );
  XNR2D1BWP12T U2257 ( .A1(n2633), .A2(n2528), .ZN(n1202) );
  OAI22D1BWP12T U2258 ( .A1(n2635), .A2(n1202), .B1(n1025), .B2(n1200), .ZN(
        mult_x_18_n915) );
  XNR2D1BWP12T U2259 ( .A1(n2609), .A2(b[6]), .ZN(n1220) );
  OAI22D1BWP12T U2260 ( .A1(n2612), .A2(n1201), .B1(n2610), .B2(n1220), .ZN(
        mult_x_18_n785) );
  OAI22D1BWP12T U2261 ( .A1(n2635), .A2(n1203), .B1(n1025), .B2(n1202), .ZN(
        mult_x_18_n916) );
  XNR2XD1BWP12T U2262 ( .A1(n2620), .A2(b[23]), .ZN(n1252) );
  OAI22D1BWP12T U2263 ( .A1(n2623), .A2(n1204), .B1(n1252), .B2(n2621), .ZN(
        mult_x_18_n929) );
  XNR2XD1BWP12T U2264 ( .A1(n2633), .A2(b[19]), .ZN(n1210) );
  OAI22D1BWP12T U2265 ( .A1(n2635), .A2(n1205), .B1(n1025), .B2(n1210), .ZN(
        mult_x_18_n904) );
  XNR2XD1BWP12T U2266 ( .A1(n2626), .A2(n2897), .ZN(n1207) );
  OAI22D1BWP12T U2267 ( .A1(n2629), .A2(n1206), .B1(n2627), .B2(n1207), .ZN(
        mult_x_18_n817) );
  XNR2XD1BWP12T U2268 ( .A1(n2626), .A2(b[11]), .ZN(n1260) );
  OAI22D1BWP12T U2269 ( .A1(n2629), .A2(n1207), .B1(n2627), .B2(n1260), .ZN(
        mult_x_18_n816) );
  OAI22D1BWP12T U2270 ( .A1(n2652), .A2(n1209), .B1(n2650), .B2(n1208), .ZN(
        mult_x_18_n962) );
  XNR2XD1BWP12T U2271 ( .A1(n2633), .A2(b[20]), .ZN(n1277) );
  OAI22D1BWP12T U2272 ( .A1(n2635), .A2(n1210), .B1(n1025), .B2(n1277), .ZN(
        mult_x_18_n903) );
  OAI22D1BWP12T U2273 ( .A1(n2646), .A2(n1212), .B1(n2644), .B2(n1211), .ZN(
        mult_x_18_n837) );
  OAI22D1BWP12T U2274 ( .A1(n2616), .A2(n1214), .B1(n2614), .B2(n1213), .ZN(
        mult_x_18_n889) );
  XNR2XD1BWP12T U2275 ( .A1(a[25]), .A2(n2639), .ZN(n1255) );
  OAI22D1BWP12T U2276 ( .A1(n2608), .A2(n1215), .B1(n2606), .B2(n1255), .ZN(
        mult_x_18_n750) );
  OAI22D1BWP12T U2277 ( .A1(n2646), .A2(n1217), .B1(n2644), .B2(n1216), .ZN(
        mult_x_18_n845) );
  IND2D1BWP12T U2278 ( .A1(n2231), .B1(n2626), .ZN(n1218) );
  OAI22D1BWP12T U2279 ( .A1(n2629), .A2(n1219), .B1(n2627), .B2(n1218), .ZN(
        mult_x_18_n721) );
  XNR2D1BWP12T U2280 ( .A1(n2609), .A2(n2605), .ZN(n1231) );
  XNR2XD1BWP12T U2281 ( .A1(n2609), .A2(b[9]), .ZN(n1283) );
  OAI22D1BWP12T U2282 ( .A1(n2612), .A2(n1231), .B1(n2610), .B2(n1283), .ZN(
        mult_x_18_n782) );
  XNR2D1BWP12T U2283 ( .A1(n2609), .A2(n2528), .ZN(n1232) );
  OAI22D1BWP12T U2284 ( .A1(n2612), .A2(n1220), .B1(n2610), .B2(n1232), .ZN(
        mult_x_18_n784) );
  XNR2D0BWP12T U2285 ( .A1(n2594), .A2(b[16]), .ZN(n1265) );
  OAI22D1BWP12T U2286 ( .A1(n2597), .A2(n1221), .B1(n1265), .B2(n2595), .ZN(
        mult_x_18_n855) );
  IND2XD0BWP12T U2287 ( .A1(n2231), .B1(n2609), .ZN(n1222) );
  OAI22D1BWP12T U2288 ( .A1(n2612), .A2(n1223), .B1(n2610), .B2(n1222), .ZN(
        mult_x_18_n719) );
  OAI22D1BWP12T U2289 ( .A1(n2601), .A2(n1225), .B1(n2599), .B2(n1224), .ZN(
        mult_x_18_n770) );
  OAI22D1BWP12T U2290 ( .A1(n2601), .A2(n1227), .B1(n2599), .B2(n1226), .ZN(
        mult_x_18_n774) );
  XNR2XD1BWP12T U2291 ( .A1(n2747), .A2(b[5]), .ZN(n1262) );
  OAI22D1BWP12T U2292 ( .A1(n2632), .A2(n1228), .B1(n1262), .B2(n2630), .ZN(
        mult_x_18_n758) );
  OAI22D1BWP12T U2293 ( .A1(n2646), .A2(n1230), .B1(n2644), .B2(n1229), .ZN(
        mult_x_18_n835) );
  OAI22D1BWP12T U2294 ( .A1(n2612), .A2(n1232), .B1(n2610), .B2(n1231), .ZN(
        mult_x_18_n783) );
  OAI22D1BWP12T U2295 ( .A1(n2638), .A2(n1234), .B1(n1233), .B2(n2636), .ZN(
        mult_x_18_n734) );
  XNR2XD1BWP12T U2296 ( .A1(a[25]), .A2(n2831), .ZN(n1254) );
  XNR2XD1BWP12T U2297 ( .A1(a[25]), .A2(n2868), .ZN(n1247) );
  OAI22D1BWP12T U2298 ( .A1(n2608), .A2(n1254), .B1(n2606), .B2(n1247), .ZN(
        mult_x_18_n748) );
  OAI22D1BWP12T U2299 ( .A1(n2652), .A2(n1236), .B1(n2650), .B2(n1235), .ZN(
        mult_x_18_n958) );
  OAI22D1BWP12T U2300 ( .A1(n2629), .A2(n1238), .B1(n2627), .B2(n1237), .ZN(
        mult_x_18_n821) );
  OAI22D1BWP12T U2301 ( .A1(n2616), .A2(n1240), .B1(n2614), .B2(n1239), .ZN(
        mult_x_18_n884) );
  OAI22D1BWP12T U2302 ( .A1(n2612), .A2(n1242), .B1(n2610), .B2(n1241), .ZN(
        mult_x_18_n789) );
  XNR2XD1BWP12T U2303 ( .A1(a[27]), .A2(n2477), .ZN(n1263) );
  XNR2XD1BWP12T U2304 ( .A1(a[27]), .A2(n2639), .ZN(n1274) );
  OAI22D1BWP12T U2305 ( .A1(n2619), .A2(n1263), .B1(n2617), .B2(n1274), .ZN(
        mult_x_18_n741) );
  XNR2XD1BWP12T U2306 ( .A1(n2725), .A2(n2605), .ZN(n1257) );
  OAI22D1BWP12T U2307 ( .A1(n2601), .A2(n1243), .B1(n2599), .B2(n1257), .ZN(
        mult_x_18_n768) );
  OAI22D1BWP12T U2308 ( .A1(n2623), .A2(n1245), .B1(n1244), .B2(n2621), .ZN(
        mult_x_18_n942) );
  OAI22D1BWP12T U2309 ( .A1(n2608), .A2(n1247), .B1(n2606), .B2(n1246), .ZN(
        mult_x_18_n747) );
  XNR2D0BWP12T U2310 ( .A1(n2643), .A2(b[15]), .ZN(n1250) );
  OAI22D1BWP12T U2311 ( .A1(n2646), .A2(n1248), .B1(n2644), .B2(n1250), .ZN(
        mult_x_18_n833) );
  XNR2D0BWP12T U2312 ( .A1(a[31]), .A2(n2231), .ZN(n1249) );
  XNR2D0BWP12T U2313 ( .A1(a[31]), .A2(n2477), .ZN(n2641) );
  OAI22D1BWP12T U2314 ( .A1(n2642), .A2(n1249), .B1(n2641), .B2(n2640), .ZN(
        mult_x_18_n730) );
  XNR2D0BWP12T U2315 ( .A1(n2643), .A2(b[16]), .ZN(n1272) );
  OAI22D1BWP12T U2316 ( .A1(n2646), .A2(n1250), .B1(n2644), .B2(n1272), .ZN(
        mult_x_18_n832) );
  XNR2XD1BWP12T U2317 ( .A1(n2679), .A2(n2598), .ZN(n1273) );
  OAI22D1BWP12T U2318 ( .A1(n2649), .A2(n1251), .B1(n1273), .B2(n2647), .ZN(
        mult_x_18_n796) );
  XNR2D0BWP12T U2319 ( .A1(n2620), .A2(b[24]), .ZN(n1270) );
  OAI22D1BWP12T U2320 ( .A1(n2623), .A2(n1252), .B1(n1270), .B2(n2621), .ZN(
        mult_x_18_n928) );
  XNR2D0BWP12T U2321 ( .A1(n2594), .A2(b[18]), .ZN(n1284) );
  OAI22D1BWP12T U2322 ( .A1(n2597), .A2(n1284), .B1(n1253), .B2(n2595), .ZN(
        mult_x_18_n852) );
  OAI22D1BWP12T U2323 ( .A1(n2608), .A2(n1255), .B1(n2606), .B2(n1254), .ZN(
        mult_x_18_n749) );
  OAI22D1BWP12T U2324 ( .A1(n2601), .A2(n1257), .B1(n2599), .B2(n1256), .ZN(
        mult_x_18_n767) );
  OAI22D1BWP12T U2325 ( .A1(n2616), .A2(n1259), .B1(n2614), .B2(n1258), .ZN(
        mult_x_18_n877) );
  XNR2XD1BWP12T U2326 ( .A1(n2626), .A2(n2598), .ZN(n1276) );
  OAI22D1BWP12T U2327 ( .A1(n2629), .A2(n1260), .B1(n2627), .B2(n1276), .ZN(
        mult_x_18_n815) );
  OAI22D1BWP12T U2328 ( .A1(n2632), .A2(n1262), .B1(n1261), .B2(n2630), .ZN(
        mult_x_18_n757) );
  XNR2XD1BWP12T U2329 ( .A1(a[27]), .A2(n2231), .ZN(n1264) );
  OAI22D1BWP12T U2330 ( .A1(n2619), .A2(n1264), .B1(n2617), .B2(n1263), .ZN(
        mult_x_18_n742) );
  XNR2D0BWP12T U2331 ( .A1(n2594), .A2(b[17]), .ZN(n1285) );
  OAI22D1BWP12T U2332 ( .A1(n2597), .A2(n1265), .B1(n1285), .B2(n2595), .ZN(
        mult_x_18_n854) );
  OAI22D1BWP12T U2333 ( .A1(n2646), .A2(n1267), .B1(n2644), .B2(n1266), .ZN(
        mult_x_18_n839) );
  XNR2D0BWP12T U2334 ( .A1(n2633), .A2(b[22]), .ZN(n1278) );
  OAI22D1BWP12T U2335 ( .A1(n2635), .A2(n1278), .B1(n1025), .B2(n1268), .ZN(
        mult_x_18_n900) );
  OAI22D1BWP12T U2336 ( .A1(n2623), .A2(n1270), .B1(n1269), .B2(n2621), .ZN(
        mult_x_18_n927) );
  OAI22D1BWP12T U2337 ( .A1(n2646), .A2(n1272), .B1(n2644), .B2(n1271), .ZN(
        mult_x_18_n831) );
  XNR2XD0BWP12T U2338 ( .A1(n2679), .A2(b[13]), .ZN(n1287) );
  OAI22D1BWP12T U2339 ( .A1(n2649), .A2(n1273), .B1(n1287), .B2(n2647), .ZN(
        mult_x_18_n795) );
  XNR2XD1BWP12T U2340 ( .A1(a[27]), .A2(n2831), .ZN(n1289) );
  OAI22D1BWP12T U2341 ( .A1(n2619), .A2(n1274), .B1(n2617), .B2(n1289), .ZN(
        mult_x_18_n740) );
  OAI22D1BWP12T U2342 ( .A1(n2629), .A2(n1276), .B1(n2627), .B2(n1275), .ZN(
        mult_x_18_n814) );
  XNR2D0BWP12T U2343 ( .A1(n2633), .A2(b[21]), .ZN(n1279) );
  OAI22D1BWP12T U2344 ( .A1(n2635), .A2(n1277), .B1(n1025), .B2(n1279), .ZN(
        mult_x_18_n902) );
  OAI22D1BWP12T U2345 ( .A1(n2635), .A2(n1279), .B1(n1025), .B2(n1278), .ZN(
        mult_x_18_n901) );
  OAI22D1BWP12T U2346 ( .A1(n2616), .A2(n1281), .B1(n2614), .B2(n1280), .ZN(
        mult_x_18_n875) );
  OAI22D1BWP12T U2347 ( .A1(n2612), .A2(n1283), .B1(n2610), .B2(n1282), .ZN(
        mult_x_18_n781) );
  OAI22D1BWP12T U2348 ( .A1(n2597), .A2(n1285), .B1(n1284), .B2(n2595), .ZN(
        mult_x_18_n853) );
  OAI22D1BWP12T U2349 ( .A1(n2649), .A2(n1287), .B1(n1286), .B2(n2647), .ZN(
        mult_x_18_n794) );
  OAI22D1BWP12T U2350 ( .A1(n2619), .A2(n1289), .B1(n2617), .B2(n1288), .ZN(
        mult_x_18_n739) );
  OAI22D1BWP12T U2351 ( .A1(n2604), .A2(n1291), .B1(n1290), .B2(n2603), .ZN(
        n1295) );
  OAI22D1BWP12T U2352 ( .A1(n2623), .A2(n1293), .B1(n1292), .B2(n2621), .ZN(
        n1294) );
  OAI22D1BWP12T U2353 ( .A1(n2604), .A2(n1297), .B1(n1296), .B2(n2603), .ZN(
        n1301) );
  OAI22D1BWP12T U2354 ( .A1(n2649), .A2(n1299), .B1(n1298), .B2(n2647), .ZN(
        n1300) );
  HA1D1BWP12T U2355 ( .A(n1301), .B(n1300), .CO(mult_x_18_n567), .S(
        mult_x_18_n568) );
  OAI22D1BWP12T U2356 ( .A1(n2604), .A2(n1303), .B1(n1302), .B2(n2603), .ZN(
        n1307) );
  CKND0BWP12T U2357 ( .I(n2679), .ZN(n1305) );
  IND2XD1BWP12T U2358 ( .A1(n2231), .B1(n2679), .ZN(n1304) );
  OAI22D1BWP12T U2359 ( .A1(n2649), .A2(n1305), .B1(n2647), .B2(n1304), .ZN(
        n1306) );
  OAI22D1BWP12T U2360 ( .A1(n2604), .A2(n1309), .B1(n1308), .B2(n2603), .ZN(
        n1313) );
  IND2D1BWP12T U2361 ( .A1(n2231), .B1(n2594), .ZN(n1310) );
  OAI22D1BWP12T U2362 ( .A1(n2597), .A2(n1311), .B1(n2595), .B2(n1310), .ZN(
        n1312) );
  HA1D0BWP12T U2363 ( .A(n1315), .B(n1314), .CO(mult_x_18_n707), .S(n448) );
  OAI22D1BWP12T U2364 ( .A1(n2604), .A2(n1325), .B1(n1324), .B2(n2603), .ZN(
        n1329) );
  OAI22D1BWP12T U2365 ( .A1(n2597), .A2(n1327), .B1(n1326), .B2(n2595), .ZN(
        n1328) );
  HA1D1BWP12T U2366 ( .A(n1329), .B(n1328), .CO(mult_x_18_n661), .S(
        mult_x_18_n662) );
  OAI22D1BWP12T U2367 ( .A1(n2604), .A2(n1331), .B1(n1330), .B2(n2603), .ZN(
        n1335) );
  OAI22D1BWP12T U2368 ( .A1(n2623), .A2(n1333), .B1(n1332), .B2(n2621), .ZN(
        n1334) );
  OAI22D1BWP12T U2369 ( .A1(n2604), .A2(n1337), .B1(n1336), .B2(n2603), .ZN(
        n1341) );
  OAI22D1BWP12T U2370 ( .A1(n2597), .A2(n1339), .B1(n1338), .B2(n2595), .ZN(
        n1340) );
  OAI22D1BWP12T U2371 ( .A1(n2604), .A2(n1343), .B1(n1342), .B2(n2603), .ZN(
        n1347) );
  OAI22D1BWP12T U2372 ( .A1(n2649), .A2(n1345), .B1(n1344), .B2(n2647), .ZN(
        n1346) );
  FA1D1BWP12T U2373 ( .A(mult_x_18_n406), .B(mult_x_18_n386), .CI(n1348), .CO(
        n2593), .S(n1740) );
  INVD1BWP12T U2374 ( .I(n1740), .ZN(n1386) );
  FA1D2BWP12T U2375 ( .A(a[30]), .B(n2291), .CI(n1349), .CO(n2660), .S(n2462)
         );
  INVD1BWP12T U2376 ( .I(n1805), .ZN(n1381) );
  HA1D0BWP12T U2377 ( .A(n2251), .B(n1351), .CO(n2665), .S(n1844) );
  CKND2D1BWP12T U2378 ( .A1(n2573), .A2(n2008), .ZN(n1357) );
  MUX2XD0BWP12T U2379 ( .I0(a[24]), .I1(n2747), .S(n2231), .Z(n1469) );
  INVD1BWP12T U2380 ( .I(n1469), .ZN(n2171) );
  MUX2NXD0BWP12T U2381 ( .I0(a[28]), .I1(a[27]), .S(n2231), .ZN(n1474) );
  TPOAI22D0BWP12T U2382 ( .A1(n1941), .A2(n2171), .B1(n1501), .B2(n1474), .ZN(
        n1353) );
  MUX2NXD0BWP12T U2383 ( .I0(n2779), .I1(n2253), .S(n2231), .ZN(n1470) );
  INVD1BWP12T U2384 ( .I(n1470), .ZN(n2172) );
  TPNR2D0BWP12T U2385 ( .A1(n1959), .A2(n2172), .ZN(n1352) );
  AOI211D0BWP12T U2386 ( .A1(a[29]), .A2(n2002), .B(n1353), .C(n1352), .ZN(
        n1354) );
  OA222D1BWP12T U2387 ( .A1(n2022), .A2(n1356), .B1(n2023), .B2(n1355), .C1(
        n2025), .C2(n1354), .Z(n2037) );
  AOI21D1BWP12T U2388 ( .A1(n1357), .A2(n2037), .B(n2964), .ZN(n1377) );
  ND2D1BWP12T U2389 ( .A1(n2932), .A2(n1920), .ZN(n1530) );
  AOI22D0BWP12T U2390 ( .A1(n2169), .A2(n2171), .B1(n2172), .B2(n2166), .ZN(
        n1359) );
  CKND2D0BWP12T U2391 ( .A1(n1474), .A2(n2170), .ZN(n1358) );
  OAI211D0BWP12T U2392 ( .A1(a[29]), .A2(n1548), .B(n1359), .C(n1358), .ZN(
        n1361) );
  NR2D0BWP12T U2393 ( .A1(n1360), .A2(a[30]), .ZN(n1814) );
  AOI211D0BWP12T U2394 ( .A1(n2769), .A2(n1361), .B(n2174), .C(n1814), .ZN(
        n1366) );
  CKND0BWP12T U2395 ( .I(n2159), .ZN(n1364) );
  AOI22D1BWP12T U2396 ( .A1(n1364), .A2(n1363), .B1(n1362), .B2(n2155), .ZN(
        n1365) );
  OA211D0BWP12T U2397 ( .A1(n2581), .A2(n2080), .B(n1366), .C(n1365), .Z(n2211) );
  CKND2D1BWP12T U2398 ( .A1(n2211), .A2(n2786), .ZN(n1375) );
  INVD1BWP12T U2399 ( .I(n2066), .ZN(n1372) );
  CKND0BWP12T U2400 ( .I(b[30]), .ZN(n2291) );
  TPNR2D0BWP12T U2401 ( .A1(n2291), .A2(n2951), .ZN(n1367) );
  AOI211XD0BWP12T U2402 ( .A1(n2291), .A2(n2948), .B(n1367), .C(n2825), .ZN(
        n1370) );
  OAI21D0BWP12T U2403 ( .A1(a[30]), .A2(n2944), .B(n2949), .ZN(n1368) );
  AOI22D0BWP12T U2404 ( .A1(n2947), .A2(n2251), .B1(n1368), .B2(b[30]), .ZN(
        n1369) );
  OAI21D0BWP12T U2405 ( .A1(n1370), .A2(n2251), .B(n1369), .ZN(n1371) );
  AOI211XD0BWP12T U2406 ( .A1(n1373), .A2(n1372), .B(n2807), .C(n1371), .ZN(
        n1374) );
  OAI211D1BWP12T U2407 ( .A1(n1849), .A2(n1530), .B(n1375), .C(n1374), .ZN(
        n1376) );
  AOI211D1BWP12T U2408 ( .A1(n1844), .A2(n2940), .B(n1377), .C(n1376), .ZN(
        n1380) );
  FA1D1BWP12T U2409 ( .A(a[30]), .B(b[30]), .CI(n1378), .CO(n2916), .S(n2397)
         );
  OAI211D2BWP12T U2410 ( .A1(n2814), .A2(n1381), .B(n1380), .C(n1379), .ZN(
        n1382) );
  TPAOI21D2BWP12T U2411 ( .A1(n2866), .A2(n2462), .B(n1382), .ZN(n1385) );
  FA1D1BWP12T U2412 ( .A(a[30]), .B(n2291), .CI(n1383), .CO(n2658), .S(n1657)
         );
  ND2D1BWP12T U2413 ( .A1(n1657), .A2(n2855), .ZN(n1384) );
  OAI211D4BWP12T U2414 ( .A1(n2822), .A2(n1386), .B(n1385), .C(n1384), .ZN(
        result[30]) );
  INVD1P75BWP12T U2415 ( .I(n1387), .ZN(n1678) );
  INVD1BWP12T U2416 ( .I(n1677), .ZN(n1388) );
  CKND2D1BWP12T U2417 ( .A1(n1388), .A2(n1676), .ZN(n1389) );
  XOR2D1BWP12T U2418 ( .A1(n1678), .A2(n1389), .Z(n1718) );
  INVD1BWP12T U2419 ( .I(n2866), .ZN(n2973) );
  INVD1BWP12T U2420 ( .I(n1396), .ZN(n1418) );
  AOI22D0BWP12T U2421 ( .A1(n1999), .A2(n2117), .B1(n2118), .B2(n1945), .ZN(
        n1402) );
  NR2D0BWP12T U2422 ( .A1(n1398), .A2(n1413), .ZN(n1399) );
  AOI22D0BWP12T U2423 ( .A1(n2002), .A2(n2120), .B1(n1400), .B2(n1399), .ZN(
        n1401) );
  ND2D1BWP12T U2424 ( .A1(n1402), .A2(n1401), .ZN(n2018) );
  CKND2D1BWP12T U2425 ( .A1(n1547), .A2(n471), .ZN(n2153) );
  INVD1BWP12T U2426 ( .I(n2153), .ZN(n1416) );
  CKND2D0BWP12T U2427 ( .A1(n2002), .A2(n1460), .ZN(n1404) );
  AOI22D0BWP12T U2428 ( .A1(n2000), .A2(n2121), .B1(n2001), .B2(n2124), .ZN(
        n1403) );
  OAI211D0BWP12T U2429 ( .A1(n1956), .A2(n1959), .B(n1404), .C(n1403), .ZN(
        n2011) );
  INVD1BWP12T U2430 ( .I(n1405), .ZN(n1830) );
  XOR2XD1BWP12T U2431 ( .A1(n1830), .A2(a[16]), .Z(n1831) );
  OAI22D0BWP12T U2432 ( .A1(n1848), .A2(n1933), .B1(n1903), .B2(n1926), .ZN(
        n1407) );
  OAI22D0BWP12T U2433 ( .A1(n1856), .A2(n1930), .B1(n1912), .B2(n2052), .ZN(
        n1406) );
  NR2D1BWP12T U2434 ( .A1(n1407), .A2(n1406), .ZN(n2063) );
  INVD1BWP12T U2435 ( .I(n2063), .ZN(n1542) );
  TPND2D0BWP12T U2436 ( .A1(n2675), .A2(n2718), .ZN(n2960) );
  AOI22D0BWP12T U2437 ( .A1(n2169), .A2(n1408), .B1(n1956), .B2(n2166), .ZN(
        n1410) );
  AOI22D0BWP12T U2438 ( .A1(n2173), .A2(n2127), .B1(n1466), .B2(n2170), .ZN(
        n1409) );
  CKND2D1BWP12T U2439 ( .A1(n1410), .A2(n1409), .ZN(n2156) );
  OAI22D0BWP12T U2440 ( .A1(n2118), .A2(n2128), .B1(n2120), .B2(n2126), .ZN(
        n1412) );
  NR2XD0BWP12T U2441 ( .A1(n2119), .A2(n2117), .ZN(n1411) );
  AOI211D1BWP12T U2442 ( .A1(n2169), .A2(n1413), .B(n1412), .C(n1411), .ZN(
        n2160) );
  CKND0BWP12T U2443 ( .I(n2160), .ZN(n1414) );
  AOI22D0BWP12T U2444 ( .A1(n2769), .A2(n2156), .B1(n1414), .B2(n2831), .ZN(
        n1415) );
  OAI211D1BWP12T U2445 ( .A1(n1416), .A2(n2870), .B(n1415), .C(n2187), .ZN(
        n2207) );
  INVD1BWP12T U2446 ( .I(n2807), .ZN(n2682) );
  AOI21D1BWP12T U2447 ( .A1(n2855), .A2(n1649), .B(n1420), .ZN(n1421) );
  IOA21D2BWP12T U2448 ( .A1(n1718), .A2(n2977), .B(n1421), .ZN(result[16]) );
  ND2D1BWP12T U2449 ( .A1(n1426), .A2(n1425), .ZN(n1427) );
  XOR2XD1BWP12T U2450 ( .A1(n1428), .A2(n1427), .Z(n1715) );
  ND2XD0BWP12T U2451 ( .A1(n1430), .A2(n1429), .ZN(n1431) );
  XNR2D1BWP12T U2452 ( .A1(n1432), .A2(n1431), .ZN(n1643) );
  INVD1BWP12T U2453 ( .I(n2454), .ZN(n1451) );
  CKND2D0BWP12T U2454 ( .A1(n1438), .A2(n1437), .ZN(n1439) );
  XNR2D1BWP12T U2455 ( .A1(n1440), .A2(n1439), .ZN(n2386) );
  AOI22D1BWP12T U2456 ( .A1(n2858), .A2(n1790), .B1(n2386), .B2(n2967), .ZN(
        n1450) );
  MAOI22D0BWP12T U2457 ( .A1(n2033), .A2(n2526), .B1(n1986), .B2(n2025), .ZN(
        n1949) );
  NR2D1BWP12T U2458 ( .A1(n1443), .A2(n2894), .ZN(n2842) );
  OAI22D0BWP12T U2459 ( .A1(n1870), .A2(n2240), .B1(n1869), .B2(n2705), .ZN(
        n1445) );
  OAI22D0BWP12T U2460 ( .A1(n1872), .A2(n2683), .B1(n1871), .B2(n2235), .ZN(
        n1444) );
  NR2D1BWP12T U2461 ( .A1(n1445), .A2(n1444), .ZN(n1883) );
  CKND2D0BWP12T U2462 ( .A1(n1883), .A2(n471), .ZN(n1447) );
  ND2XD0BWP12T U2463 ( .A1(n1881), .A2(n2639), .ZN(n1446) );
  ND2D1BWP12T U2464 ( .A1(n1447), .A2(n1446), .ZN(n1924) );
  INVD1BWP12T U2465 ( .I(n1852), .ZN(n2078) );
  INVD1BWP12T U2466 ( .I(n2155), .ZN(n2200) );
  OAI22D1BWP12T U2467 ( .A1(n2202), .A2(n1924), .B1(n2078), .B2(n2200), .ZN(
        n1884) );
  NR2D0BWP12T U2468 ( .A1(n1850), .A2(n2870), .ZN(n1886) );
  TPAOI21D0BWP12T U2469 ( .A1(n1884), .A2(n2115), .B(n2783), .ZN(n2070) );
  INVD1BWP12T U2470 ( .I(n2179), .ZN(n2534) );
  CKND2D0BWP12T U2471 ( .A1(n2534), .A2(n2831), .ZN(n1448) );
  OAI211D1BWP12T U2472 ( .A1(n2831), .A2(n2176), .B(n1448), .C(n2198), .ZN(
        n2206) );
  OAI211D1BWP12T U2473 ( .A1(n2973), .A2(n1451), .B(n1450), .C(n1449), .ZN(
        n1452) );
  AOI21D1BWP12T U2474 ( .A1(n2855), .A2(n1643), .B(n1452), .ZN(n1453) );
  IOA21D1BWP12T U2475 ( .A1(n1715), .A2(n2977), .B(n1453), .ZN(result[15]) );
  FA1D1BWP12T U2476 ( .A(mult_x_18_n448), .B(mult_x_18_n429), .CI(n1454), .CO(
        n1496), .S(n1738) );
  INVD1BWP12T U2477 ( .I(n1738), .ZN(n1495) );
  FA1D0BWP12T U2478 ( .A(a[28]), .B(n2290), .CI(n1455), .CO(n1497), .S(n2459)
         );
  ND2D1BWP12T U2479 ( .A1(n1803), .A2(n2858), .ZN(n1490) );
  FA1D2BWP12T U2480 ( .A(a[28]), .B(b[28]), .CI(n1457), .CO(n1499), .S(n2393)
         );
  ND2D1BWP12T U2481 ( .A1(n2393), .A2(n2967), .ZN(n1489) );
  OAI22D0BWP12T U2482 ( .A1(n1501), .A2(n2149), .B1(n1941), .B2(n1466), .ZN(
        n1459) );
  NR2D0BWP12T U2483 ( .A1(n1940), .A2(n2168), .ZN(n1458) );
  RCAOI211D0BWP12T U2484 ( .A1(n1460), .A2(n1999), .B(n1459), .C(n1458), .ZN(
        n2030) );
  CKND2D0BWP12T U2485 ( .A1(n1999), .A2(n1469), .ZN(n1462) );
  AOI22D0BWP12T U2486 ( .A1(n2001), .A2(n1470), .B1(n2000), .B2(n1471), .ZN(
        n1461) );
  OAI211D0BWP12T U2487 ( .A1(n1474), .A2(n1940), .B(n1462), .C(n1461), .ZN(
        n1463) );
  AOI22D0BWP12T U2488 ( .A1(n2031), .A2(n1463), .B1(n2036), .B2(n2008), .ZN(
        n1465) );
  CKND2D0BWP12T U2489 ( .A1(n2034), .A2(n2035), .ZN(n1464) );
  OAI211D0BWP12T U2490 ( .A1(n2030), .A2(n2023), .B(n1465), .C(n1464), .ZN(
        n1951) );
  AOI22D0BWP12T U2491 ( .A1(n2173), .A2(n2168), .B1(n2149), .B2(n2170), .ZN(
        n1468) );
  AOI22D0BWP12T U2492 ( .A1(n2169), .A2(n1466), .B1(n2127), .B2(n2166), .ZN(
        n1467) );
  ND2D1BWP12T U2493 ( .A1(n1468), .A2(n1467), .ZN(n2182) );
  OAI22D0BWP12T U2494 ( .A1(n1470), .A2(n2128), .B1(n1469), .B2(n2119), .ZN(
        n1473) );
  NR2D0BWP12T U2495 ( .A1(n1471), .A2(n2116), .ZN(n1472) );
  AOI211D0BWP12T U2496 ( .A1(n2173), .A2(n1474), .B(n1473), .C(n1472), .ZN(
        n1475) );
  OAI21D0BWP12T U2497 ( .A1(n1475), .A2(n2202), .B(n2115), .ZN(n1477) );
  OAI22D0BWP12T U2498 ( .A1(n2180), .A2(n2159), .B1(n2875), .B2(n2080), .ZN(
        n1476) );
  AOI211XD0BWP12T U2499 ( .A1(n2155), .A2(n2182), .B(n1477), .C(n1476), .ZN(
        n2133) );
  MOAI22D0BWP12T U2500 ( .A1(n1856), .A2(n1530), .B1(n2133), .B2(n2786), .ZN(
        n1485) );
  CKND0BWP12T U2501 ( .I(b[28]), .ZN(n2290) );
  TPNR2D0BWP12T U2502 ( .A1(n2290), .A2(n2951), .ZN(n1478) );
  AOI211XD0BWP12T U2503 ( .A1(n2290), .A2(n2948), .B(n1478), .C(n2825), .ZN(
        n1483) );
  AOI21D0BWP12T U2504 ( .A1(n1479), .A2(n2094), .B(n2095), .ZN(n2087) );
  CKND2D1BWP12T U2505 ( .A1(n2087), .A2(n2905), .ZN(n1482) );
  OAI21D0BWP12T U2506 ( .A1(a[28]), .A2(n2944), .B(n2949), .ZN(n1480) );
  AOI22D0BWP12T U2507 ( .A1(n2947), .A2(n2249), .B1(n1480), .B2(b[28]), .ZN(
        n1481) );
  OAI211D1BWP12T U2508 ( .A1(n1483), .A2(n2249), .B(n1482), .C(n1481), .ZN(
        n1484) );
  RCAOI211D0BWP12T U2509 ( .A1(n2894), .A2(n1951), .B(n1485), .C(n1484), .ZN(
        n1488) );
  HA1D1BWP12T U2510 ( .A(n2249), .B(n1486), .CO(n1500), .S(n1841) );
  ND2D1BWP12T U2511 ( .A1(n1841), .A2(n2940), .ZN(n1487) );
  ND4D1BWP12T U2512 ( .A1(n1490), .A2(n1489), .A3(n1488), .A4(n1487), .ZN(
        n1491) );
  AOI21D1BWP12T U2513 ( .A1(n2866), .A2(n2459), .B(n1491), .ZN(n1494) );
  FA1D1BWP12T U2514 ( .A(a[28]), .B(n2290), .CI(n1492), .CO(n1538), .S(n1659)
         );
  ND2D1BWP12T U2515 ( .A1(n1659), .A2(n2855), .ZN(n1493) );
  OAI211D1BWP12T U2516 ( .A1(n2822), .A2(n1495), .B(n1494), .C(n1493), .ZN(
        result[28]) );
  FA1D1BWP12T U2517 ( .A(mult_x_18_n428), .B(mult_x_18_n407), .CI(n1496), .CO(
        n1348), .S(n1739) );
  INVD1BWP12T U2518 ( .I(n1739), .ZN(n1541) );
  FA1D2BWP12T U2519 ( .A(a[29]), .B(b[29]), .CI(n1499), .CO(n1378), .S(n2396)
         );
  ND2D1BWP12T U2520 ( .A1(n2396), .A2(n2967), .ZN(n1535) );
  HA1D1BWP12T U2521 ( .A(n2248), .B(n1500), .CO(n1351), .S(n1843) );
  OAI22D0BWP12T U2522 ( .A1(n1501), .A2(n2140), .B1(n1941), .B2(n2142), .ZN(
        n1503) );
  NR2D0BWP12T U2523 ( .A1(n1959), .A2(n2141), .ZN(n1502) );
  AOI211D0BWP12T U2524 ( .A1(n1517), .A2(n2002), .B(n1503), .C(n1502), .ZN(
        n1504) );
  OAI22D0BWP12T U2525 ( .A1(n1505), .A2(n2022), .B1(n1504), .B2(n2025), .ZN(
        n1510) );
  AOI22D0BWP12T U2526 ( .A1(n2000), .A2(n1512), .B1(n2001), .B2(n1511), .ZN(
        n1507) );
  CKND2D0BWP12T U2527 ( .A1(n2002), .A2(n2143), .ZN(n1506) );
  OAI211D0BWP12T U2528 ( .A1(n1508), .A2(n1959), .B(n1507), .C(n1506), .ZN(
        n2013) );
  NR2D0BWP12T U2529 ( .A1(n2013), .A2(n2023), .ZN(n1509) );
  RCAOI211D0BWP12T U2530 ( .A1(n2008), .A2(n1947), .B(n1510), .C(n1509), .ZN(
        n2039) );
  AOI22D0BWP12T U2531 ( .A1(n1511), .A2(n2170), .B1(n2173), .B2(n2143), .ZN(
        n1515) );
  AOI22D0BWP12T U2532 ( .A1(n2166), .A2(n1513), .B1(n1512), .B2(n2169), .ZN(
        n1514) );
  ND2D1BWP12T U2533 ( .A1(n1515), .A2(n1514), .ZN(n2185) );
  OAI22D0BWP12T U2534 ( .A1(n1517), .A2(n2126), .B1(n1516), .B2(n2128), .ZN(
        n1520) );
  NR2D0BWP12T U2535 ( .A1(n1518), .A2(n2119), .ZN(n1519) );
  AOI211D0BWP12T U2536 ( .A1(n2169), .A2(n2142), .B(n1520), .C(n1519), .ZN(
        n1521) );
  OAI21D0BWP12T U2537 ( .A1(n1521), .A2(n2202), .B(n2115), .ZN(n1523) );
  OAI22D0BWP12T U2538 ( .A1(n2189), .A2(n2159), .B1(n2080), .B2(n2184), .ZN(
        n1522) );
  AOI211D1BWP12T U2539 ( .A1(n2155), .A2(n2185), .B(n1523), .C(n1522), .ZN(
        n2134) );
  AOI21D1BWP12T U2540 ( .A1(n1524), .A2(n2956), .B(n2095), .ZN(n2088) );
  AOI22D1BWP12T U2541 ( .A1(n2134), .A2(n2786), .B1(n2088), .B2(n2905), .ZN(
        n1532) );
  OAI21D0BWP12T U2542 ( .A1(a[29]), .A2(n2944), .B(n2949), .ZN(n1525) );
  AOI22D0BWP12T U2543 ( .A1(n2947), .A2(n2248), .B1(n1525), .B2(b[29]), .ZN(
        n1529) );
  CKND0BWP12T U2544 ( .I(b[29]), .ZN(n2292) );
  TPND2D0BWP12T U2545 ( .A1(n2292), .A2(n2948), .ZN(n1526) );
  OAI211D0BWP12T U2546 ( .A1(n2292), .A2(n2951), .B(n1526), .C(n2949), .ZN(
        n1527) );
  ND2XD0BWP12T U2547 ( .A1(n1527), .A2(a[29]), .ZN(n1528) );
  OA211D1BWP12T U2548 ( .A1(n1851), .A2(n1530), .B(n1529), .C(n1528), .Z(n1531) );
  OAI211D1BWP12T U2549 ( .A1(n2039), .A2(n2964), .B(n1532), .C(n1531), .ZN(
        n1533) );
  AOI21D1BWP12T U2550 ( .A1(n1843), .A2(n2940), .B(n1533), .ZN(n1534) );
  OAI211D1BWP12T U2551 ( .A1(n1536), .A2(n2814), .B(n1535), .C(n1534), .ZN(
        n1537) );
  AOI21D1BWP12T U2552 ( .A1(n2866), .A2(n2461), .B(n1537), .ZN(n1540) );
  FA1D1BWP12T U2553 ( .A(a[29]), .B(n2292), .CI(n1538), .CO(n1383), .S(n1660)
         );
  ND2D1BWP12T U2554 ( .A1(n1660), .A2(n2855), .ZN(n1539) );
  OAI211D1BWP12T U2555 ( .A1(n2822), .A2(n1541), .B(n1540), .C(n1539), .ZN(
        result[29]) );
  ND2D1BWP12T U2556 ( .A1(n1542), .A2(n2868), .ZN(n1975) );
  INVD1BWP12T U2557 ( .I(n1975), .ZN(n1555) );
  OAI22D0BWP12T U2558 ( .A1(n1870), .A2(n2869), .B1(n1869), .B2(n2532), .ZN(
        n1544) );
  OAI22D1BWP12T U2559 ( .A1(n1872), .A2(n2578), .B1(n1871), .B2(n2257), .ZN(
        n1543) );
  NR2D1BWP12T U2560 ( .A1(n1544), .A2(n1543), .ZN(n1913) );
  OAI22D0BWP12T U2561 ( .A1(n1914), .A2(n1930), .B1(n1913), .B2(n1926), .ZN(
        n1554) );
  OAI22D0BWP12T U2562 ( .A1(n1870), .A2(a[8]), .B1(n2594), .B2(n1869), .ZN(
        n1546) );
  OAI22D0BWP12T U2563 ( .A1(n2301), .A2(n1871), .B1(n1872), .B2(n2900), .ZN(
        n1545) );
  NR2D1BWP12T U2564 ( .A1(n1546), .A2(n1545), .ZN(n1910) );
  INVD1BWP12T U2565 ( .I(n1910), .ZN(n1904) );
  ND2D1BWP12T U2566 ( .A1(n1547), .A2(n1920), .ZN(n2194) );
  TPOAI21D0BWP12T U2567 ( .A1(n1904), .A2(n1933), .B(n2194), .ZN(n1553) );
  INVD1BWP12T U2568 ( .I(n1548), .ZN(n1892) );
  CKND2D0BWP12T U2569 ( .A1(n1892), .A2(n2482), .ZN(n1551) );
  CKND2D0BWP12T U2570 ( .A1(n1893), .A2(n2830), .ZN(n1550) );
  CKND2D0BWP12T U2571 ( .A1(n1894), .A2(n2303), .ZN(n1549) );
  TPAOI31D0BWP12T U2572 ( .A1(n1551), .A2(n1550), .A3(n1549), .B(n2831), .ZN(
        n1552) );
  NR3D1BWP12T U2573 ( .A1(n1554), .A2(n1553), .A3(n1552), .ZN(n1974) );
  INVD1BWP12T U2574 ( .I(n1974), .ZN(n1562) );
  AOI22D1BWP12T U2575 ( .A1(n2115), .A2(n1555), .B1(n1562), .B2(n2198), .ZN(
        n2061) );
  XNR2D0BWP12T U2576 ( .A1(n1558), .A2(n2302), .ZN(n2425) );
  INR2D0BWP12T U2577 ( .A1(n2231), .B1(n2603), .ZN(n1711) );
  CKND0BWP12T U2578 ( .I(n2951), .ZN(n2478) );
  INVD0BWP12T U2579 ( .I(n1559), .ZN(n1561) );
  INVD1BWP12T U2580 ( .I(n2061), .ZN(n1922) );
  INVD1BWP12T U2581 ( .I(n1563), .ZN(n1565) );
  ND2D1BWP12T U2582 ( .A1(n1565), .A2(n1564), .ZN(n1567) );
  XOR2XD1BWP12T U2583 ( .A1(n1567), .A2(n1566), .Z(n1712) );
  OAI22D1BWP12T U2584 ( .A1(n1870), .A2(n2257), .B1(n1869), .B2(n2550), .ZN(
        n1569) );
  OAI22D1BWP12T U2585 ( .A1(n1872), .A2(n2532), .B1(n1871), .B2(n2578), .ZN(
        n1568) );
  NR2D1BWP12T U2586 ( .A1(n1569), .A2(n1568), .ZN(n1897) );
  NR2D1BWP12T U2587 ( .A1(n1977), .A2(n2174), .ZN(n1906) );
  OAI22D1BWP12T U2588 ( .A1(n1861), .A2(n2052), .B1(n1570), .B2(n1926), .ZN(
        n1574) );
  TPAOI21D0BWP12T U2589 ( .A1(n2831), .A2(n1571), .B(n1574), .ZN(n2719) );
  ND2D1BWP12T U2590 ( .A1(n2719), .A2(n2868), .ZN(n1572) );
  RCAOI21D0BWP12T U2591 ( .A1(n1906), .A2(n1572), .B(n2058), .ZN(n2103) );
  INVD1BWP12T U2592 ( .I(n1573), .ZN(n1835) );
  INVD1BWP12T U2593 ( .I(n2535), .ZN(n2874) );
  INVD1BWP12T U2594 ( .I(n1859), .ZN(n2720) );
  AOI21D0BWP12T U2595 ( .A1(n2720), .A2(n2894), .B(n2893), .ZN(n1578) );
  INVD1BWP12T U2596 ( .I(n1575), .ZN(n2374) );
  NR2D0BWP12T U2597 ( .A1(n2284), .A2(n2951), .ZN(n1579) );
  AOI211D1BWP12T U2598 ( .A1(n2284), .A2(n2948), .B(n1579), .C(n2825), .ZN(
        n1583) );
  NR2D1BWP12T U2599 ( .A1(n2025), .A2(n2964), .ZN(n2828) );
  CKND2D0BWP12T U2600 ( .A1(n1947), .A2(n2828), .ZN(n1582) );
  OAI21D0BWP12T U2601 ( .A1(n2620), .A2(n2944), .B(n2949), .ZN(n1580) );
  AOI22D0BWP12T U2602 ( .A1(n2947), .A2(n2257), .B1(n1580), .B2(b[5]), .ZN(
        n1581) );
  INVD1BWP12T U2603 ( .I(n1584), .ZN(n1786) );
  INVD0BWP12T U2604 ( .I(n1782), .ZN(n1585) );
  NR2XD0BWP12T U2605 ( .A1(n2720), .A2(n2870), .ZN(n1978) );
  INVD1BWP12T U2606 ( .I(n1586), .ZN(n1629) );
  INVD1BWP12T U2607 ( .I(n1625), .ZN(n1587) );
  INVD1BWP12T U2608 ( .I(n1588), .ZN(n2441) );
  FA1D1BWP12T U2609 ( .A(a[26]), .B(n2774), .CI(n1591), .CO(n1654), .S(n2797)
         );
  FA1D1BWP12T U2610 ( .A(n2747), .B(n2406), .CI(n1592), .CO(n1652), .S(n2763)
         );
  FA1D0BWP12T U2611 ( .A(n2410), .B(a[20]), .CI(n1593), .CO(n1650), .S(n2937)
         );
  INVD1BWP12T U2612 ( .I(n1601), .ZN(n1603) );
  ND2D1BWP12T U2613 ( .A1(n1603), .A2(n1602), .ZN(n1605) );
  XOR2XD1BWP12T U2614 ( .A1(n1605), .A2(n1604), .Z(n2476) );
  INVD1BWP12T U2615 ( .I(n1615), .ZN(n1609) );
  AOI21D1BWP12T U2616 ( .A1(n1629), .A2(n2431), .B(n1609), .ZN(n1614) );
  INVD0BWP12T U2617 ( .I(n1610), .ZN(n1612) );
  CKND2D1BWP12T U2618 ( .A1(n1612), .A2(n1611), .ZN(n1613) );
  XOR2XD1BWP12T U2619 ( .A1(n1614), .A2(n1613), .Z(n2856) );
  ND2D1BWP12T U2620 ( .A1(n2431), .A2(n1615), .ZN(n1616) );
  XNR2D1BWP12T U2621 ( .A1(n1629), .A2(n1616), .ZN(n2824) );
  CKND0BWP12T U2622 ( .I(n1621), .ZN(n1622) );
  NR2XD0BWP12T U2623 ( .A1(n1622), .A2(n1625), .ZN(n1628) );
  CKND0BWP12T U2624 ( .I(n1623), .ZN(n1626) );
  OAI21D1BWP12T U2625 ( .A1(n1626), .A2(n1625), .B(n1624), .ZN(n1627) );
  AOI21D1BWP12T U2626 ( .A1(n1629), .A2(n1628), .B(n1627), .ZN(n1633) );
  ND2D1BWP12T U2627 ( .A1(n2419), .A2(n1631), .ZN(n1632) );
  XOR2XD1BWP12T U2628 ( .A1(n1633), .A2(n1632), .Z(n2570) );
  INVD0BWP12T U2629 ( .I(n1637), .ZN(n1638) );
  FA1D0BWP12T U2630 ( .A(n2725), .B(n2408), .CI(n1650), .CO(n769), .S(n2737)
         );
  FA1D1BWP12T U2631 ( .A(n2952), .B(a[24]), .CI(n1652), .CO(n732), .S(n2975)
         );
  FA1D1BWP12T U2632 ( .A(a[27]), .B(n2805), .CI(n1654), .CO(n1492), .S(n2818)
         );
  OR4D0BWP12T U2633 ( .A1(n2797), .A2(n1656), .A3(n1655), .A4(n2818), .Z(n1658) );
  OR4D0BWP12T U2634 ( .A1(n1660), .A2(n1659), .A3(n1658), .A4(n1657), .Z(n2470) );
  AOI21D1BWP12T U2635 ( .A1(n1670), .A2(n1669), .B(n1668), .ZN(n1673) );
  CKND2D1BWP12T U2636 ( .A1(n425), .A2(n1671), .ZN(n1672) );
  XOR2XD1BWP12T U2637 ( .A1(n1673), .A2(n1672), .Z(n2740) );
  OAI21D1BWP12T U2638 ( .A1(n1678), .A2(n1677), .B(n1676), .ZN(n1683) );
  INVD1BWP12T U2639 ( .I(n1679), .ZN(n1681) );
  ND2D1BWP12T U2640 ( .A1(n1681), .A2(n1680), .ZN(n1682) );
  INVD1BWP12T U2641 ( .I(n1696), .ZN(n1698) );
  ND2D1BWP12T U2642 ( .A1(n1698), .A2(n1697), .ZN(n1700) );
  XOR2XD1BWP12T U2643 ( .A1(n1700), .A2(n1699), .Z(n2568) );
  AOI21D1BWP12T U2644 ( .A1(n1721), .A2(n1720), .B(n1719), .ZN(n1725) );
  ND2D1BWP12T U2645 ( .A1(n1723), .A2(n1722), .ZN(n1724) );
  XOR2XD1BWP12T U2646 ( .A1(n1725), .A2(n1724), .Z(n2938) );
  INVD1BWP12T U2647 ( .I(n1730), .ZN(n1732) );
  ND2D1BWP12T U2648 ( .A1(n1732), .A2(n1731), .ZN(n1733) );
  XOR2XD1BWP12T U2649 ( .A1(n1734), .A2(n1733), .Z(n2978) );
  NR4D0BWP12T U2650 ( .A1(n1740), .A2(n1739), .A3(n1738), .A4(n1737), .ZN(
        n1741) );
  TPND2D0BWP12T U2651 ( .A1(n1742), .A2(n1741), .ZN(n2469) );
  FA1D2BWP12T U2652 ( .A(a[26]), .B(b[26]), .CI(n1743), .CO(n1800), .S(n2768)
         );
  FA1D2BWP12T U2653 ( .A(n2747), .B(b[23]), .CI(n1744), .CO(n1798), .S(n2741)
         );
  FA1D2BWP12T U2654 ( .A(a[20]), .B(b[20]), .CI(n1745), .CO(n1796), .S(n2935)
         );
  INVD1BWP12T U2655 ( .I(n1750), .ZN(n1751) );
  INVD1BWP12T U2656 ( .I(n1752), .ZN(n2347) );
  ND2D1BWP12T U2657 ( .A1(n2354), .A2(n1755), .ZN(n1757) );
  XOR2XD1BWP12T U2658 ( .A1(n1757), .A2(n1756), .Z(n2490) );
  INVD1BWP12T U2659 ( .I(n1760), .ZN(n1769) );
  INVD0BWP12T U2660 ( .I(n1768), .ZN(n1761) );
  AOI21D1BWP12T U2661 ( .A1(n1786), .A2(n1769), .B(n1761), .ZN(n1766) );
  INVD0BWP12T U2662 ( .I(n1762), .ZN(n1764) );
  CKND2D1BWP12T U2663 ( .A1(n1764), .A2(n1763), .ZN(n1765) );
  XOR2XD1BWP12T U2664 ( .A1(n1766), .A2(n1765), .Z(n2859) );
  ND2D1BWP12T U2665 ( .A1(n1769), .A2(n1768), .ZN(n1770) );
  XNR2D1BWP12T U2666 ( .A1(n1786), .A2(n1770), .ZN(n2846) );
  AOI21D1BWP12T U2667 ( .A1(n1775), .A2(n1774), .B(n1773), .ZN(n1777) );
  TPND2D0BWP12T U2668 ( .A1(n2368), .A2(n2367), .ZN(n1776) );
  XOR2XD1BWP12T U2669 ( .A1(n1777), .A2(n1776), .Z(n2561) );
  CKND0BWP12T U2670 ( .I(n1778), .ZN(n1779) );
  NR2D0BWP12T U2671 ( .A1(n1779), .A2(n1782), .ZN(n1785) );
  CKND0BWP12T U2672 ( .I(n1780), .ZN(n1783) );
  TPOAI21D0BWP12T U2673 ( .A1(n1783), .A2(n1782), .B(n1781), .ZN(n1784) );
  AOI21D1BWP12T U2674 ( .A1(n1786), .A2(n1785), .B(n1784), .ZN(n1788) );
  INVD1BWP12T U2675 ( .I(n2373), .ZN(n2351) );
  TPND2D0BWP12T U2676 ( .A1(n2351), .A2(n2372), .ZN(n1787) );
  XOR2XD1BWP12T U2677 ( .A1(n1788), .A2(n1787), .Z(n2588) );
  INVD0BWP12T U2678 ( .I(n1793), .ZN(n2338) );
  FA1D2BWP12T U2679 ( .A(n2725), .B(b[21]), .CI(n1796), .CO(n738), .S(n2715)
         );
  FA1D2BWP12T U2680 ( .A(a[24]), .B(b[24]), .CI(n1798), .CO(n700), .S(n2969)
         );
  FA1D2BWP12T U2681 ( .A(a[27]), .B(b[27]), .CI(n1800), .CO(n1456), .S(n2800)
         );
  NR4D0BWP12T U2682 ( .A1(n1805), .A2(n1804), .A3(n1803), .A4(n1802), .ZN(
        n2467) );
  NR4D0BWP12T U2683 ( .A1(a[31]), .A2(a[26]), .A3(a[27]), .A4(a[24]), .ZN(
        n1809) );
  NR4D0BWP12T U2684 ( .A1(a[29]), .A2(a[28]), .A3(a[25]), .A4(n2900), .ZN(
        n1808) );
  NR4D0BWP12T U2685 ( .A1(a[14]), .A2(n2301), .A3(a[8]), .A4(n2594), .ZN(n1807) );
  NR4D0BWP12T U2686 ( .A1(a[18]), .A2(n2626), .A3(n2643), .A4(n2308), .ZN(
        n1806) );
  ND4D1BWP12T U2687 ( .A1(n1809), .A2(n1808), .A3(n1807), .A4(n1806), .ZN(
        n1847) );
  NR4D0BWP12T U2688 ( .A1(n2747), .A2(n2679), .A3(a[16]), .A4(a[20]), .ZN(
        n1813) );
  NR4D0BWP12T U2689 ( .A1(n2620), .A2(n2871), .A3(n2830), .A4(n2482), .ZN(
        n1810) );
  AN4XD1BWP12T U2690 ( .A1(n1832), .A2(n2532), .A3(n2825), .A4(n1810), .Z(
        n1812) );
  NR4D0BWP12T U2691 ( .A1(n2609), .A2(a[22]), .A3(n2725), .A4(n2574), .ZN(
        n1811) );
  ND4D0BWP12T U2692 ( .A1(n1814), .A2(n1813), .A3(n1812), .A4(n1811), .ZN(
        n1846) );
  HA1D1BWP12T U2693 ( .A(n1816), .B(n1815), .CO(n1486), .S(n2811) );
  HA1D1BWP12T U2694 ( .A(n2779), .B(n1817), .CO(n1815), .S(n2790) );
  HA1D0BWP12T U2695 ( .A(n2946), .B(n1818), .CO(n701), .S(n2941) );
  HA1D1BWP12T U2696 ( .A(n2751), .B(n1819), .CO(n1818), .S(n2756) );
  XNR2D1BWP12T U2697 ( .A1(n1823), .A2(a[8]), .ZN(n2543) );
  HA1D0BWP12T U2698 ( .A(n1829), .B(n1828), .CO(n1838), .S(n2927) );
  XNR2XD1BWP12T U2699 ( .A1(n2482), .A2(n2603), .ZN(n2487) );
  HA1D1BWP12T U2700 ( .A(n2233), .B(n1838), .CO(n739), .S(n2731) );
  OR4D1BWP12T U2701 ( .A1(n1844), .A2(n1843), .A3(n1842), .A4(n2666), .Z(n1845) );
  OAI31D0BWP12T U2702 ( .A1(n1847), .A2(n2174), .A3(n1846), .B(n1845), .ZN(
        n2401) );
  OAI22D1BWP12T U2703 ( .A1(n1848), .A2(n2052), .B1(n1856), .B2(n1926), .ZN(
        n2961) );
  ND4D0BWP12T U2704 ( .A1(n1851), .A2(n1850), .A3(n1856), .A4(n1849), .ZN(
        n1853) );
  CKND2D1BWP12T U2705 ( .A1(n1852), .A2(n2827), .ZN(n2046) );
  OR4D0BWP12T U2706 ( .A1(n2569), .A2(n2961), .A3(n1853), .A4(n2746), .Z(n1981) );
  CKND2D1BWP12T U2707 ( .A1(n1854), .A2(n2827), .ZN(n1960) );
  INVD1BWP12T U2708 ( .I(n1960), .ZN(n2804) );
  CKND2D1BWP12T U2709 ( .A1(n2770), .A2(n2827), .ZN(n1918) );
  TPNR2D0BWP12T U2710 ( .A1(n1856), .A2(n1933), .ZN(n1857) );
  AOI21D1BWP12T U2711 ( .A1(n1858), .A2(n2827), .B(n1857), .ZN(n1969) );
  CKND2D0BWP12T U2712 ( .A1(n1969), .A2(n1859), .ZN(n1964) );
  CKND2D0BWP12T U2713 ( .A1(n1860), .A2(n2831), .ZN(n1865) );
  NR2XD0BWP12T U2714 ( .A1(n1863), .A2(n1930), .ZN(n1864) );
  AOI21D1BWP12T U2715 ( .A1(n1865), .A2(n2055), .B(n1864), .ZN(n1976) );
  NR2D0BWP12T U2716 ( .A1(n1866), .A2(n1976), .ZN(n1961) );
  INVD1BWP12T U2717 ( .I(n1866), .ZN(n1880) );
  OAI22D0BWP12T U2718 ( .A1(n1870), .A2(n2512), .B1(n1869), .B2(n1441), .ZN(
        n1868) );
  OAI22D0BWP12T U2719 ( .A1(n1872), .A2(n2241), .B1(n1871), .B2(n2242), .ZN(
        n1867) );
  NR2D1BWP12T U2720 ( .A1(n1868), .A2(n1867), .ZN(n1927) );
  OAI22D0BWP12T U2721 ( .A1(n1927), .A2(n1933), .B1(n1883), .B2(n1930), .ZN(
        n1879) );
  OAI22D0BWP12T U2722 ( .A1(n1870), .A2(n2532), .B1(n1869), .B2(n2898), .ZN(
        n1874) );
  OAI22D1BWP12T U2723 ( .A1(n1872), .A2(n2243), .B1(n1871), .B2(n2550), .ZN(
        n1873) );
  NR2D1BWP12T U2724 ( .A1(n1874), .A2(n1873), .ZN(n1925) );
  OAI21D0BWP12T U2725 ( .A1(n1925), .A2(n1926), .B(n2870), .ZN(n1878) );
  AOI22D0BWP12T U2726 ( .A1(n1892), .A2(n2871), .B1(n1891), .B2(n2830), .ZN(
        n1876) );
  AOI22D0BWP12T U2727 ( .A1(n2620), .A2(n1894), .B1(n1893), .B2(n2574), .ZN(
        n1875) );
  AOI21D0BWP12T U2728 ( .A1(n1876), .A2(n1875), .B(n2831), .ZN(n1877) );
  NR3D1BWP12T U2729 ( .A1(n1879), .A2(n1878), .A3(n1877), .ZN(n2092) );
  AOI21D1BWP12T U2730 ( .A1(n1880), .A2(n2868), .B(n2092), .ZN(n2823) );
  AOI21D1BWP12T U2731 ( .A1(n2868), .A2(n1960), .B(n2053), .ZN(n2507) );
  NR3D0BWP12T U2732 ( .A1(n2823), .A2(n2507), .A3(n1884), .ZN(n1984) );
  INR3XD0BWP12T U2733 ( .A1(n1984), .B1(n1886), .B2(n1885), .ZN(n1887) );
  OAI22D0BWP12T U2734 ( .A1(n1888), .A2(n2135), .B1(n1887), .B2(n2174), .ZN(
        n2330) );
  TPNR2D0BWP12T U2735 ( .A1(n1976), .A2(n2870), .ZN(n2496) );
  TPOAI22D0BWP12T U2736 ( .A1(n1890), .A2(n1930), .B1(n1889), .B2(n1933), .ZN(
        n1900) );
  TPAOI22D0BWP12T U2737 ( .A1(n1892), .A2(n2303), .B1(n1891), .B2(n2482), .ZN(
        n1896) );
  AOI22D0BWP12T U2738 ( .A1(n2830), .A2(n1894), .B1(n1893), .B2(n2871), .ZN(
        n1895) );
  TPAOI21D0BWP12T U2739 ( .A1(n1896), .A2(n1895), .B(n2831), .ZN(n1899) );
  TPNR2D0BWP12T U2740 ( .A1(n1897), .A2(n1926), .ZN(n1898) );
  NR3D1BWP12T U2741 ( .A1(n1900), .A2(n1899), .A3(n1898), .ZN(n2494) );
  AOI21D1BWP12T U2742 ( .A1(n2870), .A2(n2494), .B(n2174), .ZN(n2499) );
  CKND0BWP12T U2743 ( .I(n2499), .ZN(n1909) );
  OAI21D0BWP12T U2744 ( .A1(n1902), .A2(n1901), .B(n2115), .ZN(n1908) );
  CKND0BWP12T U2745 ( .I(n1978), .ZN(n1905) );
  INVD1BWP12T U2746 ( .I(n2047), .ZN(n2560) );
  AOI21D0BWP12T U2747 ( .A1(n1906), .A2(n1905), .B(n2560), .ZN(n1907) );
  OAI211D0BWP12T U2748 ( .A1(n2496), .A2(n1909), .B(n1908), .C(n1907), .ZN(
        n1923) );
  INVD1BWP12T U2749 ( .I(n1969), .ZN(n2931) );
  ND2XD0BWP12T U2750 ( .A1(n2931), .A2(n2115), .ZN(n1917) );
  AOI21D1BWP12T U2751 ( .A1(n1910), .A2(n2049), .B(n2868), .ZN(n1911) );
  TPOAI21D0BWP12T U2752 ( .A1(n1912), .A2(n1930), .B(n1911), .ZN(n1916) );
  OAI22D0BWP12T U2753 ( .A1(n1914), .A2(n1933), .B1(n1913), .B2(n2052), .ZN(
        n1915) );
  NR2D1BWP12T U2754 ( .A1(n1916), .A2(n1915), .ZN(n2872) );
  TPAOI21D0BWP12T U2755 ( .A1(n1917), .A2(n2135), .B(n2872), .ZN(n2860) );
  INVD1BWP12T U2756 ( .I(n1918), .ZN(n2895) );
  CKND2D0BWP12T U2757 ( .A1(n2895), .A2(n2115), .ZN(n1921) );
  RCAOI21D0BWP12T U2758 ( .A1(n2135), .A2(n1921), .B(n2896), .ZN(n2885) );
  NR4D0BWP12T U2759 ( .A1(n1923), .A2(n2860), .A3(n2885), .A4(n1922), .ZN(
        n1939) );
  CKND2D0BWP12T U2760 ( .A1(n2746), .A2(n2115), .ZN(n1928) );
  AOI21D0BWP12T U2761 ( .A1(n1928), .A2(n2135), .B(n2540), .ZN(n2538) );
  CKND0BWP12T U2762 ( .I(n2569), .ZN(n1935) );
  AOI211D1BWP12T U2763 ( .A1(n2868), .A2(n1935), .B(n2585), .C(n2174), .ZN(
        n2590) );
  NR4D0BWP12T U2764 ( .A1(n2538), .A2(n2590), .A3(n1936), .A4(n2495), .ZN(
        n1938) );
  ND3D0BWP12T U2765 ( .A1(n1939), .A2(n1938), .A3(n1937), .ZN(n2329) );
  TPNR2D0BWP12T U2766 ( .A1(n1940), .A2(n2121), .ZN(n1943) );
  OAI22D0BWP12T U2767 ( .A1(n1941), .A2(n2117), .B1(n1959), .B2(n2118), .ZN(
        n1942) );
  AOI211D1BWP12T U2768 ( .A1(n1945), .A2(n1944), .B(n1943), .C(n1942), .ZN(
        n1990) );
  MUX2NXD0BWP12T U2769 ( .I0(n1990), .I1(n1946), .S(n1998), .ZN(n1955) );
  NR4D0BWP12T U2770 ( .A1(n1947), .A2(n2526), .A3(n2770), .A4(n2573), .ZN(
        n1950) );
  MUX2D1BWP12T U2771 ( .I0(n1973), .I1(n1948), .S(n2017), .Z(n1965) );
  ND4D0BWP12T U2772 ( .A1(n1955), .A2(n1950), .A3(n1949), .A4(n1965), .ZN(
        n1954) );
  NR4D0BWP12T U2773 ( .A1(n1954), .A2(n1953), .A3(n1952), .A4(n1951), .ZN(
        n1968) );
  INVD1BWP12T U2774 ( .I(n1955), .ZN(n2904) );
  AOI22D0BWP12T U2775 ( .A1(n2001), .A2(n2127), .B1(n2000), .B2(n1956), .ZN(
        n1958) );
  CKND2D0BWP12T U2776 ( .A1(n2002), .A2(n2149), .ZN(n1957) );
  OAI211D0BWP12T U2777 ( .A1(n2124), .A2(n1959), .B(n1958), .C(n1957), .ZN(
        n1991) );
  ND4D0BWP12T U2778 ( .A1(n2585), .A2(n2494), .A3(n2063), .A4(n1960), .ZN(
        n1963) );
  ND3D0BWP12T U2779 ( .A1(n1961), .A2(n2540), .A3(n2872), .ZN(n1962) );
  OAI31D0BWP12T U2780 ( .A1(n1964), .A2(n1963), .A3(n1962), .B(n2870), .ZN(
        n1967) );
  INVD1BWP12T U2781 ( .I(n1965), .ZN(n2510) );
  AN4D0BWP12T U2782 ( .A1(n1968), .A2(n2772), .A3(n1967), .A4(n2802), .Z(n2112) );
  OAI22D1BWP12T U2783 ( .A1(n1970), .A2(n2025), .B1(n1969), .B2(n2872), .ZN(
        n2861) );
  NR3D0BWP12T U2784 ( .A1(n1972), .A2(n2861), .A3(n1971), .ZN(n1985) );
  ND4D0BWP12T U2785 ( .A1(n1975), .A2(n1974), .A3(n2894), .A4(n1973), .ZN(
        n1980) );
  INVD1BWP12T U2786 ( .I(n1976), .ZN(n2676) );
  OAI22D1BWP12T U2787 ( .A1(n2676), .A2(n2870), .B1(n2025), .B2(n2021), .ZN(
        n2497) );
  OAI22D1BWP12T U2788 ( .A1(n1978), .A2(n1977), .B1(n2896), .B2(n2868), .ZN(
        n1979) );
  NR4D0BWP12T U2789 ( .A1(n1981), .A2(n1980), .A3(n2497), .A4(n1979), .ZN(
        n1983) );
  ND4D0BWP12T U2790 ( .A1(n1985), .A2(n1984), .A3(n1983), .A4(n1982), .ZN(
        n2043) );
  AOI22D0BWP12T U2791 ( .A1(n1987), .A2(n2031), .B1(n1986), .B2(n1998), .ZN(
        n1988) );
  OA211D0BWP12T U2792 ( .A1(n1997), .A2(n2526), .B(n1988), .C(n2014), .Z(n2755) );
  NR2D0BWP12T U2793 ( .A1(n2755), .A2(n1989), .ZN(n1996) );
  ND4D0BWP12T U2794 ( .A1(n1996), .A2(n1995), .A3(n2708), .A4(n1994), .ZN(
        n2042) );
  OR3XD0BWP12T U2795 ( .A1(n1998), .A2(n1997), .A3(n2018), .Z(n2010) );
  CKND2D0BWP12T U2796 ( .A1(n1999), .A2(n2168), .ZN(n2005) );
  AOI22D0BWP12T U2797 ( .A1(n2001), .A2(n2167), .B1(n2000), .B2(n2149), .ZN(
        n2004) );
  CKND2D0BWP12T U2798 ( .A1(n2002), .A2(n2171), .ZN(n2003) );
  AOI31D0BWP12T U2799 ( .A1(n2005), .A2(n2004), .A3(n2003), .B(n2025), .ZN(
        n2007) );
  AOI211D0BWP12T U2800 ( .A1(n2008), .A2(n2153), .B(n2007), .C(n2006), .ZN(
        n2009) );
  OAI211D1BWP12T U2801 ( .A1(n2023), .A2(n2011), .B(n2010), .C(n2009), .ZN(
        n2965) );
  AOI22D0BWP12T U2802 ( .A1(n2031), .A2(n2013), .B1(n2012), .B2(n2508), .ZN(
        n2015) );
  OAI211D1BWP12T U2803 ( .A1(n2017), .A2(n2016), .B(n2015), .C(n2014), .ZN(
        n2717) );
  INVD1BWP12T U2804 ( .I(n2018), .ZN(n2020) );
  NR2D0BWP12T U2805 ( .A1(n2961), .A2(n2870), .ZN(n2019) );
  OA222D1BWP12T U2806 ( .A1(n2023), .A2(n2153), .B1(n2025), .B2(n2020), .C1(
        n2048), .C2(n2019), .Z(n2556) );
  OAI22D0BWP12T U2807 ( .A1(n2024), .A2(n2023), .B1(n2022), .B2(n2021), .ZN(
        n2029) );
  AOI21D0BWP12T U2808 ( .A1(n2027), .A2(n2026), .B(n2025), .ZN(n2028) );
  NR2D1BWP12T U2809 ( .A1(n2029), .A2(n2028), .ZN(n2690) );
  ND4D0BWP12T U2810 ( .A1(n2965), .A2(n2717), .A3(n2556), .A4(n2690), .ZN(
        n2041) );
  INVD1BWP12T U2811 ( .I(n2030), .ZN(n2032) );
  AOI222D1BWP12T U2812 ( .A1(n2036), .A2(n2035), .B1(n2034), .B2(n2033), .C1(
        n2032), .C2(n2031), .ZN(n2928) );
  ND4D0BWP12T U2813 ( .A1(n2039), .A2(n2928), .A3(n2038), .A4(n2037), .ZN(
        n2040) );
  NR4D0BWP12T U2814 ( .A1(n2043), .A2(n2042), .A3(n2041), .A4(n2040), .ZN(
        n2111) );
  OAI21D0BWP12T U2815 ( .A1(n2099), .A2(n471), .B(n2868), .ZN(n2044) );
  TPNR2D0BWP12T U2816 ( .A1(n2931), .A2(n2044), .ZN(n2045) );
  TPOAI31D0BWP12T U2817 ( .A1(n2872), .A2(n2174), .A3(n2045), .B(n2105), .ZN(
        n2881) );
  TPOAI21D0BWP12T U2818 ( .A1(n2046), .A2(n2068), .B(n2956), .ZN(n2743) );
  OAI211D1BWP12T U2819 ( .A1(n2048), .A2(n2099), .B(n2047), .C(n2105), .ZN(
        n2557) );
  CKND2D0BWP12T U2820 ( .A1(n2049), .A2(a[31]), .ZN(n2050) );
  OAI211D0BWP12T U2821 ( .A1(n2052), .A2(n2051), .B(n2050), .C(n2099), .ZN(
        n2083) );
  AOI21D0BWP12T U2822 ( .A1(n2115), .A2(n2083), .B(n2198), .ZN(n2054) );
  TPOAI21D0BWP12T U2823 ( .A1(n2054), .A2(n2053), .B(n2105), .ZN(n2509) );
  NR4D0BWP12T U2824 ( .A1(n2881), .A2(n2743), .A3(n2557), .A4(n2509), .ZN(
        n2062) );
  INVD1BWP12T U2825 ( .I(n2055), .ZN(n2056) );
  TPAOI21D0BWP12T U2826 ( .A1(n2831), .A2(n2057), .B(n2056), .ZN(n2674) );
  ND2D1BWP12T U2827 ( .A1(n2674), .A2(n2868), .ZN(n2059) );
  TPAOI21D0BWP12T U2828 ( .A1(n2059), .A2(n2499), .B(n2058), .ZN(n2472) );
  ND4D0BWP12T U2829 ( .A1(n2062), .A2(n2061), .A3(n2472), .A4(n2060), .ZN(
        n2075) );
  CKND0BWP12T U2830 ( .I(n2091), .ZN(n2064) );
  AN4D0BWP12T U2831 ( .A1(n2064), .A2(n2719), .A3(n2063), .A4(n2674), .Z(n2067) );
  AOI31D0BWP12T U2832 ( .A1(n2067), .A2(n2066), .A3(n2065), .B(n2068), .ZN(
        n2074) );
  OAI21D0BWP12T U2833 ( .A1(n2069), .A2(n2068), .B(n2094), .ZN(n2707) );
  ND3D0BWP12T U2834 ( .A1(n2072), .A2(n2071), .A3(n2070), .ZN(n2073) );
  NR4D0BWP12T U2835 ( .A1(n2075), .A2(n2074), .A3(n2707), .A4(n2073), .ZN(
        n2110) );
  AOI21D0BWP12T U2836 ( .A1(n2076), .A2(n2115), .B(n2198), .ZN(n2077) );
  OA21D1BWP12T U2837 ( .A1(n2077), .A2(n2585), .B(n2105), .Z(n2591) );
  ND2D1BWP12T U2838 ( .A1(n2078), .A2(n2868), .ZN(n2081) );
  AOI21D0BWP12T U2839 ( .A1(n2081), .A2(n2080), .B(n2079), .ZN(n2082) );
  TPOAI31D0BWP12T U2840 ( .A1(n2174), .A2(n2082), .A3(n2540), .B(n2105), .ZN(
        n2537) );
  TPND2D0BWP12T U2841 ( .A1(n2084), .A2(n2083), .ZN(n2803) );
  CKND2D0BWP12T U2842 ( .A1(n2084), .A2(n2961), .ZN(n2085) );
  ND4D0BWP12T U2843 ( .A1(n2803), .A2(n2905), .A3(n2310), .A4(n2085), .ZN(
        n2086) );
  NR4D0BWP12T U2844 ( .A1(n2088), .A2(n2537), .A3(n2087), .A4(n2086), .ZN(
        n2089) );
  ND3D0BWP12T U2845 ( .A1(n2090), .A2(n2591), .A3(n2089), .ZN(n2108) );
  AOI21D0BWP12T U2846 ( .A1(n2091), .A2(n2115), .B(n2198), .ZN(n2093) );
  TPOAI21D0BWP12T U2847 ( .A1(n2093), .A2(n2092), .B(n2105), .ZN(n2852) );
  AOI21D0BWP12T U2848 ( .A1(n471), .A2(n2094), .B(n2956), .ZN(n2096) );
  INVD0BWP12T U2849 ( .I(n2095), .ZN(n2100) );
  OAI21D1BWP12T U2850 ( .A1(n2096), .A2(n2931), .B(n2100), .ZN(n2933) );
  OAI21D0BWP12T U2851 ( .A1(n2101), .A2(n2782), .B(n2100), .ZN(n2102) );
  IND4D0BWP12T U2852 ( .A1(n2104), .B1(n2933), .B2(n2103), .B3(n2102), .ZN(
        n2107) );
  AOI21D0BWP12T U2853 ( .A1(n2782), .A2(n2115), .B(n2198), .ZN(n2106) );
  OAI21D1BWP12T U2854 ( .A1(n2106), .A2(n2896), .B(n2105), .ZN(n2906) );
  NR4D0BWP12T U2855 ( .A1(n2108), .A2(n2852), .A3(n2107), .A4(n2906), .ZN(
        n2109) );
  AOI22D1BWP12T U2856 ( .A1(n2112), .A2(n2111), .B1(n2110), .B2(n2109), .ZN(
        n2328) );
  IND3D0BWP12T U2857 ( .A1(n2184), .B1(n2138), .B2(n2474), .ZN(n2113) );
  NR4D0BWP12T U2858 ( .A1(n2179), .A2(n2113), .A3(n2581), .A4(n2875), .ZN(
        n2114) );
  NR2D0BWP12T U2859 ( .A1(n2114), .A2(n2135), .ZN(n2132) );
  NR2D0BWP12T U2860 ( .A1(n2164), .A2(n2831), .ZN(n2137) );
  CKND2D0BWP12T U2861 ( .A1(n2137), .A2(n2115), .ZN(n2131) );
  OAI22D0BWP12T U2862 ( .A1(n2119), .A2(n2118), .B1(n2117), .B2(n2116), .ZN(
        n2123) );
  OAI22D0BWP12T U2863 ( .A1(n2121), .A2(n2126), .B1(n2120), .B2(n2128), .ZN(
        n2122) );
  NR2D1BWP12T U2864 ( .A1(n2123), .A2(n2122), .ZN(n2163) );
  AOI22D0BWP12T U2865 ( .A1(n2169), .A2(n2125), .B1(n2124), .B2(n2166), .ZN(
        n2165) );
  CKND2D0BWP12T U2866 ( .A1(n2165), .A2(n2769), .ZN(n2129) );
  OAI22D0BWP12T U2867 ( .A1(n2128), .A2(n2127), .B1(n2149), .B2(n2126), .ZN(
        n2175) );
  OAI22D1BWP12T U2868 ( .A1(n2163), .A2(n2200), .B1(n2129), .B2(n2175), .ZN(
        n2130) );
  AOI21D0BWP12T U2869 ( .A1(n2135), .A2(n2131), .B(n2130), .ZN(n2704) );
  NR4D0BWP12T U2870 ( .A1(n2134), .A2(n2133), .A3(n2132), .A4(n2704), .ZN(
        n2162) );
  NR2XD0BWP12T U2871 ( .A1(n2160), .A2(n2831), .ZN(n2136) );
  RCAOI211D0BWP12T U2872 ( .A1(n2831), .A2(n2153), .B(n2136), .C(n2135), .ZN(
        n2546) );
  AOI211D0BWP12T U2873 ( .A1(n2198), .A2(n2137), .B(n2546), .C(n2942), .ZN(
        n2161) );
  INVD1BWP12T U2874 ( .I(n2138), .ZN(n2844) );
  AOI22D0BWP12T U2875 ( .A1(n2170), .A2(n2141), .B1(n2140), .B2(n2173), .ZN(
        n2145) );
  AOI22D0BWP12T U2876 ( .A1(n2169), .A2(n2143), .B1(n2142), .B2(n2166), .ZN(
        n2144) );
  AOI21D0BWP12T U2877 ( .A1(n2145), .A2(n2144), .B(n2202), .ZN(n2146) );
  AOI211D0BWP12T U2878 ( .A1(n2155), .A2(n2147), .B(n2174), .C(n2146), .ZN(
        n2148) );
  OAI21D0BWP12T U2879 ( .A1(n2514), .A2(n2870), .B(n2148), .ZN(n2808) );
  AOI22D0BWP12T U2880 ( .A1(n2169), .A2(n2149), .B1(n2168), .B2(n2166), .ZN(
        n2151) );
  AOI22D0BWP12T U2881 ( .A1(n2173), .A2(n2171), .B1(n2167), .B2(n2170), .ZN(
        n2150) );
  AOI21D0BWP12T U2882 ( .A1(n2151), .A2(n2150), .B(n2202), .ZN(n2152) );
  RCAOI211D0BWP12T U2883 ( .A1(n2154), .A2(n2153), .B(n2152), .C(n2174), .ZN(
        n2158) );
  TPND2D0BWP12T U2884 ( .A1(n2156), .A2(n2155), .ZN(n2157) );
  OAI211D1BWP12T U2885 ( .A1(n2160), .A2(n2159), .B(n2158), .C(n2157), .ZN(
        n2943) );
  ND4D0BWP12T U2886 ( .A1(n2162), .A2(n2161), .A3(n2808), .A4(n2943), .ZN(
        n2193) );
  MAOI22D0BWP12T U2887 ( .A1(n2177), .A2(n2769), .B1(n2176), .B2(n2827), .ZN(
        n2178) );
  OAI211D0BWP12T U2888 ( .A1(n2179), .A2(n2870), .B(n2178), .C(n2187), .ZN(
        n2744) );
  CKND0BWP12T U2889 ( .I(n2180), .ZN(n2181) );
  AOI22D0BWP12T U2890 ( .A1(n2769), .A2(n2182), .B1(n2181), .B2(n2831), .ZN(
        n2183) );
  OAI211D0BWP12T U2891 ( .A1(n2875), .A2(n2870), .B(n2183), .C(n2187), .ZN(
        n2930) );
  CKND0BWP12T U2892 ( .I(n2184), .ZN(n2186) );
  AOI22D1BWP12T U2893 ( .A1(n2868), .A2(n2186), .B1(n2185), .B2(n2769), .ZN(
        n2188) );
  OAI211D0BWP12T U2894 ( .A1(n2189), .A2(n2827), .B(n2188), .C(n2187), .ZN(
        n2728) );
  ND4D0BWP12T U2895 ( .A1(n2744), .A2(n2190), .A3(n2930), .A4(n2728), .ZN(
        n2191) );
  NR4D0BWP12T U2896 ( .A1(n2193), .A2(n2787), .A3(n2192), .A4(n2191), .ZN(
        n2326) );
  INVD1BWP12T U2897 ( .I(n2199), .ZN(n2203) );
  OAI22D0BWP12T U2898 ( .A1(n2203), .A2(n2202), .B1(n2201), .B2(n2200), .ZN(
        n2205) );
  AO211D1BWP12T U2899 ( .A1(n2868), .A2(n2474), .B(n2205), .C(n2204), .Z(n2673) );
  ND4D0BWP12T U2900 ( .A1(n2673), .A2(n2208), .A3(n2207), .A4(n2206), .ZN(
        n2212) );
  NR4D0BWP12T U2901 ( .A1(n2212), .A2(n2211), .A3(n2210), .A4(n2209), .ZN(
        n2324) );
  AOI22D1BWP12T U2902 ( .A1(n2605), .A2(a[8]), .B1(b[6]), .B2(n2574), .ZN(
        n2216) );
  AOI22D0BWP12T U2903 ( .A1(a[31]), .A2(b[31]), .B1(n2528), .B2(n2527), .ZN(
        n2215) );
  AOI22D0BWP12T U2904 ( .A1(b[13]), .A2(n2643), .B1(b[14]), .B2(a[14]), .ZN(
        n2214) );
  AOI22D0BWP12T U2905 ( .A1(b[11]), .A2(n2594), .B1(n2897), .B2(n2900), .ZN(
        n2213) );
  ND4D1BWP12T U2906 ( .A1(n2216), .A2(n2215), .A3(n2214), .A4(n2213), .ZN(
        n2322) );
  AOI22D0BWP12T U2907 ( .A1(b[26]), .A2(a[26]), .B1(n2477), .B2(n2482), .ZN(
        n2220) );
  AOI22D0BWP12T U2908 ( .A1(b[24]), .A2(a[24]), .B1(b[25]), .B2(a[25]), .ZN(
        n2219) );
  AOI22D0BWP12T U2909 ( .A1(b[5]), .A2(n2620), .B1(n2868), .B2(n2871), .ZN(
        n2218) );
  AOI22D0BWP12T U2910 ( .A1(n2831), .A2(n2830), .B1(n2639), .B2(n2303), .ZN(
        n2217) );
  ND4D1BWP12T U2911 ( .A1(n2220), .A2(n2219), .A3(n2218), .A4(n2217), .ZN(
        n2321) );
  AOI22D0BWP12T U2912 ( .A1(b[21]), .A2(n2725), .B1(b[20]), .B2(a[20]), .ZN(
        n2224) );
  AOI22D0BWP12T U2913 ( .A1(b[22]), .A2(a[22]), .B1(b[30]), .B2(a[30]), .ZN(
        n2223) );
  AOI22D0BWP12T U2914 ( .A1(b[27]), .A2(a[27]), .B1(b[29]), .B2(a[29]), .ZN(
        n2222) );
  AOI22D0BWP12T U2915 ( .A1(b[28]), .A2(a[28]), .B1(b[23]), .B2(n2747), .ZN(
        n2221) );
  ND4D1BWP12T U2916 ( .A1(n2224), .A2(n2223), .A3(n2222), .A4(n2221), .ZN(
        n2230) );
  AOI22D0BWP12T U2917 ( .A1(n2598), .A2(n2308), .B1(b[15]), .B2(n2626), .ZN(
        n2227) );
  AOI22D0BWP12T U2918 ( .A1(b[18]), .A2(a[18]), .B1(b[16]), .B2(a[16]), .ZN(
        n2226) );
  AOI22D0BWP12T U2919 ( .A1(b[19]), .A2(n2609), .B1(b[17]), .B2(n2679), .ZN(
        n2225) );
  TPND3D0BWP12T U2920 ( .A1(n2227), .A2(n2226), .A3(n2225), .ZN(n2228) );
  AO211D0BWP12T U2921 ( .A1(n2301), .A2(b[9]), .B(n2951), .C(n2228), .Z(n2229)
         );
  AO211D0BWP12T U2922 ( .A1(n2302), .A2(n2231), .B(n2230), .C(n2229), .Z(n2320) );
  AOI22D0BWP12T U2923 ( .A1(b[22]), .A2(n2232), .B1(n2751), .B2(b[23]), .ZN(
        n2239) );
  AOI22D0BWP12T U2924 ( .A1(b[20]), .A2(n2929), .B1(n2233), .B2(b[21]), .ZN(
        n2238) );
  AOI22D0BWP12T U2925 ( .A1(b[18]), .A2(n2705), .B1(n2234), .B2(b[19]), .ZN(
        n2237) );
  AOI22D0BWP12T U2926 ( .A1(b[16]), .A2(n2235), .B1(n2683), .B2(b[17]), .ZN(
        n2236) );
  ND4D1BWP12T U2927 ( .A1(n2239), .A2(n2238), .A3(n2237), .A4(n2236), .ZN(
        n2268) );
  AOI22D0BWP12T U2928 ( .A1(b[14]), .A2(n1441), .B1(n2240), .B2(b[15]), .ZN(
        n2247) );
  AOI22D0BWP12T U2929 ( .A1(n2598), .A2(n2242), .B1(n2241), .B2(b[13]), .ZN(
        n2246) );
  AOI22D0BWP12T U2930 ( .A1(n2897), .A2(n2898), .B1(n2512), .B2(b[11]), .ZN(
        n2245) );
  AOI22D1BWP12T U2931 ( .A1(n2605), .A2(n2550), .B1(n2243), .B2(b[9]), .ZN(
        n2244) );
  ND4D1BWP12T U2932 ( .A1(n2247), .A2(n2246), .A3(n2245), .A4(n2244), .ZN(
        n2267) );
  AO22XD0BWP12T U2933 ( .A1(b[28]), .A2(n2249), .B1(n2248), .B2(b[29]), .Z(
        n2250) );
  AOI211D0BWP12T U2934 ( .A1(b[30]), .A2(n2251), .B(n2250), .C(n2944), .ZN(
        n2256) );
  AOI22D0BWP12T U2935 ( .A1(b[26]), .A2(n2779), .B1(n2252), .B2(b[27]), .ZN(
        n2255) );
  AOI22D0BWP12T U2936 ( .A1(b[24]), .A2(n2946), .B1(n2253), .B2(b[25]), .ZN(
        n2254) );
  ND4D0BWP12T U2937 ( .A1(n2256), .A2(n2255), .A3(n2254), .A4(n2663), .ZN(
        n2263) );
  AOI22D1BWP12T U2938 ( .A1(b[6]), .A2(n2578), .B1(n2532), .B2(n2528), .ZN(
        n2262) );
  AOI22D0BWP12T U2939 ( .A1(n2868), .A2(n2869), .B1(n2257), .B2(b[5]), .ZN(
        n2261) );
  OAI22D0BWP12T U2940 ( .A1(n2830), .A2(n2827), .B1(n471), .B2(n2303), .ZN(
        n2259) );
  AOI211D0BWP12T U2941 ( .A1(n2477), .A2(n2481), .B(n2259), .C(n2258), .ZN(
        n2260) );
  IND4D1BWP12T U2942 ( .A1(n2263), .B1(n2262), .B2(n2261), .B3(n2260), .ZN(
        n2266) );
  OAI21D0BWP12T U2943 ( .A1(n2310), .A2(b[31]), .B(n2264), .ZN(n2265) );
  OAI31D1BWP12T U2944 ( .A1(n2268), .A2(n2267), .A3(n2266), .B(n2265), .ZN(
        n2318) );
  AOI22D0BWP12T U2945 ( .A1(a[22]), .A2(n737), .B1(n2269), .B2(a[25]), .ZN(
        n2274) );
  AOI22D0BWP12T U2946 ( .A1(a[20]), .A2(n2410), .B1(n2406), .B2(n2747), .ZN(
        n2273) );
  AOI22D0BWP12T U2947 ( .A1(a[18]), .A2(n2703), .B1(n2408), .B2(n2725), .ZN(
        n2272) );
  AOI22D0BWP12T U2948 ( .A1(a[16]), .A2(n2270), .B1(n782), .B2(n2609), .ZN(
        n2271) );
  ND4D1BWP12T U2949 ( .A1(n2274), .A2(n2273), .A3(n2272), .A4(n2271), .ZN(
        n2300) );
  AOI22D0BWP12T U2950 ( .A1(a[14]), .A2(n2275), .B1(n2678), .B2(n2679), .ZN(
        n2282) );
  AOI22D1BWP12T U2951 ( .A1(n2308), .A2(n2277), .B1(n2276), .B2(n2626), .ZN(
        n2281) );
  AOI22D0BWP12T U2952 ( .A1(n2900), .A2(n2899), .B1(n2278), .B2(n2643), .ZN(
        n2280) );
  AOI22D0BWP12T U2953 ( .A1(n2594), .A2(n2511), .B1(n2545), .B2(a[8]), .ZN(
        n2279) );
  ND4D1BWP12T U2954 ( .A1(n2282), .A2(n2281), .A3(n2280), .A4(n2279), .ZN(
        n2299) );
  AOI22D1BWP12T U2955 ( .A1(n2574), .A2(n2572), .B1(n2283), .B2(n2301), .ZN(
        n2289) );
  AOI22D0BWP12T U2956 ( .A1(n2527), .A2(n2525), .B1(n2870), .B2(n2871), .ZN(
        n2288) );
  AOI22D0BWP12T U2957 ( .A1(n2620), .A2(n2284), .B1(n471), .B2(n2303), .ZN(
        n2287) );
  AOI22D0BWP12T U2958 ( .A1(n2830), .A2(n2827), .B1(n2285), .B2(n2302), .ZN(
        n2286) );
  ND4D1BWP12T U2959 ( .A1(n2289), .A2(n2288), .A3(n2287), .A4(n2286), .ZN(
        n2298) );
  AOI22D0BWP12T U2960 ( .A1(a[30]), .A2(n2291), .B1(n2290), .B2(a[28]), .ZN(
        n2296) );
  CKND0BWP12T U2961 ( .I(b[26]), .ZN(n2774) );
  AOI22D0BWP12T U2962 ( .A1(a[26]), .A2(n2774), .B1(n2292), .B2(a[29]), .ZN(
        n2295) );
  CKND0BWP12T U2963 ( .I(b[24]), .ZN(n2952) );
  CKND0BWP12T U2964 ( .I(b[27]), .ZN(n2805) );
  AOI22D0BWP12T U2965 ( .A1(a[24]), .A2(n2952), .B1(n2805), .B2(a[27]), .ZN(
        n2294) );
  CKND2D0BWP12T U2966 ( .A1(n2483), .A2(n2482), .ZN(n2293) );
  ND4D1BWP12T U2967 ( .A1(n2296), .A2(n2295), .A3(n2294), .A4(n2293), .ZN(
        n2297) );
  NR4D0BWP12T U2968 ( .A1(n2300), .A2(n2299), .A3(n2298), .A4(n2297), .ZN(
        n2317) );
  ND4D0BWP12T U2969 ( .A1(n2301), .A2(a[8]), .A3(n2900), .A4(n2594), .ZN(n2307) );
  ND4D0BWP12T U2970 ( .A1(a[29]), .A2(a[28]), .A3(a[25]), .A4(a[24]), .ZN(
        n2306) );
  ND4D0BWP12T U2971 ( .A1(n2830), .A2(n2303), .A3(n2482), .A4(n2302), .ZN(
        n2305) );
  ND4D0BWP12T U2972 ( .A1(n2747), .A2(a[22]), .A3(n2725), .A4(a[20]), .ZN(
        n2304) );
  NR4D0BWP12T U2973 ( .A1(n2307), .A2(n2306), .A3(n2305), .A4(n2304), .ZN(
        n2316) );
  ND4D0BWP12T U2974 ( .A1(n2679), .A2(a[16]), .A3(n2643), .A4(n2308), .ZN(
        n2309) );
  NR3D0BWP12T U2975 ( .A1(n2310), .A2(n2309), .A3(n2806), .ZN(n2311) );
  ND4D0BWP12T U2976 ( .A1(n2311), .A2(a[30]), .A3(a[26]), .A4(a[27]), .ZN(
        n2314) );
  ND4D0BWP12T U2977 ( .A1(n2871), .A2(n2620), .A3(n2574), .A4(n2527), .ZN(
        n2313) );
  ND4D0BWP12T U2978 ( .A1(n2609), .A2(a[18]), .A3(a[14]), .A4(n2626), .ZN(
        n2312) );
  NR3D1BWP12T U2979 ( .A1(n2314), .A2(n2313), .A3(n2312), .ZN(n2315) );
  AOI22D1BWP12T U2980 ( .A1(n2318), .A2(n2317), .B1(n2316), .B2(n2315), .ZN(
        n2319) );
  OAI31D1BWP12T U2981 ( .A1(n2322), .A2(n2321), .A3(n2320), .B(n2319), .ZN(
        n2323) );
  AOI31D1BWP12T U2982 ( .A1(n2326), .A2(n2325), .A3(n2324), .B(n2323), .ZN(
        n2327) );
  OAI211D1BWP12T U2983 ( .A1(n2330), .A2(n2329), .B(n2328), .C(n2327), .ZN(
        n2400) );
  FA1D2BWP12T U2984 ( .A(a[27]), .B(b[27]), .CI(n2331), .CO(n1457), .S(n2801)
         );
  FA1D2BWP12T U2985 ( .A(a[26]), .B(b[26]), .CI(n2332), .CO(n2331), .S(n2791)
         );
  FA1D2BWP12T U2986 ( .A(a[24]), .B(b[24]), .CI(n2333), .CO(n727), .S(n2968)
         );
  FA1D2BWP12T U2987 ( .A(n2747), .B(b[23]), .CI(n2334), .CO(n2333), .S(n2742)
         );
  FA1D0BWP12T U2988 ( .A(a[20]), .B(b[20]), .CI(n2336), .CO(n2335), .S(n2934)
         );
  CKND2D0BWP12T U2989 ( .A1(n2338), .A2(n2337), .ZN(n2339) );
  XOR2XD1BWP12T U2990 ( .A1(n2340), .A2(n2339), .Z(n2702) );
  INVD0BWP12T U2991 ( .I(n2352), .ZN(n2354) );
  CKND2D1BWP12T U2992 ( .A1(n2354), .A2(n2353), .ZN(n2356) );
  XOR2XD1BWP12T U2993 ( .A1(n2356), .A2(n2355), .Z(n2489) );
  OR4D0BWP12T U2994 ( .A1(n2489), .A2(n2358), .A3(n2909), .A4(n2357), .Z(n2364) );
  NR4D0BWP12T U2995 ( .A1(n2365), .A2(n2587), .A3(n2364), .A4(n2838), .ZN(
        n2379) );
  NR4D0BWP12T U2996 ( .A1(n2857), .A2(n2553), .A3(n2377), .A4(n2536), .ZN(
        n2378) );
  IND3D1BWP12T U2997 ( .A1(n2380), .B1(n2379), .B2(n2378), .ZN(n2382) );
  OR4D0BWP12T U2998 ( .A1(n2892), .A2(n2506), .A3(n2382), .A4(n2381), .Z(n2384) );
  OR4D0BWP12T U2999 ( .A1(n2386), .A2(n2385), .A3(n2384), .A4(n2383), .Z(n2388) );
  OR4D0BWP12T U3000 ( .A1(n2702), .A2(n2693), .A3(n2388), .A4(n2387), .Z(n2390) );
  OR4D0BWP12T U3001 ( .A1(n2716), .A2(n2934), .A3(n2390), .A4(n2389), .Z(n2392) );
  OR4D1BWP12T U3002 ( .A1(n2968), .A2(n2742), .A3(n2392), .A4(n2391), .Z(n2394) );
  OR4D1BWP12T U3003 ( .A1(n2801), .A2(n2791), .A3(n2394), .A4(n2393), .Z(n2395) );
  NR4D0BWP12T U3004 ( .A1(n2398), .A2(n2397), .A3(n2396), .A4(n2395), .ZN(
        n2399) );
  AO211D1BWP12T U3005 ( .A1(n2603), .A2(n2401), .B(n2400), .C(n2399), .Z(n2465) );
  FA1D1BWP12T U3006 ( .A(a[27]), .B(n2805), .CI(n2402), .CO(n1455), .S(n2817)
         );
  FA1D1BWP12T U3007 ( .A(a[26]), .B(n2774), .CI(n2403), .CO(n2402), .S(n2796)
         );
  FA1D0BWP12T U3008 ( .A(n2952), .B(a[24]), .CI(n2404), .CO(n699), .S(n2939)
         );
  FA1D0BWP12T U3009 ( .A(n2747), .B(n2406), .CI(n2405), .CO(n2404), .S(n2762)
         );
  FA1D1BWP12T U3010 ( .A(n2725), .B(n2408), .CI(n2407), .CO(n736), .S(n2736)
         );
  FA1D1BWP12T U3011 ( .A(n2410), .B(a[20]), .CI(n2409), .CO(n2407), .S(n2926)
         );
  INVD0BWP12T U3012 ( .I(n2440), .ZN(n2419) );
  CKND2D1BWP12T U3013 ( .A1(n1603), .A2(n2421), .ZN(n2423) );
  XOR2XD1BWP12T U3014 ( .A1(n2423), .A2(n2422), .Z(n2491) );
  INVD0BWP12T U3015 ( .I(n2429), .ZN(n2431) );
  ND2D1BWP12T U3016 ( .A1(n1612), .A2(n2433), .ZN(n2434) );
  XNR2D1BWP12T U3017 ( .A1(n2441), .A2(n2434), .ZN(n2867) );
  INVD1BWP12T U3018 ( .I(n2445), .ZN(n2449) );
  NR4D0BWP12T U3019 ( .A1(n2463), .A2(n2462), .A3(n2461), .A4(n2460), .ZN(
        n2464) );
  AOI211D1BWP12T U3020 ( .A1(n2467), .A2(n2466), .B(n2465), .C(n2464), .ZN(
        n2468) );
  OAI211D1BWP12T U3021 ( .A1(n2471), .A2(n2470), .B(n2469), .C(n2468), .ZN(z)
         );
  MAOI22D0BWP12T U3022 ( .A1(n2473), .A2(n2977), .B1(n2472), .B2(n2957), .ZN(
        n2503) );
  INVD1BWP12T U3023 ( .I(n2474), .ZN(n2475) );
  AOI22D1BWP12T U3024 ( .A1(n2855), .A2(n2476), .B1(n2874), .B2(n2475), .ZN(
        n2502) );
  CKND0BWP12T U3025 ( .I(n2893), .ZN(n2873) );
  MUX2ND0BWP12T U3026 ( .I0(n2948), .I1(n2478), .S(n2477), .ZN(n2479) );
  AOI21D0BWP12T U3027 ( .A1(n2479), .A2(n2949), .B(n2481), .ZN(n2486) );
  AOI21D0BWP12T U3028 ( .A1(n2481), .A2(n2480), .B(n2825), .ZN(n2484) );
  OAI22D0BWP12T U3029 ( .A1(n2484), .A2(n2483), .B1(n2482), .B2(n2806), .ZN(
        n2485) );
  AO211D1BWP12T U3030 ( .A1(n2487), .A2(n2940), .B(n2486), .C(n2485), .Z(n2488) );
  TPAOI21D0BWP12T U3031 ( .A1(n2967), .A2(n2489), .B(n2488), .ZN(n2493) );
  AOI22D0BWP12T U3032 ( .A1(n2491), .A2(n2866), .B1(n2490), .B2(n2858), .ZN(
        n2492) );
  OA211D1BWP12T U3033 ( .A1(n2494), .A2(n2873), .B(n2493), .C(n2492), .Z(n2501) );
  NR2D1BWP12T U3034 ( .A1(n2496), .A2(n2495), .ZN(n2498) );
  AOI22D1BWP12T U3035 ( .A1(n2499), .A2(n2498), .B1(n2497), .B2(n2894), .ZN(
        n2500) );
  ND4D1BWP12T U3036 ( .A1(n2503), .A2(n2502), .A3(n2501), .A4(n2500), .ZN(
        result[1]) );
  CKND2D1BWP12T U3037 ( .A1(n2504), .A2(n2977), .ZN(n2521) );
  AOI22D1BWP12T U3038 ( .A1(n2967), .A2(n2506), .B1(n2505), .B2(n2940), .ZN(
        n2520) );
  NR2D1BWP12T U3039 ( .A1(n2508), .A2(n2964), .ZN(n2903) );
  AOI22D1BWP12T U3040 ( .A1(n2855), .A2(n2517), .B1(n2516), .B2(n2866), .ZN(
        n2518) );
  ND4D1BWP12T U3041 ( .A1(n2521), .A2(n2520), .A3(n2519), .A4(n2518), .ZN(
        result[11]) );
  NR2D0BWP12T U3042 ( .A1(n2525), .A2(n2951), .ZN(n2524) );
  AOI211D1BWP12T U3043 ( .A1(n2525), .A2(n2948), .B(n2524), .C(n2825), .ZN(
        n2533) );
  CKND2D1BWP12T U3044 ( .A1(n2526), .A2(n2828), .ZN(n2531) );
  TPOAI21D0BWP12T U3045 ( .A1(n2527), .A2(n2944), .B(n2949), .ZN(n2529) );
  AOI22D0BWP12T U3046 ( .A1(n2947), .A2(n2532), .B1(n2529), .B2(n2528), .ZN(
        n2530) );
  ND2D1BWP12T U3047 ( .A1(n2543), .A2(n2940), .ZN(n2555) );
  NR2D0BWP12T U3048 ( .A1(n2545), .A2(n2951), .ZN(n2544) );
  AOI211D0BWP12T U3049 ( .A1(n2545), .A2(n2948), .B(n2544), .C(n2825), .ZN(
        n2551) );
  CKND2D1BWP12T U3050 ( .A1(n2546), .A2(n2786), .ZN(n2549) );
  OAI21D0BWP12T U3051 ( .A1(a[8]), .A2(n2944), .B(n2949), .ZN(n2547) );
  AOI22D0BWP12T U3052 ( .A1(n2947), .A2(n2550), .B1(n2547), .B2(n2605), .ZN(
        n2548) );
  OAI211D1BWP12T U3053 ( .A1(n2551), .A2(n2550), .B(n2549), .C(n2548), .ZN(
        n2552) );
  AOI21D1BWP12T U3054 ( .A1(n2967), .A2(n2553), .B(n2552), .ZN(n2554) );
  OAI211D1BWP12T U3055 ( .A1(n2556), .A2(n2964), .B(n2555), .C(n2554), .ZN(
        n2566) );
  INVD1BWP12T U3056 ( .I(n2557), .ZN(n2564) );
  AOI22D0BWP12T U3057 ( .A1(n2866), .A2(n2559), .B1(n2558), .B2(n2855), .ZN(
        n2563) );
  AOI22D1BWP12T U3058 ( .A1(n2561), .A2(n2858), .B1(n2886), .B2(n2560), .ZN(
        n2562) );
  OAI211D1BWP12T U3059 ( .A1(n2564), .A2(n2957), .B(n2563), .C(n2562), .ZN(
        n2565) );
  AO211D1BWP12T U3060 ( .A1(n2567), .A2(n2977), .B(n2566), .C(n2565), .Z(
        result[8]) );
  AOI21D0BWP12T U3061 ( .A1(n2569), .A2(n2894), .B(n2893), .ZN(n2584) );
  ND2D0BWP12T U3062 ( .A1(n2570), .A2(n2855), .ZN(n2583) );
  NR2D1BWP12T U3063 ( .A1(n2572), .A2(n2951), .ZN(n2571) );
  AOI211D1BWP12T U3064 ( .A1(n2572), .A2(n2948), .B(n2571), .C(n2825), .ZN(
        n2579) );
  CKND2D1BWP12T U3065 ( .A1(n2573), .A2(n2828), .ZN(n2577) );
  OAI21D0BWP12T U3066 ( .A1(n2574), .A2(n2944), .B(n2949), .ZN(n2575) );
  AOI22D1BWP12T U3067 ( .A1(n2947), .A2(n2578), .B1(n2575), .B2(b[6]), .ZN(
        n2576) );
  OAI211D1BWP12T U3068 ( .A1(n2579), .A2(n2578), .B(n2577), .C(n2576), .ZN(
        n2580) );
  AOI21D1BWP12T U3069 ( .A1(n2581), .A2(n2874), .B(n2580), .ZN(n2582) );
  AOI22D1BWP12T U3070 ( .A1(n2858), .A2(n2588), .B1(n2587), .B2(n2967), .ZN(
        n2589) );
  CKXOR2D0BWP12T U3071 ( .A1(n2925), .A2(n2656), .Z(n2670) );
  CKND2D0BWP12T U3072 ( .A1(n2973), .A2(n2657), .ZN(n2662) );
  MUX2NXD0BWP12T U3073 ( .I0(n2662), .I1(n2922), .S(a[31]), .ZN(n2664) );
  NR2D1BWP12T U3074 ( .A1(n2664), .A2(n2663), .ZN(n2669) );
  NR2D0BWP12T U3075 ( .A1(n2665), .A2(a[31]), .ZN(n2923) );
  XNR2XD1BWP12T U3076 ( .A1(n2923), .A2(n2666), .ZN(n2667) );
  NR2D0BWP12T U3077 ( .A1(n2667), .A2(n2878), .ZN(n2668) );
  AO211D1BWP12T U3078 ( .A1(n2670), .A2(n2977), .B(n2669), .C(n2668), .Z(v) );
  ND2D1BWP12T U3079 ( .A1(n2672), .A2(n2940), .ZN(n2689) );
  INVD1BWP12T U3080 ( .I(n2673), .ZN(n2687) );
  OAI22D0BWP12T U3081 ( .A1(n2676), .A2(n2675), .B1(n2674), .B2(n2718), .ZN(
        n2686) );
  NR2D0BWP12T U3082 ( .A1(n2678), .A2(n2951), .ZN(n2677) );
  AOI211D0BWP12T U3083 ( .A1(n2678), .A2(n2948), .B(n2677), .C(n2825), .ZN(
        n2684) );
  OAI21D0BWP12T U3084 ( .A1(n2679), .A2(n2944), .B(n2949), .ZN(n2680) );
  AOI22D0BWP12T U3085 ( .A1(n2947), .A2(n2683), .B1(n2680), .B2(b[17]), .ZN(
        n2681) );
  OAI211D0BWP12T U3086 ( .A1(n2684), .A2(n2683), .B(n2682), .C(n2681), .ZN(
        n2685) );
  RCAOI211D0BWP12T U3087 ( .A1(n2687), .A2(n2786), .B(n2686), .C(n2685), .ZN(
        n2688) );
  OAI211D1BWP12T U3088 ( .A1(n2690), .A2(n2964), .B(n2689), .C(n2688), .ZN(
        n2691) );
  AOI21D1BWP12T U3089 ( .A1(n2692), .A2(n2866), .B(n2691), .ZN(n2698) );
  AOI22D1BWP12T U3090 ( .A1(n2858), .A2(n2694), .B1(n2693), .B2(n2967), .ZN(
        n2697) );
  CKND2D1BWP12T U3091 ( .A1(n2695), .A2(n2855), .ZN(n2696) );
  ND4D1BWP12T U3092 ( .A1(n2699), .A2(n2698), .A3(n2697), .A4(n2696), .ZN(
        result[17]) );
  INVD1BWP12T U3093 ( .I(n2700), .ZN(n2714) );
  CKND2D1BWP12T U3094 ( .A1(n2711), .A2(n2855), .ZN(n2712) );
  OAI211D1BWP12T U3095 ( .A1(n2822), .A2(n2714), .B(n2713), .C(n2712), .ZN(
        result[18]) );
  INVD1BWP12T U3096 ( .I(n2715), .ZN(n2734) );
  ND2D1BWP12T U3097 ( .A1(n2716), .A2(n2967), .ZN(n2733) );
  NR2D1BWP12T U3098 ( .A1(n2717), .A2(n2964), .ZN(n2730) );
  TPND2D0BWP12T U3099 ( .A1(n2408), .A2(n2948), .ZN(n2721) );
  OAI211D0BWP12T U3100 ( .A1(n2408), .A2(n2951), .B(n2721), .C(n2949), .ZN(
        n2724) );
  OAI21D0BWP12T U3101 ( .A1(n2725), .A2(n2944), .B(n2949), .ZN(n2722) );
  RCAOI211D0BWP12T U3102 ( .A1(n2725), .A2(n2724), .B(n2807), .C(n2723), .ZN(
        n2726) );
  OAI211D1BWP12T U3103 ( .A1(n2942), .A2(n2728), .B(n2727), .C(n2726), .ZN(
        n2729) );
  AOI211D1BWP12T U3104 ( .A1(n2731), .A2(n2940), .B(n2730), .C(n2729), .ZN(
        n2732) );
  OAI211D1BWP12T U3105 ( .A1(n2734), .A2(n2814), .B(n2733), .C(n2732), .ZN(
        n2735) );
  AOI21D1BWP12T U3106 ( .A1(n2866), .A2(n2736), .B(n2735), .ZN(n2739) );
  CKND2D1BWP12T U3107 ( .A1(n2737), .A2(n2855), .ZN(n2738) );
  OAI211D1BWP12T U3108 ( .A1(n2822), .A2(n427), .B(n2739), .C(n2738), .ZN(
        result[21]) );
  INVD1BWP12T U3109 ( .I(n2740), .ZN(n2766) );
  ND2D1BWP12T U3110 ( .A1(n2741), .A2(n2858), .ZN(n2760) );
  ND2D1BWP12T U3111 ( .A1(n2742), .A2(n2967), .ZN(n2759) );
  MOAI22D0BWP12T U3112 ( .A1(n2942), .A2(n2744), .B1(n2743), .B2(n2905), .ZN(
        n2754) );
  TPNR2D0BWP12T U3113 ( .A1(n2406), .A2(n2951), .ZN(n2745) );
  AOI211XD0BWP12T U3114 ( .A1(n2406), .A2(n2948), .B(n2745), .C(n2825), .ZN(
        n2752) );
  TPND2D0BWP12T U3115 ( .A1(n2746), .A2(n2932), .ZN(n2750) );
  OAI21D0BWP12T U3116 ( .A1(n2747), .A2(n2944), .B(n2949), .ZN(n2748) );
  AOI22D0BWP12T U3117 ( .A1(n2947), .A2(n2751), .B1(n2748), .B2(b[23]), .ZN(
        n2749) );
  OAI211D0BWP12T U3118 ( .A1(n2752), .A2(n2751), .B(n2750), .C(n2749), .ZN(
        n2753) );
  AOI211D1BWP12T U3119 ( .A1(n2894), .A2(n2755), .B(n2754), .C(n2753), .ZN(
        n2758) );
  ND2D1BWP12T U3120 ( .A1(n2756), .A2(n2940), .ZN(n2757) );
  ND4D1BWP12T U3121 ( .A1(n2760), .A2(n2759), .A3(n2758), .A4(n2757), .ZN(
        n2761) );
  AOI21D1BWP12T U3122 ( .A1(n2866), .A2(n2762), .B(n2761), .ZN(n2765) );
  CKND2D1BWP12T U3123 ( .A1(n2763), .A2(n2855), .ZN(n2764) );
  OAI211D1BWP12T U3124 ( .A1(n2822), .A2(n2766), .B(n2765), .C(n2764), .ZN(
        result[23]) );
  INVD1BWP12T U3125 ( .I(n2767), .ZN(n2798) );
  INVD1BWP12T U3126 ( .I(n2768), .ZN(n2794) );
  CKND2D1BWP12T U3127 ( .A1(n2770), .A2(n2769), .ZN(n2771) );
  AOI21D1BWP12T U3128 ( .A1(n2772), .A2(n2771), .B(n2964), .ZN(n2789) );
  TPNR2D0BWP12T U3129 ( .A1(n2774), .A2(n2951), .ZN(n2773) );
  RCAOI211D0BWP12T U3130 ( .A1(n2774), .A2(n2948), .B(n2773), .C(n2825), .ZN(
        n2780) );
  CKND2D0BWP12T U3131 ( .A1(n2895), .A2(n2775), .ZN(n2778) );
  OAI21D0BWP12T U3132 ( .A1(a[26]), .A2(n2944), .B(n2949), .ZN(n2776) );
  AOI22D0BWP12T U3133 ( .A1(n2947), .A2(n2779), .B1(n2776), .B2(b[26]), .ZN(
        n2777) );
  OAI211D1BWP12T U3134 ( .A1(n2780), .A2(n2779), .B(n2778), .C(n2777), .ZN(
        n2785) );
  OA21D1BWP12T U3135 ( .A1(n2783), .A2(n2782), .B(n2781), .Z(n2784) );
  AO211D1BWP12T U3136 ( .A1(n2787), .A2(n2786), .B(n2785), .C(n2784), .Z(n2788) );
  AOI211D1BWP12T U3137 ( .A1(n2790), .A2(n2940), .B(n2789), .C(n2788), .ZN(
        n2793) );
  ND2D1BWP12T U3138 ( .A1(n2791), .A2(n2967), .ZN(n2792) );
  OAI211D1BWP12T U3139 ( .A1(n2814), .A2(n2794), .B(n2793), .C(n2792), .ZN(
        n2795) );
  INVD1BWP12T U3140 ( .I(n2799), .ZN(n2821) );
  INVD1BWP12T U3141 ( .I(n2800), .ZN(n2815) );
  ND2D1BWP12T U3142 ( .A1(n2801), .A2(n2967), .ZN(n2813) );
  NR2D1BWP12T U3143 ( .A1(n2802), .A2(n2964), .ZN(n2810) );
  AOI211D1BWP12T U3144 ( .A1(n2811), .A2(n2940), .B(n2810), .C(n2809), .ZN(
        n2812) );
  OAI211D1BWP12T U3145 ( .A1(n2815), .A2(n2814), .B(n2813), .C(n2812), .ZN(
        n2816) );
  AOI21D1BWP12T U3146 ( .A1(n2866), .A2(n2817), .B(n2816), .ZN(n2820) );
  ND2D1BWP12T U3147 ( .A1(n2818), .A2(n2855), .ZN(n2819) );
  OAI211D1BWP12T U3148 ( .A1(n2822), .A2(n2821), .B(n2820), .C(n2819), .ZN(
        result[27]) );
  INVD1BWP12T U3149 ( .I(n2823), .ZN(n2841) );
  ND2D0BWP12T U3150 ( .A1(n2824), .A2(n2855), .ZN(n2840) );
  TPNR2D0BWP12T U3151 ( .A1(n2827), .A2(n2951), .ZN(n2826) );
  AOI211XD0BWP12T U3152 ( .A1(n2827), .A2(n2948), .B(n2826), .C(n2825), .ZN(
        n2836) );
  CKND2D1BWP12T U3153 ( .A1(n2829), .A2(n2828), .ZN(n2834) );
  TPOAI21D0BWP12T U3154 ( .A1(n2830), .A2(n2944), .B(n2949), .ZN(n2832) );
  AOI22D0BWP12T U3155 ( .A1(n2947), .A2(n2835), .B1(n2832), .B2(n2831), .ZN(
        n2833) );
  OAI211D1BWP12T U3156 ( .A1(n2836), .A2(n2835), .B(n2834), .C(n2833), .ZN(
        n2837) );
  AOI21D1BWP12T U3157 ( .A1(n2967), .A2(n2838), .B(n2837), .ZN(n2839) );
  OAI211D1BWP12T U3158 ( .A1(n2842), .A2(n2841), .B(n2840), .C(n2839), .ZN(
        n2851) );
  INVD1BWP12T U3159 ( .I(n2843), .ZN(n2849) );
  AOI22D1BWP12T U3160 ( .A1(n2940), .A2(n2845), .B1(n2874), .B2(n2844), .ZN(
        n2848) );
  CKND2D1BWP12T U3161 ( .A1(n2846), .A2(n2858), .ZN(n2847) );
  OAI211D1BWP12T U3162 ( .A1(n2973), .A2(n2849), .B(n2848), .C(n2847), .ZN(
        n2850) );
  AOI211D1BWP12T U3163 ( .A1(n2905), .A2(n2852), .B(n2851), .C(n2850), .ZN(
        n2853) );
  IOA21D1BWP12T U3164 ( .A1(n2854), .A2(n2977), .B(n2853), .ZN(result[3]) );
  CKND2D0BWP12T U3165 ( .A1(n2856), .A2(n2855), .ZN(n2865) );
  AOI22D0BWP12T U3166 ( .A1(n2859), .A2(n2858), .B1(n2857), .B2(n2967), .ZN(
        n2864) );
  ND2D1BWP12T U3167 ( .A1(n2860), .A2(n2886), .ZN(n2863) );
  ND2D1BWP12T U3168 ( .A1(n2861), .A2(n2894), .ZN(n2862) );
  ND4D1BWP12T U3169 ( .A1(n2865), .A2(n2864), .A3(n2863), .A4(n2862), .ZN(
        n2880) );
  ND2XD0BWP12T U3170 ( .A1(n2867), .A2(n2866), .ZN(n2877) );
  OAI211D1BWP12T U3171 ( .A1(n426), .A2(n2878), .B(n2877), .C(n2876), .ZN(
        n2879) );
  AOI211D1BWP12T U3172 ( .A1(n2905), .A2(n2881), .B(n2880), .C(n2879), .ZN(
        n2882) );
  IOA21D1BWP12T U3173 ( .A1(n2883), .A2(n2977), .B(n2882), .ZN(result[4]) );
  INVD1BWP12T U3174 ( .I(n2884), .ZN(n2891) );
  AOI22D1BWP12T U3175 ( .A1(n2887), .A2(n2940), .B1(n2886), .B2(n2885), .ZN(
        n2890) );
  CKND2D1BWP12T U3176 ( .A1(n2888), .A2(n2858), .ZN(n2889) );
  OAI211D1BWP12T U3177 ( .A1(n2973), .A2(n2891), .B(n2890), .C(n2889), .ZN(
        n2912) );
  INVD1BWP12T U3178 ( .I(n2892), .ZN(n2910) );
  ND2D1BWP12T U3179 ( .A1(n2906), .A2(n2905), .ZN(n2907) );
  OAI211D1BWP12T U3180 ( .A1(n2910), .A2(n2909), .B(n2908), .C(n2907), .ZN(
        n2911) );
  AOI211D1BWP12T U3181 ( .A1(n2855), .A2(n2913), .B(n2912), .C(n2911), .ZN(
        n2914) );
  IOA21D1BWP12T U3182 ( .A1(n2915), .A2(n2977), .B(n2914), .ZN(result[10]) );
  INVD1BWP12T U3183 ( .I(n2917), .ZN(n2920) );
  AO22D1BWP12T U3184 ( .A1(n2920), .A2(n2967), .B1(n2858), .B2(n2919), .Z(
        n2921) );
  AOI211D1BWP12T U3185 ( .A1(n2940), .A2(n2923), .B(n2922), .C(n2921), .ZN(
        n2924) );
  IOA21D1BWP12T U3186 ( .A1(n2925), .A2(n2977), .B(n2924), .ZN(c_out) );
  INVD1BWP12T U3187 ( .I(n2939), .ZN(n2972) );
  ND2D1BWP12T U3188 ( .A1(n2941), .A2(n2940), .ZN(n2963) );
  NR2D1BWP12T U3189 ( .A1(n2943), .A2(n2942), .ZN(n2959) );
  OAI21D0BWP12T U3190 ( .A1(a[24]), .A2(n2944), .B(n2949), .ZN(n2945) );
  AOI22D0BWP12T U3191 ( .A1(n2947), .A2(n2946), .B1(n2945), .B2(b[24]), .ZN(
        n2955) );
  TPND2D0BWP12T U3192 ( .A1(n2952), .A2(n2948), .ZN(n2950) );
  OAI211D0BWP12T U3193 ( .A1(n2952), .A2(n2951), .B(n2950), .C(n2949), .ZN(
        n2953) );
  CKND2D0BWP12T U3194 ( .A1(n2953), .A2(a[24]), .ZN(n2954) );
  OAI211D1BWP12T U3195 ( .A1(n2957), .A2(n2956), .B(n2955), .C(n2954), .ZN(
        n2958) );
  RCAOI211D0BWP12T U3196 ( .A1(n2961), .A2(n2960), .B(n2959), .C(n2958), .ZN(
        n2962) );
  OAI211D1BWP12T U3197 ( .A1(n2965), .A2(n2964), .B(n2963), .C(n2962), .ZN(
        n2966) );
  AOI21D1BWP12T U3198 ( .A1(n2968), .A2(n2967), .B(n2966), .ZN(n2971) );
  ND2D1BWP12T U3199 ( .A1(n2969), .A2(n2858), .ZN(n2970) );
  OAI211D1BWP12T U3200 ( .A1(n2973), .A2(n2972), .B(n2971), .C(n2970), .ZN(
        n2974) );
  AOI21D1BWP12T U3201 ( .A1(n2855), .A2(n2975), .B(n2974), .ZN(n2976) );
  IOA21D1BWP12T U3202 ( .A1(n2978), .A2(n2977), .B(n2976), .ZN(result[24]) );
  CMPE42D1BWP12T U3203 ( .A(mult_x_18_n892), .B(mult_x_18_n869), .C(
        mult_x_18_n917), .CIX(mult_x_18_n674), .D(mult_x_18_n677), .CO(
        mult_x_18_n667), .COX(mult_x_18_n666), .S(mult_x_18_n668) );
  CMPE42D1BWP12T U3204 ( .A(mult_x_18_n846), .B(mult_x_18_n867), .C(
        mult_x_18_n890), .CIX(mult_x_18_n656), .D(mult_x_18_n915), .CO(
        mult_x_18_n648), .COX(mult_x_18_n647), .S(mult_x_18_n649) );
  CMPE42D1BWP12T U3205 ( .A(mult_x_18_n843), .B(mult_x_18_n824), .C(
        mult_x_18_n631), .CIX(mult_x_18_n628), .D(mult_x_18_n619), .CO(
        mult_x_18_n613), .COX(mult_x_18_n612), .S(mult_x_18_n614) );
  CMPE42D1BWP12T U3206 ( .A(mult_x_18_n532), .B(mult_x_18_n551), .C(
        mult_x_18_n548), .CIX(mult_x_18_n541), .D(mult_x_18_n545), .CO(
        mult_x_18_n525), .COX(mult_x_18_n524), .S(mult_x_18_n526) );
  CMPE42D1BWP12T U3207 ( .A(mult_x_18_n552), .B(mult_x_18_n774), .C(
        mult_x_18_n549), .CIX(mult_x_18_n563), .D(mult_x_18_n546), .CO(
        mult_x_18_n542), .COX(mult_x_18_n541), .S(mult_x_18_n543) );
  CMPE42D1BWP12T U3208 ( .A(mult_x_18_n582), .B(mult_x_18_n789), .C(
        mult_x_18_n586), .CIX(mult_x_18_n577), .D(mult_x_18_n580), .CO(
        mult_x_18_n573), .COX(mult_x_18_n572), .S(mult_x_18_n574) );
  CMPE42D1BWP12T U3209 ( .A(mult_x_18_n772), .B(mult_x_18_n857), .C(
        mult_x_18_n785), .CIX(mult_x_18_n533), .D(mult_x_18_n520), .CO(
        mult_x_18_n511), .COX(mult_x_18_n510), .S(mult_x_18_n512) );
  CMPE42D1BWP12T U3210 ( .A(mult_x_18_n783), .B(mult_x_18_n759), .C(
        mult_x_18_n930), .CIX(mult_x_18_n494), .D(mult_x_18_n815), .CO(
        mult_x_18_n477), .COX(mult_x_18_n476), .S(mult_x_18_n478) );
  CMPE42D1BWP12T U3211 ( .A(mult_x_18_n375), .B(mult_x_18_n378), .C(
        mult_x_18_n372), .CIX(mult_x_18_n387), .D(mult_x_18_n400), .CO(
        mult_x_18_n365), .COX(mult_x_18_n364), .S(mult_x_18_n366) );
  CMPE42D1BWP12T U3212 ( .A(mult_x_18_n418), .B(mult_x_18_n421), .C(
        mult_x_18_n415), .CIX(mult_x_18_n408), .D(mult_x_18_n411), .CO(
        mult_x_18_n388), .COX(mult_x_18_n387), .S(mult_x_18_n389) );
  CMPE42D1BWP12T U3213 ( .A(mult_x_18_n463), .B(mult_x_18_n438), .C(
        mult_x_18_n457), .CIX(mult_x_18_n435), .D(mult_x_18_n460), .CO(
        mult_x_18_n431), .COX(mult_x_18_n430), .S(mult_x_18_n432) );
  CMPE42D1BWP12T U3214 ( .A(mult_x_18_n443), .B(mult_x_18_n416), .C(
        mult_x_18_n440), .CIX(mult_x_18_n434), .D(mult_x_18_n433), .CO(
        mult_x_18_n409), .COX(mult_x_18_n408), .S(mult_x_18_n410) );
  CMPE42D1BWP12T U3215 ( .A(mult_x_18_n480), .B(mult_x_18_n458), .C(
        mult_x_18_n477), .CIX(mult_x_18_n470), .D(mult_x_18_n474), .CO(
        mult_x_18_n451), .COX(mult_x_18_n450), .S(mult_x_18_n452) );
  CMPE42D1BWP12T U3216 ( .A(mult_x_18_n495), .B(mult_x_18_n481), .C(
        mult_x_18_n498), .CIX(mult_x_18_n488), .D(mult_x_18_n475), .CO(
        mult_x_18_n471), .COX(mult_x_18_n470), .S(mult_x_18_n472) );
  CMPE42D1BWP12T U3217 ( .A(mult_x_18_n738), .B(mult_x_18_n754), .C(
        mult_x_18_n850), .CIX(mult_x_18_n402), .D(mult_x_18_n745), .CO(
        mult_x_18_n371), .COX(mult_x_18_n370), .S(mult_x_18_n372) );
  CMPE42D1BWP12T U3218 ( .A(mult_x_18_n830), .B(mult_x_18_n734), .C(
        mult_x_18_n899), .CIX(mult_x_18_n414), .D(mult_x_18_n955), .CO(
        mult_x_18_n400), .COX(mult_x_18_n399), .S(mult_x_18_n401) );
  CMPE42D1BWP12T U3219 ( .A(mult_x_18_n831), .B(mult_x_18_n795), .C(
        mult_x_18_n900), .CIX(mult_x_18_n436), .D(mult_x_18_n426), .CO(
        mult_x_18_n421), .COX(mult_x_18_n420), .S(mult_x_18_n422) );
  CMPE42D1BWP12T U3220 ( .A(mult_x_18_n883), .B(mult_x_18_n775), .C(
        mult_x_18_n908), .CIX(mult_x_18_n575), .D(mult_x_18_n568), .CO(
        mult_x_18_n563), .COX(mult_x_18_n562), .S(mult_x_18_n564) );
  CMPE42D1BWP12T U3221 ( .A(mult_x_18_n838), .B(mult_x_18_n802), .C(
        mult_x_18_n907), .CIX(mult_x_18_n559), .D(mult_x_18_n963), .CO(
        mult_x_18_n548), .COX(mult_x_18_n547), .S(mult_x_18_n549) );
  CMPE42D1BWP12T U3222 ( .A(mult_x_18_n446), .B(mult_x_18_n853), .C(
        mult_x_18_n453), .CIX(mult_x_18_n441), .D(mult_x_18_n444), .CO(
        mult_x_18_n434), .COX(mult_x_18_n433), .S(mult_x_18_n435) );
  CMPE42D1BWP12T U3223 ( .A(mult_x_18_n1006), .B(mult_x_18_n871), .C(
        mult_x_18_n894), .CIX(mult_x_18_n688), .D(mult_x_18_n690), .CO(
        mult_x_18_n683), .COX(mult_x_18_n682), .S(mult_x_18_n684) );
  CMPE42D1BWP12T U3224 ( .A(mult_x_18_n928), .B(mult_x_18_n757), .C(
        mult_x_18_n813), .CIX(mult_x_18_n459), .D(mult_x_18_n901), .CO(
        mult_x_18_n440), .COX(mult_x_18_n439), .S(mult_x_18_n441) );
  CMPE42D1BWP12T U3225 ( .A(mult_x_18_n833), .B(mult_x_18_n758), .C(
        mult_x_18_n958), .CIX(mult_x_18_n473), .D(mult_x_18_n466), .CO(
        mult_x_18_n463), .COX(mult_x_18_n462), .S(mult_x_18_n464) );
  CMPE42D1BWP12T U3226 ( .A(mult_x_18_n910), .B(mult_x_18_n862), .C(
        mult_x_18_n966), .CIX(mult_x_18_n600), .D(mult_x_18_n596), .CO(
        mult_x_18_n593), .COX(mult_x_18_n592), .S(mult_x_18_n594) );
  CMPE42D1BWP12T U3227 ( .A(mult_x_18_n990), .B(mult_x_18_n743), .C(
        mult_x_18_n959), .CIX(mult_x_18_n500), .D(mult_x_18_n502), .CO(
        mult_x_18_n483), .COX(mult_x_18_n482), .S(mult_x_18_n484) );
  CMPE42D1BWP12T U3228 ( .A(mult_x_18_n566), .B(mult_x_18_n581), .C(
        mult_x_18_n564), .CIX(mult_x_18_n572), .D(mult_x_18_n561), .CO(
        mult_x_18_n557), .COX(mult_x_18_n556), .S(mult_x_18_n558) );
  CMPE42D1BWP12T U3229 ( .A(mult_x_18_n531), .B(mult_x_18_n518), .C(
        mult_x_18_n528), .CIX(mult_x_18_n524), .D(mult_x_18_n512), .CO(
        mult_x_18_n508), .COX(mult_x_18_n507), .S(mult_x_18_n509) );
  CMPE42D1BWP12T U3230 ( .A(mult_x_18_n837), .B(mult_x_18_n717), .C(
        mult_x_18_n962), .CIX(mult_x_18_n544), .D(mult_x_18_n537), .CO(
        mult_x_18_n534), .COX(mult_x_18_n533), .S(mult_x_18_n535) );
  CMPE42D1BWP12T U3231 ( .A(mult_x_18_n721), .B(mult_x_18_n826), .C(
        mult_x_18_n845), .CIX(mult_x_18_n650), .D(mult_x_18_n889), .CO(
        mult_x_18_n637), .COX(mult_x_18_n636), .S(mult_x_18_n638) );
  CMPE42D1BWP12T U3232 ( .A(mult_x_18_n879), .B(mult_x_18_n751), .C(
        mult_x_18_n904), .CIX(mult_x_18_n510), .D(mult_x_18_n503), .CO(
        mult_x_18_n498), .COX(mult_x_18_n497), .S(mult_x_18_n499) );
  CMPE42D1BWP12T U3233 ( .A(mult_x_18_n918), .B(mult_x_18_n870), .C(
        mult_x_18_n974), .CIX(mult_x_18_n679), .D(mult_x_18_n678), .CO(
        mult_x_18_n675), .COX(mult_x_18_n674), .S(mult_x_18_n676) );
  CMPE42D1BWP12T U3234 ( .A(mult_x_18_n891), .B(mult_x_18_n847), .C(
        mult_x_18_n916), .CIX(mult_x_18_n666), .D(mult_x_18_n669), .CO(
        mult_x_18_n657), .COX(mult_x_18_n656), .S(mult_x_18_n658) );
  CMPE42D1BWP12T U3235 ( .A(mult_x_18_n893), .B(mult_x_18_n945), .C(
        mult_x_18_n682), .CIX(mult_x_18_n676), .D(mult_x_18_n683), .CO(
        mult_x_18_n672), .COX(mult_x_18_n671), .S(mult_x_18_n673) );
  CMPE42D1BWP12T U3236 ( .A(mult_x_18_n851), .B(mult_x_18_n755), .C(
        mult_x_18_n746), .CIX(mult_x_18_n420), .D(mult_x_18_n766), .CO(
        mult_x_18_n394), .COX(mult_x_18_n393), .S(mult_x_18_n395) );
  CMPE42D1BWP12T U3237 ( .A(mult_x_18_n936), .B(mult_x_18_n861), .C(
        mult_x_18_n821), .CIX(mult_x_18_n592), .D(mult_x_18_n884), .CO(
        mult_x_18_n576), .COX(mult_x_18_n575), .S(mult_x_18_n577) );
  CMPE42D1BWP12T U3238 ( .A(mult_x_18_n773), .B(mult_x_18_n858), .C(
        mult_x_18_n786), .CIX(mult_x_18_n550), .D(mult_x_18_n933), .CO(
        mult_x_18_n528), .COX(mult_x_18_n527), .S(mult_x_18_n529) );
  CMPE42D1BWP12T U3239 ( .A(mult_x_18_n935), .B(mult_x_18_n788), .C(
        mult_x_18_n820), .CIX(mult_x_18_n578), .D(mult_x_18_n839), .CO(
        mult_x_18_n560), .COX(mult_x_18_n559), .S(mult_x_18_n561) );
  CMPE42D1BWP12T U3240 ( .A(mult_x_18_n825), .B(mult_x_18_n940), .C(
        mult_x_18_n844), .CIX(mult_x_18_n639), .D(mult_x_18_n632), .CO(
        mult_x_18_n626), .COX(mult_x_18_n625), .S(mult_x_18_n627) );
  CMPE42D1BWP12T U3241 ( .A(mult_x_18_n381), .B(mult_x_18_n403), .C(
        mult_x_18_n397), .CIX(mult_x_18_n390), .D(mult_x_18_n394), .CO(
        mult_x_18_n368), .COX(mult_x_18_n367), .S(mult_x_18_n369) );
  CMPE42D1BWP12T U3242 ( .A(mult_x_18_n424), .B(mult_x_18_n445), .C(
        mult_x_18_n422), .CIX(mult_x_18_n437), .D(mult_x_18_n419), .CO(
        mult_x_18_n412), .COX(mult_x_18_n411), .S(mult_x_18_n413) );
  CMPE42D1BWP12T U3243 ( .A(mult_x_18_n749), .B(mult_x_18_n854), .C(
        mult_x_18_n482), .CIX(mult_x_18_n464), .D(mult_x_18_n483), .CO(
        mult_x_18_n454), .COX(mult_x_18_n453), .S(mult_x_18_n455) );
  CMPE42D1BWP12T U3244 ( .A(mult_x_18_n818), .B(mult_x_18_n762), .C(
        mult_x_18_n881), .CIX(mult_x_18_n547), .D(mult_x_18_n906), .CO(
        mult_x_18_n531), .COX(mult_x_18_n530), .S(mult_x_18_n532) );
  CMPE42D1BWP12T U3245 ( .A(mult_x_18_n765), .B(mult_x_18_n793), .C(
        mult_x_18_n778), .CIX(mult_x_18_n399), .D(mult_x_18_n925), .CO(
        mult_x_18_n374), .COX(mult_x_18_n373), .S(mult_x_18_n375) );
  CMPE42D1BWP12T U3246 ( .A(mult_x_18_n994), .B(mult_x_18_n763), .C(
        mult_x_18_n819), .CIX(mult_x_18_n565), .D(mult_x_18_n567), .CO(
        mult_x_18_n551), .COX(mult_x_18_n550), .S(mult_x_18_n552) );
  CMPE42D1BWP12T U3247 ( .A(mult_x_18_n986), .B(mult_x_18_n731), .C(
        mult_x_18_n874), .CIX(mult_x_18_n423), .D(mult_x_18_n425), .CO(
        mult_x_18_n403), .COX(mult_x_18_n402), .S(mult_x_18_n404) );
  CMPE42D1BWP12T U3248 ( .A(mult_x_18_n829), .B(mult_x_18_n730), .C(
        mult_x_18_n954), .CIX(mult_x_18_n393), .D(mult_x_18_n383), .CO(
        mult_x_18_n380), .COX(mult_x_18_n379), .S(mult_x_18_n381) );
  CMPE42D1BWP12T U3249 ( .A(mult_x_18_n914), .B(mult_x_18_n941), .C(
        mult_x_18_n970), .CIX(mult_x_18_n647), .D(mult_x_18_n643), .CO(
        mult_x_18_n640), .COX(mult_x_18_n639), .S(mult_x_18_n641) );
  CMPE42D1BWP12T U3250 ( .A(mult_x_18_n1002), .B(mult_x_18_n827), .C(
        mult_x_18_n971), .CIX(mult_x_18_n659), .D(mult_x_18_n661), .CO(
        mult_x_18_n651), .COX(mult_x_18_n650), .S(mult_x_18_n652) );
  CMPE42D1BWP12T U3251 ( .A(mult_x_18_n404), .B(mult_x_18_n739), .C(
        mult_x_18_n401), .CIX(mult_x_18_n395), .D(mult_x_18_n398), .CO(
        mult_x_18_n391), .COX(mult_x_18_n390), .S(mult_x_18_n392) );
  CMPE42D1BWP12T U3252 ( .A(mult_x_18_n822), .B(mult_x_18_n790), .C(
        mult_x_18_n841), .CIX(mult_x_18_n603), .D(mult_x_18_n885), .CO(
        mult_x_18_n590), .COX(mult_x_18_n589), .S(mult_x_18_n591) );
  CMPE42D1BWP12T U3253 ( .A(mult_x_18_n747), .B(mult_x_18_n852), .C(
        mult_x_18_n767), .CIX(mult_x_18_n442), .D(mult_x_18_n780), .CO(
        mult_x_18_n415), .COX(mult_x_18_n414), .S(mult_x_18_n416) );
  CMPE42D1BWP12T U3254 ( .A(mult_x_18_n748), .B(mult_x_18_n741), .C(
        mult_x_18_n768), .CIX(mult_x_18_n462), .D(mult_x_18_n781), .CO(
        mult_x_18_n437), .COX(mult_x_18_n436), .S(mult_x_18_n438) );
  CMPE42D1BWP12T U3255 ( .A(mult_x_18_n769), .B(mult_x_18_n715), .C(
        mult_x_18_n782), .CIX(mult_x_18_n479), .D(mult_x_18_n929), .CO(
        mult_x_18_n457), .COX(mult_x_18_n456), .S(mult_x_18_n458) );
  CMPE42D1BWP12T U3256 ( .A(mult_x_18_n834), .B(mult_x_18_n798), .C(
        mult_x_18_n878), .CIX(mult_x_18_n497), .D(mult_x_18_n903), .CO(
        mult_x_18_n480), .COX(mult_x_18_n479), .S(mult_x_18_n481) );
  CMPE42D1BWP12T U3257 ( .A(mult_x_18_n810), .B(mult_x_18_n733), .C(
        mult_x_18_n873), .CIX(mult_x_18_n396), .D(mult_x_18_n898), .CO(
        mult_x_18_n377), .COX(mult_x_18_n376), .S(mult_x_18_n378) );
  CMPE42D1BWP12T U3258 ( .A(mult_x_18_n836), .B(mult_x_18_n800), .C(
        mult_x_18_n905), .CIX(mult_x_18_n527), .D(mult_x_18_n536), .CO(
        mult_x_18_n517), .COX(mult_x_18_n516), .S(mult_x_18_n518) );
  CMPE42D1BWP12T U3259 ( .A(mult_x_18_n814), .B(mult_x_18_n742), .C(
        mult_x_18_n877), .CIX(mult_x_18_n476), .D(mult_x_18_n902), .CO(
        mult_x_18_n460), .COX(mult_x_18_n459), .S(mult_x_18_n461) );
  CMPE42D1BWP12T U3260 ( .A(mult_x_18_n369), .B(mult_x_18_n391), .C(
        mult_x_18_n366), .CIX(mult_x_18_n384), .D(mult_x_18_n388), .CO(
        mult_x_18_n362), .COX(mult_x_18_n361), .S(mult_x_18_n363) );
  CMPE42D1BWP12T U3261 ( .A(mult_x_18_n412), .B(mult_x_18_n392), .C(
        mult_x_18_n389), .CIX(mult_x_18_n405), .D(mult_x_18_n409), .CO(
        mult_x_18_n385), .COX(mult_x_18_n384), .S(mult_x_18_n386) );
  CMPE42D1BWP12T U3262 ( .A(mult_x_18_n413), .B(mult_x_18_n430), .C(
        mult_x_18_n410), .CIX(mult_x_18_n427), .D(mult_x_18_n431), .CO(
        mult_x_18_n406), .COX(mult_x_18_n405), .S(mult_x_18_n407) );
  CMPE42D1BWP12T U3263 ( .A(mult_x_18_n450), .B(mult_x_18_n454), .C(
        mult_x_18_n432), .CIX(mult_x_18_n447), .D(mult_x_18_n451), .CO(
        mult_x_18_n428), .COX(mult_x_18_n427), .S(mult_x_18_n429) );
  CMPE42D1BWP12T U3264 ( .A(mult_x_18_n937), .B(mult_x_18_n719), .C(
        mult_x_18_n606), .CIX(mult_x_18_n594), .D(mult_x_18_n607), .CO(
        mult_x_18_n587), .COX(mult_x_18_n586), .S(mult_x_18_n588) );
  CMPE42D1BWP12T U3265 ( .A(mult_x_18_n784), .B(mult_x_18_n771), .C(
        mult_x_18_n519), .CIX(mult_x_18_n516), .D(mult_x_18_n501), .CO(
        mult_x_18_n492), .COX(mult_x_18_n491), .S(mult_x_18_n493) );
  CMPE42D1BWP12T U3266 ( .A(mult_x_18_n927), .B(mult_x_18_n740), .C(
        mult_x_18_n812), .CIX(mult_x_18_n439), .D(mult_x_18_n875), .CO(
        mult_x_18_n418), .COX(mult_x_18_n417), .S(mult_x_18_n419) );
  CMPE42D1BWP12T U3267 ( .A(mult_x_18_n750), .B(mult_x_18_n855), .C(
        mult_x_18_n770), .CIX(mult_x_18_n484), .D(mult_x_18_n491), .CO(
        mult_x_18_n474), .COX(mult_x_18_n473), .S(mult_x_18_n475) );
  CMPE42D1BWP12T U3268 ( .A(mult_x_18_n840), .B(mult_x_18_n804), .C(
        mult_x_18_n909), .CIX(mult_x_18_n589), .D(mult_x_18_n595), .CO(
        mult_x_18_n579), .COX(mult_x_18_n578), .S(mult_x_18_n580) );
  CMPE42D1BWP12T U3269 ( .A(mult_x_18_n832), .B(mult_x_18_n796), .C(
        mult_x_18_n957), .CIX(mult_x_18_n456), .D(mult_x_18_n465), .CO(
        mult_x_18_n443), .COX(mult_x_18_n442), .S(mult_x_18_n444) );
  CMPE42D1BWP12T U3270 ( .A(mult_x_18_n779), .B(mult_x_18_n794), .C(
        mult_x_18_n926), .CIX(mult_x_18_n417), .D(mult_x_18_n811), .CO(
        mult_x_18_n397), .COX(mult_x_18_n396), .S(mult_x_18_n398) );
  CMPE42D1BWP12T U3271 ( .A(mult_x_18_n787), .B(mult_x_18_n859), .C(
        mult_x_18_n934), .CIX(mult_x_18_n562), .D(mult_x_18_n882), .CO(
        mult_x_18_n545), .COX(mult_x_18_n544), .S(mult_x_18_n546) );
  CMPE42D1BWP12T U3272 ( .A(mult_x_18_n492), .B(mult_x_18_n478), .C(
        mult_x_18_n472), .CIX(mult_x_18_n485), .D(mult_x_18_n489), .CO(
        mult_x_18_n468), .COX(mult_x_18_n467), .S(mult_x_18_n469) );
  CMPE42D1BWP12T U3273 ( .A(mult_x_18_n576), .B(mult_x_18_n579), .C(
        mult_x_18_n573), .CIX(mult_x_18_n558), .D(mult_x_18_n569), .CO(
        mult_x_18_n554), .COX(mult_x_18_n553), .S(mult_x_18_n555) );
  CMPE42D1BWP12T U3274 ( .A(mult_x_18_n590), .B(mult_x_18_n593), .C(
        mult_x_18_n587), .CIX(mult_x_18_n574), .D(mult_x_18_n583), .CO(
        mult_x_18_n570), .COX(mult_x_18_n569), .S(mult_x_18_n571) );
  CMPE42D1BWP12T U3275 ( .A(mult_x_18_n455), .B(mult_x_18_n461), .C(
        mult_x_18_n452), .CIX(mult_x_18_n467), .D(mult_x_18_n471), .CO(
        mult_x_18_n448), .COX(mult_x_18_n447), .S(mult_x_18_n449) );
  CMPE42D1BWP12T U3276 ( .A(mult_x_18_n641), .B(mult_x_18_n651), .C(
        mult_x_18_n638), .CIX(mult_x_18_n644), .D(mult_x_18_n648), .CO(
        mult_x_18_n634), .COX(mult_x_18_n633), .S(mult_x_18_n635) );
  CMPE42D1BWP12T U3277 ( .A(mult_x_18_n640), .B(mult_x_18_n630), .C(
        mult_x_18_n637), .CIX(mult_x_18_n633), .D(mult_x_18_n627), .CO(
        mult_x_18_n623), .COX(mult_x_18_n622), .S(mult_x_18_n624) );
  CMPE42D1BWP12T U3278 ( .A(mult_x_18_n556), .B(mult_x_18_n560), .C(
        mult_x_18_n543), .CIX(mult_x_18_n553), .D(mult_x_18_n557), .CO(
        mult_x_18_n539), .COX(mult_x_18_n538), .S(mult_x_18_n540) );
  CMPE42D1BWP12T U3279 ( .A(mult_x_18_n529), .B(mult_x_18_n535), .C(
        mult_x_18_n542), .CIX(mult_x_18_n538), .D(mult_x_18_n526), .CO(
        mult_x_18_n522), .COX(mult_x_18_n521), .S(mult_x_18_n523) );
  CMPE42D1BWP12T U3280 ( .A(mult_x_18_n534), .B(mult_x_18_n515), .C(
        mult_x_18_n525), .CIX(mult_x_18_n521), .D(mult_x_18_n509), .CO(
        mult_x_18_n505), .COX(mult_x_18_n504), .S(mult_x_18_n506) );
endmodule


module top7 ( clock, reset, stall_from_instructionfetch, decoder_pc_update, 
        MEM_MEMCTRL_from_mem_data, MEMCTRL_MEM_to_mem_read_enable, 
        MEMCTRL_MEM_to_mem_write_enable, MEMCTRL_MEM_to_mem_mem_enable, 
        MEMCTRL_MEM_to_mem_address, MEMCTRL_MEM_to_mem_data );
  input [15:0] MEM_MEMCTRL_from_mem_data;
  output [11:0] MEMCTRL_MEM_to_mem_address;
  output [15:0] MEMCTRL_MEM_to_mem_data;
  input clock, reset, stall_from_instructionfetch;
  output decoder_pc_update, MEMCTRL_MEM_to_mem_read_enable,
         MEMCTRL_MEM_to_mem_write_enable, MEMCTRL_MEM_to_mem_mem_enable;
  wire   ALU_OUT_n, ALU_OUT_c, ALU_OUT_z, ALU_OUT_v, ALU_IN_c, MEMCTRL_load_in,
         n3, n4, memory_interface_inst1_fsm_state_3_,
         memory_interface_inst1_fsm_state_2_,
         memory_interface_inst1_fsm_state_1_,
         memory_interface_inst1_fsm_state_0_, memory_interface_inst1_fsm_N32,
         memory_interface_inst1_fsm_N33, memory_interface_inst1_fsm_N34,
         memory_interface_inst1_fsm_N35,
         memory_interface_inst1_delayed_is_signed,
         memory_interface_inst1_delay_addr_for_adder_0_,
         memory_interface_inst1_delay_addr_for_adder_1_,
         memory_interface_inst1_delay_addr_for_adder_2_,
         memory_interface_inst1_delay_addr_for_adder_3_,
         memory_interface_inst1_delay_addr_for_adder_4_,
         memory_interface_inst1_delay_addr_for_adder_5_,
         memory_interface_inst1_delay_addr_for_adder_6_,
         memory_interface_inst1_delay_addr_for_adder_7_,
         memory_interface_inst1_delay_addr_for_adder_8_,
         memory_interface_inst1_delay_addr_for_adder_9_,
         memory_interface_inst1_delay_addr_for_adder_10_,
         memory_interface_inst1_delay_addr_for_adder_11_,
         register_file_inst1_n2648, register_file_inst1_n2647,
         register_file_inst1_n2646, register_file_inst1_n2645,
         register_file_inst1_n2644, register_file_inst1_n2643,
         register_file_inst1_n2642, register_file_inst1_n2641,
         register_file_inst1_n2640, register_file_inst1_n2639,
         register_file_inst1_n2638, register_file_inst1_n2637,
         register_file_inst1_n2636, register_file_inst1_n2635,
         register_file_inst1_n2634, register_file_inst1_n2633,
         register_file_inst1_n2632, register_file_inst1_n2631,
         register_file_inst1_n2630, register_file_inst1_n2629,
         register_file_inst1_n2628, register_file_inst1_n2627,
         register_file_inst1_n2626, register_file_inst1_n2625,
         register_file_inst1_n2624, register_file_inst1_n2623,
         register_file_inst1_n2622, register_file_inst1_n2621,
         register_file_inst1_n2620, register_file_inst1_n2619,
         register_file_inst1_n2618, register_file_inst1_n2617,
         register_file_inst1_n2616, register_file_inst1_n2615,
         register_file_inst1_n2614, register_file_inst1_n2613,
         register_file_inst1_n2612, register_file_inst1_n2611,
         register_file_inst1_n2610, register_file_inst1_n2609,
         register_file_inst1_n2608, register_file_inst1_n2607,
         register_file_inst1_n2606, register_file_inst1_n2605,
         register_file_inst1_n2604, register_file_inst1_n2603,
         register_file_inst1_n2602, register_file_inst1_n2601,
         register_file_inst1_n2600, register_file_inst1_n2599,
         register_file_inst1_n2598, register_file_inst1_n2597,
         register_file_inst1_n2596, register_file_inst1_n2595,
         register_file_inst1_n2594, register_file_inst1_n2593,
         register_file_inst1_n2592, register_file_inst1_n2591,
         register_file_inst1_n2590, register_file_inst1_n2589,
         register_file_inst1_n2588, register_file_inst1_n2587,
         register_file_inst1_n2586, register_file_inst1_n2585,
         register_file_inst1_n2584, register_file_inst1_n2583,
         register_file_inst1_n2582, register_file_inst1_n2581,
         register_file_inst1_n2580, register_file_inst1_n2579,
         register_file_inst1_n2578, register_file_inst1_n2577,
         register_file_inst1_n2576, register_file_inst1_n2575,
         register_file_inst1_n2574, register_file_inst1_n2573,
         register_file_inst1_n2572, register_file_inst1_n2571,
         register_file_inst1_n2570, register_file_inst1_n2569,
         register_file_inst1_n2568, register_file_inst1_n2567,
         register_file_inst1_n2566, register_file_inst1_n2565,
         register_file_inst1_n2564, register_file_inst1_n2563,
         register_file_inst1_n2562, register_file_inst1_n2561,
         register_file_inst1_n2560, register_file_inst1_n2559,
         register_file_inst1_n2558, register_file_inst1_n2557,
         register_file_inst1_n2556, register_file_inst1_n2555,
         register_file_inst1_n2554, register_file_inst1_n2553,
         register_file_inst1_n2552, register_file_inst1_n2551,
         register_file_inst1_n2550, register_file_inst1_n2549,
         register_file_inst1_n2548, register_file_inst1_n2547,
         register_file_inst1_n2546, register_file_inst1_n2545,
         register_file_inst1_n2544, register_file_inst1_n2543,
         register_file_inst1_n2542, register_file_inst1_n2541,
         register_file_inst1_n2540, register_file_inst1_n2539,
         register_file_inst1_n2538, register_file_inst1_n2537,
         register_file_inst1_n2536, register_file_inst1_n2535,
         register_file_inst1_n2534, register_file_inst1_n2533,
         register_file_inst1_n2532, register_file_inst1_n2531,
         register_file_inst1_n2530, register_file_inst1_n2529,
         register_file_inst1_n2528, register_file_inst1_n2527,
         register_file_inst1_n2526, register_file_inst1_n2525,
         register_file_inst1_n2524, register_file_inst1_n2523,
         register_file_inst1_n2522, register_file_inst1_n2521,
         register_file_inst1_n2520, register_file_inst1_n2519,
         register_file_inst1_n2518, register_file_inst1_n2517,
         register_file_inst1_n2516, register_file_inst1_n2515,
         register_file_inst1_n2514, register_file_inst1_n2513,
         register_file_inst1_n2512, register_file_inst1_n2511,
         register_file_inst1_n2510, register_file_inst1_n2509,
         register_file_inst1_n2508, register_file_inst1_n2507,
         register_file_inst1_n2506, register_file_inst1_n2505,
         register_file_inst1_n2504, register_file_inst1_n2503,
         register_file_inst1_n2502, register_file_inst1_n2501,
         register_file_inst1_n2500, register_file_inst1_n2499,
         register_file_inst1_n2498, register_file_inst1_n2497,
         register_file_inst1_n2496, register_file_inst1_n2495,
         register_file_inst1_n2494, register_file_inst1_n2493,
         register_file_inst1_n2492, register_file_inst1_n2491,
         register_file_inst1_n2490, register_file_inst1_n2489,
         register_file_inst1_n2488, register_file_inst1_n2487,
         register_file_inst1_n2486, register_file_inst1_n2485,
         register_file_inst1_n2484, register_file_inst1_n2483,
         register_file_inst1_n2482, register_file_inst1_n2481,
         register_file_inst1_n2480, register_file_inst1_n2479,
         register_file_inst1_n2478, register_file_inst1_n2477,
         register_file_inst1_n2476, register_file_inst1_n2475,
         register_file_inst1_n2474, register_file_inst1_n2473,
         register_file_inst1_n2472, register_file_inst1_n2471,
         register_file_inst1_n2470, register_file_inst1_n2469,
         register_file_inst1_n2468, register_file_inst1_n2467,
         register_file_inst1_n2466, register_file_inst1_n2465,
         register_file_inst1_n2464, register_file_inst1_n2463,
         register_file_inst1_n2462, register_file_inst1_n2461,
         register_file_inst1_n2460, register_file_inst1_n2459,
         register_file_inst1_n2458, register_file_inst1_n2457,
         register_file_inst1_n2456, register_file_inst1_n2455,
         register_file_inst1_n2454, register_file_inst1_n2453,
         register_file_inst1_n2452, register_file_inst1_n2451,
         register_file_inst1_n2450, register_file_inst1_n2449,
         register_file_inst1_n2448, register_file_inst1_n2447,
         register_file_inst1_n2446, register_file_inst1_n2445,
         register_file_inst1_n2444, register_file_inst1_n2443,
         register_file_inst1_n2442, register_file_inst1_n2441,
         register_file_inst1_n2440, register_file_inst1_n2439,
         register_file_inst1_n2438, register_file_inst1_n2437,
         register_file_inst1_n2436, register_file_inst1_n2435,
         register_file_inst1_n2434, register_file_inst1_n2433,
         register_file_inst1_n2432, register_file_inst1_n2431,
         register_file_inst1_n2430, register_file_inst1_n2429,
         register_file_inst1_n2428, register_file_inst1_n2427,
         register_file_inst1_n2426, register_file_inst1_n2425,
         register_file_inst1_n2424, register_file_inst1_n2423,
         register_file_inst1_n2422, register_file_inst1_n2421,
         register_file_inst1_n2420, register_file_inst1_n2419,
         register_file_inst1_n2418, register_file_inst1_n2417,
         register_file_inst1_n2416, register_file_inst1_n2415,
         register_file_inst1_n2414, register_file_inst1_n2413,
         register_file_inst1_n2412, register_file_inst1_n2411,
         register_file_inst1_n2410, register_file_inst1_n2409,
         register_file_inst1_n2408, register_file_inst1_n2407,
         register_file_inst1_n2406, register_file_inst1_n2405,
         register_file_inst1_n2404, register_file_inst1_n2403,
         register_file_inst1_n2402, register_file_inst1_n2401,
         register_file_inst1_n2400, register_file_inst1_n2399,
         register_file_inst1_n2398, register_file_inst1_n2397,
         register_file_inst1_n2396, register_file_inst1_n2395,
         register_file_inst1_n2394, register_file_inst1_n2393,
         register_file_inst1_n2392, register_file_inst1_n2391,
         register_file_inst1_n2390, register_file_inst1_n2389,
         register_file_inst1_n2388, register_file_inst1_n2387,
         register_file_inst1_n2386, register_file_inst1_n2385,
         register_file_inst1_n2384, register_file_inst1_n2383,
         register_file_inst1_n2382, register_file_inst1_n2381,
         register_file_inst1_n2380, register_file_inst1_n2379,
         register_file_inst1_n2378, register_file_inst1_n2377,
         register_file_inst1_n2376, register_file_inst1_n2375,
         register_file_inst1_n2374, register_file_inst1_n2373,
         register_file_inst1_n2372, register_file_inst1_n2371,
         register_file_inst1_n2370, register_file_inst1_n2369,
         register_file_inst1_n2368, register_file_inst1_n2367,
         register_file_inst1_n2366, register_file_inst1_n2365,
         register_file_inst1_n2364, register_file_inst1_n2363,
         register_file_inst1_n2362, register_file_inst1_n2361,
         register_file_inst1_n2360, register_file_inst1_n2359,
         register_file_inst1_n2358, register_file_inst1_n2357,
         register_file_inst1_n2356, register_file_inst1_n2355,
         register_file_inst1_n2354, register_file_inst1_n2353,
         register_file_inst1_n2352, register_file_inst1_n2351,
         register_file_inst1_n2350, register_file_inst1_n2349,
         register_file_inst1_n2348, register_file_inst1_n2347,
         register_file_inst1_n2346, register_file_inst1_n2345,
         register_file_inst1_n2344, register_file_inst1_n2343,
         register_file_inst1_n2342, register_file_inst1_n2341,
         register_file_inst1_n2340, register_file_inst1_n2339,
         register_file_inst1_n2338, register_file_inst1_n2337,
         register_file_inst1_n2336, register_file_inst1_n2335,
         register_file_inst1_n2334, register_file_inst1_n2333,
         register_file_inst1_n2332, register_file_inst1_n2331,
         register_file_inst1_n2330, register_file_inst1_n2329,
         register_file_inst1_n2328, register_file_inst1_n2327,
         register_file_inst1_n2326, register_file_inst1_n2325,
         register_file_inst1_n2324, register_file_inst1_n2323,
         register_file_inst1_n2322, register_file_inst1_n2321,
         register_file_inst1_n2320, register_file_inst1_n2319,
         register_file_inst1_n2318, register_file_inst1_n2317,
         register_file_inst1_n2316, register_file_inst1_n2315,
         register_file_inst1_n2314, register_file_inst1_n2313,
         register_file_inst1_n2312, register_file_inst1_n2311,
         register_file_inst1_n2310, register_file_inst1_n2309,
         register_file_inst1_n2308, register_file_inst1_n2307,
         register_file_inst1_n2306, register_file_inst1_n2305,
         register_file_inst1_n2304, register_file_inst1_n2303,
         register_file_inst1_n2302, register_file_inst1_n2301,
         register_file_inst1_n2300, register_file_inst1_n2299,
         register_file_inst1_n2298, register_file_inst1_n2297,
         register_file_inst1_n2296, register_file_inst1_n2295,
         register_file_inst1_n2294, register_file_inst1_n2293,
         register_file_inst1_n2292, register_file_inst1_n2291,
         register_file_inst1_n2290, register_file_inst1_n2289,
         register_file_inst1_n2288, register_file_inst1_n2287,
         register_file_inst1_n2286, register_file_inst1_n2285,
         register_file_inst1_n2284, register_file_inst1_n2283,
         register_file_inst1_n2282, register_file_inst1_n2281,
         register_file_inst1_n2280, register_file_inst1_n2279,
         register_file_inst1_n2278, register_file_inst1_n2277,
         register_file_inst1_n2276, register_file_inst1_n2275,
         register_file_inst1_n2274, register_file_inst1_n2273,
         register_file_inst1_n2272, register_file_inst1_n2271,
         register_file_inst1_n2270, register_file_inst1_n2269,
         register_file_inst1_n2268, register_file_inst1_n2267,
         register_file_inst1_n2266, register_file_inst1_n2265,
         register_file_inst1_n2264, register_file_inst1_n2263,
         register_file_inst1_n2262, register_file_inst1_n2261,
         register_file_inst1_n2260, register_file_inst1_n2259,
         register_file_inst1_n2258, register_file_inst1_n2257,
         register_file_inst1_n2256, register_file_inst1_n2255,
         register_file_inst1_n2254, register_file_inst1_n2253,
         register_file_inst1_n2252, register_file_inst1_n2251,
         register_file_inst1_n2250, register_file_inst1_n2249,
         register_file_inst1_n2248, register_file_inst1_n2247,
         register_file_inst1_n2246, register_file_inst1_n2245,
         register_file_inst1_n2244, register_file_inst1_n2243,
         register_file_inst1_n2242, register_file_inst1_n2241,
         register_file_inst1_n2240, register_file_inst1_n2239,
         register_file_inst1_n2238, register_file_inst1_n2237,
         register_file_inst1_n2236, register_file_inst1_n2235,
         register_file_inst1_n2234, register_file_inst1_n2233,
         register_file_inst1_n2232, register_file_inst1_n2231,
         register_file_inst1_n2230, register_file_inst1_n2229,
         register_file_inst1_n2228, register_file_inst1_n2227,
         register_file_inst1_n2226, register_file_inst1_n2225,
         register_file_inst1_n2224, register_file_inst1_n2223,
         register_file_inst1_n2222, register_file_inst1_n2221,
         register_file_inst1_n2220, register_file_inst1_n2219,
         register_file_inst1_n2218, register_file_inst1_n2217,
         register_file_inst1_n2216, register_file_inst1_n2215,
         register_file_inst1_n2214, register_file_inst1_n2213,
         register_file_inst1_n2212, register_file_inst1_n2211,
         register_file_inst1_n2210, register_file_inst1_n2209,
         register_file_inst1_n2208, register_file_inst1_n2207,
         register_file_inst1_n2206, register_file_inst1_n2205,
         register_file_inst1_n2204, register_file_inst1_n2203,
         register_file_inst1_n2202, register_file_inst1_n2201,
         register_file_inst1_n2200, register_file_inst1_n2199,
         register_file_inst1_n2198, register_file_inst1_n2197,
         register_file_inst1_n2196, register_file_inst1_n2195,
         register_file_inst1_n2194, register_file_inst1_n2193,
         register_file_inst1_n2192, register_file_inst1_n2191,
         register_file_inst1_n2190, register_file_inst1_n2189,
         register_file_inst1_n2188, register_file_inst1_n2187,
         register_file_inst1_n2186, register_file_inst1_n2185,
         register_file_inst1_n2184, register_file_inst1_n2183,
         register_file_inst1_n2182, register_file_inst1_n2181,
         register_file_inst1_n2180, register_file_inst1_n2179,
         register_file_inst1_n2178, register_file_inst1_n2177,
         register_file_inst1_n2176, register_file_inst1_n2175,
         register_file_inst1_n2174, register_file_inst1_n2173,
         register_file_inst1_n2172, register_file_inst1_n2171,
         register_file_inst1_n2170, register_file_inst1_n2169,
         register_file_inst1_n2168, register_file_inst1_n2167,
         register_file_inst1_n2166, register_file_inst1_n2165,
         register_file_inst1_n2164, register_file_inst1_n2163,
         register_file_inst1_n2162, register_file_inst1_n2161,
         register_file_inst1_n2160, register_file_inst1_n2159,
         register_file_inst1_n2158, register_file_inst1_n2157,
         register_file_inst1_n2156, register_file_inst1_n2155,
         register_file_inst1_n2154, register_file_inst1_n2153,
         register_file_inst1_n2152, register_file_inst1_n2151,
         register_file_inst1_n2150, register_file_inst1_n2149,
         register_file_inst1_n2148, register_file_inst1_n2147,
         register_file_inst1_n2146, register_file_inst1_n2145,
         register_file_inst1_n2144, register_file_inst1_n2143,
         register_file_inst1_n2142, register_file_inst1_n2141,
         register_file_inst1_n2140, register_file_inst1_n2139,
         register_file_inst1_n2138, register_file_inst1_n2136,
         register_file_inst1_pc_write_in_0_,
         register_file_inst1_pc_write_in_1_,
         register_file_inst1_pc_write_in_3_,
         register_file_inst1_pc_write_in_5_,
         register_file_inst1_pc_write_in_7_,
         register_file_inst1_pc_write_in_11_,
         register_file_inst1_pc_write_in_12_,
         register_file_inst1_pc_write_in_13_,
         register_file_inst1_pc_write_in_14_,
         register_file_inst1_pc_write_in_15_, register_file_inst1_tmp1_0_,
         register_file_inst1_tmp1_1_, register_file_inst1_tmp1_2_,
         register_file_inst1_tmp1_3_, register_file_inst1_tmp1_4_,
         register_file_inst1_tmp1_5_, register_file_inst1_tmp1_6_,
         register_file_inst1_tmp1_7_, register_file_inst1_tmp1_8_,
         register_file_inst1_tmp1_9_, register_file_inst1_tmp1_10_,
         register_file_inst1_tmp1_11_, register_file_inst1_tmp1_12_,
         register_file_inst1_tmp1_13_, register_file_inst1_tmp1_14_,
         register_file_inst1_tmp1_15_, register_file_inst1_tmp1_16_,
         register_file_inst1_tmp1_17_, register_file_inst1_tmp1_18_,
         register_file_inst1_tmp1_19_, register_file_inst1_tmp1_20_,
         register_file_inst1_tmp1_21_, register_file_inst1_tmp1_22_,
         register_file_inst1_tmp1_23_, register_file_inst1_tmp1_24_,
         register_file_inst1_tmp1_25_, register_file_inst1_tmp1_26_,
         register_file_inst1_tmp1_27_, register_file_inst1_tmp1_28_,
         register_file_inst1_tmp1_29_, register_file_inst1_tmp1_30_,
         register_file_inst1_tmp1_31_, register_file_inst1_lr_0_,
         register_file_inst1_lr_1_, register_file_inst1_lr_2_,
         register_file_inst1_lr_3_, register_file_inst1_lr_4_,
         register_file_inst1_lr_5_, register_file_inst1_lr_6_,
         register_file_inst1_lr_7_, register_file_inst1_lr_8_,
         register_file_inst1_lr_9_, register_file_inst1_lr_10_,
         register_file_inst1_lr_11_, register_file_inst1_lr_12_,
         register_file_inst1_lr_13_, register_file_inst1_lr_14_,
         register_file_inst1_lr_15_, register_file_inst1_lr_16_,
         register_file_inst1_lr_17_, register_file_inst1_lr_18_,
         register_file_inst1_lr_19_, register_file_inst1_lr_20_,
         register_file_inst1_lr_21_, register_file_inst1_lr_22_,
         register_file_inst1_lr_23_, register_file_inst1_lr_24_,
         register_file_inst1_lr_25_, register_file_inst1_lr_26_,
         register_file_inst1_lr_27_, register_file_inst1_lr_28_,
         register_file_inst1_lr_29_, register_file_inst1_lr_30_,
         register_file_inst1_lr_31_, register_file_inst1_r12_0_,
         register_file_inst1_r12_1_, register_file_inst1_r12_2_,
         register_file_inst1_r12_3_, register_file_inst1_r12_4_,
         register_file_inst1_r12_5_, register_file_inst1_r12_6_,
         register_file_inst1_r12_7_, register_file_inst1_r12_8_,
         register_file_inst1_r12_9_, register_file_inst1_r12_10_,
         register_file_inst1_r12_11_, register_file_inst1_r12_12_,
         register_file_inst1_r12_13_, register_file_inst1_r12_14_,
         register_file_inst1_r12_15_, register_file_inst1_r12_16_,
         register_file_inst1_r12_17_, register_file_inst1_r12_18_,
         register_file_inst1_r12_19_, register_file_inst1_r12_20_,
         register_file_inst1_r12_21_, register_file_inst1_r12_22_,
         register_file_inst1_r12_23_, register_file_inst1_r12_24_,
         register_file_inst1_r12_25_, register_file_inst1_r12_26_,
         register_file_inst1_r12_27_, register_file_inst1_r12_28_,
         register_file_inst1_r12_29_, register_file_inst1_r12_30_,
         register_file_inst1_r12_31_, register_file_inst1_r11_0_,
         register_file_inst1_r11_1_, register_file_inst1_r11_2_,
         register_file_inst1_r11_3_, register_file_inst1_r11_4_,
         register_file_inst1_r11_5_, register_file_inst1_r11_6_,
         register_file_inst1_r11_7_, register_file_inst1_r11_8_,
         register_file_inst1_r11_9_, register_file_inst1_r11_10_,
         register_file_inst1_r11_11_, register_file_inst1_r11_12_,
         register_file_inst1_r11_13_, register_file_inst1_r11_14_,
         register_file_inst1_r11_15_, register_file_inst1_r11_16_,
         register_file_inst1_r11_17_, register_file_inst1_r11_18_,
         register_file_inst1_r11_19_, register_file_inst1_r11_20_,
         register_file_inst1_r11_21_, register_file_inst1_r11_22_,
         register_file_inst1_r11_23_, register_file_inst1_r11_24_,
         register_file_inst1_r11_25_, register_file_inst1_r11_26_,
         register_file_inst1_r11_27_, register_file_inst1_r11_28_,
         register_file_inst1_r11_29_, register_file_inst1_r11_30_,
         register_file_inst1_r11_31_, register_file_inst1_r10_0_,
         register_file_inst1_r10_1_, register_file_inst1_r10_2_,
         register_file_inst1_r10_3_, register_file_inst1_r10_4_,
         register_file_inst1_r10_5_, register_file_inst1_r10_6_,
         register_file_inst1_r10_7_, register_file_inst1_r10_8_,
         register_file_inst1_r10_9_, register_file_inst1_r10_10_,
         register_file_inst1_r10_11_, register_file_inst1_r10_12_,
         register_file_inst1_r10_13_, register_file_inst1_r10_14_,
         register_file_inst1_r10_15_, register_file_inst1_r10_16_,
         register_file_inst1_r10_17_, register_file_inst1_r10_18_,
         register_file_inst1_r10_19_, register_file_inst1_r10_20_,
         register_file_inst1_r10_21_, register_file_inst1_r10_22_,
         register_file_inst1_r10_23_, register_file_inst1_r10_24_,
         register_file_inst1_r10_25_, register_file_inst1_r10_26_,
         register_file_inst1_r10_27_, register_file_inst1_r10_28_,
         register_file_inst1_r10_29_, register_file_inst1_r10_30_,
         register_file_inst1_r10_31_, register_file_inst1_r9_0_,
         register_file_inst1_r9_1_, register_file_inst1_r9_2_,
         register_file_inst1_r9_3_, register_file_inst1_r9_4_,
         register_file_inst1_r9_5_, register_file_inst1_r9_6_,
         register_file_inst1_r9_7_, register_file_inst1_r9_8_,
         register_file_inst1_r9_9_, register_file_inst1_r9_10_,
         register_file_inst1_r9_11_, register_file_inst1_r9_12_,
         register_file_inst1_r9_13_, register_file_inst1_r9_14_,
         register_file_inst1_r9_15_, register_file_inst1_r9_16_,
         register_file_inst1_r9_17_, register_file_inst1_r9_18_,
         register_file_inst1_r9_19_, register_file_inst1_r9_20_,
         register_file_inst1_r9_21_, register_file_inst1_r9_22_,
         register_file_inst1_r9_23_, register_file_inst1_r9_24_,
         register_file_inst1_r9_25_, register_file_inst1_r9_26_,
         register_file_inst1_r9_27_, register_file_inst1_r9_28_,
         register_file_inst1_r9_29_, register_file_inst1_r9_30_,
         register_file_inst1_r9_31_, register_file_inst1_r8_0_,
         register_file_inst1_r8_1_, register_file_inst1_r8_2_,
         register_file_inst1_r8_3_, register_file_inst1_r8_4_,
         register_file_inst1_r8_5_, register_file_inst1_r8_6_,
         register_file_inst1_r8_7_, register_file_inst1_r8_8_,
         register_file_inst1_r8_9_, register_file_inst1_r8_10_,
         register_file_inst1_r8_11_, register_file_inst1_r8_12_,
         register_file_inst1_r8_13_, register_file_inst1_r8_14_,
         register_file_inst1_r8_15_, register_file_inst1_r8_16_,
         register_file_inst1_r8_17_, register_file_inst1_r8_18_,
         register_file_inst1_r8_19_, register_file_inst1_r8_20_,
         register_file_inst1_r8_21_, register_file_inst1_r8_22_,
         register_file_inst1_r8_23_, register_file_inst1_r8_24_,
         register_file_inst1_r8_25_, register_file_inst1_r8_26_,
         register_file_inst1_r8_27_, register_file_inst1_r8_28_,
         register_file_inst1_r8_29_, register_file_inst1_r8_30_,
         register_file_inst1_r8_31_, register_file_inst1_r7_0_,
         register_file_inst1_r7_1_, register_file_inst1_r7_2_,
         register_file_inst1_r7_3_, register_file_inst1_r7_4_,
         register_file_inst1_r7_5_, register_file_inst1_r7_6_,
         register_file_inst1_r7_7_, register_file_inst1_r7_8_,
         register_file_inst1_r7_9_, register_file_inst1_r7_10_,
         register_file_inst1_r7_11_, register_file_inst1_r7_12_,
         register_file_inst1_r7_13_, register_file_inst1_r7_14_,
         register_file_inst1_r7_15_, register_file_inst1_r7_16_,
         register_file_inst1_r7_17_, register_file_inst1_r7_18_,
         register_file_inst1_r7_19_, register_file_inst1_r7_20_,
         register_file_inst1_r7_21_, register_file_inst1_r7_22_,
         register_file_inst1_r7_23_, register_file_inst1_r7_24_,
         register_file_inst1_r7_25_, register_file_inst1_r7_26_,
         register_file_inst1_r7_27_, register_file_inst1_r7_28_,
         register_file_inst1_r7_29_, register_file_inst1_r7_30_,
         register_file_inst1_r7_31_, register_file_inst1_r6_0_,
         register_file_inst1_r6_1_, register_file_inst1_r6_2_,
         register_file_inst1_r6_3_, register_file_inst1_r6_4_,
         register_file_inst1_r6_5_, register_file_inst1_r6_6_,
         register_file_inst1_r6_7_, register_file_inst1_r6_8_,
         register_file_inst1_r6_9_, register_file_inst1_r6_10_,
         register_file_inst1_r6_11_, register_file_inst1_r6_12_,
         register_file_inst1_r6_13_, register_file_inst1_r6_14_,
         register_file_inst1_r6_15_, register_file_inst1_r6_16_,
         register_file_inst1_r6_17_, register_file_inst1_r6_18_,
         register_file_inst1_r6_19_, register_file_inst1_r6_20_,
         register_file_inst1_r6_21_, register_file_inst1_r6_22_,
         register_file_inst1_r6_23_, register_file_inst1_r6_24_,
         register_file_inst1_r6_25_, register_file_inst1_r6_26_,
         register_file_inst1_r6_27_, register_file_inst1_r6_28_,
         register_file_inst1_r6_29_, register_file_inst1_r6_30_,
         register_file_inst1_r6_31_, register_file_inst1_r5_0_,
         register_file_inst1_r5_1_, register_file_inst1_r5_2_,
         register_file_inst1_r5_3_, register_file_inst1_r5_4_,
         register_file_inst1_r5_5_, register_file_inst1_r5_6_,
         register_file_inst1_r5_7_, register_file_inst1_r5_8_,
         register_file_inst1_r5_9_, register_file_inst1_r5_10_,
         register_file_inst1_r5_11_, register_file_inst1_r5_12_,
         register_file_inst1_r5_13_, register_file_inst1_r5_14_,
         register_file_inst1_r5_15_, register_file_inst1_r5_16_,
         register_file_inst1_r5_17_, register_file_inst1_r5_18_,
         register_file_inst1_r5_19_, register_file_inst1_r5_20_,
         register_file_inst1_r5_21_, register_file_inst1_r5_22_,
         register_file_inst1_r5_23_, register_file_inst1_r5_24_,
         register_file_inst1_r5_25_, register_file_inst1_r5_26_,
         register_file_inst1_r5_27_, register_file_inst1_r5_28_,
         register_file_inst1_r5_29_, register_file_inst1_r5_30_,
         register_file_inst1_r5_31_, register_file_inst1_r4_0_,
         register_file_inst1_r4_1_, register_file_inst1_r4_2_,
         register_file_inst1_r4_3_, register_file_inst1_r4_4_,
         register_file_inst1_r4_5_, register_file_inst1_r4_6_,
         register_file_inst1_r4_7_, register_file_inst1_r4_8_,
         register_file_inst1_r4_9_, register_file_inst1_r4_10_,
         register_file_inst1_r4_11_, register_file_inst1_r4_12_,
         register_file_inst1_r4_13_, register_file_inst1_r4_14_,
         register_file_inst1_r4_15_, register_file_inst1_r4_16_,
         register_file_inst1_r4_17_, register_file_inst1_r4_18_,
         register_file_inst1_r4_19_, register_file_inst1_r4_20_,
         register_file_inst1_r4_21_, register_file_inst1_r4_22_,
         register_file_inst1_r4_23_, register_file_inst1_r4_24_,
         register_file_inst1_r4_25_, register_file_inst1_r4_26_,
         register_file_inst1_r4_27_, register_file_inst1_r4_28_,
         register_file_inst1_r4_29_, register_file_inst1_r4_30_,
         register_file_inst1_r4_31_, register_file_inst1_r3_0_,
         register_file_inst1_r3_1_, register_file_inst1_r3_2_,
         register_file_inst1_r3_3_, register_file_inst1_r3_4_,
         register_file_inst1_r3_5_, register_file_inst1_r3_6_,
         register_file_inst1_r3_7_, register_file_inst1_r3_8_,
         register_file_inst1_r3_9_, register_file_inst1_r3_10_,
         register_file_inst1_r3_11_, register_file_inst1_r3_12_,
         register_file_inst1_r3_13_, register_file_inst1_r3_14_,
         register_file_inst1_r3_15_, register_file_inst1_r3_16_,
         register_file_inst1_r3_17_, register_file_inst1_r3_18_,
         register_file_inst1_r3_19_, register_file_inst1_r3_20_,
         register_file_inst1_r3_21_, register_file_inst1_r3_22_,
         register_file_inst1_r3_23_, register_file_inst1_r3_24_,
         register_file_inst1_r3_25_, register_file_inst1_r3_26_,
         register_file_inst1_r3_27_, register_file_inst1_r3_28_,
         register_file_inst1_r3_29_, register_file_inst1_r3_30_,
         register_file_inst1_r3_31_, register_file_inst1_r2_0_,
         register_file_inst1_r2_1_, register_file_inst1_r2_2_,
         register_file_inst1_r2_3_, register_file_inst1_r2_4_,
         register_file_inst1_r2_5_, register_file_inst1_r2_6_,
         register_file_inst1_r2_7_, register_file_inst1_r2_8_,
         register_file_inst1_r2_9_, register_file_inst1_r2_10_,
         register_file_inst1_r2_11_, register_file_inst1_r2_12_,
         register_file_inst1_r2_13_, register_file_inst1_r2_14_,
         register_file_inst1_r2_15_, register_file_inst1_r2_16_,
         register_file_inst1_r2_17_, register_file_inst1_r2_18_,
         register_file_inst1_r2_19_, register_file_inst1_r2_20_,
         register_file_inst1_r2_21_, register_file_inst1_r2_22_,
         register_file_inst1_r2_23_, register_file_inst1_r2_24_,
         register_file_inst1_r2_25_, register_file_inst1_r2_26_,
         register_file_inst1_r2_27_, register_file_inst1_r2_28_,
         register_file_inst1_r2_29_, register_file_inst1_r2_30_,
         register_file_inst1_r2_31_, register_file_inst1_r1_0_,
         register_file_inst1_r1_1_, register_file_inst1_r1_2_,
         register_file_inst1_r1_3_, register_file_inst1_r1_4_,
         register_file_inst1_r1_5_, register_file_inst1_r1_6_,
         register_file_inst1_r1_7_, register_file_inst1_r1_8_,
         register_file_inst1_r1_9_, register_file_inst1_r1_10_,
         register_file_inst1_r1_11_, register_file_inst1_r1_12_,
         register_file_inst1_r1_13_, register_file_inst1_r1_14_,
         register_file_inst1_r1_15_, register_file_inst1_r1_16_,
         register_file_inst1_r1_17_, register_file_inst1_r1_18_,
         register_file_inst1_r1_19_, register_file_inst1_r1_20_,
         register_file_inst1_r1_21_, register_file_inst1_r1_22_,
         register_file_inst1_r1_23_, register_file_inst1_r1_24_,
         register_file_inst1_r1_25_, register_file_inst1_r1_26_,
         register_file_inst1_r1_27_, register_file_inst1_r1_28_,
         register_file_inst1_r1_29_, register_file_inst1_r1_30_,
         register_file_inst1_r1_31_, register_file_inst1_r0_0_,
         register_file_inst1_r0_1_, register_file_inst1_r0_2_,
         register_file_inst1_r0_3_, register_file_inst1_r0_4_,
         register_file_inst1_r0_5_, register_file_inst1_r0_6_,
         register_file_inst1_r0_7_, register_file_inst1_r0_8_,
         register_file_inst1_r0_9_, register_file_inst1_r0_10_,
         register_file_inst1_r0_11_, register_file_inst1_r0_12_,
         register_file_inst1_r0_13_, register_file_inst1_r0_14_,
         register_file_inst1_r0_15_, register_file_inst1_r0_16_,
         register_file_inst1_r0_17_, register_file_inst1_r0_18_,
         register_file_inst1_r0_19_, register_file_inst1_r0_20_,
         register_file_inst1_r0_21_, register_file_inst1_r0_22_,
         register_file_inst1_r0_23_, register_file_inst1_r0_24_,
         register_file_inst1_r0_25_, register_file_inst1_r0_26_,
         register_file_inst1_r0_27_, register_file_inst1_r0_28_,
         register_file_inst1_r0_29_, register_file_inst1_r0_30_,
         register_file_inst1_r0_31_, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333;
  wire   [31:0] ALU_MISC_OUT_result;
  wire   [31:0] STACK_RF_next_sp;
  wire   [31:0] RF_ALU_STACK_operand_a;
  wire   [31:0] RF_ALU_operand_b;
  wire   [31:0] RF_MEMCTRL_data_reg;
  wire   [12:2] RF_MEMCTRL_address_reg;
  wire   [11:0] MEMCTRL_IN_address;
  wire   [15:0] memory_interface_inst1_delay_first_two_bytes_out;
  wire   [31:0] memory_interface_inst1_delay_data_in32;
  wire   [11:0] memory_interface_inst1_delay_addr_single;
  wire   [3:0] register_file_inst1_cpsrin;
  wire   [30:2] register_file_inst1_pc_write_in_plus_two;
  wire   [31:0] register_file_inst1_spin;
  tri   clock;
  tri   reset;
  tri   stall_from_instructionfetch;
  tri   decoder_pc_update;
  tri   DEC_CPSR_update_flag_n;
  tri   RF_OUT_n;
  tri   DEC_CPSR_update_flag_c;
  tri   RF_OUT_c;
  tri   DEC_CPSR_update_flag_z;
  tri   RF_OUT_z;
  tri   DEC_CPSR_update_flag_v;
  tri   RF_OUT_v;
  tri   [31:0] IF_DEC_instruction;
  tri   IF_DEC_instruction_valid;
  tri   MEMCTRL_write_finished;
  tri   MEMCTRL_read_finished;
  tri   [4:0] DEC_RF_operand_a;
  tri   [4:0] DEC_RF_operand_b;
  tri   [31:0] DEC_RF_offset_a;
  tri   [31:0] DEC_RF_offset_b;
  tri   [4:0] DEC_ALU_alu_opcode;
  tri   [4:0] DEC_RF_alu_stack_write_to_reg;
  tri   DEC_RF_alu_stack_write_to_reg_enable;
  tri   [4:0] DEC_RF_memory_write_to_reg;
  tri   DEC_RF_memory_write_to_reg_enable;
  tri   [4:0] DEC_RF_memory_store_data_reg;
  tri   [4:0] DEC_RF_memory_store_address_reg;
  tri   DEC_MISC_OUT_memory_address_source_is_reg;
  tri   [1:0] DEC_MEMCTRL_load_store_width;
  tri   DEC_MEMCTRL_memorycontroller_sign_extend;
  tri   DEC_MEMCTRL_CTRL_memory_load_request;
  tri   DEC_MEMCTRL_CTRL_memory_store_request;
  tri   DEC_IF_stall_to_instructionfetch;
  tri   [15:0] MEMCTRL_RF_IF_data_in;
  tri   [31:0] IF_RF_incremented_pc_out;
  tri   IF_RF_incremented_pc_write_enable;
  tri   [31:0] RF_pc_out;
  tri   IF_memory_load_req;
  tri   [11:0] IF_instruction_memory_address;

  irdecode irdecode_inst1 ( .clock(clock), .reset(reset), .instruction(
        IF_DEC_instruction), .flag_n(RF_OUT_n), .flag_z(RF_OUT_z), .flag_c(
        RF_OUT_c), .flag_v(RF_OUT_v), .stall_from_instructionfetch(
        stall_from_instructionfetch), .instruction_valid(
        IF_DEC_instruction_valid), .memory_write_finished(
        MEMCTRL_write_finished), .memory_read_finished(MEMCTRL_read_finished), 
        .operand_a(DEC_RF_operand_a), .operand_b(DEC_RF_operand_b), .offset_a(
        DEC_RF_offset_a), .offset_b(DEC_RF_offset_b), .alu_opcode(
        DEC_ALU_alu_opcode), .update_flag_n(DEC_CPSR_update_flag_n), 
        .update_flag_z(DEC_CPSR_update_flag_z), .update_flag_c(
        DEC_CPSR_update_flag_c), .update_flag_v(DEC_CPSR_update_flag_v), 
        .alu_stack_write_to_reg(DEC_RF_alu_stack_write_to_reg), 
        .alu_stack_write_to_reg_enable(DEC_RF_alu_stack_write_to_reg_enable), 
        .memory_write_to_reg(DEC_RF_memory_write_to_reg), 
        .memory_write_to_reg_enable(DEC_RF_memory_write_to_reg_enable), 
        .memory_store_data_reg(DEC_RF_memory_store_data_reg), 
        .memory_store_address_reg(DEC_RF_memory_store_address_reg), 
        .memory_address_source_is_reg(
        DEC_MISC_OUT_memory_address_source_is_reg), .load_store_width(
        DEC_MEMCTRL_load_store_width), .memorycontroller_sign_extend(
        DEC_MEMCTRL_memorycontroller_sign_extend), .memory_load_request(
        DEC_MEMCTRL_CTRL_memory_load_request), .memory_store_request(
        DEC_MEMCTRL_CTRL_memory_store_request), .stall_to_instructionfetch(
        DEC_IF_stall_to_instructionfetch), .decoder_pc_update(
        decoder_pc_update) );
  ALU_VARIABLE ALU_VARIABLE_inst1 ( .a(RF_ALU_STACK_operand_a), .b(
        RF_ALU_operand_b), .op(DEC_ALU_alu_opcode[3:0]), .c_in(ALU_IN_c), 
        .result(ALU_MISC_OUT_result), .c_out(ALU_OUT_c), .z(ALU_OUT_z), .n(
        ALU_OUT_n), .v(ALU_OUT_v) );
  Instruction_Fetch Instruction_Fetch_inst1 ( .clk(clock), .reset(reset), 
        .stall_decoder_in(DEC_IF_stall_to_instructionfetch), 
        .memory_output_valid(MEMCTRL_read_finished), .current_pc_in(RF_pc_out), 
        .instruction_in(MEMCTRL_RF_IF_data_in), .memory_load_request(
        IF_memory_load_req), .incremented_pc_write_enable(
        IF_RF_incremented_pc_write_enable), .memory_address(
        IF_instruction_memory_address), .incremented_pc_out(
        IF_RF_incremented_pc_out), .instruction_out(IF_DEC_instruction), 
        .instruction_valid(IF_DEC_instruction_valid) );
  DFQD1BWP12T memory_interface_inst1_delayed_is_signed_reg ( .D(
        DEC_MEMCTRL_memorycontroller_sign_extend), .CP(clock), .Q(
        memory_interface_inst1_delayed_is_signed) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_0_ ( .D(
        MEMCTRL_IN_address[0]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[0]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_2_ ( .D(
        MEMCTRL_IN_address[2]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_3_ ( .D(
        MEMCTRL_IN_address[3]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_4_ ( .D(
        MEMCTRL_IN_address[4]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[4]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_5_ ( .D(
        MEMCTRL_IN_address[5]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[5]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_6_ ( .D(
        MEMCTRL_IN_address[6]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_7_ ( .D(
        MEMCTRL_IN_address[7]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_8_ ( .D(
        MEMCTRL_IN_address[8]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_9_ ( .D(
        MEMCTRL_IN_address[9]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_10_ ( .D(
        MEMCTRL_IN_address[10]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_11_ ( .D(
        MEMCTRL_IN_address[11]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[11]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_0_ ( .D(
        MEMCTRL_IN_address[0]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_0_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_2_ ( .D(
        MEMCTRL_IN_address[2]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_2_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_3_ ( .D(
        MEMCTRL_IN_address[3]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_3_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_4_ ( .D(
        MEMCTRL_IN_address[4]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_4_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_5_ ( .D(
        MEMCTRL_IN_address[5]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_5_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_6_ ( .D(
        MEMCTRL_IN_address[6]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_6_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_7_ ( .D(
        MEMCTRL_IN_address[7]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_7_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_8_ ( .D(
        MEMCTRL_IN_address[8]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_8_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_9_ ( .D(
        MEMCTRL_IN_address[9]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_9_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_10_ ( .D(
        MEMCTRL_IN_address[10]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_10_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_11_ ( .D(
        MEMCTRL_IN_address[11]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_11_) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_0_ ( .D(
        MEM_MEMCTRL_from_mem_data[8]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[0]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_1_ ( .D(
        MEM_MEMCTRL_from_mem_data[9]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[1]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_2_ ( .D(
        MEM_MEMCTRL_from_mem_data[10]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_3_ ( .D(
        MEM_MEMCTRL_from_mem_data[11]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_4_ ( .D(
        MEM_MEMCTRL_from_mem_data[12]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[4]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_5_ ( .D(
        MEM_MEMCTRL_from_mem_data[13]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[5]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_6_ ( .D(
        MEM_MEMCTRL_from_mem_data[14]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_7_ ( .D(
        MEM_MEMCTRL_from_mem_data[15]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_8_ ( .D(
        MEM_MEMCTRL_from_mem_data[0]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_9_ ( .D(
        MEM_MEMCTRL_from_mem_data[1]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_10_ ( .D(
        MEM_MEMCTRL_from_mem_data[2]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_11_ ( .D(
        MEM_MEMCTRL_from_mem_data[3]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[11]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_12_ ( .D(
        MEM_MEMCTRL_from_mem_data[4]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[12]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_13_ ( .D(
        MEM_MEMCTRL_from_mem_data[5]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[13]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_14_ ( .D(
        MEM_MEMCTRL_from_mem_data[6]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[14]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_15_ ( .D(
        MEM_MEMCTRL_from_mem_data[7]), .CP(clock), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[15]) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_2_ ( .D(register_file_inst1_n2139), 
        .CP(clock), .Q(register_file_inst1_tmp1_2_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_3_ ( .D(register_file_inst1_n2140), 
        .CP(clock), .Q(register_file_inst1_tmp1_3_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_4_ ( .D(register_file_inst1_n2141), 
        .CP(clock), .Q(register_file_inst1_tmp1_4_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_5_ ( .D(register_file_inst1_n2142), 
        .CP(clock), .Q(register_file_inst1_tmp1_5_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_6_ ( .D(register_file_inst1_n2143), 
        .CP(clock), .Q(register_file_inst1_tmp1_6_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_7_ ( .D(register_file_inst1_n2144), 
        .CP(clock), .Q(register_file_inst1_tmp1_7_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_8_ ( .D(register_file_inst1_n2145), 
        .CP(clock), .Q(register_file_inst1_tmp1_8_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_9_ ( .D(register_file_inst1_n2146), 
        .CP(clock), .Q(register_file_inst1_tmp1_9_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_10_ ( .D(register_file_inst1_n2147), 
        .CP(clock), .Q(register_file_inst1_tmp1_10_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_11_ ( .D(register_file_inst1_n2148), 
        .CP(clock), .Q(register_file_inst1_tmp1_11_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_12_ ( .D(register_file_inst1_n2149), 
        .CP(clock), .Q(register_file_inst1_tmp1_12_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_13_ ( .D(register_file_inst1_n2150), 
        .CP(clock), .Q(register_file_inst1_tmp1_13_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_14_ ( .D(register_file_inst1_n2151), 
        .CP(clock), .Q(register_file_inst1_tmp1_14_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_15_ ( .D(register_file_inst1_n2152), 
        .CP(clock), .Q(register_file_inst1_tmp1_15_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_16_ ( .D(register_file_inst1_n2153), 
        .CP(clock), .Q(register_file_inst1_tmp1_16_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_17_ ( .D(register_file_inst1_n2154), 
        .CP(clock), .Q(register_file_inst1_tmp1_17_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_18_ ( .D(register_file_inst1_n2155), 
        .CP(clock), .Q(register_file_inst1_tmp1_18_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_19_ ( .D(register_file_inst1_n2156), 
        .CP(clock), .Q(register_file_inst1_tmp1_19_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_20_ ( .D(register_file_inst1_n2157), 
        .CP(clock), .Q(register_file_inst1_tmp1_20_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_21_ ( .D(register_file_inst1_n2158), 
        .CP(clock), .Q(register_file_inst1_tmp1_21_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_22_ ( .D(register_file_inst1_n2159), 
        .CP(clock), .Q(register_file_inst1_tmp1_22_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_23_ ( .D(register_file_inst1_n2160), 
        .CP(clock), .Q(register_file_inst1_tmp1_23_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_24_ ( .D(register_file_inst1_n2161), 
        .CP(clock), .Q(register_file_inst1_tmp1_24_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_25_ ( .D(register_file_inst1_n2162), 
        .CP(clock), .Q(register_file_inst1_tmp1_25_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_26_ ( .D(register_file_inst1_n2163), 
        .CP(clock), .Q(register_file_inst1_tmp1_26_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_27_ ( .D(register_file_inst1_n2164), 
        .CP(clock), .Q(register_file_inst1_tmp1_27_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_28_ ( .D(register_file_inst1_n2165), 
        .CP(clock), .Q(register_file_inst1_tmp1_28_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_29_ ( .D(register_file_inst1_n2166), 
        .CP(clock), .Q(register_file_inst1_tmp1_29_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_30_ ( .D(register_file_inst1_n2167), 
        .CP(clock), .Q(register_file_inst1_tmp1_30_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_31_ ( .D(register_file_inst1_n2168), 
        .CP(clock), .Q(register_file_inst1_tmp1_31_) );
  DFQD1BWP12T register_file_inst1_cpsr_reg_0_ ( .D(
        register_file_inst1_cpsrin[0]), .CP(clock), .Q(RF_OUT_v) );
  DFQD1BWP12T register_file_inst1_cpsr_reg_1_ ( .D(
        register_file_inst1_cpsrin[1]), .CP(clock), .Q(RF_OUT_z) );
  DFQD1BWP12T register_file_inst1_cpsr_reg_2_ ( .D(
        register_file_inst1_cpsrin[2]), .CP(clock), .Q(RF_OUT_c) );
  DFQD1BWP12T register_file_inst1_cpsr_reg_3_ ( .D(
        register_file_inst1_cpsrin[3]), .CP(clock), .Q(RF_OUT_n) );
  DFQD1BWP12T register_file_inst1_pc_reg_0_ ( .D(register_file_inst1_n2169), 
        .CP(clock), .Q(RF_pc_out[0]) );
  DFQD1BWP12T register_file_inst1_pc_reg_2_ ( .D(register_file_inst1_n2171), 
        .CP(clock), .Q(RF_pc_out[2]) );
  DFQD1BWP12T register_file_inst1_pc_reg_3_ ( .D(register_file_inst1_n2172), 
        .CP(clock), .Q(RF_pc_out[3]) );
  DFQD1BWP12T register_file_inst1_pc_reg_4_ ( .D(register_file_inst1_n2173), 
        .CP(clock), .Q(RF_pc_out[4]) );
  DFQD1BWP12T register_file_inst1_pc_reg_5_ ( .D(register_file_inst1_n2174), 
        .CP(clock), .Q(RF_pc_out[5]) );
  DFQD1BWP12T register_file_inst1_pc_reg_6_ ( .D(register_file_inst1_n2175), 
        .CP(clock), .Q(RF_pc_out[6]) );
  DFQD1BWP12T register_file_inst1_pc_reg_7_ ( .D(register_file_inst1_n2176), 
        .CP(clock), .Q(RF_pc_out[7]) );
  DFQD1BWP12T register_file_inst1_pc_reg_8_ ( .D(register_file_inst1_n2177), 
        .CP(clock), .Q(RF_pc_out[8]) );
  DFQD1BWP12T register_file_inst1_pc_reg_9_ ( .D(register_file_inst1_n2178), 
        .CP(clock), .Q(RF_pc_out[9]) );
  DFQD1BWP12T register_file_inst1_pc_reg_10_ ( .D(register_file_inst1_n2179), 
        .CP(clock), .Q(RF_pc_out[10]) );
  DFQD1BWP12T register_file_inst1_pc_reg_11_ ( .D(register_file_inst1_n2180), 
        .CP(clock), .Q(RF_pc_out[11]) );
  DFQD1BWP12T register_file_inst1_pc_reg_12_ ( .D(register_file_inst1_n2181), 
        .CP(clock), .Q(RF_pc_out[12]) );
  DFQD1BWP12T register_file_inst1_pc_reg_13_ ( .D(register_file_inst1_n2182), 
        .CP(clock), .Q(RF_pc_out[13]) );
  DFQD1BWP12T register_file_inst1_pc_reg_14_ ( .D(register_file_inst1_n2183), 
        .CP(clock), .Q(RF_pc_out[14]) );
  DFQD1BWP12T register_file_inst1_pc_reg_15_ ( .D(register_file_inst1_n2184), 
        .CP(clock), .Q(RF_pc_out[15]) );
  DFQD1BWP12T register_file_inst1_pc_reg_16_ ( .D(register_file_inst1_n2185), 
        .CP(clock), .Q(RF_pc_out[16]) );
  DFQD1BWP12T register_file_inst1_pc_reg_17_ ( .D(register_file_inst1_n2186), 
        .CP(clock), .Q(RF_pc_out[17]) );
  DFQD1BWP12T register_file_inst1_pc_reg_18_ ( .D(register_file_inst1_n2187), 
        .CP(clock), .Q(RF_pc_out[18]) );
  DFQD1BWP12T register_file_inst1_pc_reg_19_ ( .D(register_file_inst1_n2188), 
        .CP(clock), .Q(RF_pc_out[19]) );
  DFQD1BWP12T register_file_inst1_pc_reg_20_ ( .D(register_file_inst1_n2189), 
        .CP(clock), .Q(RF_pc_out[20]) );
  DFQD1BWP12T register_file_inst1_pc_reg_21_ ( .D(register_file_inst1_n2190), 
        .CP(clock), .Q(RF_pc_out[21]) );
  DFQD1BWP12T register_file_inst1_pc_reg_22_ ( .D(register_file_inst1_n2191), 
        .CP(clock), .Q(RF_pc_out[22]) );
  DFQD1BWP12T register_file_inst1_pc_reg_23_ ( .D(register_file_inst1_n2192), 
        .CP(clock), .Q(RF_pc_out[23]) );
  DFQD1BWP12T register_file_inst1_pc_reg_24_ ( .D(register_file_inst1_n2193), 
        .CP(clock), .Q(RF_pc_out[24]) );
  DFQD1BWP12T register_file_inst1_pc_reg_25_ ( .D(register_file_inst1_n2194), 
        .CP(clock), .Q(RF_pc_out[25]) );
  DFQD1BWP12T register_file_inst1_pc_reg_26_ ( .D(register_file_inst1_n2195), 
        .CP(clock), .Q(RF_pc_out[26]) );
  DFQD1BWP12T register_file_inst1_pc_reg_27_ ( .D(register_file_inst1_n2196), 
        .CP(clock), .Q(RF_pc_out[27]) );
  DFQD1BWP12T register_file_inst1_pc_reg_28_ ( .D(register_file_inst1_n2197), 
        .CP(clock), .Q(RF_pc_out[28]) );
  DFQD1BWP12T register_file_inst1_pc_reg_29_ ( .D(register_file_inst1_n2198), 
        .CP(clock), .Q(RF_pc_out[29]) );
  DFQD1BWP12T register_file_inst1_pc_reg_30_ ( .D(register_file_inst1_n2199), 
        .CP(clock), .Q(RF_pc_out[30]) );
  DFQD1BWP12T register_file_inst1_pc_reg_31_ ( .D(register_file_inst1_n2200), 
        .CP(clock), .Q(RF_pc_out[31]) );
  DFQD1BWP12T register_file_inst1_sp_reg_5_ ( .D(register_file_inst1_spin[5]), 
        .CP(clock), .Q(STACK_RF_next_sp[5]) );
  DFQD1BWP12T register_file_inst1_sp_reg_6_ ( .D(register_file_inst1_spin[6]), 
        .CP(clock), .Q(STACK_RF_next_sp[6]) );
  DFQD1BWP12T register_file_inst1_sp_reg_7_ ( .D(register_file_inst1_spin[7]), 
        .CP(clock), .Q(STACK_RF_next_sp[7]) );
  DFQD1BWP12T register_file_inst1_sp_reg_8_ ( .D(register_file_inst1_spin[8]), 
        .CP(clock), .Q(STACK_RF_next_sp[8]) );
  DFQD1BWP12T register_file_inst1_sp_reg_9_ ( .D(register_file_inst1_spin[9]), 
        .CP(clock), .Q(STACK_RF_next_sp[9]) );
  DFQD1BWP12T register_file_inst1_sp_reg_10_ ( .D(register_file_inst1_spin[10]), .CP(clock), .Q(STACK_RF_next_sp[10]) );
  DFQD1BWP12T register_file_inst1_sp_reg_11_ ( .D(register_file_inst1_spin[11]), .CP(clock), .Q(STACK_RF_next_sp[11]) );
  DFQD1BWP12T register_file_inst1_sp_reg_12_ ( .D(register_file_inst1_spin[12]), .CP(clock), .Q(STACK_RF_next_sp[12]) );
  DFQD1BWP12T register_file_inst1_sp_reg_13_ ( .D(register_file_inst1_spin[13]), .CP(clock), .Q(STACK_RF_next_sp[13]) );
  DFQD1BWP12T register_file_inst1_sp_reg_14_ ( .D(register_file_inst1_spin[14]), .CP(clock), .Q(STACK_RF_next_sp[14]) );
  DFQD1BWP12T register_file_inst1_sp_reg_15_ ( .D(register_file_inst1_spin[15]), .CP(clock), .Q(STACK_RF_next_sp[15]) );
  DFQD1BWP12T register_file_inst1_sp_reg_16_ ( .D(register_file_inst1_spin[16]), .CP(clock), .Q(STACK_RF_next_sp[16]) );
  DFQD1BWP12T register_file_inst1_sp_reg_17_ ( .D(register_file_inst1_spin[17]), .CP(clock), .Q(STACK_RF_next_sp[17]) );
  DFQD1BWP12T register_file_inst1_sp_reg_18_ ( .D(register_file_inst1_spin[18]), .CP(clock), .Q(STACK_RF_next_sp[18]) );
  DFQD1BWP12T register_file_inst1_sp_reg_19_ ( .D(register_file_inst1_spin[19]), .CP(clock), .Q(STACK_RF_next_sp[19]) );
  DFQD1BWP12T register_file_inst1_sp_reg_20_ ( .D(register_file_inst1_spin[20]), .CP(clock), .Q(STACK_RF_next_sp[20]) );
  DFQD1BWP12T register_file_inst1_sp_reg_21_ ( .D(register_file_inst1_spin[21]), .CP(clock), .Q(STACK_RF_next_sp[21]) );
  DFQD1BWP12T register_file_inst1_sp_reg_22_ ( .D(register_file_inst1_spin[22]), .CP(clock), .Q(STACK_RF_next_sp[22]) );
  DFQD1BWP12T register_file_inst1_sp_reg_23_ ( .D(register_file_inst1_spin[23]), .CP(clock), .Q(STACK_RF_next_sp[23]) );
  DFQD1BWP12T register_file_inst1_sp_reg_24_ ( .D(register_file_inst1_spin[24]), .CP(clock), .Q(STACK_RF_next_sp[24]) );
  DFQD1BWP12T register_file_inst1_sp_reg_25_ ( .D(register_file_inst1_spin[25]), .CP(clock), .Q(STACK_RF_next_sp[25]) );
  DFQD1BWP12T register_file_inst1_sp_reg_26_ ( .D(register_file_inst1_spin[26]), .CP(clock), .Q(STACK_RF_next_sp[26]) );
  DFQD1BWP12T register_file_inst1_sp_reg_27_ ( .D(register_file_inst1_spin[27]), .CP(clock), .Q(STACK_RF_next_sp[27]) );
  DFQD1BWP12T register_file_inst1_sp_reg_28_ ( .D(register_file_inst1_spin[28]), .CP(clock), .Q(STACK_RF_next_sp[28]) );
  DFQD1BWP12T register_file_inst1_sp_reg_29_ ( .D(register_file_inst1_spin[29]), .CP(clock), .Q(STACK_RF_next_sp[29]) );
  DFQD1BWP12T register_file_inst1_sp_reg_30_ ( .D(register_file_inst1_spin[30]), .CP(clock), .Q(STACK_RF_next_sp[30]) );
  DFQD1BWP12T register_file_inst1_sp_reg_31_ ( .D(register_file_inst1_spin[31]), .CP(clock), .Q(STACK_RF_next_sp[31]) );
  DFQD1BWP12T register_file_inst1_lr_reg_0_ ( .D(register_file_inst1_n2201), 
        .CP(clock), .Q(register_file_inst1_lr_0_) );
  DFQD1BWP12T register_file_inst1_lr_reg_2_ ( .D(register_file_inst1_n2203), 
        .CP(clock), .Q(register_file_inst1_lr_2_) );
  DFQD1BWP12T register_file_inst1_lr_reg_3_ ( .D(register_file_inst1_n2204), 
        .CP(clock), .Q(register_file_inst1_lr_3_) );
  DFQD1BWP12T register_file_inst1_lr_reg_4_ ( .D(register_file_inst1_n2205), 
        .CP(clock), .Q(register_file_inst1_lr_4_) );
  DFQD1BWP12T register_file_inst1_lr_reg_5_ ( .D(register_file_inst1_n2206), 
        .CP(clock), .Q(register_file_inst1_lr_5_) );
  DFQD1BWP12T register_file_inst1_lr_reg_6_ ( .D(register_file_inst1_n2207), 
        .CP(clock), .Q(register_file_inst1_lr_6_) );
  DFQD1BWP12T register_file_inst1_lr_reg_7_ ( .D(register_file_inst1_n2208), 
        .CP(clock), .Q(register_file_inst1_lr_7_) );
  DFQD1BWP12T register_file_inst1_lr_reg_8_ ( .D(register_file_inst1_n2209), 
        .CP(clock), .Q(register_file_inst1_lr_8_) );
  DFQD1BWP12T register_file_inst1_lr_reg_9_ ( .D(register_file_inst1_n2210), 
        .CP(clock), .Q(register_file_inst1_lr_9_) );
  DFQD1BWP12T register_file_inst1_lr_reg_10_ ( .D(register_file_inst1_n2211), 
        .CP(clock), .Q(register_file_inst1_lr_10_) );
  DFQD1BWP12T register_file_inst1_lr_reg_11_ ( .D(register_file_inst1_n2212), 
        .CP(clock), .Q(register_file_inst1_lr_11_) );
  DFQD1BWP12T register_file_inst1_lr_reg_12_ ( .D(register_file_inst1_n2213), 
        .CP(clock), .Q(register_file_inst1_lr_12_) );
  DFQD1BWP12T register_file_inst1_lr_reg_13_ ( .D(register_file_inst1_n2214), 
        .CP(clock), .Q(register_file_inst1_lr_13_) );
  DFQD1BWP12T register_file_inst1_lr_reg_14_ ( .D(register_file_inst1_n2215), 
        .CP(clock), .Q(register_file_inst1_lr_14_) );
  DFQD1BWP12T register_file_inst1_lr_reg_15_ ( .D(register_file_inst1_n2216), 
        .CP(clock), .Q(register_file_inst1_lr_15_) );
  DFQD1BWP12T register_file_inst1_lr_reg_16_ ( .D(register_file_inst1_n2217), 
        .CP(clock), .Q(register_file_inst1_lr_16_) );
  DFQD1BWP12T register_file_inst1_lr_reg_17_ ( .D(register_file_inst1_n2218), 
        .CP(clock), .Q(register_file_inst1_lr_17_) );
  DFQD1BWP12T register_file_inst1_lr_reg_18_ ( .D(register_file_inst1_n2219), 
        .CP(clock), .Q(register_file_inst1_lr_18_) );
  DFQD1BWP12T register_file_inst1_lr_reg_19_ ( .D(register_file_inst1_n2220), 
        .CP(clock), .Q(register_file_inst1_lr_19_) );
  DFQD1BWP12T register_file_inst1_lr_reg_20_ ( .D(register_file_inst1_n2221), 
        .CP(clock), .Q(register_file_inst1_lr_20_) );
  DFQD1BWP12T register_file_inst1_lr_reg_21_ ( .D(register_file_inst1_n2222), 
        .CP(clock), .Q(register_file_inst1_lr_21_) );
  DFQD1BWP12T register_file_inst1_lr_reg_22_ ( .D(register_file_inst1_n2223), 
        .CP(clock), .Q(register_file_inst1_lr_22_) );
  DFQD1BWP12T register_file_inst1_lr_reg_23_ ( .D(register_file_inst1_n2224), 
        .CP(clock), .Q(register_file_inst1_lr_23_) );
  DFQD1BWP12T register_file_inst1_lr_reg_24_ ( .D(register_file_inst1_n2225), 
        .CP(clock), .Q(register_file_inst1_lr_24_) );
  DFQD1BWP12T register_file_inst1_lr_reg_25_ ( .D(register_file_inst1_n2226), 
        .CP(clock), .Q(register_file_inst1_lr_25_) );
  DFQD1BWP12T register_file_inst1_lr_reg_26_ ( .D(register_file_inst1_n2227), 
        .CP(clock), .Q(register_file_inst1_lr_26_) );
  DFQD1BWP12T register_file_inst1_lr_reg_27_ ( .D(register_file_inst1_n2228), 
        .CP(clock), .Q(register_file_inst1_lr_27_) );
  DFQD1BWP12T register_file_inst1_lr_reg_28_ ( .D(register_file_inst1_n2229), 
        .CP(clock), .Q(register_file_inst1_lr_28_) );
  DFQD1BWP12T register_file_inst1_lr_reg_29_ ( .D(register_file_inst1_n2230), 
        .CP(clock), .Q(register_file_inst1_lr_29_) );
  DFQD1BWP12T register_file_inst1_lr_reg_30_ ( .D(register_file_inst1_n2231), 
        .CP(clock), .Q(register_file_inst1_lr_30_) );
  DFQD1BWP12T register_file_inst1_lr_reg_31_ ( .D(register_file_inst1_n2232), 
        .CP(clock), .Q(register_file_inst1_lr_31_) );
  DFQD1BWP12T register_file_inst1_r12_reg_2_ ( .D(register_file_inst1_n2235), 
        .CP(clock), .Q(register_file_inst1_r12_2_) );
  DFQD1BWP12T register_file_inst1_r12_reg_3_ ( .D(register_file_inst1_n2236), 
        .CP(clock), .Q(register_file_inst1_r12_3_) );
  DFQD1BWP12T register_file_inst1_r12_reg_4_ ( .D(register_file_inst1_n2237), 
        .CP(clock), .Q(register_file_inst1_r12_4_) );
  DFQD1BWP12T register_file_inst1_r12_reg_5_ ( .D(register_file_inst1_n2238), 
        .CP(clock), .Q(register_file_inst1_r12_5_) );
  DFQD1BWP12T register_file_inst1_r12_reg_6_ ( .D(register_file_inst1_n2239), 
        .CP(clock), .Q(register_file_inst1_r12_6_) );
  DFQD1BWP12T register_file_inst1_r12_reg_7_ ( .D(register_file_inst1_n2240), 
        .CP(clock), .Q(register_file_inst1_r12_7_) );
  DFQD1BWP12T register_file_inst1_r12_reg_8_ ( .D(register_file_inst1_n2241), 
        .CP(clock), .Q(register_file_inst1_r12_8_) );
  DFQD1BWP12T register_file_inst1_r12_reg_9_ ( .D(register_file_inst1_n2242), 
        .CP(clock), .Q(register_file_inst1_r12_9_) );
  DFQD1BWP12T register_file_inst1_r12_reg_10_ ( .D(register_file_inst1_n2243), 
        .CP(clock), .Q(register_file_inst1_r12_10_) );
  DFQD1BWP12T register_file_inst1_r12_reg_11_ ( .D(register_file_inst1_n2244), 
        .CP(clock), .Q(register_file_inst1_r12_11_) );
  DFQD1BWP12T register_file_inst1_r12_reg_12_ ( .D(register_file_inst1_n2245), 
        .CP(clock), .Q(register_file_inst1_r12_12_) );
  DFQD1BWP12T register_file_inst1_r12_reg_13_ ( .D(register_file_inst1_n2246), 
        .CP(clock), .Q(register_file_inst1_r12_13_) );
  DFQD1BWP12T register_file_inst1_r12_reg_14_ ( .D(register_file_inst1_n2247), 
        .CP(clock), .Q(register_file_inst1_r12_14_) );
  DFQD1BWP12T register_file_inst1_r12_reg_15_ ( .D(register_file_inst1_n2248), 
        .CP(clock), .Q(register_file_inst1_r12_15_) );
  DFQD1BWP12T register_file_inst1_r12_reg_16_ ( .D(register_file_inst1_n2249), 
        .CP(clock), .Q(register_file_inst1_r12_16_) );
  DFQD1BWP12T register_file_inst1_r12_reg_17_ ( .D(register_file_inst1_n2250), 
        .CP(clock), .Q(register_file_inst1_r12_17_) );
  DFQD1BWP12T register_file_inst1_r12_reg_18_ ( .D(register_file_inst1_n2251), 
        .CP(clock), .Q(register_file_inst1_r12_18_) );
  DFQD1BWP12T register_file_inst1_r12_reg_19_ ( .D(register_file_inst1_n2252), 
        .CP(clock), .Q(register_file_inst1_r12_19_) );
  DFQD1BWP12T register_file_inst1_r12_reg_20_ ( .D(register_file_inst1_n2253), 
        .CP(clock), .Q(register_file_inst1_r12_20_) );
  DFQD1BWP12T register_file_inst1_r12_reg_21_ ( .D(register_file_inst1_n2254), 
        .CP(clock), .Q(register_file_inst1_r12_21_) );
  DFQD1BWP12T register_file_inst1_r12_reg_22_ ( .D(register_file_inst1_n2255), 
        .CP(clock), .Q(register_file_inst1_r12_22_) );
  DFQD1BWP12T register_file_inst1_r12_reg_23_ ( .D(register_file_inst1_n2256), 
        .CP(clock), .Q(register_file_inst1_r12_23_) );
  DFQD1BWP12T register_file_inst1_r12_reg_24_ ( .D(register_file_inst1_n2257), 
        .CP(clock), .Q(register_file_inst1_r12_24_) );
  DFQD1BWP12T register_file_inst1_r12_reg_25_ ( .D(register_file_inst1_n2258), 
        .CP(clock), .Q(register_file_inst1_r12_25_) );
  DFQD1BWP12T register_file_inst1_r12_reg_26_ ( .D(register_file_inst1_n2259), 
        .CP(clock), .Q(register_file_inst1_r12_26_) );
  DFQD1BWP12T register_file_inst1_r12_reg_27_ ( .D(register_file_inst1_n2260), 
        .CP(clock), .Q(register_file_inst1_r12_27_) );
  DFQD1BWP12T register_file_inst1_r12_reg_28_ ( .D(register_file_inst1_n2261), 
        .CP(clock), .Q(register_file_inst1_r12_28_) );
  DFQD1BWP12T register_file_inst1_r12_reg_29_ ( .D(register_file_inst1_n2262), 
        .CP(clock), .Q(register_file_inst1_r12_29_) );
  DFQD1BWP12T register_file_inst1_r12_reg_30_ ( .D(register_file_inst1_n2263), 
        .CP(clock), .Q(register_file_inst1_r12_30_) );
  DFQD1BWP12T register_file_inst1_r12_reg_31_ ( .D(register_file_inst1_n2264), 
        .CP(clock), .Q(register_file_inst1_r12_31_) );
  DFQD1BWP12T register_file_inst1_r11_reg_0_ ( .D(register_file_inst1_n2265), 
        .CP(clock), .Q(register_file_inst1_r11_0_) );
  DFQD1BWP12T register_file_inst1_r11_reg_2_ ( .D(register_file_inst1_n2267), 
        .CP(clock), .Q(register_file_inst1_r11_2_) );
  DFQD1BWP12T register_file_inst1_r11_reg_3_ ( .D(register_file_inst1_n2268), 
        .CP(clock), .Q(register_file_inst1_r11_3_) );
  DFQD1BWP12T register_file_inst1_r11_reg_4_ ( .D(register_file_inst1_n2269), 
        .CP(clock), .Q(register_file_inst1_r11_4_) );
  DFQD1BWP12T register_file_inst1_r11_reg_5_ ( .D(register_file_inst1_n2270), 
        .CP(clock), .Q(register_file_inst1_r11_5_) );
  DFQD1BWP12T register_file_inst1_r11_reg_6_ ( .D(register_file_inst1_n2271), 
        .CP(clock), .Q(register_file_inst1_r11_6_) );
  DFQD1BWP12T register_file_inst1_r11_reg_7_ ( .D(register_file_inst1_n2272), 
        .CP(clock), .Q(register_file_inst1_r11_7_) );
  DFQD1BWP12T register_file_inst1_r11_reg_8_ ( .D(register_file_inst1_n2273), 
        .CP(clock), .Q(register_file_inst1_r11_8_) );
  DFQD1BWP12T register_file_inst1_r11_reg_9_ ( .D(register_file_inst1_n2274), 
        .CP(clock), .Q(register_file_inst1_r11_9_) );
  DFQD1BWP12T register_file_inst1_r11_reg_10_ ( .D(register_file_inst1_n2275), 
        .CP(clock), .Q(register_file_inst1_r11_10_) );
  DFQD1BWP12T register_file_inst1_r11_reg_11_ ( .D(register_file_inst1_n2276), 
        .CP(clock), .Q(register_file_inst1_r11_11_) );
  DFQD1BWP12T register_file_inst1_r11_reg_12_ ( .D(register_file_inst1_n2277), 
        .CP(clock), .Q(register_file_inst1_r11_12_) );
  DFQD1BWP12T register_file_inst1_r11_reg_13_ ( .D(register_file_inst1_n2278), 
        .CP(clock), .Q(register_file_inst1_r11_13_) );
  DFQD1BWP12T register_file_inst1_r11_reg_14_ ( .D(register_file_inst1_n2279), 
        .CP(clock), .Q(register_file_inst1_r11_14_) );
  DFQD1BWP12T register_file_inst1_r11_reg_15_ ( .D(register_file_inst1_n2280), 
        .CP(clock), .Q(register_file_inst1_r11_15_) );
  DFQD1BWP12T register_file_inst1_r11_reg_16_ ( .D(register_file_inst1_n2281), 
        .CP(clock), .Q(register_file_inst1_r11_16_) );
  DFQD1BWP12T register_file_inst1_r11_reg_17_ ( .D(register_file_inst1_n2282), 
        .CP(clock), .Q(register_file_inst1_r11_17_) );
  DFQD1BWP12T register_file_inst1_r11_reg_18_ ( .D(register_file_inst1_n2283), 
        .CP(clock), .Q(register_file_inst1_r11_18_) );
  DFQD1BWP12T register_file_inst1_r11_reg_19_ ( .D(register_file_inst1_n2284), 
        .CP(clock), .Q(register_file_inst1_r11_19_) );
  DFQD1BWP12T register_file_inst1_r11_reg_20_ ( .D(register_file_inst1_n2285), 
        .CP(clock), .Q(register_file_inst1_r11_20_) );
  DFQD1BWP12T register_file_inst1_r11_reg_21_ ( .D(register_file_inst1_n2286), 
        .CP(clock), .Q(register_file_inst1_r11_21_) );
  DFQD1BWP12T register_file_inst1_r11_reg_22_ ( .D(register_file_inst1_n2287), 
        .CP(clock), .Q(register_file_inst1_r11_22_) );
  DFQD1BWP12T register_file_inst1_r11_reg_23_ ( .D(register_file_inst1_n2288), 
        .CP(clock), .Q(register_file_inst1_r11_23_) );
  DFQD1BWP12T register_file_inst1_r11_reg_24_ ( .D(register_file_inst1_n2289), 
        .CP(clock), .Q(register_file_inst1_r11_24_) );
  DFQD1BWP12T register_file_inst1_r11_reg_25_ ( .D(register_file_inst1_n2290), 
        .CP(clock), .Q(register_file_inst1_r11_25_) );
  DFQD1BWP12T register_file_inst1_r11_reg_26_ ( .D(register_file_inst1_n2291), 
        .CP(clock), .Q(register_file_inst1_r11_26_) );
  DFQD1BWP12T register_file_inst1_r11_reg_27_ ( .D(register_file_inst1_n2292), 
        .CP(clock), .Q(register_file_inst1_r11_27_) );
  DFQD1BWP12T register_file_inst1_r11_reg_28_ ( .D(register_file_inst1_n2293), 
        .CP(clock), .Q(register_file_inst1_r11_28_) );
  DFQD1BWP12T register_file_inst1_r11_reg_29_ ( .D(register_file_inst1_n2294), 
        .CP(clock), .Q(register_file_inst1_r11_29_) );
  DFQD1BWP12T register_file_inst1_r11_reg_30_ ( .D(register_file_inst1_n2295), 
        .CP(clock), .Q(register_file_inst1_r11_30_) );
  DFQD1BWP12T register_file_inst1_r11_reg_31_ ( .D(register_file_inst1_n2296), 
        .CP(clock), .Q(register_file_inst1_r11_31_) );
  DFQD1BWP12T register_file_inst1_r10_reg_0_ ( .D(register_file_inst1_n2297), 
        .CP(clock), .Q(register_file_inst1_r10_0_) );
  DFQD1BWP12T register_file_inst1_r10_reg_2_ ( .D(register_file_inst1_n2299), 
        .CP(clock), .Q(register_file_inst1_r10_2_) );
  DFQD1BWP12T register_file_inst1_r10_reg_3_ ( .D(register_file_inst1_n2300), 
        .CP(clock), .Q(register_file_inst1_r10_3_) );
  DFQD1BWP12T register_file_inst1_r10_reg_4_ ( .D(register_file_inst1_n2301), 
        .CP(clock), .Q(register_file_inst1_r10_4_) );
  DFQD1BWP12T register_file_inst1_r10_reg_5_ ( .D(register_file_inst1_n2302), 
        .CP(clock), .Q(register_file_inst1_r10_5_) );
  DFQD1BWP12T register_file_inst1_r10_reg_6_ ( .D(register_file_inst1_n2303), 
        .CP(clock), .Q(register_file_inst1_r10_6_) );
  DFQD1BWP12T register_file_inst1_r10_reg_7_ ( .D(register_file_inst1_n2304), 
        .CP(clock), .Q(register_file_inst1_r10_7_) );
  DFQD1BWP12T register_file_inst1_r10_reg_8_ ( .D(register_file_inst1_n2305), 
        .CP(clock), .Q(register_file_inst1_r10_8_) );
  DFQD1BWP12T register_file_inst1_r10_reg_9_ ( .D(register_file_inst1_n2306), 
        .CP(clock), .Q(register_file_inst1_r10_9_) );
  DFQD1BWP12T register_file_inst1_r10_reg_10_ ( .D(register_file_inst1_n2307), 
        .CP(clock), .Q(register_file_inst1_r10_10_) );
  DFQD1BWP12T register_file_inst1_r10_reg_11_ ( .D(register_file_inst1_n2308), 
        .CP(clock), .Q(register_file_inst1_r10_11_) );
  DFQD1BWP12T register_file_inst1_r10_reg_12_ ( .D(register_file_inst1_n2309), 
        .CP(clock), .Q(register_file_inst1_r10_12_) );
  DFQD1BWP12T register_file_inst1_r10_reg_13_ ( .D(register_file_inst1_n2310), 
        .CP(clock), .Q(register_file_inst1_r10_13_) );
  DFQD1BWP12T register_file_inst1_r10_reg_14_ ( .D(register_file_inst1_n2311), 
        .CP(clock), .Q(register_file_inst1_r10_14_) );
  DFQD1BWP12T register_file_inst1_r10_reg_15_ ( .D(register_file_inst1_n2312), 
        .CP(clock), .Q(register_file_inst1_r10_15_) );
  DFQD1BWP12T register_file_inst1_r10_reg_16_ ( .D(register_file_inst1_n2313), 
        .CP(clock), .Q(register_file_inst1_r10_16_) );
  DFQD1BWP12T register_file_inst1_r10_reg_17_ ( .D(register_file_inst1_n2314), 
        .CP(clock), .Q(register_file_inst1_r10_17_) );
  DFQD1BWP12T register_file_inst1_r10_reg_18_ ( .D(register_file_inst1_n2315), 
        .CP(clock), .Q(register_file_inst1_r10_18_) );
  DFQD1BWP12T register_file_inst1_r10_reg_19_ ( .D(register_file_inst1_n2316), 
        .CP(clock), .Q(register_file_inst1_r10_19_) );
  DFQD1BWP12T register_file_inst1_r10_reg_20_ ( .D(register_file_inst1_n2317), 
        .CP(clock), .Q(register_file_inst1_r10_20_) );
  DFQD1BWP12T register_file_inst1_r10_reg_21_ ( .D(register_file_inst1_n2318), 
        .CP(clock), .Q(register_file_inst1_r10_21_) );
  DFQD1BWP12T register_file_inst1_r10_reg_22_ ( .D(register_file_inst1_n2319), 
        .CP(clock), .Q(register_file_inst1_r10_22_) );
  DFQD1BWP12T register_file_inst1_r10_reg_23_ ( .D(register_file_inst1_n2320), 
        .CP(clock), .Q(register_file_inst1_r10_23_) );
  DFQD1BWP12T register_file_inst1_r10_reg_24_ ( .D(register_file_inst1_n2321), 
        .CP(clock), .Q(register_file_inst1_r10_24_) );
  DFQD1BWP12T register_file_inst1_r10_reg_25_ ( .D(register_file_inst1_n2322), 
        .CP(clock), .Q(register_file_inst1_r10_25_) );
  DFQD1BWP12T register_file_inst1_r10_reg_26_ ( .D(register_file_inst1_n2323), 
        .CP(clock), .Q(register_file_inst1_r10_26_) );
  DFQD1BWP12T register_file_inst1_r10_reg_27_ ( .D(register_file_inst1_n2324), 
        .CP(clock), .Q(register_file_inst1_r10_27_) );
  DFQD1BWP12T register_file_inst1_r10_reg_28_ ( .D(register_file_inst1_n2325), 
        .CP(clock), .Q(register_file_inst1_r10_28_) );
  DFQD1BWP12T register_file_inst1_r10_reg_29_ ( .D(register_file_inst1_n2326), 
        .CP(clock), .Q(register_file_inst1_r10_29_) );
  DFQD1BWP12T register_file_inst1_r10_reg_30_ ( .D(register_file_inst1_n2327), 
        .CP(clock), .Q(register_file_inst1_r10_30_) );
  DFQD1BWP12T register_file_inst1_r10_reg_31_ ( .D(register_file_inst1_n2328), 
        .CP(clock), .Q(register_file_inst1_r10_31_) );
  DFQD1BWP12T register_file_inst1_r9_reg_2_ ( .D(register_file_inst1_n2331), 
        .CP(clock), .Q(register_file_inst1_r9_2_) );
  DFQD1BWP12T register_file_inst1_r9_reg_3_ ( .D(register_file_inst1_n2332), 
        .CP(clock), .Q(register_file_inst1_r9_3_) );
  DFQD1BWP12T register_file_inst1_r9_reg_4_ ( .D(register_file_inst1_n2333), 
        .CP(clock), .Q(register_file_inst1_r9_4_) );
  DFQD1BWP12T register_file_inst1_r9_reg_5_ ( .D(register_file_inst1_n2334), 
        .CP(clock), .Q(register_file_inst1_r9_5_) );
  DFQD1BWP12T register_file_inst1_r9_reg_6_ ( .D(register_file_inst1_n2335), 
        .CP(clock), .Q(register_file_inst1_r9_6_) );
  DFQD1BWP12T register_file_inst1_r9_reg_7_ ( .D(register_file_inst1_n2336), 
        .CP(clock), .Q(register_file_inst1_r9_7_) );
  DFQD1BWP12T register_file_inst1_r9_reg_8_ ( .D(register_file_inst1_n2337), 
        .CP(clock), .Q(register_file_inst1_r9_8_) );
  DFQD1BWP12T register_file_inst1_r9_reg_9_ ( .D(register_file_inst1_n2338), 
        .CP(clock), .Q(register_file_inst1_r9_9_) );
  DFQD1BWP12T register_file_inst1_r9_reg_10_ ( .D(register_file_inst1_n2339), 
        .CP(clock), .Q(register_file_inst1_r9_10_) );
  DFQD1BWP12T register_file_inst1_r9_reg_11_ ( .D(register_file_inst1_n2340), 
        .CP(clock), .Q(register_file_inst1_r9_11_) );
  DFQD1BWP12T register_file_inst1_r9_reg_12_ ( .D(register_file_inst1_n2341), 
        .CP(clock), .Q(register_file_inst1_r9_12_) );
  DFQD1BWP12T register_file_inst1_r9_reg_13_ ( .D(register_file_inst1_n2342), 
        .CP(clock), .Q(register_file_inst1_r9_13_) );
  DFQD1BWP12T register_file_inst1_r9_reg_14_ ( .D(register_file_inst1_n2343), 
        .CP(clock), .Q(register_file_inst1_r9_14_) );
  DFQD1BWP12T register_file_inst1_r9_reg_15_ ( .D(register_file_inst1_n2344), 
        .CP(clock), .Q(register_file_inst1_r9_15_) );
  DFQD1BWP12T register_file_inst1_r9_reg_16_ ( .D(register_file_inst1_n2345), 
        .CP(clock), .Q(register_file_inst1_r9_16_) );
  DFQD1BWP12T register_file_inst1_r9_reg_17_ ( .D(register_file_inst1_n2346), 
        .CP(clock), .Q(register_file_inst1_r9_17_) );
  DFQD1BWP12T register_file_inst1_r9_reg_18_ ( .D(register_file_inst1_n2347), 
        .CP(clock), .Q(register_file_inst1_r9_18_) );
  DFQD1BWP12T register_file_inst1_r9_reg_19_ ( .D(register_file_inst1_n2348), 
        .CP(clock), .Q(register_file_inst1_r9_19_) );
  DFQD1BWP12T register_file_inst1_r9_reg_20_ ( .D(register_file_inst1_n2349), 
        .CP(clock), .Q(register_file_inst1_r9_20_) );
  DFQD1BWP12T register_file_inst1_r9_reg_21_ ( .D(register_file_inst1_n2350), 
        .CP(clock), .Q(register_file_inst1_r9_21_) );
  DFQD1BWP12T register_file_inst1_r9_reg_22_ ( .D(register_file_inst1_n2351), 
        .CP(clock), .Q(register_file_inst1_r9_22_) );
  DFQD1BWP12T register_file_inst1_r9_reg_23_ ( .D(register_file_inst1_n2352), 
        .CP(clock), .Q(register_file_inst1_r9_23_) );
  DFQD1BWP12T register_file_inst1_r9_reg_24_ ( .D(register_file_inst1_n2353), 
        .CP(clock), .Q(register_file_inst1_r9_24_) );
  DFQD1BWP12T register_file_inst1_r9_reg_25_ ( .D(register_file_inst1_n2354), 
        .CP(clock), .Q(register_file_inst1_r9_25_) );
  DFQD1BWP12T register_file_inst1_r9_reg_26_ ( .D(register_file_inst1_n2355), 
        .CP(clock), .Q(register_file_inst1_r9_26_) );
  DFQD1BWP12T register_file_inst1_r9_reg_27_ ( .D(register_file_inst1_n2356), 
        .CP(clock), .Q(register_file_inst1_r9_27_) );
  DFQD1BWP12T register_file_inst1_r9_reg_28_ ( .D(register_file_inst1_n2357), 
        .CP(clock), .Q(register_file_inst1_r9_28_) );
  DFQD1BWP12T register_file_inst1_r9_reg_29_ ( .D(register_file_inst1_n2358), 
        .CP(clock), .Q(register_file_inst1_r9_29_) );
  DFQD1BWP12T register_file_inst1_r9_reg_30_ ( .D(register_file_inst1_n2359), 
        .CP(clock), .Q(register_file_inst1_r9_30_) );
  DFQD1BWP12T register_file_inst1_r9_reg_31_ ( .D(register_file_inst1_n2360), 
        .CP(clock), .Q(register_file_inst1_r9_31_) );
  DFQD1BWP12T register_file_inst1_r8_reg_2_ ( .D(register_file_inst1_n2363), 
        .CP(clock), .Q(register_file_inst1_r8_2_) );
  DFQD1BWP12T register_file_inst1_r8_reg_3_ ( .D(register_file_inst1_n2364), 
        .CP(clock), .Q(register_file_inst1_r8_3_) );
  DFQD1BWP12T register_file_inst1_r8_reg_4_ ( .D(register_file_inst1_n2365), 
        .CP(clock), .Q(register_file_inst1_r8_4_) );
  DFQD1BWP12T register_file_inst1_r8_reg_5_ ( .D(register_file_inst1_n2366), 
        .CP(clock), .Q(register_file_inst1_r8_5_) );
  DFQD1BWP12T register_file_inst1_r8_reg_6_ ( .D(register_file_inst1_n2367), 
        .CP(clock), .Q(register_file_inst1_r8_6_) );
  DFQD1BWP12T register_file_inst1_r8_reg_7_ ( .D(register_file_inst1_n2368), 
        .CP(clock), .Q(register_file_inst1_r8_7_) );
  DFQD1BWP12T register_file_inst1_r8_reg_8_ ( .D(register_file_inst1_n2369), 
        .CP(clock), .Q(register_file_inst1_r8_8_) );
  DFQD1BWP12T register_file_inst1_r8_reg_9_ ( .D(register_file_inst1_n2370), 
        .CP(clock), .Q(register_file_inst1_r8_9_) );
  DFQD1BWP12T register_file_inst1_r8_reg_10_ ( .D(register_file_inst1_n2371), 
        .CP(clock), .Q(register_file_inst1_r8_10_) );
  DFQD1BWP12T register_file_inst1_r8_reg_11_ ( .D(register_file_inst1_n2372), 
        .CP(clock), .Q(register_file_inst1_r8_11_) );
  DFQD1BWP12T register_file_inst1_r8_reg_12_ ( .D(register_file_inst1_n2373), 
        .CP(clock), .Q(register_file_inst1_r8_12_) );
  DFQD1BWP12T register_file_inst1_r8_reg_13_ ( .D(register_file_inst1_n2374), 
        .CP(clock), .Q(register_file_inst1_r8_13_) );
  DFQD1BWP12T register_file_inst1_r8_reg_14_ ( .D(register_file_inst1_n2375), 
        .CP(clock), .Q(register_file_inst1_r8_14_) );
  DFQD1BWP12T register_file_inst1_r8_reg_15_ ( .D(register_file_inst1_n2376), 
        .CP(clock), .Q(register_file_inst1_r8_15_) );
  DFQD1BWP12T register_file_inst1_r8_reg_16_ ( .D(register_file_inst1_n2377), 
        .CP(clock), .Q(register_file_inst1_r8_16_) );
  DFQD1BWP12T register_file_inst1_r8_reg_17_ ( .D(register_file_inst1_n2378), 
        .CP(clock), .Q(register_file_inst1_r8_17_) );
  DFQD1BWP12T register_file_inst1_r8_reg_18_ ( .D(register_file_inst1_n2379), 
        .CP(clock), .Q(register_file_inst1_r8_18_) );
  DFQD1BWP12T register_file_inst1_r8_reg_19_ ( .D(register_file_inst1_n2380), 
        .CP(clock), .Q(register_file_inst1_r8_19_) );
  DFQD1BWP12T register_file_inst1_r8_reg_20_ ( .D(register_file_inst1_n2381), 
        .CP(clock), .Q(register_file_inst1_r8_20_) );
  DFQD1BWP12T register_file_inst1_r8_reg_21_ ( .D(register_file_inst1_n2382), 
        .CP(clock), .Q(register_file_inst1_r8_21_) );
  DFQD1BWP12T register_file_inst1_r8_reg_22_ ( .D(register_file_inst1_n2383), 
        .CP(clock), .Q(register_file_inst1_r8_22_) );
  DFQD1BWP12T register_file_inst1_r8_reg_23_ ( .D(register_file_inst1_n2384), 
        .CP(clock), .Q(register_file_inst1_r8_23_) );
  DFQD1BWP12T register_file_inst1_r8_reg_24_ ( .D(register_file_inst1_n2385), 
        .CP(clock), .Q(register_file_inst1_r8_24_) );
  DFQD1BWP12T register_file_inst1_r8_reg_25_ ( .D(register_file_inst1_n2386), 
        .CP(clock), .Q(register_file_inst1_r8_25_) );
  DFQD1BWP12T register_file_inst1_r8_reg_26_ ( .D(register_file_inst1_n2387), 
        .CP(clock), .Q(register_file_inst1_r8_26_) );
  DFQD1BWP12T register_file_inst1_r8_reg_27_ ( .D(register_file_inst1_n2388), 
        .CP(clock), .Q(register_file_inst1_r8_27_) );
  DFQD1BWP12T register_file_inst1_r8_reg_28_ ( .D(register_file_inst1_n2389), 
        .CP(clock), .Q(register_file_inst1_r8_28_) );
  DFQD1BWP12T register_file_inst1_r8_reg_29_ ( .D(register_file_inst1_n2390), 
        .CP(clock), .Q(register_file_inst1_r8_29_) );
  DFQD1BWP12T register_file_inst1_r8_reg_30_ ( .D(register_file_inst1_n2391), 
        .CP(clock), .Q(register_file_inst1_r8_30_) );
  DFQD1BWP12T register_file_inst1_r8_reg_31_ ( .D(register_file_inst1_n2392), 
        .CP(clock), .Q(register_file_inst1_r8_31_) );
  DFQD1BWP12T register_file_inst1_r7_reg_0_ ( .D(register_file_inst1_n2393), 
        .CP(clock), .Q(register_file_inst1_r7_0_) );
  DFQD1BWP12T register_file_inst1_r7_reg_2_ ( .D(register_file_inst1_n2395), 
        .CP(clock), .Q(register_file_inst1_r7_2_) );
  DFQD1BWP12T register_file_inst1_r7_reg_4_ ( .D(register_file_inst1_n2397), 
        .CP(clock), .Q(register_file_inst1_r7_4_) );
  DFQD1BWP12T register_file_inst1_r7_reg_5_ ( .D(register_file_inst1_n2398), 
        .CP(clock), .Q(register_file_inst1_r7_5_) );
  DFQD1BWP12T register_file_inst1_r7_reg_6_ ( .D(register_file_inst1_n2399), 
        .CP(clock), .Q(register_file_inst1_r7_6_) );
  DFQD1BWP12T register_file_inst1_r7_reg_7_ ( .D(register_file_inst1_n2400), 
        .CP(clock), .Q(register_file_inst1_r7_7_) );
  DFQD1BWP12T register_file_inst1_r7_reg_8_ ( .D(register_file_inst1_n2401), 
        .CP(clock), .Q(register_file_inst1_r7_8_) );
  DFQD1BWP12T register_file_inst1_r7_reg_9_ ( .D(register_file_inst1_n2402), 
        .CP(clock), .Q(register_file_inst1_r7_9_) );
  DFQD1BWP12T register_file_inst1_r7_reg_10_ ( .D(register_file_inst1_n2403), 
        .CP(clock), .Q(register_file_inst1_r7_10_) );
  DFQD1BWP12T register_file_inst1_r7_reg_11_ ( .D(register_file_inst1_n2404), 
        .CP(clock), .Q(register_file_inst1_r7_11_) );
  DFQD1BWP12T register_file_inst1_r7_reg_12_ ( .D(register_file_inst1_n2405), 
        .CP(clock), .Q(register_file_inst1_r7_12_) );
  DFQD1BWP12T register_file_inst1_r7_reg_13_ ( .D(register_file_inst1_n2406), 
        .CP(clock), .Q(register_file_inst1_r7_13_) );
  DFQD1BWP12T register_file_inst1_r7_reg_14_ ( .D(register_file_inst1_n2407), 
        .CP(clock), .Q(register_file_inst1_r7_14_) );
  DFQD1BWP12T register_file_inst1_r7_reg_15_ ( .D(register_file_inst1_n2408), 
        .CP(clock), .Q(register_file_inst1_r7_15_) );
  DFQD1BWP12T register_file_inst1_r7_reg_16_ ( .D(register_file_inst1_n2409), 
        .CP(clock), .Q(register_file_inst1_r7_16_) );
  DFQD1BWP12T register_file_inst1_r7_reg_17_ ( .D(register_file_inst1_n2410), 
        .CP(clock), .Q(register_file_inst1_r7_17_) );
  DFQD1BWP12T register_file_inst1_r7_reg_18_ ( .D(register_file_inst1_n2411), 
        .CP(clock), .Q(register_file_inst1_r7_18_) );
  DFQD1BWP12T register_file_inst1_r7_reg_19_ ( .D(register_file_inst1_n2412), 
        .CP(clock), .Q(register_file_inst1_r7_19_) );
  DFQD1BWP12T register_file_inst1_r7_reg_20_ ( .D(register_file_inst1_n2413), 
        .CP(clock), .Q(register_file_inst1_r7_20_) );
  DFQD1BWP12T register_file_inst1_r7_reg_21_ ( .D(register_file_inst1_n2414), 
        .CP(clock), .Q(register_file_inst1_r7_21_) );
  DFQD1BWP12T register_file_inst1_r7_reg_22_ ( .D(register_file_inst1_n2415), 
        .CP(clock), .Q(register_file_inst1_r7_22_) );
  DFQD1BWP12T register_file_inst1_r7_reg_23_ ( .D(register_file_inst1_n2416), 
        .CP(clock), .Q(register_file_inst1_r7_23_) );
  DFQD1BWP12T register_file_inst1_r7_reg_24_ ( .D(register_file_inst1_n2417), 
        .CP(clock), .Q(register_file_inst1_r7_24_) );
  DFQD1BWP12T register_file_inst1_r7_reg_25_ ( .D(register_file_inst1_n2418), 
        .CP(clock), .Q(register_file_inst1_r7_25_) );
  DFQD1BWP12T register_file_inst1_r7_reg_26_ ( .D(register_file_inst1_n2419), 
        .CP(clock), .Q(register_file_inst1_r7_26_) );
  DFQD1BWP12T register_file_inst1_r7_reg_27_ ( .D(register_file_inst1_n2420), 
        .CP(clock), .Q(register_file_inst1_r7_27_) );
  DFQD1BWP12T register_file_inst1_r7_reg_28_ ( .D(register_file_inst1_n2421), 
        .CP(clock), .Q(register_file_inst1_r7_28_) );
  DFQD1BWP12T register_file_inst1_r7_reg_29_ ( .D(register_file_inst1_n2422), 
        .CP(clock), .Q(register_file_inst1_r7_29_) );
  DFQD1BWP12T register_file_inst1_r7_reg_30_ ( .D(register_file_inst1_n2423), 
        .CP(clock), .Q(register_file_inst1_r7_30_) );
  DFQD1BWP12T register_file_inst1_r7_reg_31_ ( .D(register_file_inst1_n2424), 
        .CP(clock), .Q(register_file_inst1_r7_31_) );
  DFQD1BWP12T register_file_inst1_r6_reg_0_ ( .D(register_file_inst1_n2425), 
        .CP(clock), .Q(register_file_inst1_r6_0_) );
  DFQD1BWP12T register_file_inst1_r6_reg_2_ ( .D(register_file_inst1_n2427), 
        .CP(clock), .Q(register_file_inst1_r6_2_) );
  DFQD1BWP12T register_file_inst1_r6_reg_3_ ( .D(register_file_inst1_n2428), 
        .CP(clock), .Q(register_file_inst1_r6_3_) );
  DFQD1BWP12T register_file_inst1_r6_reg_4_ ( .D(register_file_inst1_n2429), 
        .CP(clock), .Q(register_file_inst1_r6_4_) );
  DFQD1BWP12T register_file_inst1_r6_reg_6_ ( .D(register_file_inst1_n2431), 
        .CP(clock), .Q(register_file_inst1_r6_6_) );
  DFQD1BWP12T register_file_inst1_r6_reg_7_ ( .D(register_file_inst1_n2432), 
        .CP(clock), .Q(register_file_inst1_r6_7_) );
  DFQD1BWP12T register_file_inst1_r6_reg_8_ ( .D(register_file_inst1_n2433), 
        .CP(clock), .Q(register_file_inst1_r6_8_) );
  DFQD1BWP12T register_file_inst1_r6_reg_9_ ( .D(register_file_inst1_n2434), 
        .CP(clock), .Q(register_file_inst1_r6_9_) );
  DFQD1BWP12T register_file_inst1_r6_reg_10_ ( .D(register_file_inst1_n2435), 
        .CP(clock), .Q(register_file_inst1_r6_10_) );
  DFQD1BWP12T register_file_inst1_r6_reg_11_ ( .D(register_file_inst1_n2436), 
        .CP(clock), .Q(register_file_inst1_r6_11_) );
  DFQD1BWP12T register_file_inst1_r6_reg_12_ ( .D(register_file_inst1_n2437), 
        .CP(clock), .Q(register_file_inst1_r6_12_) );
  DFQD1BWP12T register_file_inst1_r6_reg_13_ ( .D(register_file_inst1_n2438), 
        .CP(clock), .Q(register_file_inst1_r6_13_) );
  DFQD1BWP12T register_file_inst1_r6_reg_14_ ( .D(register_file_inst1_n2439), 
        .CP(clock), .Q(register_file_inst1_r6_14_) );
  DFQD1BWP12T register_file_inst1_r6_reg_15_ ( .D(register_file_inst1_n2440), 
        .CP(clock), .Q(register_file_inst1_r6_15_) );
  DFQD1BWP12T register_file_inst1_r6_reg_16_ ( .D(register_file_inst1_n2441), 
        .CP(clock), .Q(register_file_inst1_r6_16_) );
  DFQD1BWP12T register_file_inst1_r6_reg_17_ ( .D(register_file_inst1_n2442), 
        .CP(clock), .Q(register_file_inst1_r6_17_) );
  DFQD1BWP12T register_file_inst1_r6_reg_18_ ( .D(register_file_inst1_n2443), 
        .CP(clock), .Q(register_file_inst1_r6_18_) );
  DFQD1BWP12T register_file_inst1_r6_reg_19_ ( .D(register_file_inst1_n2444), 
        .CP(clock), .Q(register_file_inst1_r6_19_) );
  DFQD1BWP12T register_file_inst1_r6_reg_20_ ( .D(register_file_inst1_n2445), 
        .CP(clock), .Q(register_file_inst1_r6_20_) );
  DFQD1BWP12T register_file_inst1_r6_reg_21_ ( .D(register_file_inst1_n2446), 
        .CP(clock), .Q(register_file_inst1_r6_21_) );
  DFQD1BWP12T register_file_inst1_r6_reg_22_ ( .D(register_file_inst1_n2447), 
        .CP(clock), .Q(register_file_inst1_r6_22_) );
  DFQD1BWP12T register_file_inst1_r6_reg_23_ ( .D(register_file_inst1_n2448), 
        .CP(clock), .Q(register_file_inst1_r6_23_) );
  DFQD1BWP12T register_file_inst1_r6_reg_24_ ( .D(register_file_inst1_n2449), 
        .CP(clock), .Q(register_file_inst1_r6_24_) );
  DFQD1BWP12T register_file_inst1_r6_reg_25_ ( .D(register_file_inst1_n2450), 
        .CP(clock), .Q(register_file_inst1_r6_25_) );
  DFQD1BWP12T register_file_inst1_r6_reg_26_ ( .D(register_file_inst1_n2451), 
        .CP(clock), .Q(register_file_inst1_r6_26_) );
  DFQD1BWP12T register_file_inst1_r6_reg_27_ ( .D(register_file_inst1_n2452), 
        .CP(clock), .Q(register_file_inst1_r6_27_) );
  DFQD1BWP12T register_file_inst1_r6_reg_28_ ( .D(register_file_inst1_n2453), 
        .CP(clock), .Q(register_file_inst1_r6_28_) );
  DFQD1BWP12T register_file_inst1_r6_reg_29_ ( .D(register_file_inst1_n2454), 
        .CP(clock), .Q(register_file_inst1_r6_29_) );
  DFQD1BWP12T register_file_inst1_r6_reg_30_ ( .D(register_file_inst1_n2455), 
        .CP(clock), .Q(register_file_inst1_r6_30_) );
  DFQD1BWP12T register_file_inst1_r6_reg_31_ ( .D(register_file_inst1_n2456), 
        .CP(clock), .Q(register_file_inst1_r6_31_) );
  DFQD1BWP12T register_file_inst1_r5_reg_0_ ( .D(register_file_inst1_n2457), 
        .CP(clock), .Q(register_file_inst1_r5_0_) );
  DFQD1BWP12T register_file_inst1_r5_reg_2_ ( .D(register_file_inst1_n2459), 
        .CP(clock), .Q(register_file_inst1_r5_2_) );
  DFQD1BWP12T register_file_inst1_r5_reg_3_ ( .D(register_file_inst1_n2460), 
        .CP(clock), .Q(register_file_inst1_r5_3_) );
  DFQD1BWP12T register_file_inst1_r5_reg_4_ ( .D(register_file_inst1_n2461), 
        .CP(clock), .Q(register_file_inst1_r5_4_) );
  DFQD1BWP12T register_file_inst1_r5_reg_5_ ( .D(register_file_inst1_n2462), 
        .CP(clock), .Q(register_file_inst1_r5_5_) );
  DFQD1BWP12T register_file_inst1_r5_reg_6_ ( .D(register_file_inst1_n2463), 
        .CP(clock), .Q(register_file_inst1_r5_6_) );
  DFQD1BWP12T register_file_inst1_r5_reg_7_ ( .D(register_file_inst1_n2464), 
        .CP(clock), .Q(register_file_inst1_r5_7_) );
  DFQD1BWP12T register_file_inst1_r5_reg_8_ ( .D(register_file_inst1_n2465), 
        .CP(clock), .Q(register_file_inst1_r5_8_) );
  DFQD1BWP12T register_file_inst1_r5_reg_9_ ( .D(register_file_inst1_n2466), 
        .CP(clock), .Q(register_file_inst1_r5_9_) );
  DFQD1BWP12T register_file_inst1_r5_reg_10_ ( .D(register_file_inst1_n2467), 
        .CP(clock), .Q(register_file_inst1_r5_10_) );
  DFQD1BWP12T register_file_inst1_r5_reg_11_ ( .D(register_file_inst1_n2468), 
        .CP(clock), .Q(register_file_inst1_r5_11_) );
  DFQD1BWP12T register_file_inst1_r5_reg_12_ ( .D(register_file_inst1_n2469), 
        .CP(clock), .Q(register_file_inst1_r5_12_) );
  DFQD1BWP12T register_file_inst1_r5_reg_13_ ( .D(register_file_inst1_n2470), 
        .CP(clock), .Q(register_file_inst1_r5_13_) );
  DFQD1BWP12T register_file_inst1_r5_reg_14_ ( .D(register_file_inst1_n2471), 
        .CP(clock), .Q(register_file_inst1_r5_14_) );
  DFQD1BWP12T register_file_inst1_r5_reg_15_ ( .D(register_file_inst1_n2472), 
        .CP(clock), .Q(register_file_inst1_r5_15_) );
  DFQD1BWP12T register_file_inst1_r5_reg_16_ ( .D(register_file_inst1_n2473), 
        .CP(clock), .Q(register_file_inst1_r5_16_) );
  DFQD1BWP12T register_file_inst1_r5_reg_17_ ( .D(register_file_inst1_n2474), 
        .CP(clock), .Q(register_file_inst1_r5_17_) );
  DFQD1BWP12T register_file_inst1_r5_reg_18_ ( .D(register_file_inst1_n2475), 
        .CP(clock), .Q(register_file_inst1_r5_18_) );
  DFQD1BWP12T register_file_inst1_r5_reg_19_ ( .D(register_file_inst1_n2476), 
        .CP(clock), .Q(register_file_inst1_r5_19_) );
  DFQD1BWP12T register_file_inst1_r5_reg_20_ ( .D(register_file_inst1_n2477), 
        .CP(clock), .Q(register_file_inst1_r5_20_) );
  DFQD1BWP12T register_file_inst1_r5_reg_21_ ( .D(register_file_inst1_n2478), 
        .CP(clock), .Q(register_file_inst1_r5_21_) );
  DFQD1BWP12T register_file_inst1_r5_reg_22_ ( .D(register_file_inst1_n2479), 
        .CP(clock), .Q(register_file_inst1_r5_22_) );
  DFQD1BWP12T register_file_inst1_r5_reg_23_ ( .D(register_file_inst1_n2480), 
        .CP(clock), .Q(register_file_inst1_r5_23_) );
  DFQD1BWP12T register_file_inst1_r5_reg_24_ ( .D(register_file_inst1_n2481), 
        .CP(clock), .Q(register_file_inst1_r5_24_) );
  DFQD1BWP12T register_file_inst1_r5_reg_25_ ( .D(register_file_inst1_n2482), 
        .CP(clock), .Q(register_file_inst1_r5_25_) );
  DFQD1BWP12T register_file_inst1_r5_reg_26_ ( .D(register_file_inst1_n2483), 
        .CP(clock), .Q(register_file_inst1_r5_26_) );
  DFQD1BWP12T register_file_inst1_r5_reg_27_ ( .D(register_file_inst1_n2484), 
        .CP(clock), .Q(register_file_inst1_r5_27_) );
  DFQD1BWP12T register_file_inst1_r5_reg_28_ ( .D(register_file_inst1_n2485), 
        .CP(clock), .Q(register_file_inst1_r5_28_) );
  DFQD1BWP12T register_file_inst1_r5_reg_29_ ( .D(register_file_inst1_n2486), 
        .CP(clock), .Q(register_file_inst1_r5_29_) );
  DFQD1BWP12T register_file_inst1_r5_reg_30_ ( .D(register_file_inst1_n2487), 
        .CP(clock), .Q(register_file_inst1_r5_30_) );
  DFQD1BWP12T register_file_inst1_r5_reg_31_ ( .D(register_file_inst1_n2488), 
        .CP(clock), .Q(register_file_inst1_r5_31_) );
  DFQD1BWP12T register_file_inst1_r4_reg_0_ ( .D(register_file_inst1_n2489), 
        .CP(clock), .Q(register_file_inst1_r4_0_) );
  DFQD1BWP12T register_file_inst1_r4_reg_2_ ( .D(register_file_inst1_n2491), 
        .CP(clock), .Q(register_file_inst1_r4_2_) );
  DFQD1BWP12T register_file_inst1_r4_reg_3_ ( .D(register_file_inst1_n2492), 
        .CP(clock), .Q(register_file_inst1_r4_3_) );
  DFQD1BWP12T register_file_inst1_r4_reg_4_ ( .D(register_file_inst1_n2493), 
        .CP(clock), .Q(register_file_inst1_r4_4_) );
  DFQD1BWP12T register_file_inst1_r4_reg_5_ ( .D(register_file_inst1_n2494), 
        .CP(clock), .Q(register_file_inst1_r4_5_) );
  DFQD1BWP12T register_file_inst1_r4_reg_6_ ( .D(register_file_inst1_n2495), 
        .CP(clock), .Q(register_file_inst1_r4_6_) );
  DFQD1BWP12T register_file_inst1_r4_reg_7_ ( .D(register_file_inst1_n2496), 
        .CP(clock), .Q(register_file_inst1_r4_7_) );
  DFQD1BWP12T register_file_inst1_r4_reg_8_ ( .D(register_file_inst1_n2497), 
        .CP(clock), .Q(register_file_inst1_r4_8_) );
  DFQD1BWP12T register_file_inst1_r4_reg_9_ ( .D(register_file_inst1_n2498), 
        .CP(clock), .Q(register_file_inst1_r4_9_) );
  DFQD1BWP12T register_file_inst1_r4_reg_10_ ( .D(register_file_inst1_n2499), 
        .CP(clock), .Q(register_file_inst1_r4_10_) );
  DFQD1BWP12T register_file_inst1_r4_reg_11_ ( .D(register_file_inst1_n2500), 
        .CP(clock), .Q(register_file_inst1_r4_11_) );
  DFQD1BWP12T register_file_inst1_r4_reg_12_ ( .D(register_file_inst1_n2501), 
        .CP(clock), .Q(register_file_inst1_r4_12_) );
  DFQD1BWP12T register_file_inst1_r4_reg_13_ ( .D(register_file_inst1_n2502), 
        .CP(clock), .Q(register_file_inst1_r4_13_) );
  DFQD1BWP12T register_file_inst1_r4_reg_14_ ( .D(register_file_inst1_n2503), 
        .CP(clock), .Q(register_file_inst1_r4_14_) );
  DFQD1BWP12T register_file_inst1_r4_reg_15_ ( .D(register_file_inst1_n2504), 
        .CP(clock), .Q(register_file_inst1_r4_15_) );
  DFQD1BWP12T register_file_inst1_r4_reg_16_ ( .D(register_file_inst1_n2505), 
        .CP(clock), .Q(register_file_inst1_r4_16_) );
  DFQD1BWP12T register_file_inst1_r4_reg_17_ ( .D(register_file_inst1_n2506), 
        .CP(clock), .Q(register_file_inst1_r4_17_) );
  DFQD1BWP12T register_file_inst1_r4_reg_18_ ( .D(register_file_inst1_n2507), 
        .CP(clock), .Q(register_file_inst1_r4_18_) );
  DFQD1BWP12T register_file_inst1_r4_reg_19_ ( .D(register_file_inst1_n2508), 
        .CP(clock), .Q(register_file_inst1_r4_19_) );
  DFQD1BWP12T register_file_inst1_r4_reg_20_ ( .D(register_file_inst1_n2509), 
        .CP(clock), .Q(register_file_inst1_r4_20_) );
  DFQD1BWP12T register_file_inst1_r4_reg_21_ ( .D(register_file_inst1_n2510), 
        .CP(clock), .Q(register_file_inst1_r4_21_) );
  DFQD1BWP12T register_file_inst1_r4_reg_22_ ( .D(register_file_inst1_n2511), 
        .CP(clock), .Q(register_file_inst1_r4_22_) );
  DFQD1BWP12T register_file_inst1_r4_reg_23_ ( .D(register_file_inst1_n2512), 
        .CP(clock), .Q(register_file_inst1_r4_23_) );
  DFQD1BWP12T register_file_inst1_r4_reg_24_ ( .D(register_file_inst1_n2513), 
        .CP(clock), .Q(register_file_inst1_r4_24_) );
  DFQD1BWP12T register_file_inst1_r4_reg_25_ ( .D(register_file_inst1_n2514), 
        .CP(clock), .Q(register_file_inst1_r4_25_) );
  DFQD1BWP12T register_file_inst1_r4_reg_26_ ( .D(register_file_inst1_n2515), 
        .CP(clock), .Q(register_file_inst1_r4_26_) );
  DFQD1BWP12T register_file_inst1_r4_reg_27_ ( .D(register_file_inst1_n2516), 
        .CP(clock), .Q(register_file_inst1_r4_27_) );
  DFQD1BWP12T register_file_inst1_r4_reg_28_ ( .D(register_file_inst1_n2517), 
        .CP(clock), .Q(register_file_inst1_r4_28_) );
  DFQD1BWP12T register_file_inst1_r4_reg_29_ ( .D(register_file_inst1_n2518), 
        .CP(clock), .Q(register_file_inst1_r4_29_) );
  DFQD1BWP12T register_file_inst1_r4_reg_30_ ( .D(register_file_inst1_n2519), 
        .CP(clock), .Q(register_file_inst1_r4_30_) );
  DFQD1BWP12T register_file_inst1_r4_reg_31_ ( .D(register_file_inst1_n2520), 
        .CP(clock), .Q(register_file_inst1_r4_31_) );
  DFQD1BWP12T register_file_inst1_r3_reg_0_ ( .D(register_file_inst1_n2521), 
        .CP(clock), .Q(register_file_inst1_r3_0_) );
  DFQD1BWP12T register_file_inst1_r3_reg_2_ ( .D(register_file_inst1_n2523), 
        .CP(clock), .Q(register_file_inst1_r3_2_) );
  DFQD1BWP12T register_file_inst1_r3_reg_3_ ( .D(register_file_inst1_n2524), 
        .CP(clock), .Q(register_file_inst1_r3_3_) );
  DFQD1BWP12T register_file_inst1_r3_reg_4_ ( .D(register_file_inst1_n2525), 
        .CP(clock), .Q(register_file_inst1_r3_4_) );
  DFQD1BWP12T register_file_inst1_r3_reg_5_ ( .D(register_file_inst1_n2526), 
        .CP(clock), .Q(register_file_inst1_r3_5_) );
  DFQD1BWP12T register_file_inst1_r3_reg_6_ ( .D(register_file_inst1_n2527), 
        .CP(clock), .Q(register_file_inst1_r3_6_) );
  DFQD1BWP12T register_file_inst1_r3_reg_7_ ( .D(register_file_inst1_n2528), 
        .CP(clock), .Q(register_file_inst1_r3_7_) );
  DFQD1BWP12T register_file_inst1_r3_reg_8_ ( .D(register_file_inst1_n2529), 
        .CP(clock), .Q(register_file_inst1_r3_8_) );
  DFQD1BWP12T register_file_inst1_r3_reg_10_ ( .D(register_file_inst1_n2531), 
        .CP(clock), .Q(register_file_inst1_r3_10_) );
  DFQD1BWP12T register_file_inst1_r3_reg_11_ ( .D(register_file_inst1_n2532), 
        .CP(clock), .Q(register_file_inst1_r3_11_) );
  DFQD1BWP12T register_file_inst1_r3_reg_12_ ( .D(register_file_inst1_n2533), 
        .CP(clock), .Q(register_file_inst1_r3_12_) );
  DFQD1BWP12T register_file_inst1_r3_reg_13_ ( .D(register_file_inst1_n2534), 
        .CP(clock), .Q(register_file_inst1_r3_13_) );
  DFQD1BWP12T register_file_inst1_r3_reg_14_ ( .D(register_file_inst1_n2535), 
        .CP(clock), .Q(register_file_inst1_r3_14_) );
  DFQD1BWP12T register_file_inst1_r3_reg_15_ ( .D(register_file_inst1_n2536), 
        .CP(clock), .Q(register_file_inst1_r3_15_) );
  DFQD1BWP12T register_file_inst1_r3_reg_16_ ( .D(register_file_inst1_n2537), 
        .CP(clock), .Q(register_file_inst1_r3_16_) );
  DFQD1BWP12T register_file_inst1_r3_reg_17_ ( .D(register_file_inst1_n2538), 
        .CP(clock), .Q(register_file_inst1_r3_17_) );
  DFQD1BWP12T register_file_inst1_r3_reg_18_ ( .D(register_file_inst1_n2539), 
        .CP(clock), .Q(register_file_inst1_r3_18_) );
  DFQD1BWP12T register_file_inst1_r3_reg_19_ ( .D(register_file_inst1_n2540), 
        .CP(clock), .Q(register_file_inst1_r3_19_) );
  DFQD1BWP12T register_file_inst1_r3_reg_20_ ( .D(register_file_inst1_n2541), 
        .CP(clock), .Q(register_file_inst1_r3_20_) );
  DFQD1BWP12T register_file_inst1_r3_reg_21_ ( .D(register_file_inst1_n2542), 
        .CP(clock), .Q(register_file_inst1_r3_21_) );
  DFQD1BWP12T register_file_inst1_r3_reg_22_ ( .D(register_file_inst1_n2543), 
        .CP(clock), .Q(register_file_inst1_r3_22_) );
  DFQD1BWP12T register_file_inst1_r3_reg_23_ ( .D(register_file_inst1_n2544), 
        .CP(clock), .Q(register_file_inst1_r3_23_) );
  DFQD1BWP12T register_file_inst1_r3_reg_24_ ( .D(register_file_inst1_n2545), 
        .CP(clock), .Q(register_file_inst1_r3_24_) );
  DFQD1BWP12T register_file_inst1_r3_reg_25_ ( .D(register_file_inst1_n2546), 
        .CP(clock), .Q(register_file_inst1_r3_25_) );
  DFQD1BWP12T register_file_inst1_r3_reg_26_ ( .D(register_file_inst1_n2547), 
        .CP(clock), .Q(register_file_inst1_r3_26_) );
  DFQD1BWP12T register_file_inst1_r3_reg_27_ ( .D(register_file_inst1_n2548), 
        .CP(clock), .Q(register_file_inst1_r3_27_) );
  DFQD1BWP12T register_file_inst1_r3_reg_28_ ( .D(register_file_inst1_n2549), 
        .CP(clock), .Q(register_file_inst1_r3_28_) );
  DFQD1BWP12T register_file_inst1_r3_reg_29_ ( .D(register_file_inst1_n2550), 
        .CP(clock), .Q(register_file_inst1_r3_29_) );
  DFQD1BWP12T register_file_inst1_r3_reg_30_ ( .D(register_file_inst1_n2551), 
        .CP(clock), .Q(register_file_inst1_r3_30_) );
  DFQD1BWP12T register_file_inst1_r3_reg_31_ ( .D(register_file_inst1_n2552), 
        .CP(clock), .Q(register_file_inst1_r3_31_) );
  DFQD1BWP12T register_file_inst1_r2_reg_2_ ( .D(register_file_inst1_n2555), 
        .CP(clock), .Q(register_file_inst1_r2_2_) );
  DFQD1BWP12T register_file_inst1_r2_reg_3_ ( .D(register_file_inst1_n2556), 
        .CP(clock), .Q(register_file_inst1_r2_3_) );
  DFQD1BWP12T register_file_inst1_r2_reg_4_ ( .D(register_file_inst1_n2557), 
        .CP(clock), .Q(register_file_inst1_r2_4_) );
  DFQD1BWP12T register_file_inst1_r2_reg_5_ ( .D(register_file_inst1_n2558), 
        .CP(clock), .Q(register_file_inst1_r2_5_) );
  DFQD1BWP12T register_file_inst1_r2_reg_6_ ( .D(register_file_inst1_n2559), 
        .CP(clock), .Q(register_file_inst1_r2_6_) );
  DFQD1BWP12T register_file_inst1_r2_reg_7_ ( .D(register_file_inst1_n2560), 
        .CP(clock), .Q(register_file_inst1_r2_7_) );
  DFQD1BWP12T register_file_inst1_r2_reg_8_ ( .D(register_file_inst1_n2561), 
        .CP(clock), .Q(register_file_inst1_r2_8_) );
  DFQD1BWP12T register_file_inst1_r2_reg_9_ ( .D(register_file_inst1_n2562), 
        .CP(clock), .Q(register_file_inst1_r2_9_) );
  DFQD1BWP12T register_file_inst1_r2_reg_10_ ( .D(register_file_inst1_n2563), 
        .CP(clock), .Q(register_file_inst1_r2_10_) );
  DFQD1BWP12T register_file_inst1_r2_reg_11_ ( .D(register_file_inst1_n2564), 
        .CP(clock), .Q(register_file_inst1_r2_11_) );
  DFQD1BWP12T register_file_inst1_r2_reg_12_ ( .D(register_file_inst1_n2565), 
        .CP(clock), .Q(register_file_inst1_r2_12_) );
  DFQD1BWP12T register_file_inst1_r2_reg_13_ ( .D(register_file_inst1_n2566), 
        .CP(clock), .Q(register_file_inst1_r2_13_) );
  DFQD1BWP12T register_file_inst1_r2_reg_14_ ( .D(register_file_inst1_n2567), 
        .CP(clock), .Q(register_file_inst1_r2_14_) );
  DFQD1BWP12T register_file_inst1_r2_reg_15_ ( .D(register_file_inst1_n2568), 
        .CP(clock), .Q(register_file_inst1_r2_15_) );
  DFQD1BWP12T register_file_inst1_r2_reg_16_ ( .D(register_file_inst1_n2569), 
        .CP(clock), .Q(register_file_inst1_r2_16_) );
  DFQD1BWP12T register_file_inst1_r2_reg_17_ ( .D(register_file_inst1_n2570), 
        .CP(clock), .Q(register_file_inst1_r2_17_) );
  DFQD1BWP12T register_file_inst1_r2_reg_18_ ( .D(register_file_inst1_n2571), 
        .CP(clock), .Q(register_file_inst1_r2_18_) );
  DFQD1BWP12T register_file_inst1_r2_reg_19_ ( .D(register_file_inst1_n2572), 
        .CP(clock), .Q(register_file_inst1_r2_19_) );
  DFQD1BWP12T register_file_inst1_r2_reg_20_ ( .D(register_file_inst1_n2573), 
        .CP(clock), .Q(register_file_inst1_r2_20_) );
  DFQD1BWP12T register_file_inst1_r2_reg_21_ ( .D(register_file_inst1_n2574), 
        .CP(clock), .Q(register_file_inst1_r2_21_) );
  DFQD1BWP12T register_file_inst1_r2_reg_22_ ( .D(register_file_inst1_n2575), 
        .CP(clock), .Q(register_file_inst1_r2_22_) );
  DFQD1BWP12T register_file_inst1_r2_reg_23_ ( .D(register_file_inst1_n2576), 
        .CP(clock), .Q(register_file_inst1_r2_23_) );
  DFQD1BWP12T register_file_inst1_r2_reg_24_ ( .D(register_file_inst1_n2577), 
        .CP(clock), .Q(register_file_inst1_r2_24_) );
  DFQD1BWP12T register_file_inst1_r2_reg_25_ ( .D(register_file_inst1_n2578), 
        .CP(clock), .Q(register_file_inst1_r2_25_) );
  DFQD1BWP12T register_file_inst1_r2_reg_26_ ( .D(register_file_inst1_n2579), 
        .CP(clock), .Q(register_file_inst1_r2_26_) );
  DFQD1BWP12T register_file_inst1_r2_reg_27_ ( .D(register_file_inst1_n2580), 
        .CP(clock), .Q(register_file_inst1_r2_27_) );
  DFQD1BWP12T register_file_inst1_r2_reg_28_ ( .D(register_file_inst1_n2581), 
        .CP(clock), .Q(register_file_inst1_r2_28_) );
  DFQD1BWP12T register_file_inst1_r2_reg_29_ ( .D(register_file_inst1_n2582), 
        .CP(clock), .Q(register_file_inst1_r2_29_) );
  DFQD1BWP12T register_file_inst1_r2_reg_30_ ( .D(register_file_inst1_n2583), 
        .CP(clock), .Q(register_file_inst1_r2_30_) );
  DFQD1BWP12T register_file_inst1_r2_reg_31_ ( .D(register_file_inst1_n2584), 
        .CP(clock), .Q(register_file_inst1_r2_31_) );
  DFQD1BWP12T register_file_inst1_r1_reg_0_ ( .D(register_file_inst1_n2585), 
        .CP(clock), .Q(register_file_inst1_r1_0_) );
  DFQD1BWP12T register_file_inst1_r1_reg_2_ ( .D(register_file_inst1_n2587), 
        .CP(clock), .Q(register_file_inst1_r1_2_) );
  DFQD1BWP12T register_file_inst1_r1_reg_3_ ( .D(register_file_inst1_n2588), 
        .CP(clock), .Q(register_file_inst1_r1_3_) );
  DFQD1BWP12T register_file_inst1_r1_reg_4_ ( .D(register_file_inst1_n2589), 
        .CP(clock), .Q(register_file_inst1_r1_4_) );
  DFQD1BWP12T register_file_inst1_r1_reg_5_ ( .D(register_file_inst1_n2590), 
        .CP(clock), .Q(register_file_inst1_r1_5_) );
  DFQD1BWP12T register_file_inst1_r1_reg_6_ ( .D(register_file_inst1_n2591), 
        .CP(clock), .Q(register_file_inst1_r1_6_) );
  DFQD1BWP12T register_file_inst1_r1_reg_7_ ( .D(register_file_inst1_n2592), 
        .CP(clock), .Q(register_file_inst1_r1_7_) );
  DFQD1BWP12T register_file_inst1_r1_reg_8_ ( .D(register_file_inst1_n2593), 
        .CP(clock), .Q(register_file_inst1_r1_8_) );
  DFQD1BWP12T register_file_inst1_r1_reg_9_ ( .D(register_file_inst1_n2594), 
        .CP(clock), .Q(register_file_inst1_r1_9_) );
  DFQD1BWP12T register_file_inst1_r1_reg_10_ ( .D(register_file_inst1_n2595), 
        .CP(clock), .Q(register_file_inst1_r1_10_) );
  DFQD1BWP12T register_file_inst1_r1_reg_11_ ( .D(register_file_inst1_n2596), 
        .CP(clock), .Q(register_file_inst1_r1_11_) );
  DFQD1BWP12T register_file_inst1_r1_reg_12_ ( .D(register_file_inst1_n2597), 
        .CP(clock), .Q(register_file_inst1_r1_12_) );
  DFQD1BWP12T register_file_inst1_r1_reg_13_ ( .D(register_file_inst1_n2598), 
        .CP(clock), .Q(register_file_inst1_r1_13_) );
  DFQD1BWP12T register_file_inst1_r1_reg_14_ ( .D(register_file_inst1_n2599), 
        .CP(clock), .Q(register_file_inst1_r1_14_) );
  DFQD1BWP12T register_file_inst1_r1_reg_15_ ( .D(register_file_inst1_n2600), 
        .CP(clock), .Q(register_file_inst1_r1_15_) );
  DFQD1BWP12T register_file_inst1_r1_reg_16_ ( .D(register_file_inst1_n2601), 
        .CP(clock), .Q(register_file_inst1_r1_16_) );
  DFQD1BWP12T register_file_inst1_r1_reg_17_ ( .D(register_file_inst1_n2602), 
        .CP(clock), .Q(register_file_inst1_r1_17_) );
  DFQD1BWP12T register_file_inst1_r1_reg_18_ ( .D(register_file_inst1_n2603), 
        .CP(clock), .Q(register_file_inst1_r1_18_) );
  DFQD1BWP12T register_file_inst1_r1_reg_19_ ( .D(register_file_inst1_n2604), 
        .CP(clock), .Q(register_file_inst1_r1_19_) );
  DFQD1BWP12T register_file_inst1_r1_reg_20_ ( .D(register_file_inst1_n2605), 
        .CP(clock), .Q(register_file_inst1_r1_20_) );
  DFQD1BWP12T register_file_inst1_r1_reg_21_ ( .D(register_file_inst1_n2606), 
        .CP(clock), .Q(register_file_inst1_r1_21_) );
  DFQD1BWP12T register_file_inst1_r1_reg_22_ ( .D(register_file_inst1_n2607), 
        .CP(clock), .Q(register_file_inst1_r1_22_) );
  DFQD1BWP12T register_file_inst1_r1_reg_23_ ( .D(register_file_inst1_n2608), 
        .CP(clock), .Q(register_file_inst1_r1_23_) );
  DFQD1BWP12T register_file_inst1_r1_reg_24_ ( .D(register_file_inst1_n2609), 
        .CP(clock), .Q(register_file_inst1_r1_24_) );
  DFQD1BWP12T register_file_inst1_r1_reg_25_ ( .D(register_file_inst1_n2610), 
        .CP(clock), .Q(register_file_inst1_r1_25_) );
  DFQD1BWP12T register_file_inst1_r1_reg_26_ ( .D(register_file_inst1_n2611), 
        .CP(clock), .Q(register_file_inst1_r1_26_) );
  DFQD1BWP12T register_file_inst1_r1_reg_27_ ( .D(register_file_inst1_n2612), 
        .CP(clock), .Q(register_file_inst1_r1_27_) );
  DFQD1BWP12T register_file_inst1_r1_reg_28_ ( .D(register_file_inst1_n2613), 
        .CP(clock), .Q(register_file_inst1_r1_28_) );
  DFQD1BWP12T register_file_inst1_r1_reg_29_ ( .D(register_file_inst1_n2614), 
        .CP(clock), .Q(register_file_inst1_r1_29_) );
  DFQD1BWP12T register_file_inst1_r1_reg_30_ ( .D(register_file_inst1_n2615), 
        .CP(clock), .Q(register_file_inst1_r1_30_) );
  DFQD1BWP12T register_file_inst1_r1_reg_31_ ( .D(register_file_inst1_n2616), 
        .CP(clock), .Q(register_file_inst1_r1_31_) );
  DFQD1BWP12T register_file_inst1_r0_reg_0_ ( .D(register_file_inst1_n2617), 
        .CP(clock), .Q(register_file_inst1_r0_0_) );
  DFQD1BWP12T register_file_inst1_r0_reg_2_ ( .D(register_file_inst1_n2619), 
        .CP(clock), .Q(register_file_inst1_r0_2_) );
  DFQD1BWP12T register_file_inst1_r0_reg_3_ ( .D(register_file_inst1_n2620), 
        .CP(clock), .Q(register_file_inst1_r0_3_) );
  DFQD1BWP12T register_file_inst1_r0_reg_4_ ( .D(register_file_inst1_n2621), 
        .CP(clock), .Q(register_file_inst1_r0_4_) );
  DFQD1BWP12T register_file_inst1_r0_reg_5_ ( .D(register_file_inst1_n2622), 
        .CP(clock), .Q(register_file_inst1_r0_5_) );
  DFQD1BWP12T register_file_inst1_r0_reg_6_ ( .D(register_file_inst1_n2623), 
        .CP(clock), .Q(register_file_inst1_r0_6_) );
  DFQD1BWP12T register_file_inst1_r0_reg_7_ ( .D(register_file_inst1_n2624), 
        .CP(clock), .Q(register_file_inst1_r0_7_) );
  DFQD1BWP12T register_file_inst1_r0_reg_8_ ( .D(register_file_inst1_n2625), 
        .CP(clock), .Q(register_file_inst1_r0_8_) );
  DFQD1BWP12T register_file_inst1_r0_reg_9_ ( .D(register_file_inst1_n2626), 
        .CP(clock), .Q(register_file_inst1_r0_9_) );
  DFQD1BWP12T register_file_inst1_r0_reg_10_ ( .D(register_file_inst1_n2627), 
        .CP(clock), .Q(register_file_inst1_r0_10_) );
  DFQD1BWP12T register_file_inst1_r0_reg_11_ ( .D(register_file_inst1_n2628), 
        .CP(clock), .Q(register_file_inst1_r0_11_) );
  DFQD1BWP12T register_file_inst1_r0_reg_12_ ( .D(register_file_inst1_n2629), 
        .CP(clock), .Q(register_file_inst1_r0_12_) );
  DFQD1BWP12T register_file_inst1_r0_reg_13_ ( .D(register_file_inst1_n2630), 
        .CP(clock), .Q(register_file_inst1_r0_13_) );
  DFQD1BWP12T register_file_inst1_r0_reg_14_ ( .D(register_file_inst1_n2631), 
        .CP(clock), .Q(register_file_inst1_r0_14_) );
  DFQD1BWP12T register_file_inst1_r0_reg_15_ ( .D(register_file_inst1_n2632), 
        .CP(clock), .Q(register_file_inst1_r0_15_) );
  DFQD1BWP12T register_file_inst1_r0_reg_16_ ( .D(register_file_inst1_n2633), 
        .CP(clock), .Q(register_file_inst1_r0_16_) );
  DFQD1BWP12T register_file_inst1_r0_reg_17_ ( .D(register_file_inst1_n2634), 
        .CP(clock), .Q(register_file_inst1_r0_17_) );
  DFQD1BWP12T register_file_inst1_r0_reg_18_ ( .D(register_file_inst1_n2635), 
        .CP(clock), .Q(register_file_inst1_r0_18_) );
  DFQD1BWP12T register_file_inst1_r0_reg_19_ ( .D(register_file_inst1_n2636), 
        .CP(clock), .Q(register_file_inst1_r0_19_) );
  DFQD1BWP12T register_file_inst1_r0_reg_20_ ( .D(register_file_inst1_n2637), 
        .CP(clock), .Q(register_file_inst1_r0_20_) );
  DFQD1BWP12T register_file_inst1_r0_reg_21_ ( .D(register_file_inst1_n2638), 
        .CP(clock), .Q(register_file_inst1_r0_21_) );
  DFQD1BWP12T register_file_inst1_r0_reg_22_ ( .D(register_file_inst1_n2639), 
        .CP(clock), .Q(register_file_inst1_r0_22_) );
  DFQD1BWP12T register_file_inst1_r0_reg_23_ ( .D(register_file_inst1_n2640), 
        .CP(clock), .Q(register_file_inst1_r0_23_) );
  DFQD1BWP12T register_file_inst1_r0_reg_24_ ( .D(register_file_inst1_n2641), 
        .CP(clock), .Q(register_file_inst1_r0_24_) );
  DFQD1BWP12T register_file_inst1_r0_reg_25_ ( .D(register_file_inst1_n2642), 
        .CP(clock), .Q(register_file_inst1_r0_25_) );
  DFQD1BWP12T register_file_inst1_r0_reg_26_ ( .D(register_file_inst1_n2643), 
        .CP(clock), .Q(register_file_inst1_r0_26_) );
  DFQD1BWP12T register_file_inst1_r0_reg_27_ ( .D(register_file_inst1_n2644), 
        .CP(clock), .Q(register_file_inst1_r0_27_) );
  DFQD1BWP12T register_file_inst1_r0_reg_28_ ( .D(register_file_inst1_n2645), 
        .CP(clock), .Q(register_file_inst1_r0_28_) );
  DFQD1BWP12T register_file_inst1_r0_reg_29_ ( .D(register_file_inst1_n2646), 
        .CP(clock), .Q(register_file_inst1_r0_29_) );
  DFQD1BWP12T register_file_inst1_r0_reg_30_ ( .D(register_file_inst1_n2647), 
        .CP(clock), .Q(register_file_inst1_r0_30_) );
  DFQD1BWP12T register_file_inst1_r0_reg_31_ ( .D(register_file_inst1_n2648), 
        .CP(clock), .Q(register_file_inst1_r0_31_) );
  DFQD1BWP12T register_file_inst1_r7_reg_3_ ( .D(register_file_inst1_n2396), 
        .CP(clock), .Q(register_file_inst1_r7_3_) );
  DFQD1BWP12T register_file_inst1_r6_reg_5_ ( .D(register_file_inst1_n2430), 
        .CP(clock), .Q(register_file_inst1_r6_5_) );
  AO222D1BWP12T U12 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[11]), .B1(RF_MEMCTRL_address_reg[12]), 
        .B2(n3), .C1(ALU_MISC_OUT_result[12]), .C2(n4), .Z(
        MEMCTRL_IN_address[11]) );
  AO222D1BWP12T U15 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[8]), .B1(n4), .B2(ALU_MISC_OUT_result[9]), .C1(RF_MEMCTRL_address_reg[9]), .C2(n3), .Z(MEMCTRL_IN_address[8]) );
  AO222D1BWP12T U16 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[7]), .B1(n4), .B2(ALU_MISC_OUT_result[8]), .C1(RF_MEMCTRL_address_reg[8]), .C2(n3), .Z(MEMCTRL_IN_address[7]) );
  AO222D1BWP12T U14 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[9]), .B1(n4), .B2(
        ALU_MISC_OUT_result[10]), .C1(RF_MEMCTRL_address_reg[10]), .C2(n3), 
        .Z(MEMCTRL_IN_address[9]) );
  AO222D1BWP12T U17 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[6]), .B1(n4), .B2(ALU_MISC_OUT_result[7]), .C1(RF_MEMCTRL_address_reg[7]), .C2(n3), .Z(MEMCTRL_IN_address[6]) );
  AO222D1BWP12T U18 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[5]), .B1(n4), .B2(ALU_MISC_OUT_result[6]), .C1(RF_MEMCTRL_address_reg[6]), .C2(n3), .Z(MEMCTRL_IN_address[5]) );
  AO222D1BWP12T U19 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[4]), .B1(n4), .B2(ALU_MISC_OUT_result[5]), .C1(RF_MEMCTRL_address_reg[5]), .C2(n3), .Z(MEMCTRL_IN_address[4]) );
  AO222D1BWP12T U20 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[3]), .B1(n4), .B2(ALU_MISC_OUT_result[4]), .C1(RF_MEMCTRL_address_reg[4]), .C2(n3), .Z(MEMCTRL_IN_address[3]) );
  AO222D1BWP12T U21 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[2]), .B1(n4), .B2(ALU_MISC_OUT_result[3]), .C1(RF_MEMCTRL_address_reg[3]), .C2(n3), .Z(MEMCTRL_IN_address[2]) );
  AO222D1BWP12T U22 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[1]), .B1(n4), .B2(ALU_MISC_OUT_result[2]), .C1(RF_MEMCTRL_address_reg[2]), .C2(n3), .Z(MEMCTRL_IN_address[1]) );
  AO222D1BWP12T U13 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[10]), .B1(n4), .B2(
        ALU_MISC_OUT_result[11]), .C1(RF_MEMCTRL_address_reg[11]), .C2(n3), 
        .Z(MEMCTRL_IN_address[10]) );
  OR2XD1BWP12T U24 ( .A1(IF_memory_load_req), .A2(
        DEC_MEMCTRL_CTRL_memory_load_request), .Z(MEMCTRL_load_in) );
  CKAN2D1BWP12T U23 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[0]), .Z(MEMCTRL_IN_address[0]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_0_ ( .D(
        RF_MEMCTRL_data_reg[0]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[0]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_31_ ( .D(
        RF_MEMCTRL_data_reg[31]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[31]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_25_ ( .D(
        RF_MEMCTRL_data_reg[25]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[25]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_28_ ( .D(
        RF_MEMCTRL_data_reg[28]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[28]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_26_ ( .D(
        RF_MEMCTRL_data_reg[26]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[26]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_30_ ( .D(
        RF_MEMCTRL_data_reg[30]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[30]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_24_ ( .D(
        RF_MEMCTRL_data_reg[24]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[24]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_7_ ( .D(
        RF_MEMCTRL_data_reg[7]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_4_ ( .D(
        RF_MEMCTRL_data_reg[4]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[4]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_3_ ( .D(
        RF_MEMCTRL_data_reg[3]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_2_ ( .D(
        RF_MEMCTRL_data_reg[2]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_29_ ( .D(
        RF_MEMCTRL_data_reg[29]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[29]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_27_ ( .D(
        RF_MEMCTRL_data_reg[27]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[27]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_8_ ( .D(
        RF_MEMCTRL_data_reg[8]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_1_ ( .D(
        RF_MEMCTRL_data_reg[1]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[1]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_14_ ( .D(
        RF_MEMCTRL_data_reg[14]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[14]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_13_ ( .D(
        RF_MEMCTRL_data_reg[13]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[13]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_15_ ( .D(
        RF_MEMCTRL_data_reg[15]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[15]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_17_ ( .D(
        RF_MEMCTRL_data_reg[17]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[17]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_19_ ( .D(
        RF_MEMCTRL_data_reg[19]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[19]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_23_ ( .D(
        RF_MEMCTRL_data_reg[23]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[23]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_5_ ( .D(
        RF_MEMCTRL_data_reg[5]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[5]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_12_ ( .D(
        RF_MEMCTRL_data_reg[12]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[12]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_11_ ( .D(
        RF_MEMCTRL_data_reg[11]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[11]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_10_ ( .D(
        RF_MEMCTRL_data_reg[10]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_9_ ( .D(
        RF_MEMCTRL_data_reg[9]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_6_ ( .D(
        RF_MEMCTRL_data_reg[6]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_20_ ( .D(
        RF_MEMCTRL_data_reg[20]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[20]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_21_ ( .D(
        RF_MEMCTRL_data_reg[21]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[21]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_22_ ( .D(
        RF_MEMCTRL_data_reg[22]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[22]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_18_ ( .D(
        RF_MEMCTRL_data_reg[18]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[18]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_16_ ( .D(
        RF_MEMCTRL_data_reg[16]), .CP(clock), .Q(
        memory_interface_inst1_delay_data_in32[16]) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_2_ ( .D(
        memory_interface_inst1_fsm_N34), .CP(clock), .Q(
        memory_interface_inst1_fsm_state_2_) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_1_ ( .D(
        memory_interface_inst1_fsm_N33), .CP(clock), .Q(
        memory_interface_inst1_fsm_state_1_) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_3_ ( .D(
        memory_interface_inst1_fsm_N35), .CP(clock), .Q(
        memory_interface_inst1_fsm_state_3_) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_0_ ( .D(
        memory_interface_inst1_fsm_N32), .CP(clock), .Q(
        memory_interface_inst1_fsm_state_0_) );
  DFQD1BWP12T register_file_inst1_sp_reg_1_ ( .D(register_file_inst1_spin[1]), 
        .CP(clock), .Q(STACK_RF_next_sp[1]) );
  DFQD1BWP12T register_file_inst1_pc_reg_1_ ( .D(register_file_inst1_n2170), 
        .CP(clock), .Q(RF_pc_out[1]) );
  DFQD1BWP12T register_file_inst1_sp_reg_2_ ( .D(register_file_inst1_spin[2]), 
        .CP(clock), .Q(STACK_RF_next_sp[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_single_reg_1_ ( .D(
        MEMCTRL_IN_address[1]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_single[1]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_1_ ( .D(
        MEMCTRL_IN_address[1]), .CP(clock), .Q(
        memory_interface_inst1_delay_addr_for_adder_1_) );
  DFQD1BWP12T register_file_inst1_r12_reg_1_ ( .D(register_file_inst1_n2234), 
        .CP(clock), .Q(register_file_inst1_r12_1_) );
  DFQD1BWP12T register_file_inst1_r8_reg_1_ ( .D(register_file_inst1_n2362), 
        .CP(clock), .Q(register_file_inst1_r8_1_) );
  DFQD1BWP12T register_file_inst1_r9_reg_1_ ( .D(register_file_inst1_n2330), 
        .CP(clock), .Q(register_file_inst1_r9_1_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_1_ ( .D(register_file_inst1_n2138), 
        .CP(clock), .Q(register_file_inst1_tmp1_1_) );
  DFQD1BWP12T register_file_inst1_r11_reg_1_ ( .D(register_file_inst1_n2266), 
        .CP(clock), .Q(register_file_inst1_r11_1_) );
  DFQD1BWP12T register_file_inst1_r2_reg_1_ ( .D(register_file_inst1_n2554), 
        .CP(clock), .Q(register_file_inst1_r2_1_) );
  DFQD1BWP12T register_file_inst1_r3_reg_1_ ( .D(register_file_inst1_n2522), 
        .CP(clock), .Q(register_file_inst1_r3_1_) );
  DFQD1BWP12T register_file_inst1_r10_reg_1_ ( .D(register_file_inst1_n2298), 
        .CP(clock), .Q(register_file_inst1_r10_1_) );
  DFQD1BWP12T register_file_inst1_r4_reg_1_ ( .D(register_file_inst1_n2490), 
        .CP(clock), .Q(register_file_inst1_r4_1_) );
  DFQD1BWP12T register_file_inst1_r0_reg_1_ ( .D(register_file_inst1_n2618), 
        .CP(clock), .Q(register_file_inst1_r0_1_) );
  DFQD1BWP12T register_file_inst1_lr_reg_1_ ( .D(register_file_inst1_n2202), 
        .CP(clock), .Q(register_file_inst1_lr_1_) );
  DFQD1BWP12T register_file_inst1_r7_reg_1_ ( .D(register_file_inst1_n2394), 
        .CP(clock), .Q(register_file_inst1_r7_1_) );
  DFQD1BWP12T register_file_inst1_r5_reg_1_ ( .D(register_file_inst1_n2458), 
        .CP(clock), .Q(register_file_inst1_r5_1_) );
  DFQD1BWP12T register_file_inst1_r1_reg_1_ ( .D(register_file_inst1_n2586), 
        .CP(clock), .Q(register_file_inst1_r1_1_) );
  DFQD1BWP12T register_file_inst1_r6_reg_1_ ( .D(register_file_inst1_n2426), 
        .CP(clock), .Q(register_file_inst1_r6_1_) );
  DFQD1BWP12T register_file_inst1_sp_reg_4_ ( .D(register_file_inst1_spin[4]), 
        .CP(clock), .Q(STACK_RF_next_sp[4]) );
  DFQD1BWP12T register_file_inst1_sp_reg_0_ ( .D(register_file_inst1_spin[0]), 
        .CP(clock), .Q(STACK_RF_next_sp[0]) );
  DFQD1BWP12T register_file_inst1_sp_reg_3_ ( .D(register_file_inst1_spin[3]), 
        .CP(clock), .Q(STACK_RF_next_sp[3]) );
  DFQD1BWP12T register_file_inst1_r2_reg_0_ ( .D(register_file_inst1_n2553), 
        .CP(clock), .Q(register_file_inst1_r2_0_) );
  DFQD1BWP12T register_file_inst1_r12_reg_0_ ( .D(register_file_inst1_n2233), 
        .CP(clock), .Q(register_file_inst1_r12_0_) );
  DFQD1BWP12T register_file_inst1_r8_reg_0_ ( .D(register_file_inst1_n2361), 
        .CP(clock), .Q(register_file_inst1_r8_0_) );
  DFQD1BWP12T register_file_inst1_r9_reg_0_ ( .D(register_file_inst1_n2329), 
        .CP(clock), .Q(register_file_inst1_r9_0_) );
  DFQD1BWP12T register_file_inst1_tmp1_reg_0_ ( .D(register_file_inst1_n2136), 
        .CP(clock), .Q(register_file_inst1_tmp1_0_) );
  DFQD1BWP12T register_file_inst1_r3_reg_9_ ( .D(register_file_inst1_n2530), 
        .CP(clock), .Q(register_file_inst1_r3_9_) );
  TIELBWP12T U25 ( .ZN(n6) );
  INVD1BWP12T U26 ( .I(n6), .ZN(MEMCTRL_MEM_to_mem_mem_enable) );
  OAI22D1BWP12T U27 ( .A1(n1822), .A2(n1861), .B1(n1817), .B2(n1859), .ZN(
        n1735) );
  NR4D0BWP12T U28 ( .A1(n1677), .A2(n1676), .A3(n1675), .A4(n1674), .ZN(n1683)
         );
  NR2D1BWP12T U29 ( .A1(n2311), .A2(n2314), .ZN(n850) );
  NR2D1BWP12T U30 ( .A1(n289), .A2(n2314), .ZN(n1948) );
  NR2D1BWP12T U31 ( .A1(n2307), .A2(n2314), .ZN(n852) );
  NR2D1BWP12T U32 ( .A1(n2307), .A2(n2308), .ZN(n1947) );
  NR2D1BWP12T U33 ( .A1(n2309), .A2(n2308), .ZN(n1932) );
  NR2D1BWP12T U34 ( .A1(n284), .A2(n2311), .ZN(n845) );
  NR2D1BWP12T U35 ( .A1(n2311), .A2(n2310), .ZN(n844) );
  NR2D1BWP12T U36 ( .A1(n2310), .A2(n2309), .ZN(n841) );
  NR2D1BWP12T U37 ( .A1(n284), .A2(n289), .ZN(n843) );
  NR2D1BWP12T U38 ( .A1(n2310), .A2(n2307), .ZN(n839) );
  INVD1BWP12T U39 ( .I(DEC_RF_memory_store_data_reg[4]), .ZN(n2306) );
  INVD1BWP12T U40 ( .I(register_file_inst1_r7_5_), .ZN(n1703) );
  MUX2D1BWP12T U41 ( .I0(MEMCTRL_RF_IF_data_in[14]), .I1(
        ALU_MISC_OUT_result[14]), .S(n2277), .Z(
        register_file_inst1_pc_write_in_14_) );
  MUX2D1BWP12T U42 ( .I0(MEMCTRL_RF_IF_data_in[12]), .I1(
        ALU_MISC_OUT_result[12]), .S(n2277), .Z(
        register_file_inst1_pc_write_in_12_) );
  TPNR2D1BWP12T U43 ( .A1(n210), .A2(n16), .ZN(n917) );
  INVD1BWP12T U44 ( .I(ALU_MISC_OUT_result[31]), .ZN(n1103) );
  INVD1BWP12T U45 ( .I(ALU_MISC_OUT_result[27]), .ZN(n503) );
  INVD1BWP12T U46 ( .I(ALU_MISC_OUT_result[23]), .ZN(n511) );
  RCIAO21D0BWP12T U47 ( .A1(n2328), .A2(n885), .B(n500), .ZN(n989) );
  INVD1BWP12T U48 ( .I(ALU_MISC_OUT_result[21]), .ZN(n513) );
  INVD1BWP12T U49 ( .I(ALU_MISC_OUT_result[18]), .ZN(n218) );
  RCIAO21D0BWP12T U50 ( .A1(n2331), .A2(n885), .B(n500), .ZN(n967) );
  INVD1BWP12T U51 ( .I(MEMCTRL_RF_IF_data_in[15]), .ZN(n2135) );
  INVD1BWP12T U52 ( .I(MEMCTRL_RF_IF_data_in[14]), .ZN(n2132) );
  INVD1BWP12T U53 ( .I(MEMCTRL_RF_IF_data_in[13]), .ZN(n2129) );
  INVD1BWP12T U54 ( .I(MEMCTRL_RF_IF_data_in[12]), .ZN(n2126) );
  INVD1BWP12T U55 ( .I(MEMCTRL_RF_IF_data_in[11]), .ZN(n2123) );
  INVD1BWP12T U56 ( .I(MEMCTRL_RF_IF_data_in[10]), .ZN(n2120) );
  INVD1BWP12T U57 ( .I(MEMCTRL_RF_IF_data_in[9]), .ZN(n2117) );
  INVD1BWP12T U58 ( .I(MEMCTRL_RF_IF_data_in[8]), .ZN(n2115) );
  INVD1BWP12T U59 ( .I(n1928), .ZN(n1835) );
  NR2D1BWP12T U60 ( .A1(n2090), .A2(n2092), .ZN(n1868) );
  NR2D1BWP12T U61 ( .A1(n2090), .A2(n2094), .ZN(n1867) );
  INVD1BWP12T U62 ( .I(n1873), .ZN(n1742) );
  NR2D1BWP12T U63 ( .A1(n2181), .A2(n2176), .ZN(n1911) );
  NR2D1BWP12T U64 ( .A1(n28), .A2(n2176), .ZN(n1910) );
  ND2D1BWP12T U65 ( .A1(n30), .A2(n27), .ZN(n1903) );
  IND2D1BWP12T U66 ( .A1(n28), .B1(n31), .ZN(n1901) );
  IND2D1BWP12T U67 ( .A1(n2181), .B1(n31), .ZN(n1905) );
  NR2D1BWP12T U68 ( .A1(n107), .A2(n2093), .ZN(n1942) );
  NR2D1BWP12T U69 ( .A1(n2089), .A2(n2096), .ZN(n1941) );
  NR2D1BWP12T U70 ( .A1(n106), .A2(n2179), .ZN(n1946) );
  NR2D1BWP12T U71 ( .A1(n2175), .A2(n2182), .ZN(n1945) );
  ND3D0BWP12T U72 ( .A1(n2289), .A2(memory_interface_inst1_delayed_is_signed), 
        .A3(MEM_MEMCTRL_from_mem_data[7]), .ZN(n7) );
  CKND0BWP12T U73 ( .I(n2251), .ZN(n8) );
  AOI211D0BWP12T U74 ( .A1(n2288), .A2(
        memory_interface_inst1_delayed_is_signed), .B(n772), .C(n8), .ZN(n9)
         );
  MUX2ND0BWP12T U75 ( .I0(n2327), .I1(n7), .S(n9), .ZN(n500) );
  INVD1BWP12T U76 ( .I(ALU_MISC_OUT_result[26]), .ZN(n505) );
  INR2D0BWP12T U77 ( .A1(n2251), .B1(n2289), .ZN(n886) );
  INVD1BWP12T U78 ( .I(ALU_MISC_OUT_result[25]), .ZN(n507) );
  OR3D0BWP12T U79 ( .A1(memory_interface_inst1_fsm_state_1_), .A2(
        memory_interface_inst1_fsm_state_3_), .A3(
        memory_interface_inst1_fsm_state_2_), .Z(n498) );
  IND3D1BWP12T U80 ( .A1(n136), .B1(n2293), .B2(n1095), .ZN(n1093) );
  INVD1BWP12T U81 ( .I(ALU_MISC_OUT_result[20]), .ZN(n516) );
  INR2D0BWP12T U82 ( .A1(n634), .B1(n633), .ZN(n763) );
  IND3D1BWP12T U83 ( .A1(n118), .B1(n2293), .B2(n1092), .ZN(n1090) );
  IND2D0BWP12T U84 ( .A1(n137), .B1(n1980), .ZN(n1075) );
  IND2D0BWP12T U85 ( .A1(memory_interface_inst1_delayed_is_signed), .B1(n2288), 
        .ZN(n10) );
  ND4D0BWP12T U86 ( .A1(n885), .A2(n2327), .A3(n886), .A4(n10), .ZN(n2267) );
  INR3D0BWP12T U87 ( .A1(n772), .B1(n2332), .B2(MEMCTRL_load_in), .ZN(n862) );
  IND3D1BWP12T U88 ( .A1(n69), .B1(n2293), .B2(n1089), .ZN(n1086) );
  IND3D1BWP12T U89 ( .A1(n123), .B1(n2293), .B2(n1098), .ZN(n1096) );
  IND3D1BWP12T U90 ( .A1(n73), .B1(n2293), .B2(n74), .ZN(n1068) );
  NR3D0BWP12T U91 ( .A1(memory_interface_inst1_fsm_state_0_), .A2(
        memory_interface_inst1_fsm_state_3_), .A3(n2250), .ZN(n2288) );
  INR2D0BWP12T U92 ( .A1(n2276), .B1(n1973), .ZN(n161) );
  IND2D0BWP12T U93 ( .A1(n145), .B1(n1970), .ZN(n1079) );
  IND2D0BWP12T U94 ( .A1(n148), .B1(n1971), .ZN(n1071) );
  MAOI22D0BWP12T U95 ( .A1(n2277), .A2(ALU_MISC_OUT_result[31]), .B1(n2277), 
        .B2(n1101), .ZN(n519) );
  IND2D0BWP12T U96 ( .A1(n886), .B1(n885), .ZN(n2269) );
  AN3D0BWP12T U97 ( .A1(memory_interface_inst1_fsm_state_2_), .A2(n2247), .A3(
        n617), .Z(n501) );
  IND2D0BWP12T U98 ( .A1(n2093), .B1(n76), .ZN(n1871) );
  XNR2XD0BWP12T U99 ( .A1(n1016), .A2(n1015), .ZN(
        register_file_inst1_pc_write_in_plus_two[22]) );
  CKND2D2BWP12T U100 ( .A1(n1014), .A2(n1015), .ZN(n1017) );
  CKND2D2BWP12T U101 ( .A1(n130), .A2(register_file_inst1_pc_write_in_11_), 
        .ZN(n109) );
  OR4D2BWP12T U102 ( .A1(n1489), .A2(n1488), .A3(n1487), .A4(n1486), .Z(
        RF_ALU_operand_b[6]) );
  MUX2D1BWP12T U103 ( .I0(n507), .I1(n506), .S(n514), .Z(n11) );
  MUX2D1BWP12T U104 ( .I0(n503), .I1(n502), .S(n514), .Z(n12) );
  ND2D1BWP12T U105 ( .A1(n49), .A2(n48), .ZN(RF_ALU_STACK_operand_a[14]) );
  MUX2D1BWP12T U106 ( .I0(n1030), .I1(n1031), .S(n514), .Z(n13) );
  MUX2D1BWP12T U107 ( .I0(n970), .I1(n971), .S(n514), .Z(n14) );
  OR4XD1BWP12T U108 ( .A1(n592), .A2(n591), .A3(n590), .A4(n589), .Z(
        RF_ALU_STACK_operand_a[26]) );
  OR4XD1BWP12T U109 ( .A1(n557), .A2(n556), .A3(n555), .A4(n554), .Z(
        RF_ALU_operand_b[21]) );
  OR4XD1BWP12T U110 ( .A1(n579), .A2(n578), .A3(n577), .A4(n576), .Z(
        RF_ALU_STACK_operand_a[24]) );
  OR4XD1BWP12T U111 ( .A1(n566), .A2(n565), .A3(n564), .A4(n563), .Z(
        RF_ALU_operand_b[22]) );
  OR4XD1BWP12T U112 ( .A1(n602), .A2(n601), .A3(n600), .A4(n599), .Z(
        RF_ALU_STACK_operand_a[22]) );
  MUX2ND0BWP12T U113 ( .I0(MEMCTRL_RF_IF_data_in[2]), .I1(
        ALU_MISC_OUT_result[2]), .S(n2277), .ZN(n15) );
  MUX2ND0BWP12T U114 ( .I0(MEMCTRL_RF_IF_data_in[4]), .I1(
        ALU_MISC_OUT_result[4]), .S(n2277), .ZN(n16) );
  OR4XD1BWP12T U115 ( .A1(n545), .A2(n544), .A3(n543), .A4(n542), .Z(
        RF_ALU_operand_b[20]) );
  MUX2ND0BWP12T U116 ( .I0(MEMCTRL_RF_IF_data_in[8]), .I1(
        ALU_MISC_OUT_result[8]), .S(n2277), .ZN(n17) );
  INVD1BWP12T U117 ( .I(register_file_inst1_pc_write_in_7_), .ZN(n18) );
  INVD1BWP12T U118 ( .I(register_file_inst1_pc_write_in_1_), .ZN(n226) );
  NR2XD1BWP12T U119 ( .A1(n15), .A2(n226), .ZN(n894) );
  TPND2D1BWP12T U120 ( .A1(register_file_inst1_pc_write_in_3_), .A2(n894), 
        .ZN(n210) );
  TPND2D1BWP12T U121 ( .A1(register_file_inst1_pc_write_in_5_), .A2(n917), 
        .ZN(n195) );
  TPNR2D1BWP12T U122 ( .A1(n1930), .A2(n195), .ZN(n59) );
  XNR2XD1BWP12T U123 ( .A1(n18), .A2(n59), .ZN(
        register_file_inst1_pc_write_in_plus_two[7]) );
  INVD1BWP12T U124 ( .I(register_file_inst1_r11_22_), .ZN(n593) );
  INVD1BWP12T U125 ( .I(n161), .ZN(n19) );
  OAI211D1BWP12T U126 ( .A1(n2279), .A2(n1974), .B(n2293), .C(n19), .ZN(n1021)
         );
  OR3D1BWP12T U127 ( .A1(n161), .A2(n1975), .A3(n2279), .Z(n1020) );
  INVD1BWP12T U128 ( .I(MEM_MEMCTRL_from_mem_data[14]), .ZN(n2328) );
  NR2D1BWP12T U129 ( .A1(memory_interface_inst1_fsm_state_1_), .A2(
        memory_interface_inst1_fsm_state_0_), .ZN(n617) );
  INVD1BWP12T U130 ( .I(memory_interface_inst1_fsm_state_3_), .ZN(n2247) );
  INVD1BWP12T U131 ( .I(n501), .ZN(n885) );
  INVD1BWP12T U132 ( .I(n498), .ZN(n2289) );
  INVD1BWP12T U133 ( .I(MEM_MEMCTRL_from_mem_data[15]), .ZN(n2327) );
  INR2D1BWP12T U134 ( .A1(memory_interface_inst1_fsm_state_1_), .B1(
        memory_interface_inst1_fsm_state_2_), .ZN(n858) );
  INVD1BWP12T U135 ( .I(n858), .ZN(n2250) );
  INVD1BWP12T U136 ( .I(memory_interface_inst1_fsm_state_0_), .ZN(n499) );
  INR2D1BWP12T U137 ( .A1(n499), .B1(n498), .ZN(n772) );
  ND2D1BWP12T U138 ( .A1(n2276), .A2(n1976), .ZN(n1019) );
  INVD3BWP12T U139 ( .I(ALU_MISC_OUT_result[22]), .ZN(n988) );
  OAI222D0BWP12T U140 ( .A1(n593), .A2(n1021), .B1(n1020), .B2(n989), .C1(
        n1019), .C2(n988), .ZN(register_file_inst1_n2287) );
  INVD1BWP12T U141 ( .I(register_file_inst1_r12_4_), .ZN(n1668) );
  ND2D1BWP12T U142 ( .A1(n2303), .A2(n2175), .ZN(n28) );
  NR2D1BWP12T U143 ( .A1(n28), .A2(n2178), .ZN(n1915) );
  INVD1BWP12T U144 ( .I(n1915), .ZN(n1798) );
  INVD1BWP12T U145 ( .I(STACK_RF_next_sp[4]), .ZN(n20) );
  NR2D1BWP12T U146 ( .A1(n2178), .A2(n2181), .ZN(n1914) );
  INVD1BWP12T U147 ( .I(n1914), .ZN(n1796) );
  OAI22D1BWP12T U148 ( .A1(n1668), .A2(n1798), .B1(n20), .B2(n1796), .ZN(n24)
         );
  NR2D1BWP12T U149 ( .A1(n2181), .A2(n2183), .ZN(n1937) );
  INVD1BWP12T U150 ( .I(n1937), .ZN(n1802) );
  INVD1BWP12T U151 ( .I(register_file_inst1_r0_4_), .ZN(n255) );
  ND2D1BWP12T U152 ( .A1(n2302), .A2(n2175), .ZN(n106) );
  NR2D1BWP12T U153 ( .A1(n106), .A2(n2176), .ZN(n1938) );
  INVD1BWP12T U154 ( .I(n1938), .ZN(n1800) );
  OAI22D1BWP12T U155 ( .A1(n2190), .A2(n1802), .B1(n255), .B2(n1800), .ZN(n23)
         );
  CKND1BWP12T U156 ( .I(register_file_inst1_lr_4_), .ZN(n1671) );
  NR2D1BWP12T U157 ( .A1(n28), .A2(n2183), .ZN(n1917) );
  INVD1BWP12T U158 ( .I(n1917), .ZN(n1805) );
  INVD1BWP12T U159 ( .I(register_file_inst1_r3_4_), .ZN(n1669) );
  NR2D1BWP12T U160 ( .A1(n2179), .A2(n2180), .ZN(n1916) );
  INVD1BWP12T U161 ( .I(n1916), .ZN(n1803) );
  OAI22D1BWP12T U162 ( .A1(n1671), .A2(n1805), .B1(n1669), .B2(n1803), .ZN(n22) );
  CKND1BWP12T U163 ( .I(register_file_inst1_r1_4_), .ZN(n254) );
  NR2D1BWP12T U164 ( .A1(n2176), .A2(n2180), .ZN(n1919) );
  INVD1BWP12T U165 ( .I(n1919), .ZN(n1809) );
  INVD1BWP12T U166 ( .I(register_file_inst1_r7_4_), .ZN(n250) );
  NR2D1BWP12T U167 ( .A1(n2183), .A2(n2180), .ZN(n1918) );
  INVD1BWP12T U168 ( .I(n1918), .ZN(n1807) );
  OAI22D1BWP12T U169 ( .A1(n254), .A2(n1809), .B1(n250), .B2(n1807), .ZN(n21)
         );
  NR4D0BWP12T U170 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n37) );
  CKND2D1BWP12T U171 ( .A1(register_file_inst1_r9_4_), .A2(n1911), .ZN(n26) );
  CKND2D1BWP12T U172 ( .A1(register_file_inst1_r8_4_), .A2(n1910), .ZN(n25) );
  ND3D1BWP12T U173 ( .A1(n2191), .A2(n26), .A3(n25), .ZN(n35) );
  INVD1BWP12T U174 ( .I(register_file_inst1_r4_4_), .ZN(n1670) );
  INVD1BWP12T U175 ( .I(n2178), .ZN(n30) );
  INVD1BWP12T U176 ( .I(n106), .ZN(n27) );
  CKND1BWP12T U177 ( .I(register_file_inst1_r10_4_), .ZN(n1672) );
  INVD1BWP12T U178 ( .I(n2179), .ZN(n31) );
  OAI22D1BWP12T U179 ( .A1(n1670), .A2(n1903), .B1(n1672), .B2(n1901), .ZN(n34) );
  INVD1BWP12T U180 ( .I(register_file_inst1_r5_4_), .ZN(n256) );
  INVD1BWP12T U181 ( .I(n2180), .ZN(n29) );
  ND2D2BWP12T U182 ( .A1(n30), .A2(n29), .ZN(n1907) );
  CKND1BWP12T U183 ( .I(register_file_inst1_r11_4_), .ZN(n249) );
  OAI22D1BWP12T U184 ( .A1(n256), .A2(n1907), .B1(n249), .B2(n1905), .ZN(n33)
         );
  INVD1BWP12T U185 ( .I(register_file_inst1_tmp1_4_), .ZN(n252) );
  INVD1BWP12T U186 ( .I(n2244), .ZN(n1823) );
  INVD1BWP12T U187 ( .I(register_file_inst1_r6_4_), .ZN(n1673) );
  NR2D1BWP12T U188 ( .A1(n2183), .A2(n106), .ZN(n1909) );
  INVD1BWP12T U189 ( .I(n1909), .ZN(n1821) );
  OAI22D1BWP12T U190 ( .A1(n252), .A2(n1823), .B1(n1673), .B2(n1821), .ZN(n32)
         );
  NR4D0BWP12T U191 ( .A1(n35), .A2(n34), .A3(n33), .A4(n32), .ZN(n36) );
  ND2D1BWP12T U192 ( .A1(n37), .A2(n36), .ZN(RF_ALU_STACK_operand_a[4]) );
  TPND2D0BWP12T U193 ( .A1(n501), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[5]), .ZN(n2272) );
  TPND2D0BWP12T U194 ( .A1(n501), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[4]), .ZN(n2273) );
  INVD1BWP12T U195 ( .I(register_file_inst1_r12_14_), .ZN(n232) );
  INVD1BWP12T U196 ( .I(STACK_RF_next_sp[14]), .ZN(n227) );
  OAI22D1BWP12T U197 ( .A1(n232), .A2(n1798), .B1(n227), .B2(n1796), .ZN(n41)
         );
  INVD1BWP12T U198 ( .I(register_file_inst1_r0_14_), .ZN(n234) );
  OAI22D1BWP12T U199 ( .A1(n2210), .A2(n1802), .B1(n234), .B2(n1800), .ZN(n40)
         );
  INVD1BWP12T U200 ( .I(register_file_inst1_lr_14_), .ZN(n231) );
  INVD1BWP12T U201 ( .I(register_file_inst1_r3_14_), .ZN(n221) );
  OAI22D1BWP12T U202 ( .A1(n231), .A2(n1805), .B1(n221), .B2(n1803), .ZN(n39)
         );
  INVD1BWP12T U203 ( .I(register_file_inst1_r1_14_), .ZN(n1254) );
  INVD1BWP12T U204 ( .I(register_file_inst1_r7_14_), .ZN(n1256) );
  OAI22D1BWP12T U205 ( .A1(n1254), .A2(n1809), .B1(n1256), .B2(n1807), .ZN(n38) );
  NR4D0BWP12T U206 ( .A1(n41), .A2(n40), .A3(n39), .A4(n38), .ZN(n49) );
  CKND2D1BWP12T U207 ( .A1(register_file_inst1_r9_14_), .A2(n1911), .ZN(n43)
         );
  CKND2D1BWP12T U208 ( .A1(register_file_inst1_r8_14_), .A2(n1910), .ZN(n42)
         );
  ND3D1BWP12T U209 ( .A1(n2211), .A2(n43), .A3(n42), .ZN(n47) );
  INVD1BWP12T U210 ( .I(register_file_inst1_r4_14_), .ZN(n230) );
  INVD1BWP12T U211 ( .I(register_file_inst1_r10_14_), .ZN(n220) );
  OAI22D1BWP12T U212 ( .A1(n230), .A2(n1903), .B1(n220), .B2(n1901), .ZN(n46)
         );
  INVD1BWP12T U213 ( .I(register_file_inst1_r5_14_), .ZN(n223) );
  INVD1BWP12T U214 ( .I(register_file_inst1_r11_14_), .ZN(n1253) );
  OAI22D1BWP12T U215 ( .A1(n223), .A2(n1907), .B1(n1253), .B2(n1905), .ZN(n45)
         );
  INVD1BWP12T U216 ( .I(register_file_inst1_tmp1_14_), .ZN(n228) );
  INVD1BWP12T U217 ( .I(register_file_inst1_r6_14_), .ZN(n225) );
  OAI22D1BWP12T U218 ( .A1(n228), .A2(n1823), .B1(n225), .B2(n1821), .ZN(n44)
         );
  NR4D0BWP12T U219 ( .A1(n47), .A2(n46), .A3(n45), .A4(n44), .ZN(n48) );
  INVD1BWP12T U220 ( .I(register_file_inst1_r4_30_), .ZN(n1048) );
  INVD1BWP12T U221 ( .I(register_file_inst1_r10_30_), .ZN(n1041) );
  OAI22D1BWP12T U222 ( .A1(n1048), .A2(n1903), .B1(n1041), .B2(n1901), .ZN(n58) );
  INVD1BWP12T U223 ( .I(register_file_inst1_r5_30_), .ZN(n1042) );
  INVD1BWP12T U224 ( .I(register_file_inst1_r11_30_), .ZN(n1617) );
  OAI22D1BWP12T U225 ( .A1(n1042), .A2(n1907), .B1(n1617), .B2(n1905), .ZN(n57) );
  AOI22D1BWP12T U226 ( .A1(register_file_inst1_tmp1_30_), .A2(n2244), .B1(
        register_file_inst1_r6_30_), .B2(n1909), .ZN(n51) );
  AOI22D1BWP12T U227 ( .A1(register_file_inst1_r9_30_), .A2(n1911), .B1(
        register_file_inst1_r8_30_), .B2(n1910), .ZN(n50) );
  ND3D1BWP12T U228 ( .A1(n51), .A2(n50), .A3(n2242), .ZN(n56) );
  AOI22D1BWP12T U229 ( .A1(register_file_inst1_r12_30_), .A2(n1915), .B1(
        STACK_RF_next_sp[30]), .B2(n1914), .ZN(n54) );
  AOI22D1BWP12T U230 ( .A1(register_file_inst1_lr_30_), .A2(n1917), .B1(
        register_file_inst1_r3_30_), .B2(n1916), .ZN(n53) );
  AOI22D0BWP12T U231 ( .A1(register_file_inst1_r1_30_), .A2(n1919), .B1(
        register_file_inst1_r7_30_), .B2(n1918), .ZN(n52) );
  ND4D1BWP12T U232 ( .A1(n54), .A2(n2243), .A3(n53), .A4(n52), .ZN(n55) );
  OR4D1BWP12T U233 ( .A1(n58), .A2(n57), .A3(n56), .A4(n55), .Z(
        RF_ALU_STACK_operand_a[30]) );
  ND2D1BWP12T U234 ( .A1(n2316), .A2(n2315), .ZN(n289) );
  OR2D1BWP12T U235 ( .A1(n2311), .A2(n2308), .Z(n745) );
  INVD1BWP12T U236 ( .I(n745), .ZN(n1927) );
  TPND2D0BWP12T U237 ( .A1(n2293), .A2(n1960), .ZN(n1962) );
  INVD1BWP12T U238 ( .I(MEM_MEMCTRL_from_mem_data[3]), .ZN(n2261) );
  INVD1BWP12T U239 ( .I(MEM_MEMCTRL_from_mem_data[4]), .ZN(n2259) );
  INVD1BWP12T U240 ( .I(MEM_MEMCTRL_from_mem_data[5]), .ZN(n2257) );
  INVD1BWP12T U241 ( .I(MEM_MEMCTRL_from_mem_data[0]), .ZN(n2268) );
  INVD1BWP12T U242 ( .I(MEM_MEMCTRL_from_mem_data[7]), .ZN(n2253) );
  INVD1BWP12T U243 ( .I(MEM_MEMCTRL_from_mem_data[1]), .ZN(n2265) );
  INVD1BWP12T U244 ( .I(MEM_MEMCTRL_from_mem_data[6]), .ZN(n2255) );
  INVD1BWP12T U245 ( .I(MEM_MEMCTRL_from_mem_data[2]), .ZN(n2263) );
  INVD1BWP12T U246 ( .I(register_file_inst1_pc_write_in_13_), .ZN(n62) );
  TPNR2D1BWP12T U247 ( .A1(n1931), .A2(n17), .ZN(n60) );
  TPND2D1BWP12T U248 ( .A1(register_file_inst1_pc_write_in_7_), .A2(n59), .ZN(
        n972) );
  INVD1P75BWP12T U249 ( .I(n972), .ZN(n974) );
  TPND2D2BWP12T U250 ( .A1(n60), .A2(n974), .ZN(n155) );
  NR2XD1BWP12T U251 ( .A1(n155), .A2(n1929), .ZN(n130) );
  INVD1BWP12T U252 ( .I(n109), .ZN(n993) );
  CKND2D1BWP12T U253 ( .A1(register_file_inst1_pc_write_in_12_), .A2(n993), 
        .ZN(n61) );
  CKXOR2D1BWP12T U254 ( .A1(n62), .A2(n61), .Z(
        register_file_inst1_pc_write_in_plus_two[13]) );
  CKND0BWP12T U255 ( .I(register_file_inst1_r6_20_), .ZN(n65) );
  ND2D1BWP12T U256 ( .A1(n1968), .A2(n2083), .ZN(n1043) );
  NR2D1BWP12T U257 ( .A1(n2278), .A2(n1969), .ZN(n64) );
  INVD0BWP12T U258 ( .I(n64), .ZN(n63) );
  ND3D1BWP12T U259 ( .A1(n2293), .A2(n1043), .A3(n63), .ZN(n1045) );
  ND3D1BWP12T U260 ( .A1(n64), .A2(n2293), .A3(n1043), .ZN(n1044) );
  INVD1BWP12T U261 ( .I(MEM_MEMCTRL_from_mem_data[12]), .ZN(n2330) );
  IAO21D1BWP12T U262 ( .A1(n2330), .A2(n885), .B(n500), .ZN(n515) );
  OAI222D0BWP12T U263 ( .A1(n65), .A2(n1045), .B1(n1044), .B2(n515), .C1(n1043), .C2(n516), .ZN(register_file_inst1_n2445) );
  CKND0BWP12T U264 ( .I(register_file_inst1_lr_20_), .ZN(n68) );
  ND2D1BWP12T U265 ( .A1(n2083), .A2(n1981), .ZN(n1085) );
  ND2D1BWP12T U266 ( .A1(n2300), .A2(n2298), .ZN(n147) );
  NR2D1BWP12T U267 ( .A1(n2278), .A2(n147), .ZN(n67) );
  INVD0BWP12T U268 ( .I(n67), .ZN(n66) );
  ND3D1BWP12T U269 ( .A1(n2293), .A2(n1085), .A3(n66), .ZN(n1082) );
  ND3D1BWP12T U270 ( .A1(n67), .A2(n2293), .A3(n1085), .ZN(n1084) );
  OAI222D0BWP12T U271 ( .A1(n68), .A2(n1082), .B1(n1084), .B2(n515), .C1(n1085), .C2(n516), .ZN(register_file_inst1_n2221) );
  CKND0BWP12T U272 ( .I(register_file_inst1_r0_20_), .ZN(n70) );
  ND2D1BWP12T U273 ( .A1(n1979), .A2(n1968), .ZN(n1089) );
  ND2D1BWP12T U274 ( .A1(n1972), .A2(n1963), .ZN(n144) );
  NR2D1BWP12T U275 ( .A1(n144), .A2(n1969), .ZN(n69) );
  ND3D1BWP12T U276 ( .A1(n69), .A2(n2293), .A3(n1089), .ZN(n1088) );
  OAI222D0BWP12T U277 ( .A1(n70), .A2(n1086), .B1(n1088), .B2(n515), .C1(n1089), .C2(n516), .ZN(register_file_inst1_n2637) );
  CKND0BWP12T U278 ( .I(STACK_RF_next_sp[20]), .ZN(n72) );
  NR2D1BWP12T U279 ( .A1(n2279), .A2(n1977), .ZN(n71) );
  INVD1BWP12T U280 ( .I(n71), .ZN(n215) );
  ND2D1BWP12T U281 ( .A1(n1978), .A2(n215), .ZN(n1037) );
  ND2D1BWP12T U282 ( .A1(n1978), .A2(n71), .ZN(n1102) );
  NR2D1BWP12T U283 ( .A1(n1964), .A2(n1962), .ZN(n149) );
  ND2D1BWP12T U284 ( .A1(n2276), .A2(n149), .ZN(n1104) );
  OAI222D0BWP12T U285 ( .A1(n72), .A2(n1037), .B1(n1102), .B2(n515), .C1(n1104), .C2(n516), .ZN(register_file_inst1_spin[20]) );
  NR2D1BWP12T U286 ( .A1(n147), .A2(n1975), .ZN(n73) );
  INVD1BWP12T U287 ( .I(n1973), .ZN(n139) );
  CKND2D1BWP12T U288 ( .A1(n1981), .A2(n139), .ZN(n74) );
  ND2D1BWP12T U289 ( .A1(n73), .A2(n74), .ZN(n1069) );
  INVD1BWP12T U290 ( .I(ALU_MISC_OUT_result[4]), .ZN(n257) );
  ND2D1BWP12T U291 ( .A1(n1981), .A2(n1976), .ZN(n1070) );
  OAI222D0BWP12T U292 ( .A1(n2105), .A2(n1069), .B1(n257), .B2(n1070), .C1(
        n1068), .C2(n1672), .ZN(register_file_inst1_n2301) );
  INVD1BWP12T U293 ( .I(MEM_MEMCTRL_from_mem_data[13]), .ZN(n2329) );
  INVD1BWP12T U294 ( .I(register_file_inst1_r1_19_), .ZN(n1532) );
  INVD1BWP12T U295 ( .I(n2097), .ZN(n77) );
  INVD1BWP12T U296 ( .I(n2092), .ZN(n75) );
  ND2D1BWP12T U297 ( .A1(n77), .A2(n75), .ZN(n1873) );
  INVD1BWP12T U298 ( .I(register_file_inst1_r11_19_), .ZN(n1541) );
  INVD1BWP12T U299 ( .I(n2094), .ZN(n76) );
  OAI22D1BWP12T U300 ( .A1(n1532), .A2(n1873), .B1(n1541), .B2(n1871), .ZN(n86) );
  INVD1BWP12T U301 ( .I(register_file_inst1_r7_19_), .ZN(n1531) );
  CKND1BWP12T U302 ( .I(n2088), .ZN(n2095) );
  ND2D1BWP12T U303 ( .A1(n75), .A2(n2095), .ZN(n1877) );
  INVD1BWP12T U304 ( .I(register_file_inst1_r9_19_), .ZN(n969) );
  ND2D1BWP12T U305 ( .A1(n77), .A2(n76), .ZN(n1875) );
  OAI22D1BWP12T U306 ( .A1(n1531), .A2(n1877), .B1(n969), .B2(n1875), .ZN(n85)
         );
  ND2D1BWP12T U307 ( .A1(n2304), .A2(n2089), .ZN(n107) );
  NR2D1BWP12T U308 ( .A1(n2097), .A2(n107), .ZN(n1633) );
  AOI22D1BWP12T U309 ( .A1(register_file_inst1_tmp1_19_), .A2(n1835), .B1(
        register_file_inst1_r0_19_), .B2(n1633), .ZN(n79) );
  AOI22D1BWP12T U310 ( .A1(register_file_inst1_r5_19_), .A2(n1868), .B1(
        STACK_RF_next_sp[19]), .B2(n1867), .ZN(n78) );
  ND3D1BWP12T U311 ( .A1(n79), .A2(n78), .A3(n2144), .ZN(n84) );
  ND2D1BWP12T U312 ( .A1(n2305), .A2(n2089), .ZN(n105) );
  NR2D1BWP12T U313 ( .A1(n105), .A2(n2090), .ZN(n1659) );
  NR2D1BWP12T U314 ( .A1(n2097), .A2(n105), .ZN(n1838) );
  AOI22D1BWP12T U315 ( .A1(register_file_inst1_r12_19_), .A2(n1659), .B1(
        register_file_inst1_r8_19_), .B2(n1838), .ZN(n82) );
  NR2D1BWP12T U316 ( .A1(n2090), .A2(n107), .ZN(n1595) );
  NR2D1BWP12T U317 ( .A1(n2093), .A2(n2092), .ZN(n1839) );
  AOI22D1BWP12T U318 ( .A1(register_file_inst1_r4_19_), .A2(n1595), .B1(
        register_file_inst1_r3_19_), .B2(n1839), .ZN(n81) );
  NR2D1BWP12T U319 ( .A1(n107), .A2(n2088), .ZN(n1596) );
  NR2D1BWP12T U320 ( .A1(n105), .A2(n2093), .ZN(n1840) );
  AOI22D1BWP12T U321 ( .A1(register_file_inst1_r6_19_), .A2(n1596), .B1(
        register_file_inst1_r10_19_), .B2(n1840), .ZN(n80) );
  ND4D1BWP12T U322 ( .A1(n82), .A2(n81), .A3(n2145), .A4(n80), .ZN(n83) );
  OR4D1BWP12T U323 ( .A1(n86), .A2(n85), .A3(n84), .A4(n83), .Z(
        RF_ALU_operand_b[19]) );
  INVD1BWP12T U324 ( .I(register_file_inst1_r1_23_), .ZN(n193) );
  INVD1BWP12T U325 ( .I(register_file_inst1_r11_23_), .ZN(n1890) );
  OAI22D1BWP12T U326 ( .A1(n193), .A2(n1873), .B1(n1890), .B2(n1871), .ZN(n95)
         );
  INVD1BWP12T U327 ( .I(register_file_inst1_r7_23_), .ZN(n190) );
  INVD1BWP12T U328 ( .I(register_file_inst1_r9_23_), .ZN(n183) );
  OAI22D1BWP12T U329 ( .A1(n190), .A2(n1877), .B1(n183), .B2(n1875), .ZN(n94)
         );
  AOI22D1BWP12T U330 ( .A1(register_file_inst1_tmp1_23_), .A2(n1835), .B1(
        register_file_inst1_r0_23_), .B2(n1633), .ZN(n88) );
  AOI22D1BWP12T U331 ( .A1(register_file_inst1_r5_23_), .A2(n1868), .B1(
        STACK_RF_next_sp[23]), .B2(n1867), .ZN(n87) );
  ND3D1BWP12T U332 ( .A1(n88), .A2(n87), .A3(n2152), .ZN(n93) );
  AOI22D1BWP12T U333 ( .A1(register_file_inst1_r12_23_), .A2(n1659), .B1(
        register_file_inst1_r8_23_), .B2(n1838), .ZN(n91) );
  AOI22D1BWP12T U334 ( .A1(register_file_inst1_r4_23_), .A2(n1595), .B1(
        register_file_inst1_r3_23_), .B2(n1839), .ZN(n90) );
  AOI22D1BWP12T U335 ( .A1(register_file_inst1_r6_23_), .A2(n1596), .B1(
        register_file_inst1_r10_23_), .B2(n1840), .ZN(n89) );
  ND4D1BWP12T U336 ( .A1(n91), .A2(n90), .A3(n2153), .A4(n89), .ZN(n92) );
  OR4D1BWP12T U337 ( .A1(n95), .A2(n94), .A3(n93), .A4(n92), .Z(
        RF_ALU_operand_b[23]) );
  INR2XD0BWP12T U338 ( .A1(memory_interface_inst1_fsm_state_0_), .B1(n2247), 
        .ZN(n614) );
  CKND2D0BWP12T U339 ( .A1(n858), .A2(n614), .ZN(n621) );
  INVD1BWP12T U340 ( .I(n621), .ZN(n618) );
  AOI211D1BWP12T U341 ( .A1(n862), .A2(n1953), .B(n1951), .C(n618), .ZN(n1952)
         );
  INVD1BWP12T U342 ( .I(register_file_inst1_r1_24_), .ZN(n171) );
  INVD1BWP12T U343 ( .I(register_file_inst1_r11_24_), .ZN(n569) );
  INVD1BWP12T U344 ( .I(n1871), .ZN(n1741) );
  OAI22D1BWP12T U345 ( .A1(n171), .A2(n1873), .B1(n569), .B2(n1871), .ZN(n104)
         );
  INVD1BWP12T U346 ( .I(register_file_inst1_r7_24_), .ZN(n175) );
  INVD1BWP12T U347 ( .I(register_file_inst1_r9_24_), .ZN(n174) );
  INVD1BWP12T U348 ( .I(n1875), .ZN(n1743) );
  OAI22D1BWP12T U349 ( .A1(n175), .A2(n1877), .B1(n174), .B2(n1875), .ZN(n103)
         );
  AOI22D1BWP12T U350 ( .A1(register_file_inst1_tmp1_24_), .A2(n1835), .B1(
        register_file_inst1_r0_24_), .B2(n1633), .ZN(n97) );
  AOI22D1BWP12T U351 ( .A1(register_file_inst1_r5_24_), .A2(n1868), .B1(
        STACK_RF_next_sp[24]), .B2(n1867), .ZN(n96) );
  ND3D1BWP12T U352 ( .A1(n97), .A2(n96), .A3(n2154), .ZN(n102) );
  INVD1BWP12T U353 ( .I(n1659), .ZN(n1850) );
  AOI22D1BWP12T U354 ( .A1(register_file_inst1_r12_24_), .A2(n1659), .B1(
        register_file_inst1_r8_24_), .B2(n1838), .ZN(n100) );
  INVD1BWP12T U355 ( .I(n1595), .ZN(n1854) );
  AOI22D1BWP12T U356 ( .A1(register_file_inst1_r4_24_), .A2(n1595), .B1(
        register_file_inst1_r3_24_), .B2(n1839), .ZN(n99) );
  INVD1BWP12T U357 ( .I(n1596), .ZN(n1861) );
  AOI22D1BWP12T U358 ( .A1(register_file_inst1_r6_24_), .A2(n1596), .B1(
        register_file_inst1_r10_24_), .B2(n1840), .ZN(n98) );
  ND4D1BWP12T U359 ( .A1(n100), .A2(n99), .A3(n2155), .A4(n98), .ZN(n101) );
  OR4D1BWP12T U360 ( .A1(n104), .A2(n103), .A3(n102), .A4(n101), .Z(
        RF_ALU_operand_b[24]) );
  CKND2D0BWP12T U361 ( .A1(n501), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[15]), .ZN(n2252) );
  CKND2D0BWP12T U362 ( .A1(n501), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[0]), .ZN(n2274) );
  NR2D1BWP12T U363 ( .A1(n105), .A2(n2088), .ZN(n1943) );
  INVD4BWP12T U364 ( .I(ALU_MISC_OUT_result[19]), .ZN(n970) );
  AOI21D1BWP12T U365 ( .A1(n501), .A2(MEM_MEMCTRL_from_mem_data[11]), .B(n500), 
        .ZN(n971) );
  ND2D1BWP12T U366 ( .A1(n2276), .A2(n2275), .ZN(n514) );
  AOI21D1BWP12T U367 ( .A1(n501), .A2(MEM_MEMCTRL_from_mem_data[10]), .B(n500), 
        .ZN(n219) );
  MUX2ND4BWP12T U368 ( .I0(n218), .I1(n219), .S(n514), .ZN(n995) );
  INVD1BWP12T U369 ( .I(n514), .ZN(n2277) );
  AOI21D1BWP12T U370 ( .A1(n501), .A2(MEM_MEMCTRL_from_mem_data[9]), .B(n500), 
        .ZN(n217) );
  CKND2D1BWP12T U371 ( .A1(ALU_MISC_OUT_result[17]), .A2(n2277), .ZN(n108) );
  OA21D1BWP12T U372 ( .A1(n2277), .A2(n217), .B(n108), .Z(n112) );
  INVD3BWP12T U373 ( .I(ALU_MISC_OUT_result[16]), .ZN(n966) );
  INVD1BWP12T U374 ( .I(MEM_MEMCTRL_from_mem_data[8]), .ZN(n2331) );
  MUX2NXD0BWP12T U375 ( .I0(n966), .I1(n967), .S(n514), .ZN(n113) );
  INVD1BWP12T U376 ( .I(register_file_inst1_pc_write_in_15_), .ZN(n117) );
  TPND2D1BWP12T U377 ( .A1(register_file_inst1_pc_write_in_13_), .A2(
        register_file_inst1_pc_write_in_12_), .ZN(n110) );
  NR2XD1BWP12T U378 ( .A1(n110), .A2(n109), .ZN(n991) );
  TPND2D1BWP12T U379 ( .A1(n991), .A2(register_file_inst1_pc_write_in_14_), 
        .ZN(n116) );
  NR2XD1BWP12T U380 ( .A1(n117), .A2(n116), .ZN(n114) );
  TPND2D1BWP12T U381 ( .A1(n113), .A2(n114), .ZN(n111) );
  NR2XD1BWP12T U382 ( .A1(n112), .A2(n111), .ZN(n996) );
  TPND2D1BWP12T U383 ( .A1(n995), .A2(n996), .ZN(n517) );
  XOR2XD1BWP12T U384 ( .A1(n14), .A2(n517), .Z(
        register_file_inst1_pc_write_in_plus_two[19]) );
  XOR2XD1BWP12T U385 ( .A1(n112), .A2(n111), .Z(
        register_file_inst1_pc_write_in_plus_two[17]) );
  INVD1BWP12T U386 ( .I(n113), .ZN(n115) );
  XNR2XD1BWP12T U387 ( .A1(n115), .A2(n114), .ZN(
        register_file_inst1_pc_write_in_plus_two[16]) );
  XOR2XD1BWP12T U388 ( .A1(n117), .A2(n116), .Z(
        register_file_inst1_pc_write_in_plus_two[15]) );
  INVD1BWP12T U389 ( .I(register_file_inst1_r4_27_), .ZN(n1565) );
  ND2D1BWP12T U390 ( .A1(n149), .A2(n1968), .ZN(n1092) );
  NR2D1BWP12T U391 ( .A1(n1977), .A2(n1969), .ZN(n118) );
  ND3D1BWP12T U392 ( .A1(n118), .A2(n2293), .A3(n1092), .ZN(n1091) );
  AOI21D1BWP12T U393 ( .A1(n501), .A2(MEM_MEMCTRL_from_mem_data[3]), .B(n500), 
        .ZN(n502) );
  OAI222D0BWP12T U394 ( .A1(n1565), .A2(n1090), .B1(n1091), .B2(n502), .C1(
        n1092), .C2(n503), .ZN(register_file_inst1_n2516) );
  CKND0BWP12T U395 ( .I(STACK_RF_next_sp[27]), .ZN(n119) );
  ND2D1BWP12T U396 ( .A1(n1978), .A2(n215), .ZN(n1099) );
  OAI222D0BWP12T U397 ( .A1(n119), .A2(n1099), .B1(n1102), .B2(n502), .C1(
        n1104), .C2(n503), .ZN(register_file_inst1_spin[27]) );
  CKND0BWP12T U398 ( .I(register_file_inst1_tmp1_27_), .ZN(n122) );
  INR3D0BWP12T U399 ( .A1(n2300), .B1(n2278), .B2(n2298), .ZN(n121) );
  CKND0BWP12T U400 ( .I(n121), .ZN(n120) );
  ND3D1BWP12T U401 ( .A1(n2293), .A2(n2168), .A3(n120), .ZN(n1027) );
  ND3D1BWP12T U402 ( .A1(n121), .A2(n2293), .A3(n2168), .ZN(n1026) );
  OAI222D0BWP12T U403 ( .A1(n122), .A2(n1027), .B1(n1026), .B2(n502), .C1(
        n2168), .C2(n503), .ZN(register_file_inst1_n2164) );
  INVD1BWP12T U404 ( .I(register_file_inst1_r5_27_), .ZN(n1567) );
  NR2D1BWP12T U405 ( .A1(n2082), .A2(n1965), .ZN(n134) );
  ND2D1BWP12T U406 ( .A1(n134), .A2(n149), .ZN(n1098) );
  ND2D1BWP12T U407 ( .A1(n2301), .A2(n2299), .ZN(n135) );
  NR2D1BWP12T U408 ( .A1(n135), .A2(n1977), .ZN(n123) );
  ND3D1BWP12T U409 ( .A1(n123), .A2(n2293), .A3(n1098), .ZN(n1097) );
  OAI222D0BWP12T U410 ( .A1(n1567), .A2(n1096), .B1(n1097), .B2(n502), .C1(
        n1098), .C2(n503), .ZN(register_file_inst1_n2484) );
  CKND0BWP12T U411 ( .I(register_file_inst1_r6_27_), .ZN(n124) );
  OAI222D0BWP12T U412 ( .A1(n124), .A2(n1045), .B1(n1044), .B2(n502), .C1(
        n1043), .C2(n503), .ZN(register_file_inst1_n2452) );
  CKND0BWP12T U413 ( .I(register_file_inst1_r3_27_), .ZN(n128) );
  TPND2D0BWP12T U414 ( .A1(n134), .A2(n139), .ZN(n126) );
  NR2D1BWP12T U415 ( .A1(n135), .A2(n1975), .ZN(n127) );
  CKND0BWP12T U416 ( .I(n127), .ZN(n125) );
  ND3D1BWP12T U417 ( .A1(n2293), .A2(n126), .A3(n125), .ZN(n1064) );
  ND2D1BWP12T U418 ( .A1(n127), .A2(n126), .ZN(n1066) );
  ND2D1BWP12T U419 ( .A1(n134), .A2(n1976), .ZN(n1067) );
  OAI222D0BWP12T U420 ( .A1(n128), .A2(n1064), .B1(n1066), .B2(n502), .C1(
        n1067), .C2(n503), .ZN(register_file_inst1_n2548) );
  CKND0BWP12T U421 ( .I(register_file_inst1_r0_27_), .ZN(n129) );
  OAI222D0BWP12T U422 ( .A1(n129), .A2(n1086), .B1(n1088), .B2(n502), .C1(
        n1089), .C2(n503), .ZN(register_file_inst1_n2644) );
  INVD1BWP12T U423 ( .I(register_file_inst1_pc_write_in_11_), .ZN(n131) );
  XNR2XD1BWP12T U424 ( .A1(n131), .A2(n130), .ZN(
        register_file_inst1_pc_write_in_plus_two[11]) );
  INVD1BWP12T U425 ( .I(register_file_inst1_r7_27_), .ZN(n488) );
  ND2D1BWP12T U426 ( .A1(n134), .A2(n2083), .ZN(n1049) );
  NR2D1BWP12T U427 ( .A1(n2278), .A2(n135), .ZN(n133) );
  INVD0BWP12T U428 ( .I(n133), .ZN(n132) );
  ND3D1BWP12T U429 ( .A1(n2293), .A2(n1049), .A3(n132), .ZN(n1051) );
  ND3D1BWP12T U430 ( .A1(n133), .A2(n2293), .A3(n1049), .ZN(n1050) );
  OAI222D0BWP12T U431 ( .A1(n488), .A2(n1051), .B1(n1050), .B2(n502), .C1(
        n1049), .C2(n503), .ZN(register_file_inst1_n2420) );
  INVD1BWP12T U432 ( .I(register_file_inst1_r1_27_), .ZN(n486) );
  ND2D1BWP12T U433 ( .A1(n134), .A2(n1979), .ZN(n1095) );
  NR2D1BWP12T U434 ( .A1(n135), .A2(n144), .ZN(n136) );
  ND3D1BWP12T U435 ( .A1(n136), .A2(n2293), .A3(n1095), .ZN(n1094) );
  OAI222D0BWP12T U436 ( .A1(n486), .A2(n1093), .B1(n1094), .B2(n502), .C1(
        n1095), .C2(n503), .ZN(register_file_inst1_n2612) );
  INVD1BWP12T U437 ( .I(register_file_inst1_r10_27_), .ZN(n1564) );
  OAI222D0BWP12T U438 ( .A1(n1564), .A2(n1068), .B1(n1069), .B2(n502), .C1(
        n1070), .C2(n503), .ZN(register_file_inst1_n2324) );
  INVD1BWP12T U439 ( .I(register_file_inst1_r11_27_), .ZN(n1566) );
  OAI222D0BWP12T U440 ( .A1(n1566), .A2(n1021), .B1(n1020), .B2(n502), .C1(
        n1019), .C2(n503), .ZN(register_file_inst1_n2292) );
  CKND0BWP12T U441 ( .I(register_file_inst1_r8_27_), .ZN(n138) );
  NR2D1BWP12T U442 ( .A1(n144), .A2(n147), .ZN(n137) );
  ND2D1BWP12T U443 ( .A1(n1980), .A2(n137), .ZN(n1077) );
  ND2D1BWP12T U444 ( .A1(n1979), .A2(n1981), .ZN(n1078) );
  OAI222D0BWP12T U445 ( .A1(n138), .A2(n1075), .B1(n1077), .B2(n502), .C1(
        n1078), .C2(n503), .ZN(register_file_inst1_n2388) );
  CKND0BWP12T U446 ( .I(register_file_inst1_r2_27_), .ZN(n143) );
  CKND2D1BWP12T U447 ( .A1(n1968), .A2(n139), .ZN(n141) );
  NR2D1BWP12T U448 ( .A1(n1969), .A2(n1975), .ZN(n142) );
  CKND0BWP12T U449 ( .I(n142), .ZN(n140) );
  ND3D1BWP12T U450 ( .A1(n2293), .A2(n141), .A3(n140), .ZN(n1060) );
  ND2D1BWP12T U451 ( .A1(n142), .A2(n141), .ZN(n1062) );
  ND2D1BWP12T U452 ( .A1(n1968), .A2(n1976), .ZN(n1063) );
  OAI222D0BWP12T U453 ( .A1(n143), .A2(n1060), .B1(n1062), .B2(n502), .C1(
        n1063), .C2(n503), .ZN(register_file_inst1_n2580) );
  INVD1BWP12T U454 ( .I(register_file_inst1_r9_27_), .ZN(n487) );
  NR2D1BWP12T U455 ( .A1(n2279), .A2(n144), .ZN(n145) );
  ND2D1BWP12T U456 ( .A1(n1970), .A2(n145), .ZN(n1080) );
  ND2D1BWP12T U457 ( .A1(n2276), .A2(n1979), .ZN(n1081) );
  OAI222D0BWP12T U458 ( .A1(n487), .A2(n1079), .B1(n1080), .B2(n502), .C1(
        n1081), .C2(n503), .ZN(register_file_inst1_n2356) );
  CKND0BWP12T U459 ( .I(register_file_inst1_lr_27_), .ZN(n146) );
  OAI222D0BWP12T U460 ( .A1(n146), .A2(n1082), .B1(n1084), .B2(n502), .C1(
        n1085), .C2(n503), .ZN(register_file_inst1_n2228) );
  CKND0BWP12T U461 ( .I(register_file_inst1_r12_27_), .ZN(n150) );
  NR2D1BWP12T U462 ( .A1(n1977), .A2(n147), .ZN(n148) );
  ND2D1BWP12T U463 ( .A1(n1971), .A2(n148), .ZN(n1073) );
  ND2D1BWP12T U464 ( .A1(n149), .A2(n1981), .ZN(n1074) );
  OAI222D0BWP12T U465 ( .A1(n150), .A2(n1071), .B1(n1073), .B2(n502), .C1(
        n1074), .C2(n503), .ZN(register_file_inst1_n2260) );
  INVD1BWP12T U466 ( .I(register_file_inst1_r9_26_), .ZN(n466) );
  AOI21D1BWP12T U467 ( .A1(n501), .A2(MEM_MEMCTRL_from_mem_data[2]), .B(n500), 
        .ZN(n504) );
  OAI222D0BWP12T U468 ( .A1(n466), .A2(n1079), .B1(n1080), .B2(n504), .C1(
        n1081), .C2(n505), .ZN(register_file_inst1_n2355) );
  CKND0BWP12T U469 ( .I(register_file_inst1_r12_26_), .ZN(n151) );
  OAI222D0BWP12T U470 ( .A1(n151), .A2(n1071), .B1(n1073), .B2(n504), .C1(
        n1074), .C2(n505), .ZN(register_file_inst1_n2259) );
  INVD1BWP12T U471 ( .I(register_file_inst1_r5_26_), .ZN(n583) );
  OAI222D0BWP12T U472 ( .A1(n583), .A2(n1096), .B1(n1097), .B2(n504), .C1(
        n1098), .C2(n505), .ZN(register_file_inst1_n2483) );
  CKND0BWP12T U473 ( .I(STACK_RF_next_sp[26]), .ZN(n152) );
  OAI222D0BWP12T U474 ( .A1(n152), .A2(n1037), .B1(n1102), .B2(n504), .C1(
        n1104), .C2(n505), .ZN(register_file_inst1_spin[26]) );
  INVD1BWP12T U475 ( .I(register_file_inst1_r7_26_), .ZN(n467) );
  OAI222D0BWP12T U476 ( .A1(n467), .A2(n1051), .B1(n1050), .B2(n504), .C1(
        n1049), .C2(n505), .ZN(register_file_inst1_n2419) );
  INVD1BWP12T U477 ( .I(register_file_inst1_r10_26_), .ZN(n580) );
  OAI222D0BWP12T U478 ( .A1(n580), .A2(n1068), .B1(n1069), .B2(n504), .C1(
        n1070), .C2(n505), .ZN(register_file_inst1_n2323) );
  CKND0BWP12T U479 ( .I(register_file_inst1_r6_26_), .ZN(n153) );
  OAI222D0BWP12T U480 ( .A1(n153), .A2(n1045), .B1(n1044), .B2(n504), .C1(
        n1043), .C2(n505), .ZN(register_file_inst1_n2451) );
  CKND0BWP12T U481 ( .I(register_file_inst1_r0_26_), .ZN(n154) );
  OAI222D0BWP12T U482 ( .A1(n154), .A2(n1086), .B1(n1088), .B2(n504), .C1(
        n1089), .C2(n505), .ZN(register_file_inst1_n2643) );
  XOR2XD1BWP12T U483 ( .A1(n155), .A2(n1929), .Z(
        register_file_inst1_pc_write_in_plus_two[10]) );
  CKND0BWP12T U484 ( .I(register_file_inst1_r2_26_), .ZN(n156) );
  OAI222D0BWP12T U485 ( .A1(n156), .A2(n1060), .B1(n1062), .B2(n504), .C1(
        n1063), .C2(n505), .ZN(register_file_inst1_n2579) );
  CKND0BWP12T U486 ( .I(register_file_inst1_lr_26_), .ZN(n157) );
  OAI222D0BWP12T U487 ( .A1(n157), .A2(n1082), .B1(n1084), .B2(n504), .C1(
        n1085), .C2(n505), .ZN(register_file_inst1_n2227) );
  CKND0BWP12T U488 ( .I(register_file_inst1_tmp1_26_), .ZN(n158) );
  OAI222D0BWP12T U489 ( .A1(n158), .A2(n1027), .B1(n1026), .B2(n504), .C1(
        n2168), .C2(n505), .ZN(register_file_inst1_n2163) );
  INVD1BWP12T U490 ( .I(register_file_inst1_r4_26_), .ZN(n581) );
  OAI222D0BWP12T U491 ( .A1(n581), .A2(n1090), .B1(n1091), .B2(n504), .C1(
        n1092), .C2(n505), .ZN(register_file_inst1_n2515) );
  INVD1BWP12T U492 ( .I(register_file_inst1_r1_26_), .ZN(n465) );
  OAI222D0BWP12T U493 ( .A1(n465), .A2(n1093), .B1(n1094), .B2(n504), .C1(
        n1095), .C2(n505), .ZN(register_file_inst1_n2611) );
  CKND0BWP12T U494 ( .I(register_file_inst1_r8_26_), .ZN(n159) );
  OAI222D0BWP12T U495 ( .A1(n159), .A2(n1075), .B1(n1077), .B2(n504), .C1(
        n1078), .C2(n505), .ZN(register_file_inst1_n2387) );
  CKND0BWP12T U496 ( .I(register_file_inst1_r3_26_), .ZN(n160) );
  OAI222D0BWP12T U497 ( .A1(n160), .A2(n1064), .B1(n1066), .B2(n504), .C1(
        n1067), .C2(n505), .ZN(register_file_inst1_n2547) );
  INVD1BWP12T U498 ( .I(register_file_inst1_r11_26_), .ZN(n582) );
  OR3D1BWP12T U499 ( .A1(n161), .A2(n1975), .A3(n2279), .Z(n964) );
  OAI222D0BWP12T U500 ( .A1(n582), .A2(n1021), .B1(n964), .B2(n504), .C1(n1019), .C2(n505), .ZN(register_file_inst1_n2291) );
  CKND0BWP12T U501 ( .I(register_file_inst1_r2_25_), .ZN(n162) );
  AOI21D1BWP12T U502 ( .A1(n501), .A2(MEM_MEMCTRL_from_mem_data[1]), .B(n500), 
        .ZN(n506) );
  OAI222D0BWP12T U503 ( .A1(n162), .A2(n1060), .B1(n1062), .B2(n506), .C1(
        n1063), .C2(n507), .ZN(register_file_inst1_n2578) );
  INVD1BWP12T U504 ( .I(register_file_inst1_r9_25_), .ZN(n432) );
  OAI222D0BWP12T U505 ( .A1(n432), .A2(n1079), .B1(n1080), .B2(n506), .C1(
        n1081), .C2(n507), .ZN(register_file_inst1_n2354) );
  INVD1BWP12T U506 ( .I(register_file_inst1_r7_25_), .ZN(n433) );
  OAI222D0BWP12T U507 ( .A1(n433), .A2(n1051), .B1(n1050), .B2(n506), .C1(
        n1049), .C2(n507), .ZN(register_file_inst1_n2418) );
  INVD1BWP12T U508 ( .I(register_file_inst1_r10_25_), .ZN(n1551) );
  OAI222D0BWP12T U509 ( .A1(n1551), .A2(n1068), .B1(n1069), .B2(n506), .C1(
        n1070), .C2(n507), .ZN(register_file_inst1_n2322) );
  INVD1BWP12T U510 ( .I(register_file_inst1_r4_25_), .ZN(n1552) );
  OAI222D0BWP12T U511 ( .A1(n1552), .A2(n1090), .B1(n1091), .B2(n506), .C1(
        n1092), .C2(n507), .ZN(register_file_inst1_n2514) );
  CKND0BWP12T U512 ( .I(register_file_inst1_r12_25_), .ZN(n163) );
  OAI222D0BWP12T U513 ( .A1(n163), .A2(n1071), .B1(n1073), .B2(n506), .C1(
        n1074), .C2(n507), .ZN(register_file_inst1_n2258) );
  INVD1BWP12T U514 ( .I(register_file_inst1_r1_25_), .ZN(n431) );
  OAI222D0BWP12T U515 ( .A1(n431), .A2(n1093), .B1(n1094), .B2(n506), .C1(
        n1095), .C2(n507), .ZN(register_file_inst1_n2610) );
  CKND0BWP12T U516 ( .I(register_file_inst1_tmp1_25_), .ZN(n164) );
  OAI222D0BWP12T U517 ( .A1(n164), .A2(n1027), .B1(n1026), .B2(n506), .C1(
        n2168), .C2(n507), .ZN(register_file_inst1_n2162) );
  CKND0BWP12T U518 ( .I(register_file_inst1_r0_25_), .ZN(n165) );
  OAI222D0BWP12T U519 ( .A1(n165), .A2(n1086), .B1(n1088), .B2(n506), .C1(
        n1089), .C2(n507), .ZN(register_file_inst1_n2642) );
  INVD1BWP12T U520 ( .I(register_file_inst1_r11_25_), .ZN(n1553) );
  OAI222D0BWP12T U521 ( .A1(n1553), .A2(n1021), .B1(n1020), .B2(n506), .C1(
        n1019), .C2(n507), .ZN(register_file_inst1_n2290) );
  CKND0BWP12T U522 ( .I(register_file_inst1_r6_25_), .ZN(n166) );
  OAI222D0BWP12T U523 ( .A1(n166), .A2(n1045), .B1(n1044), .B2(n506), .C1(
        n1043), .C2(n507), .ZN(register_file_inst1_n2450) );
  CKND0BWP12T U524 ( .I(register_file_inst1_r3_25_), .ZN(n167) );
  OAI222D0BWP12T U525 ( .A1(n167), .A2(n1064), .B1(n1066), .B2(n506), .C1(
        n1067), .C2(n507), .ZN(register_file_inst1_n2546) );
  INVD1BWP12T U526 ( .I(register_file_inst1_r5_25_), .ZN(n1554) );
  OAI222D0BWP12T U527 ( .A1(n1554), .A2(n1096), .B1(n1097), .B2(n506), .C1(
        n1098), .C2(n507), .ZN(register_file_inst1_n2482) );
  CKND0BWP12T U528 ( .I(register_file_inst1_lr_25_), .ZN(n168) );
  OAI222D0BWP12T U529 ( .A1(n168), .A2(n1082), .B1(n1084), .B2(n506), .C1(
        n1085), .C2(n507), .ZN(register_file_inst1_n2226) );
  CKND0BWP12T U530 ( .I(register_file_inst1_r8_25_), .ZN(n169) );
  OAI222D0BWP12T U531 ( .A1(n169), .A2(n1075), .B1(n1077), .B2(n506), .C1(
        n1078), .C2(n507), .ZN(register_file_inst1_n2386) );
  CKND0BWP12T U532 ( .I(STACK_RF_next_sp[25]), .ZN(n170) );
  OAI222D0BWP12T U533 ( .A1(n170), .A2(n1099), .B1(n1102), .B2(n506), .C1(
        n1104), .C2(n507), .ZN(register_file_inst1_spin[25]) );
  AOI21D1BWP12T U534 ( .A1(n501), .A2(MEM_MEMCTRL_from_mem_data[0]), .B(n500), 
        .ZN(n508) );
  INVD2BWP12T U535 ( .I(ALU_MISC_OUT_result[24]), .ZN(n509) );
  OAI222D0BWP12T U536 ( .A1(n171), .A2(n1093), .B1(n1094), .B2(n508), .C1(
        n1095), .C2(n509), .ZN(register_file_inst1_n2609) );
  CKND0BWP12T U537 ( .I(register_file_inst1_r12_24_), .ZN(n172) );
  OAI222D0BWP12T U538 ( .A1(n172), .A2(n1071), .B1(n1073), .B2(n508), .C1(
        n1074), .C2(n509), .ZN(register_file_inst1_n2257) );
  CKND0BWP12T U539 ( .I(register_file_inst1_r0_24_), .ZN(n173) );
  OAI222D0BWP12T U540 ( .A1(n173), .A2(n1086), .B1(n1088), .B2(n508), .C1(
        n1089), .C2(n509), .ZN(register_file_inst1_n2641) );
  OAI222D0BWP12T U541 ( .A1(n174), .A2(n1079), .B1(n1080), .B2(n508), .C1(
        n1081), .C2(n509), .ZN(register_file_inst1_n2353) );
  OAI222D0BWP12T U542 ( .A1(n175), .A2(n1051), .B1(n1050), .B2(n508), .C1(
        n1049), .C2(n509), .ZN(register_file_inst1_n2417) );
  CKND0BWP12T U543 ( .I(register_file_inst1_r6_24_), .ZN(n176) );
  OAI222D0BWP12T U544 ( .A1(n176), .A2(n1045), .B1(n1044), .B2(n508), .C1(
        n1043), .C2(n509), .ZN(register_file_inst1_n2449) );
  CKND0BWP12T U545 ( .I(register_file_inst1_r3_24_), .ZN(n177) );
  OAI222D0BWP12T U546 ( .A1(n177), .A2(n1064), .B1(n1066), .B2(n508), .C1(
        n1067), .C2(n509), .ZN(register_file_inst1_n2545) );
  INVD1BWP12T U547 ( .I(register_file_inst1_r10_24_), .ZN(n567) );
  OAI222D0BWP12T U548 ( .A1(n567), .A2(n1068), .B1(n1069), .B2(n508), .C1(
        n1070), .C2(n509), .ZN(register_file_inst1_n2321) );
  CKND0BWP12T U549 ( .I(register_file_inst1_r8_24_), .ZN(n178) );
  OAI222D0BWP12T U550 ( .A1(n178), .A2(n1075), .B1(n1077), .B2(n508), .C1(
        n1078), .C2(n509), .ZN(register_file_inst1_n2385) );
  CKND0BWP12T U551 ( .I(register_file_inst1_tmp1_24_), .ZN(n179) );
  OAI222D0BWP12T U552 ( .A1(n179), .A2(n1027), .B1(n1026), .B2(n508), .C1(
        n2168), .C2(n509), .ZN(register_file_inst1_n2161) );
  CKND0BWP12T U553 ( .I(register_file_inst1_r2_24_), .ZN(n180) );
  OAI222D0BWP12T U554 ( .A1(n180), .A2(n1060), .B1(n1062), .B2(n508), .C1(
        n1063), .C2(n509), .ZN(register_file_inst1_n2577) );
  OAI222D0BWP12T U555 ( .A1(n569), .A2(n1021), .B1(n964), .B2(n508), .C1(n1019), .C2(n509), .ZN(register_file_inst1_n2289) );
  INVD1BWP12T U556 ( .I(register_file_inst1_r5_24_), .ZN(n570) );
  OAI222D0BWP12T U557 ( .A1(n570), .A2(n1096), .B1(n1097), .B2(n508), .C1(
        n1098), .C2(n509), .ZN(register_file_inst1_n2481) );
  CKND0BWP12T U558 ( .I(STACK_RF_next_sp[24]), .ZN(n181) );
  OAI222D0BWP12T U559 ( .A1(n181), .A2(n1099), .B1(n1102), .B2(n508), .C1(
        n1104), .C2(n509), .ZN(register_file_inst1_spin[24]) );
  CKND0BWP12T U560 ( .I(register_file_inst1_lr_24_), .ZN(n182) );
  OAI222D0BWP12T U561 ( .A1(n182), .A2(n1082), .B1(n1084), .B2(n508), .C1(
        n1085), .C2(n509), .ZN(register_file_inst1_n2225) );
  INVD1BWP12T U562 ( .I(register_file_inst1_r4_24_), .ZN(n568) );
  OAI222D0BWP12T U563 ( .A1(n568), .A2(n1090), .B1(n1091), .B2(n508), .C1(
        n1092), .C2(n509), .ZN(register_file_inst1_n2513) );
  IAO21D1BWP12T U564 ( .A1(n2327), .A2(n885), .B(n500), .ZN(n510) );
  OAI222D0BWP12T U565 ( .A1(n183), .A2(n1079), .B1(n1080), .B2(n510), .C1(
        n1081), .C2(n511), .ZN(register_file_inst1_n2352) );
  OAI222D0BWP12T U566 ( .A1(n1890), .A2(n1021), .B1(n964), .B2(n510), .C1(
        n1019), .C2(n511), .ZN(register_file_inst1_n2288) );
  CKND0BWP12T U567 ( .I(STACK_RF_next_sp[23]), .ZN(n184) );
  OAI222D0BWP12T U568 ( .A1(n184), .A2(n1037), .B1(n1102), .B2(n510), .C1(
        n1104), .C2(n511), .ZN(register_file_inst1_spin[23]) );
  INVD1BWP12T U569 ( .I(register_file_inst1_r10_23_), .ZN(n1888) );
  OAI222D0BWP12T U570 ( .A1(n1888), .A2(n1068), .B1(n1069), .B2(n510), .C1(
        n1070), .C2(n511), .ZN(register_file_inst1_n2320) );
  CKND0BWP12T U571 ( .I(register_file_inst1_r8_23_), .ZN(n185) );
  OAI222D0BWP12T U572 ( .A1(n185), .A2(n1075), .B1(n1077), .B2(n510), .C1(
        n1078), .C2(n511), .ZN(register_file_inst1_n2384) );
  CKND0BWP12T U573 ( .I(register_file_inst1_r0_23_), .ZN(n186) );
  OAI222D0BWP12T U574 ( .A1(n186), .A2(n1086), .B1(n1088), .B2(n510), .C1(
        n1089), .C2(n511), .ZN(register_file_inst1_n2640) );
  CKND0BWP12T U575 ( .I(register_file_inst1_lr_23_), .ZN(n187) );
  OAI222D0BWP12T U576 ( .A1(n187), .A2(n1082), .B1(n1084), .B2(n510), .C1(
        n1085), .C2(n511), .ZN(register_file_inst1_n2224) );
  CKND0BWP12T U577 ( .I(register_file_inst1_r2_23_), .ZN(n188) );
  OAI222D0BWP12T U578 ( .A1(n188), .A2(n1060), .B1(n1062), .B2(n510), .C1(
        n1063), .C2(n511), .ZN(register_file_inst1_n2576) );
  CKND0BWP12T U579 ( .I(register_file_inst1_r12_23_), .ZN(n189) );
  OAI222D0BWP12T U580 ( .A1(n189), .A2(n1071), .B1(n1073), .B2(n510), .C1(
        n1074), .C2(n511), .ZN(register_file_inst1_n2256) );
  OAI222D0BWP12T U581 ( .A1(n190), .A2(n1051), .B1(n1050), .B2(n510), .C1(
        n1049), .C2(n511), .ZN(register_file_inst1_n2416) );
  INVD1BWP12T U582 ( .I(register_file_inst1_r5_23_), .ZN(n1891) );
  OAI222D0BWP12T U583 ( .A1(n1891), .A2(n1096), .B1(n1097), .B2(n510), .C1(
        n1098), .C2(n511), .ZN(register_file_inst1_n2480) );
  CKND0BWP12T U584 ( .I(register_file_inst1_tmp1_23_), .ZN(n191) );
  OAI222D0BWP12T U585 ( .A1(n191), .A2(n1027), .B1(n1026), .B2(n510), .C1(
        n2168), .C2(n511), .ZN(register_file_inst1_n2160) );
  CKND0BWP12T U586 ( .I(register_file_inst1_r6_23_), .ZN(n192) );
  OAI222D0BWP12T U587 ( .A1(n192), .A2(n1045), .B1(n1044), .B2(n510), .C1(
        n1043), .C2(n511), .ZN(register_file_inst1_n2448) );
  OAI222D0BWP12T U588 ( .A1(n193), .A2(n1093), .B1(n1094), .B2(n510), .C1(
        n1095), .C2(n511), .ZN(register_file_inst1_n2608) );
  INVD1BWP12T U589 ( .I(register_file_inst1_r4_23_), .ZN(n1889) );
  OAI222D0BWP12T U590 ( .A1(n1889), .A2(n1090), .B1(n1091), .B2(n510), .C1(
        n1092), .C2(n511), .ZN(register_file_inst1_n2512) );
  CKND0BWP12T U591 ( .I(register_file_inst1_r3_23_), .ZN(n194) );
  OAI222D0BWP12T U592 ( .A1(n194), .A2(n1064), .B1(n1066), .B2(n510), .C1(
        n1067), .C2(n511), .ZN(register_file_inst1_n2544) );
  XOR2XD1BWP12T U593 ( .A1(n1930), .A2(n195), .Z(
        register_file_inst1_pc_write_in_plus_two[6]) );
  CKND0BWP12T U594 ( .I(register_file_inst1_lr_21_), .ZN(n196) );
  IAO21D1BWP12T U595 ( .A1(n2329), .A2(n885), .B(n500), .ZN(n512) );
  OAI222D0BWP12T U596 ( .A1(n196), .A2(n1082), .B1(n1084), .B2(n512), .C1(
        n1085), .C2(n513), .ZN(register_file_inst1_n2222) );
  INVD1BWP12T U597 ( .I(register_file_inst1_r7_21_), .ZN(n548) );
  OAI222D0BWP12T U598 ( .A1(n548), .A2(n1051), .B1(n1050), .B2(n512), .C1(
        n1049), .C2(n513), .ZN(register_file_inst1_n2414) );
  CKND0BWP12T U599 ( .I(register_file_inst1_tmp1_21_), .ZN(n197) );
  OAI222D0BWP12T U600 ( .A1(n197), .A2(n1027), .B1(n1026), .B2(n512), .C1(
        n2168), .C2(n513), .ZN(register_file_inst1_n2158) );
  CKND0BWP12T U601 ( .I(register_file_inst1_r6_21_), .ZN(n198) );
  OAI222D0BWP12T U602 ( .A1(n198), .A2(n1045), .B1(n1044), .B2(n512), .C1(
        n1043), .C2(n513), .ZN(register_file_inst1_n2446) );
  INVD1BWP12T U603 ( .I(register_file_inst1_r11_21_), .ZN(n1906) );
  OAI222D0BWP12T U604 ( .A1(n1906), .A2(n1021), .B1(n964), .B2(n512), .C1(
        n1019), .C2(n513), .ZN(register_file_inst1_n2286) );
  CKND0BWP12T U605 ( .I(register_file_inst1_r2_21_), .ZN(n199) );
  OAI222D0BWP12T U606 ( .A1(n199), .A2(n1060), .B1(n1062), .B2(n512), .C1(
        n1063), .C2(n513), .ZN(register_file_inst1_n2574) );
  INVD1BWP12T U607 ( .I(register_file_inst1_r5_21_), .ZN(n1908) );
  OAI222D0BWP12T U608 ( .A1(n1908), .A2(n1096), .B1(n1097), .B2(n512), .C1(
        n1098), .C2(n513), .ZN(register_file_inst1_n2478) );
  INVD1BWP12T U609 ( .I(register_file_inst1_lr_19_), .ZN(n1530) );
  OAI222D1BWP12T U610 ( .A1(n1530), .A2(n1082), .B1(n1084), .B2(n971), .C1(
        n1085), .C2(n970), .ZN(register_file_inst1_n2220) );
  INVD1BWP12T U611 ( .I(register_file_inst1_r9_21_), .ZN(n547) );
  OAI222D0BWP12T U612 ( .A1(n547), .A2(n1079), .B1(n1080), .B2(n512), .C1(
        n1081), .C2(n513), .ZN(register_file_inst1_n2350) );
  CKND0BWP12T U613 ( .I(register_file_inst1_r3_21_), .ZN(n200) );
  OAI222D0BWP12T U614 ( .A1(n200), .A2(n1064), .B1(n1066), .B2(n512), .C1(
        n1067), .C2(n513), .ZN(register_file_inst1_n2542) );
  INVD1BWP12T U615 ( .I(register_file_inst1_r1_21_), .ZN(n546) );
  OAI222D0BWP12T U616 ( .A1(n546), .A2(n1093), .B1(n1094), .B2(n512), .C1(
        n1095), .C2(n513), .ZN(register_file_inst1_n2606) );
  CKND0BWP12T U617 ( .I(STACK_RF_next_sp[21]), .ZN(n201) );
  OAI222D0BWP12T U618 ( .A1(n201), .A2(n1099), .B1(n1102), .B2(n512), .C1(
        n1104), .C2(n513), .ZN(register_file_inst1_spin[21]) );
  CKND0BWP12T U619 ( .I(register_file_inst1_r12_21_), .ZN(n202) );
  OAI222D0BWP12T U620 ( .A1(n202), .A2(n1071), .B1(n1073), .B2(n512), .C1(
        n1074), .C2(n513), .ZN(register_file_inst1_n2254) );
  CKND0BWP12T U621 ( .I(register_file_inst1_r8_21_), .ZN(n203) );
  OAI222D0BWP12T U622 ( .A1(n203), .A2(n1075), .B1(n1077), .B2(n512), .C1(
        n1078), .C2(n513), .ZN(register_file_inst1_n2382) );
  CKND0BWP12T U623 ( .I(register_file_inst1_r0_21_), .ZN(n204) );
  OAI222D0BWP12T U624 ( .A1(n204), .A2(n1086), .B1(n1088), .B2(n512), .C1(
        n1089), .C2(n513), .ZN(register_file_inst1_n2638) );
  INVD1BWP12T U625 ( .I(register_file_inst1_r10_21_), .ZN(n1902) );
  OAI222D0BWP12T U626 ( .A1(n1902), .A2(n1068), .B1(n1069), .B2(n512), .C1(
        n1070), .C2(n513), .ZN(register_file_inst1_n2318) );
  INVD1BWP12T U627 ( .I(register_file_inst1_r4_21_), .ZN(n1904) );
  OAI222D0BWP12T U628 ( .A1(n1904), .A2(n1090), .B1(n1091), .B2(n512), .C1(
        n1092), .C2(n513), .ZN(register_file_inst1_n2510) );
  INVD1BWP12T U629 ( .I(register_file_inst1_r9_18_), .ZN(n1137) );
  OAI222D0BWP12T U630 ( .A1(n1137), .A2(n1079), .B1(n1080), .B2(n219), .C1(
        n1081), .C2(n218), .ZN(register_file_inst1_n2347) );
  INVD1BWP12T U631 ( .I(register_file_inst1_r12_17_), .ZN(n1159) );
  INVD1BWP12T U632 ( .I(ALU_MISC_OUT_result[17]), .ZN(n216) );
  OAI222D0BWP12T U633 ( .A1(n1159), .A2(n1071), .B1(n1073), .B2(n217), .C1(
        n1074), .C2(n216), .ZN(register_file_inst1_n2250) );
  INVD1BWP12T U634 ( .I(STACK_RF_next_sp[17]), .ZN(n1158) );
  OAI222D0BWP12T U635 ( .A1(n1158), .A2(n1099), .B1(n1102), .B2(n217), .C1(
        n1104), .C2(n216), .ZN(register_file_inst1_spin[17]) );
  INVD1BWP12T U636 ( .I(register_file_inst1_r9_17_), .ZN(n1148) );
  OAI222D0BWP12T U637 ( .A1(n1148), .A2(n1079), .B1(n1080), .B2(n217), .C1(
        n1081), .C2(n216), .ZN(register_file_inst1_n2346) );
  CKND0BWP12T U638 ( .I(register_file_inst1_r8_18_), .ZN(n205) );
  OAI222D0BWP12T U639 ( .A1(n205), .A2(n1075), .B1(n1077), .B2(n219), .C1(
        n1078), .C2(n218), .ZN(register_file_inst1_n2379) );
  INVD1BWP12T U640 ( .I(register_file_inst1_r4_20_), .ZN(n522) );
  OAI222D0BWP12T U641 ( .A1(n522), .A2(n1090), .B1(n1091), .B2(n515), .C1(
        n1092), .C2(n516), .ZN(register_file_inst1_n2509) );
  CKND0BWP12T U642 ( .I(register_file_inst1_tmp1_20_), .ZN(n206) );
  OAI222D0BWP12T U643 ( .A1(n206), .A2(n1027), .B1(n1026), .B2(n515), .C1(
        n2168), .C2(n516), .ZN(register_file_inst1_n2157) );
  INVD1BWP12T U644 ( .I(register_file_inst1_r11_18_), .ZN(n1135) );
  OAI222D0BWP12T U645 ( .A1(n1135), .A2(n1021), .B1(n964), .B2(n219), .C1(
        n1019), .C2(n218), .ZN(register_file_inst1_n2283) );
  INVD1BWP12T U646 ( .I(register_file_inst1_r5_20_), .ZN(n523) );
  OAI222D0BWP12T U647 ( .A1(n523), .A2(n1096), .B1(n1097), .B2(n515), .C1(
        n1098), .C2(n516), .ZN(register_file_inst1_n2477) );
  INVD1BWP12T U648 ( .I(register_file_inst1_r4_18_), .ZN(n1125) );
  OAI222D0BWP12T U649 ( .A1(n1125), .A2(n1090), .B1(n1091), .B2(n219), .C1(
        n1092), .C2(n218), .ZN(register_file_inst1_n2507) );
  INVD1BWP12T U650 ( .I(register_file_inst1_lr_18_), .ZN(n1117) );
  OAI222D0BWP12T U651 ( .A1(n1117), .A2(n1082), .B1(n1084), .B2(n219), .C1(
        n1085), .C2(n218), .ZN(register_file_inst1_n2219) );
  INVD1BWP12T U652 ( .I(register_file_inst1_r4_17_), .ZN(n1172) );
  OAI222D0BWP12T U653 ( .A1(n1172), .A2(n1090), .B1(n1091), .B2(n217), .C1(
        n1092), .C2(n216), .ZN(register_file_inst1_n2506) );
  INVD1BWP12T U654 ( .I(register_file_inst1_tmp1_18_), .ZN(n1128) );
  OAI222D0BWP12T U655 ( .A1(n1128), .A2(n1027), .B1(n1026), .B2(n219), .C1(
        n2168), .C2(n218), .ZN(register_file_inst1_n2155) );
  CKND0BWP12T U656 ( .I(register_file_inst1_r8_20_), .ZN(n207) );
  OAI222D0BWP12T U657 ( .A1(n207), .A2(n1075), .B1(n1077), .B2(n515), .C1(
        n1078), .C2(n516), .ZN(register_file_inst1_n2381) );
  INVD1BWP12T U658 ( .I(register_file_inst1_tmp1_17_), .ZN(n1176) );
  OAI222D0BWP12T U659 ( .A1(n1176), .A2(n1027), .B1(n1026), .B2(n217), .C1(
        n2168), .C2(n216), .ZN(register_file_inst1_n2154) );
  INVD1BWP12T U660 ( .I(register_file_inst1_r7_17_), .ZN(n1163) );
  OAI222D0BWP12T U661 ( .A1(n1163), .A2(n1051), .B1(n1050), .B2(n217), .C1(
        n1049), .C2(n216), .ZN(register_file_inst1_n2410) );
  INVD1BWP12T U662 ( .I(register_file_inst1_r0_18_), .ZN(n1115) );
  OAI222D0BWP12T U663 ( .A1(n1115), .A2(n1086), .B1(n1088), .B2(n219), .C1(
        n1089), .C2(n218), .ZN(register_file_inst1_n2635) );
  INVD1BWP12T U664 ( .I(register_file_inst1_r10_17_), .ZN(n1171) );
  OAI222D0BWP12T U665 ( .A1(n1171), .A2(n1068), .B1(n1069), .B2(n217), .C1(
        n1070), .C2(n216), .ZN(register_file_inst1_n2314) );
  INVD1BWP12T U666 ( .I(register_file_inst1_r0_17_), .ZN(n1160) );
  OAI222D0BWP12T U667 ( .A1(n1160), .A2(n1086), .B1(n1088), .B2(n217), .C1(
        n1089), .C2(n216), .ZN(register_file_inst1_n2634) );
  INVD1BWP12T U668 ( .I(register_file_inst1_lr_17_), .ZN(n1162) );
  OAI222D0BWP12T U669 ( .A1(n1162), .A2(n1082), .B1(n1084), .B2(n217), .C1(
        n1085), .C2(n216), .ZN(register_file_inst1_n2218) );
  INVD1BWP12T U670 ( .I(register_file_inst1_r10_18_), .ZN(n1124) );
  OAI222D0BWP12T U671 ( .A1(n1124), .A2(n1068), .B1(n1069), .B2(n219), .C1(
        n1070), .C2(n218), .ZN(register_file_inst1_n2315) );
  INVD1BWP12T U672 ( .I(register_file_inst1_r11_17_), .ZN(n1173) );
  OAI222D0BWP12T U673 ( .A1(n1173), .A2(n1021), .B1(n1020), .B2(n217), .C1(
        n1019), .C2(n216), .ZN(register_file_inst1_n2282) );
  INVD1BWP12T U674 ( .I(register_file_inst1_r7_18_), .ZN(n1138) );
  OAI222D0BWP12T U675 ( .A1(n1138), .A2(n1051), .B1(n1050), .B2(n219), .C1(
        n1049), .C2(n218), .ZN(register_file_inst1_n2411) );
  INVD1BWP12T U676 ( .I(register_file_inst1_r7_20_), .ZN(n536) );
  OAI222D0BWP12T U677 ( .A1(n536), .A2(n1051), .B1(n1050), .B2(n515), .C1(
        n1049), .C2(n516), .ZN(register_file_inst1_n2413) );
  INVD1BWP12T U678 ( .I(register_file_inst1_r10_20_), .ZN(n521) );
  OAI222D0BWP12T U679 ( .A1(n521), .A2(n1068), .B1(n1069), .B2(n515), .C1(
        n1070), .C2(n516), .ZN(register_file_inst1_n2317) );
  CKND0BWP12T U680 ( .I(register_file_inst1_r8_17_), .ZN(n208) );
  OAI222D0BWP12T U681 ( .A1(n208), .A2(n1075), .B1(n1077), .B2(n217), .C1(
        n1078), .C2(n216), .ZN(register_file_inst1_n2378) );
  INVD1BWP12T U682 ( .I(register_file_inst1_r1_17_), .ZN(n1164) );
  OAI222D0BWP12T U683 ( .A1(n1164), .A2(n1093), .B1(n1094), .B2(n217), .C1(
        n1095), .C2(n216), .ZN(register_file_inst1_n2602) );
  INVD1BWP12T U684 ( .I(register_file_inst1_r3_17_), .ZN(n1161) );
  OAI222D0BWP12T U685 ( .A1(n1161), .A2(n1064), .B1(n1066), .B2(n217), .C1(
        n1067), .C2(n216), .ZN(register_file_inst1_n2538) );
  INVD1BWP12T U686 ( .I(register_file_inst1_r11_20_), .ZN(n533) );
  OAI222D0BWP12T U687 ( .A1(n533), .A2(n1021), .B1(n1020), .B2(n515), .C1(
        n1019), .C2(n516), .ZN(register_file_inst1_n2285) );
  CKND0BWP12T U688 ( .I(register_file_inst1_r12_20_), .ZN(n209) );
  OAI222D0BWP12T U689 ( .A1(n209), .A2(n1071), .B1(n1073), .B2(n515), .C1(
        n1074), .C2(n516), .ZN(register_file_inst1_n2253) );
  INVD1BWP12T U690 ( .I(register_file_inst1_r9_20_), .ZN(n535) );
  OAI222D0BWP12T U691 ( .A1(n535), .A2(n1079), .B1(n1080), .B2(n515), .C1(
        n1081), .C2(n516), .ZN(register_file_inst1_n2349) );
  CKXOR2D1BWP12T U692 ( .A1(n16), .A2(n210), .Z(
        register_file_inst1_pc_write_in_plus_two[4]) );
  CKND0BWP12T U693 ( .I(register_file_inst1_r3_20_), .ZN(n211) );
  OAI222D0BWP12T U694 ( .A1(n211), .A2(n1064), .B1(n1066), .B2(n515), .C1(
        n1067), .C2(n516), .ZN(register_file_inst1_n2541) );
  CKND0BWP12T U695 ( .I(register_file_inst1_r2_17_), .ZN(n212) );
  OAI222D0BWP12T U696 ( .A1(n212), .A2(n1060), .B1(n1062), .B2(n217), .C1(
        n1063), .C2(n216), .ZN(register_file_inst1_n2570) );
  INVD1BWP12T U697 ( .I(register_file_inst1_r12_18_), .ZN(n1114) );
  OAI222D0BWP12T U698 ( .A1(n1114), .A2(n1071), .B1(n1073), .B2(n219), .C1(
        n1074), .C2(n218), .ZN(register_file_inst1_n2251) );
  INVD1BWP12T U699 ( .I(register_file_inst1_r1_20_), .ZN(n534) );
  OAI222D0BWP12T U700 ( .A1(n534), .A2(n1093), .B1(n1094), .B2(n515), .C1(
        n1095), .C2(n516), .ZN(register_file_inst1_n2605) );
  INVD1BWP12T U701 ( .I(register_file_inst1_r3_18_), .ZN(n1116) );
  OAI222D0BWP12T U702 ( .A1(n1116), .A2(n1064), .B1(n1066), .B2(n219), .C1(
        n1067), .C2(n218), .ZN(register_file_inst1_n2539) );
  CKND0BWP12T U703 ( .I(register_file_inst1_r2_20_), .ZN(n213) );
  OAI222D0BWP12T U704 ( .A1(n213), .A2(n1060), .B1(n1062), .B2(n515), .C1(
        n1063), .C2(n516), .ZN(register_file_inst1_n2573) );
  INVD1BWP12T U705 ( .I(register_file_inst1_r6_17_), .ZN(n1175) );
  OAI222D0BWP12T U706 ( .A1(n1175), .A2(n1045), .B1(n1044), .B2(n217), .C1(
        n1043), .C2(n216), .ZN(register_file_inst1_n2442) );
  CKND0BWP12T U707 ( .I(register_file_inst1_r2_18_), .ZN(n214) );
  OAI222D0BWP12T U708 ( .A1(n214), .A2(n1060), .B1(n1062), .B2(n219), .C1(
        n1063), .C2(n218), .ZN(register_file_inst1_n2571) );
  INVD1BWP12T U709 ( .I(STACK_RF_next_sp[18]), .ZN(n1113) );
  ND2D1BWP12T U710 ( .A1(n1978), .A2(n215), .ZN(n975) );
  OAI222D0BWP12T U711 ( .A1(n1113), .A2(n975), .B1(n1102), .B2(n219), .C1(
        n1104), .C2(n218), .ZN(register_file_inst1_spin[18]) );
  INVD1BWP12T U712 ( .I(register_file_inst1_r1_18_), .ZN(n1136) );
  OAI222D0BWP12T U713 ( .A1(n1136), .A2(n1093), .B1(n1094), .B2(n219), .C1(
        n1095), .C2(n218), .ZN(register_file_inst1_n2603) );
  INVD1BWP12T U714 ( .I(register_file_inst1_r5_18_), .ZN(n1126) );
  OAI222D0BWP12T U715 ( .A1(n1126), .A2(n1096), .B1(n1097), .B2(n219), .C1(
        n1098), .C2(n218), .ZN(register_file_inst1_n2475) );
  INVD1BWP12T U716 ( .I(register_file_inst1_r5_17_), .ZN(n1174) );
  OAI222D0BWP12T U717 ( .A1(n1174), .A2(n1096), .B1(n1097), .B2(n217), .C1(
        n1098), .C2(n216), .ZN(register_file_inst1_n2474) );
  INVD1BWP12T U718 ( .I(register_file_inst1_r6_18_), .ZN(n1127) );
  OAI222D0BWP12T U719 ( .A1(n1127), .A2(n1045), .B1(n1044), .B2(n219), .C1(
        n1043), .C2(n218), .ZN(register_file_inst1_n2443) );
  INVD1BWP12T U720 ( .I(ALU_MISC_OUT_result[14]), .ZN(n233) );
  OAI222D0BWP12T U721 ( .A1(n1254), .A2(n1093), .B1(n233), .B2(n1095), .C1(
        n2132), .C2(n1094), .ZN(register_file_inst1_n2599) );
  OAI222D0BWP12T U722 ( .A1(n1256), .A2(n1051), .B1(n233), .B2(n1049), .C1(
        n2132), .C2(n1050), .ZN(register_file_inst1_n2407) );
  INVD1BWP12T U723 ( .I(register_file_inst1_r6_15_), .ZN(n1245) );
  INVD1BWP12T U724 ( .I(ALU_MISC_OUT_result[15]), .ZN(n236) );
  OAI222D0BWP12T U725 ( .A1(n1245), .A2(n1045), .B1(n236), .B2(n1043), .C1(
        n2135), .C2(n1044), .ZN(register_file_inst1_n2440) );
  OAI222D0BWP12T U726 ( .A1(n2132), .A2(n1069), .B1(n233), .B2(n1070), .C1(
        n1068), .C2(n220), .ZN(register_file_inst1_n2311) );
  OAI222D0BWP12T U727 ( .A1(n2132), .A2(n1066), .B1(n233), .B2(n1067), .C1(
        n1064), .C2(n221), .ZN(register_file_inst1_n2535) );
  CKND0BWP12T U728 ( .I(register_file_inst1_r2_15_), .ZN(n222) );
  OAI222D0BWP12T U729 ( .A1(n2135), .A2(n1062), .B1(n236), .B2(n1063), .C1(
        n1060), .C2(n222), .ZN(register_file_inst1_n2568) );
  INVD1BWP12T U730 ( .I(register_file_inst1_r10_15_), .ZN(n1241) );
  OAI222D0BWP12T U731 ( .A1(n2135), .A2(n1069), .B1(n236), .B2(n1070), .C1(
        n1068), .C2(n1241), .ZN(register_file_inst1_n2312) );
  INVD1BWP12T U732 ( .I(register_file_inst1_r3_15_), .ZN(n1231) );
  OAI222D0BWP12T U733 ( .A1(n2135), .A2(n1066), .B1(n236), .B2(n1067), .C1(
        n1064), .C2(n1231), .ZN(register_file_inst1_n2536) );
  INVD1BWP12T U734 ( .I(register_file_inst1_tmp1_15_), .ZN(n1246) );
  OAI222D0BWP12T U735 ( .A1(n2135), .A2(n1026), .B1(n236), .B2(n2168), .C1(
        n1027), .C2(n1246), .ZN(register_file_inst1_n2152) );
  INVD1BWP12T U736 ( .I(register_file_inst1_r7_15_), .ZN(n1233) );
  OAI222D0BWP12T U737 ( .A1(n1233), .A2(n1051), .B1(n236), .B2(n1049), .C1(
        n2135), .C2(n1050), .ZN(register_file_inst1_n2408) );
  OAI222D0BWP12T U738 ( .A1(n223), .A2(n1096), .B1(n233), .B2(n1098), .C1(
        n2132), .C2(n1097), .ZN(register_file_inst1_n2471) );
  CKND0BWP12T U739 ( .I(register_file_inst1_r2_14_), .ZN(n224) );
  OAI222D0BWP12T U740 ( .A1(n2132), .A2(n1062), .B1(n233), .B2(n1063), .C1(
        n1060), .C2(n224), .ZN(register_file_inst1_n2567) );
  INVD1BWP12T U741 ( .I(register_file_inst1_r1_15_), .ZN(n1234) );
  OAI222D0BWP12T U742 ( .A1(n1234), .A2(n1093), .B1(n236), .B2(n1095), .C1(
        n2135), .C2(n1094), .ZN(register_file_inst1_n2600) );
  OAI222D0BWP12T U743 ( .A1(n225), .A2(n1045), .B1(n233), .B2(n1043), .C1(
        n2132), .C2(n1044), .ZN(register_file_inst1_n2439) );
  INVD1BWP12T U744 ( .I(register_file_inst1_r5_15_), .ZN(n1244) );
  OAI222D0BWP12T U745 ( .A1(n1244), .A2(n1096), .B1(n236), .B2(n1098), .C1(
        n2135), .C2(n1097), .ZN(register_file_inst1_n2472) );
  XOR2XD1BWP12T U746 ( .A1(n15), .A2(n226), .Z(
        register_file_inst1_pc_write_in_plus_two[2]) );
  OAI222D0BWP12T U747 ( .A1(n227), .A2(n1099), .B1(n233), .B2(n1104), .C1(
        n2132), .C2(n1102), .ZN(register_file_inst1_spin[14]) );
  OAI222D0BWP12T U748 ( .A1(n2132), .A2(n1020), .B1(n233), .B2(n1019), .C1(
        n1021), .C2(n1253), .ZN(register_file_inst1_n2279) );
  INVD1BWP12T U749 ( .I(register_file_inst1_r9_14_), .ZN(n1255) );
  OAI222D0BWP12T U750 ( .A1(n1255), .A2(n1079), .B1(n233), .B2(n1081), .C1(
        n2132), .C2(n1080), .ZN(register_file_inst1_n2343) );
  INVD1BWP12T U751 ( .I(register_file_inst1_r11_15_), .ZN(n1243) );
  OAI222D0BWP12T U752 ( .A1(n2135), .A2(n1020), .B1(n236), .B2(n1019), .C1(
        n1021), .C2(n1243), .ZN(register_file_inst1_n2280) );
  OAI222D0BWP12T U753 ( .A1(n2132), .A2(n1026), .B1(n233), .B2(n2168), .C1(
        n1027), .C2(n228), .ZN(register_file_inst1_n2151) );
  INVD1BWP12T U754 ( .I(register_file_inst1_r12_15_), .ZN(n1229) );
  OAI222D0BWP12T U755 ( .A1(n1229), .A2(n1071), .B1(n236), .B2(n1074), .C1(
        n2135), .C2(n1073), .ZN(register_file_inst1_n2248) );
  CKND0BWP12T U756 ( .I(register_file_inst1_r8_14_), .ZN(n229) );
  OAI222D0BWP12T U757 ( .A1(n229), .A2(n1075), .B1(n233), .B2(n1078), .C1(
        n2132), .C2(n1077), .ZN(register_file_inst1_n2375) );
  INVD1BWP12T U758 ( .I(register_file_inst1_r9_15_), .ZN(n1218) );
  OAI222D0BWP12T U759 ( .A1(n1218), .A2(n1079), .B1(n236), .B2(n1081), .C1(
        n2135), .C2(n1080), .ZN(register_file_inst1_n2344) );
  OAI222D0BWP12T U760 ( .A1(n230), .A2(n1090), .B1(n233), .B2(n1092), .C1(
        n2132), .C2(n1091), .ZN(register_file_inst1_n2503) );
  OAI222D0BWP12T U761 ( .A1(n231), .A2(n1082), .B1(n233), .B2(n1085), .C1(
        n2132), .C2(n1084), .ZN(register_file_inst1_n2215) );
  INVD1BWP12T U762 ( .I(register_file_inst1_r4_15_), .ZN(n1242) );
  OAI222D0BWP12T U763 ( .A1(n1242), .A2(n1090), .B1(n236), .B2(n1092), .C1(
        n2135), .C2(n1091), .ZN(register_file_inst1_n2504) );
  INVD1BWP12T U764 ( .I(register_file_inst1_lr_15_), .ZN(n1232) );
  OAI222D0BWP12T U765 ( .A1(n1232), .A2(n1082), .B1(n236), .B2(n1085), .C1(
        n2135), .C2(n1084), .ZN(register_file_inst1_n2216) );
  OAI222D0BWP12T U766 ( .A1(n232), .A2(n1071), .B1(n233), .B2(n1074), .C1(
        n2132), .C2(n1073), .ZN(register_file_inst1_n2247) );
  OAI222D0BWP12T U767 ( .A1(n234), .A2(n1086), .B1(n233), .B2(n1089), .C1(
        n2132), .C2(n1088), .ZN(register_file_inst1_n2631) );
  CKND0BWP12T U768 ( .I(register_file_inst1_r8_15_), .ZN(n235) );
  OAI222D0BWP12T U769 ( .A1(n235), .A2(n1075), .B1(n236), .B2(n1078), .C1(
        n2135), .C2(n1077), .ZN(register_file_inst1_n2376) );
  INVD1BWP12T U770 ( .I(register_file_inst1_r0_15_), .ZN(n1230) );
  OAI222D0BWP12T U771 ( .A1(n1230), .A2(n1086), .B1(n236), .B2(n1089), .C1(
        n2135), .C2(n1088), .ZN(register_file_inst1_n2632) );
  INVD1BWP12T U772 ( .I(STACK_RF_next_sp[15]), .ZN(n1228) );
  OAI222D0BWP12T U773 ( .A1(n1228), .A2(n975), .B1(n236), .B2(n1104), .C1(
        n2135), .C2(n1102), .ZN(register_file_inst1_spin[15]) );
  INVD1BWP12T U774 ( .I(ALU_MISC_OUT_result[2]), .ZN(n239) );
  INVD1BWP12T U775 ( .I(register_file_inst1_r3_2_), .ZN(n1804) );
  OAI222D0BWP12T U776 ( .A1(n2101), .A2(n1066), .B1(n239), .B2(n1067), .C1(
        n1064), .C2(n1804), .ZN(register_file_inst1_n2523) );
  TPOAI21D0BWP12T U777 ( .A1(n239), .A2(n1104), .B(n1991), .ZN(
        register_file_inst1_spin[2]) );
  INVD1BWP12T U778 ( .I(register_file_inst1_tmp1_2_), .ZN(n1824) );
  OAI222D0BWP12T U779 ( .A1(n2101), .A2(n1026), .B1(n239), .B2(n2168), .C1(
        n1027), .C2(n1824), .ZN(register_file_inst1_n2139) );
  INVD1BWP12T U780 ( .I(register_file_inst1_r8_2_), .ZN(n1734) );
  OAI222D0BWP12T U781 ( .A1(n1734), .A2(n1075), .B1(n239), .B2(n1078), .C1(
        n2101), .C2(n1077), .ZN(register_file_inst1_n2363) );
  INVD1BWP12T U782 ( .I(register_file_inst1_r7_2_), .ZN(n1808) );
  OAI222D0BWP12T U783 ( .A1(n1808), .A2(n1051), .B1(n239), .B2(n1049), .C1(
        n2101), .C2(n1050), .ZN(register_file_inst1_n2395) );
  INVD1BWP12T U784 ( .I(register_file_inst1_r4_2_), .ZN(n1818) );
  OAI222D0BWP12T U785 ( .A1(n1818), .A2(n1090), .B1(n239), .B2(n1092), .C1(
        n2101), .C2(n1091), .ZN(register_file_inst1_n2491) );
  INVD1BWP12T U786 ( .I(register_file_inst1_r5_2_), .ZN(n1820) );
  OAI222D0BWP12T U787 ( .A1(n1820), .A2(n1096), .B1(n239), .B2(n1098), .C1(
        n2101), .C2(n1097), .ZN(register_file_inst1_n2459) );
  INVD1BWP12T U788 ( .I(register_file_inst1_lr_2_), .ZN(n1806) );
  OAI222D0BWP12T U789 ( .A1(n1806), .A2(n1082), .B1(n239), .B2(n1085), .C1(
        n2101), .C2(n1084), .ZN(register_file_inst1_n2203) );
  CKND0BWP12T U790 ( .I(register_file_inst1_r2_2_), .ZN(n237) );
  OAI222D0BWP12T U791 ( .A1(n2101), .A2(n1062), .B1(n239), .B2(n1063), .C1(
        n1060), .C2(n237), .ZN(register_file_inst1_n2555) );
  INVD1BWP12T U792 ( .I(register_file_inst1_r12_2_), .ZN(n1799) );
  OAI222D0BWP12T U793 ( .A1(n1799), .A2(n1071), .B1(n239), .B2(n1074), .C1(
        n2101), .C2(n1073), .ZN(register_file_inst1_n2235) );
  INVD1BWP12T U794 ( .I(register_file_inst1_r11_2_), .ZN(n1819) );
  OAI222D0BWP12T U795 ( .A1(n2101), .A2(n964), .B1(n239), .B2(n1019), .C1(
        n1021), .C2(n1819), .ZN(register_file_inst1_n2267) );
  INVD1BWP12T U796 ( .I(register_file_inst1_r1_2_), .ZN(n1810) );
  OAI222D0BWP12T U797 ( .A1(n1810), .A2(n1093), .B1(n239), .B2(n1095), .C1(
        n2101), .C2(n1094), .ZN(register_file_inst1_n2587) );
  INVD1BWP12T U798 ( .I(register_file_inst1_r6_2_), .ZN(n1822) );
  OAI222D0BWP12T U799 ( .A1(n1822), .A2(n1045), .B1(n239), .B2(n1043), .C1(
        n2101), .C2(n1044), .ZN(register_file_inst1_n2427) );
  CKND1BWP12T U800 ( .I(register_file_inst1_r10_2_), .ZN(n1817) );
  OAI222D0BWP12T U801 ( .A1(n2101), .A2(n1069), .B1(n239), .B2(n1070), .C1(
        n1068), .C2(n1817), .ZN(register_file_inst1_n2299) );
  CKND0BWP12T U802 ( .I(register_file_inst1_r9_2_), .ZN(n238) );
  OAI222D0BWP12T U803 ( .A1(n238), .A2(n1079), .B1(n239), .B2(n1081), .C1(
        n2101), .C2(n1080), .ZN(register_file_inst1_n2331) );
  INVD1BWP12T U804 ( .I(register_file_inst1_r0_2_), .ZN(n1801) );
  OAI222D0BWP12T U805 ( .A1(n1801), .A2(n1086), .B1(n239), .B2(n1089), .C1(
        n2101), .C2(n1088), .ZN(register_file_inst1_n2619) );
  INVD1BWP12T U806 ( .I(ALU_MISC_OUT_result[12]), .ZN(n245) );
  CKND0BWP12T U807 ( .I(register_file_inst1_r2_12_), .ZN(n240) );
  OAI222D0BWP12T U808 ( .A1(n2126), .A2(n1062), .B1(n245), .B2(n1063), .C1(
        n1060), .C2(n240), .ZN(register_file_inst1_n2565) );
  INVD1BWP12T U809 ( .I(ALU_MISC_OUT_result[11]), .ZN(n247) );
  CKND0BWP12T U810 ( .I(register_file_inst1_r2_11_), .ZN(n241) );
  OAI222D0BWP12T U811 ( .A1(n2123), .A2(n1062), .B1(n247), .B2(n1063), .C1(
        n1060), .C2(n241), .ZN(register_file_inst1_n2564) );
  INVD1BWP12T U812 ( .I(register_file_inst1_r0_11_), .ZN(n1432) );
  OAI222D0BWP12T U813 ( .A1(n1432), .A2(n1086), .B1(n247), .B2(n1089), .C1(
        n2123), .C2(n1088), .ZN(register_file_inst1_n2628) );
  INVD1BWP12T U814 ( .I(register_file_inst1_r5_11_), .ZN(n1446) );
  OAI222D0BWP12T U815 ( .A1(n1446), .A2(n1096), .B1(n247), .B2(n1098), .C1(
        n2123), .C2(n1097), .ZN(register_file_inst1_n2468) );
  INVD1BWP12T U816 ( .I(ALU_MISC_OUT_result[13]), .ZN(n246) );
  INVD1BWP12T U817 ( .I(register_file_inst1_tmp1_13_), .ZN(n1294) );
  OAI222D0BWP12T U818 ( .A1(n2129), .A2(n1026), .B1(n246), .B2(n2168), .C1(
        n1027), .C2(n1294), .ZN(register_file_inst1_n2150) );
  CKND0BWP12T U819 ( .I(register_file_inst1_r2_13_), .ZN(n242) );
  OAI222D0BWP12T U820 ( .A1(n2129), .A2(n1062), .B1(n246), .B2(n1063), .C1(
        n1060), .C2(n242), .ZN(register_file_inst1_n2566) );
  INVD1BWP12T U821 ( .I(register_file_inst1_r9_11_), .ZN(n1420) );
  OAI222D0BWP12T U822 ( .A1(n1420), .A2(n1079), .B1(n247), .B2(n1081), .C1(
        n2123), .C2(n1080), .ZN(register_file_inst1_n2340) );
  INVD1BWP12T U823 ( .I(register_file_inst1_r0_13_), .ZN(n1278) );
  OAI222D0BWP12T U824 ( .A1(n1278), .A2(n1086), .B1(n246), .B2(n1089), .C1(
        n2129), .C2(n1088), .ZN(register_file_inst1_n2630) );
  INVD1BWP12T U825 ( .I(register_file_inst1_r9_12_), .ZN(n1325) );
  OAI222D0BWP12T U826 ( .A1(n1325), .A2(n1079), .B1(n245), .B2(n1081), .C1(
        n2126), .C2(n1080), .ZN(register_file_inst1_n2341) );
  INVD1BWP12T U827 ( .I(register_file_inst1_r11_13_), .ZN(n1291) );
  OAI222D0BWP12T U828 ( .A1(n2129), .A2(n964), .B1(n246), .B2(n1019), .C1(
        n1021), .C2(n1291), .ZN(register_file_inst1_n2278) );
  INVD1BWP12T U829 ( .I(register_file_inst1_r9_13_), .ZN(n1266) );
  OAI222D0BWP12T U830 ( .A1(n1266), .A2(n1079), .B1(n246), .B2(n1081), .C1(
        n2129), .C2(n1080), .ZN(register_file_inst1_n2342) );
  INVD1BWP12T U831 ( .I(register_file_inst1_r12_12_), .ZN(n1302) );
  OAI222D0BWP12T U832 ( .A1(n1302), .A2(n1071), .B1(n245), .B2(n1074), .C1(
        n2126), .C2(n1073), .ZN(register_file_inst1_n2245) );
  TPOAI21D0BWP12T U833 ( .A1(n245), .A2(n1104), .B(n2008), .ZN(
        register_file_inst1_spin[12]) );
  INVD1BWP12T U834 ( .I(register_file_inst1_tmp1_12_), .ZN(n1316) );
  OAI222D0BWP12T U835 ( .A1(n2126), .A2(n1026), .B1(n245), .B2(n2168), .C1(
        n1027), .C2(n1316), .ZN(register_file_inst1_n2149) );
  INVD1BWP12T U836 ( .I(register_file_inst1_r5_12_), .ZN(n1314) );
  OAI222D0BWP12T U837 ( .A1(n1314), .A2(n1096), .B1(n245), .B2(n1098), .C1(
        n2126), .C2(n1097), .ZN(register_file_inst1_n2469) );
  INVD1BWP12T U838 ( .I(register_file_inst1_r11_12_), .ZN(n1323) );
  OAI222D0BWP12T U839 ( .A1(n2126), .A2(n964), .B1(n245), .B2(n1019), .C1(
        n1021), .C2(n1323), .ZN(register_file_inst1_n2277) );
  INVD1BWP12T U840 ( .I(register_file_inst1_r6_11_), .ZN(n1447) );
  OAI222D0BWP12T U841 ( .A1(n1447), .A2(n1045), .B1(n247), .B2(n1043), .C1(
        n2123), .C2(n1044), .ZN(register_file_inst1_n2436) );
  INVD1BWP12T U842 ( .I(register_file_inst1_r11_11_), .ZN(n1445) );
  OAI222D0BWP12T U843 ( .A1(n2123), .A2(n1020), .B1(n247), .B2(n1019), .C1(
        n1021), .C2(n1445), .ZN(register_file_inst1_n2276) );
  INVD1BWP12T U844 ( .I(register_file_inst1_r0_12_), .ZN(n1303) );
  OAI222D0BWP12T U845 ( .A1(n1303), .A2(n1086), .B1(n245), .B2(n1089), .C1(
        n2126), .C2(n1088), .ZN(register_file_inst1_n2629) );
  INVD1BWP12T U846 ( .I(register_file_inst1_r12_11_), .ZN(n1431) );
  OAI222D0BWP12T U847 ( .A1(n1431), .A2(n1071), .B1(n247), .B2(n1074), .C1(
        n2123), .C2(n1073), .ZN(register_file_inst1_n2244) );
  INVD1BWP12T U848 ( .I(register_file_inst1_r6_12_), .ZN(n1315) );
  OAI222D0BWP12T U849 ( .A1(n1315), .A2(n1045), .B1(n245), .B2(n1043), .C1(
        n2126), .C2(n1044), .ZN(register_file_inst1_n2437) );
  INVD1BWP12T U850 ( .I(register_file_inst1_r6_13_), .ZN(n1293) );
  OAI222D0BWP12T U851 ( .A1(n1293), .A2(n1045), .B1(n246), .B2(n1043), .C1(
        n2129), .C2(n1044), .ZN(register_file_inst1_n2438) );
  INVD1BWP12T U852 ( .I(STACK_RF_next_sp[13]), .ZN(n1276) );
  OAI222D0BWP12T U853 ( .A1(n1276), .A2(n1037), .B1(n246), .B2(n1104), .C1(
        n2129), .C2(n1102), .ZN(register_file_inst1_spin[13]) );
  INVD1BWP12T U854 ( .I(register_file_inst1_r5_13_), .ZN(n1292) );
  OAI222D0BWP12T U855 ( .A1(n1292), .A2(n1096), .B1(n246), .B2(n1098), .C1(
        n2129), .C2(n1097), .ZN(register_file_inst1_n2470) );
  INVD1BWP12T U856 ( .I(register_file_inst1_r12_13_), .ZN(n1277) );
  OAI222D0BWP12T U857 ( .A1(n1277), .A2(n1071), .B1(n246), .B2(n1074), .C1(
        n2129), .C2(n1073), .ZN(register_file_inst1_n2246) );
  INVD1BWP12T U858 ( .I(register_file_inst1_r10_13_), .ZN(n1289) );
  OAI222D0BWP12T U859 ( .A1(n2129), .A2(n1069), .B1(n246), .B2(n1070), .C1(
        n1068), .C2(n1289), .ZN(register_file_inst1_n2310) );
  INVD1BWP12T U860 ( .I(register_file_inst1_lr_13_), .ZN(n1280) );
  OAI222D0BWP12T U861 ( .A1(n1280), .A2(n1082), .B1(n246), .B2(n1085), .C1(
        n2129), .C2(n1084), .ZN(register_file_inst1_n2214) );
  CKND0BWP12T U862 ( .I(register_file_inst1_r8_12_), .ZN(n243) );
  OAI222D0BWP12T U863 ( .A1(n243), .A2(n1075), .B1(n245), .B2(n1078), .C1(
        n2126), .C2(n1077), .ZN(register_file_inst1_n2373) );
  INVD1BWP12T U864 ( .I(register_file_inst1_r4_11_), .ZN(n1444) );
  OAI222D0BWP12T U865 ( .A1(n1444), .A2(n1090), .B1(n247), .B2(n1092), .C1(
        n2123), .C2(n1091), .ZN(register_file_inst1_n2500) );
  INVD1BWP12T U866 ( .I(register_file_inst1_r4_12_), .ZN(n1313) );
  OAI222D0BWP12T U867 ( .A1(n1313), .A2(n1090), .B1(n245), .B2(n1092), .C1(
        n2126), .C2(n1091), .ZN(register_file_inst1_n2501) );
  INVD1BWP12T U868 ( .I(register_file_inst1_r10_12_), .ZN(n1312) );
  OAI222D0BWP12T U869 ( .A1(n2126), .A2(n1069), .B1(n245), .B2(n1070), .C1(
        n1068), .C2(n1312), .ZN(register_file_inst1_n2309) );
  INVD1BWP12T U870 ( .I(register_file_inst1_lr_11_), .ZN(n1434) );
  OAI222D0BWP12T U871 ( .A1(n1434), .A2(n1082), .B1(n247), .B2(n1085), .C1(
        n2123), .C2(n1084), .ZN(register_file_inst1_n2212) );
  INVD1BWP12T U872 ( .I(register_file_inst1_r3_13_), .ZN(n1279) );
  OAI222D0BWP12T U873 ( .A1(n2129), .A2(n1066), .B1(n246), .B2(n1067), .C1(
        n1064), .C2(n1279), .ZN(register_file_inst1_n2534) );
  TPOAI21D0BWP12T U874 ( .A1(n247), .A2(n1104), .B(n2011), .ZN(
        register_file_inst1_spin[11]) );
  INVD1BWP12T U875 ( .I(register_file_inst1_r3_11_), .ZN(n1433) );
  OAI222D0BWP12T U876 ( .A1(n2123), .A2(n1066), .B1(n247), .B2(n1067), .C1(
        n1064), .C2(n1433), .ZN(register_file_inst1_n2532) );
  INVD1BWP12T U877 ( .I(register_file_inst1_r10_11_), .ZN(n1443) );
  OAI222D0BWP12T U878 ( .A1(n2123), .A2(n1069), .B1(n247), .B2(n1070), .C1(
        n1068), .C2(n1443), .ZN(register_file_inst1_n2308) );
  INVD1BWP12T U879 ( .I(register_file_inst1_r7_11_), .ZN(n1435) );
  OAI222D0BWP12T U880 ( .A1(n1435), .A2(n1051), .B1(n247), .B2(n1049), .C1(
        n2123), .C2(n1050), .ZN(register_file_inst1_n2404) );
  INVD1BWP12T U881 ( .I(register_file_inst1_r3_12_), .ZN(n1304) );
  OAI222D0BWP12T U882 ( .A1(n2126), .A2(n1066), .B1(n245), .B2(n1067), .C1(
        n1064), .C2(n1304), .ZN(register_file_inst1_n2533) );
  INVD1BWP12T U883 ( .I(register_file_inst1_lr_12_), .ZN(n1305) );
  OAI222D0BWP12T U884 ( .A1(n1305), .A2(n1082), .B1(n245), .B2(n1085), .C1(
        n2126), .C2(n1084), .ZN(register_file_inst1_n2213) );
  INVD1BWP12T U885 ( .I(register_file_inst1_r1_11_), .ZN(n1436) );
  OAI222D0BWP12T U886 ( .A1(n1436), .A2(n1093), .B1(n247), .B2(n1095), .C1(
        n2123), .C2(n1094), .ZN(register_file_inst1_n2596) );
  INVD1BWP12T U887 ( .I(register_file_inst1_tmp1_11_), .ZN(n1448) );
  OAI222D0BWP12T U888 ( .A1(n2123), .A2(n1026), .B1(n247), .B2(n2168), .C1(
        n1027), .C2(n1448), .ZN(register_file_inst1_n2148) );
  CKND0BWP12T U889 ( .I(register_file_inst1_r8_13_), .ZN(n244) );
  OAI222D0BWP12T U890 ( .A1(n244), .A2(n1075), .B1(n246), .B2(n1078), .C1(
        n2129), .C2(n1077), .ZN(register_file_inst1_n2374) );
  INVD1BWP12T U891 ( .I(register_file_inst1_r4_13_), .ZN(n1290) );
  OAI222D0BWP12T U892 ( .A1(n1290), .A2(n1090), .B1(n246), .B2(n1092), .C1(
        n2129), .C2(n1091), .ZN(register_file_inst1_n2502) );
  INVD1BWP12T U893 ( .I(register_file_inst1_r7_13_), .ZN(n1281) );
  OAI222D0BWP12T U894 ( .A1(n1281), .A2(n1051), .B1(n246), .B2(n1049), .C1(
        n2129), .C2(n1050), .ZN(register_file_inst1_n2406) );
  INVD1BWP12T U895 ( .I(register_file_inst1_r1_12_), .ZN(n1324) );
  OAI222D0BWP12T U896 ( .A1(n1324), .A2(n1093), .B1(n245), .B2(n1095), .C1(
        n2126), .C2(n1094), .ZN(register_file_inst1_n2597) );
  INVD1BWP12T U897 ( .I(register_file_inst1_r7_12_), .ZN(n1326) );
  OAI222D0BWP12T U898 ( .A1(n1326), .A2(n1051), .B1(n245), .B2(n1049), .C1(
        n2126), .C2(n1050), .ZN(register_file_inst1_n2405) );
  INVD1BWP12T U899 ( .I(register_file_inst1_r1_13_), .ZN(n1282) );
  OAI222D0BWP12T U900 ( .A1(n1282), .A2(n1093), .B1(n246), .B2(n1095), .C1(
        n2129), .C2(n1094), .ZN(register_file_inst1_n2598) );
  CKND0BWP12T U901 ( .I(register_file_inst1_r8_11_), .ZN(n248) );
  OAI222D0BWP12T U902 ( .A1(n248), .A2(n1075), .B1(n247), .B2(n1078), .C1(
        n2123), .C2(n1077), .ZN(register_file_inst1_n2372) );
  OAI222D0BWP12T U903 ( .A1(n2105), .A2(n1020), .B1(n257), .B2(n1019), .C1(
        n1021), .C2(n249), .ZN(register_file_inst1_n2269) );
  OAI222D0BWP12T U904 ( .A1(n250), .A2(n1051), .B1(n257), .B2(n1049), .C1(
        n2105), .C2(n1050), .ZN(register_file_inst1_n2397) );
  CKND0BWP12T U905 ( .I(register_file_inst1_r9_4_), .ZN(n251) );
  OAI222D0BWP12T U906 ( .A1(n251), .A2(n1079), .B1(n257), .B2(n1081), .C1(
        n2105), .C2(n1080), .ZN(register_file_inst1_n2333) );
  INVD1BWP12T U907 ( .I(register_file_inst1_r8_4_), .ZN(n1667) );
  OAI222D0BWP12T U908 ( .A1(n1667), .A2(n1075), .B1(n257), .B2(n1078), .C1(
        n2105), .C2(n1077), .ZN(register_file_inst1_n2365) );
  OAI222D0BWP12T U909 ( .A1(n1668), .A2(n1071), .B1(n257), .B2(n1074), .C1(
        n2105), .C2(n1073), .ZN(register_file_inst1_n2237) );
  TPOAI21D0BWP12T U910 ( .A1(n257), .A2(n1104), .B(n2029), .ZN(
        register_file_inst1_spin[4]) );
  OAI222D0BWP12T U911 ( .A1(n1671), .A2(n1082), .B1(n257), .B2(n1085), .C1(
        n2105), .C2(n1084), .ZN(register_file_inst1_n2205) );
  OAI222D0BWP12T U912 ( .A1(n2105), .A2(n1026), .B1(n257), .B2(n2168), .C1(
        n1027), .C2(n252), .ZN(register_file_inst1_n2141) );
  CKND0BWP12T U913 ( .I(register_file_inst1_r2_4_), .ZN(n253) );
  OAI222D0BWP12T U914 ( .A1(n2105), .A2(n1062), .B1(n257), .B2(n1063), .C1(
        n1060), .C2(n253), .ZN(register_file_inst1_n2557) );
  OAI222D0BWP12T U915 ( .A1(n1670), .A2(n1090), .B1(n257), .B2(n1092), .C1(
        n2105), .C2(n1091), .ZN(register_file_inst1_n2493) );
  OAI222D0BWP12T U916 ( .A1(n254), .A2(n1093), .B1(n257), .B2(n1095), .C1(
        n2105), .C2(n1094), .ZN(register_file_inst1_n2589) );
  OAI222D0BWP12T U917 ( .A1(n2105), .A2(n1066), .B1(n257), .B2(n1067), .C1(
        n1064), .C2(n1669), .ZN(register_file_inst1_n2525) );
  OAI222D0BWP12T U918 ( .A1(n255), .A2(n1086), .B1(n257), .B2(n1089), .C1(
        n2105), .C2(n1088), .ZN(register_file_inst1_n2621) );
  OAI222D0BWP12T U919 ( .A1(n256), .A2(n1096), .B1(n257), .B2(n1098), .C1(
        n2105), .C2(n1097), .ZN(register_file_inst1_n2461) );
  OAI222D0BWP12T U920 ( .A1(n1673), .A2(n1045), .B1(n257), .B2(n1043), .C1(
        n2105), .C2(n1044), .ZN(register_file_inst1_n2429) );
  INVD1BWP12T U921 ( .I(ALU_MISC_OUT_result[6]), .ZN(n271) );
  TPOAI21D0BWP12T U922 ( .A1(n271), .A2(n1104), .B(n2026), .ZN(
        register_file_inst1_spin[6]) );
  INVD1BWP12T U923 ( .I(register_file_inst1_r4_10_), .ZN(n455) );
  INVD1BWP12T U924 ( .I(ALU_MISC_OUT_result[10]), .ZN(n274) );
  OAI222D0BWP12T U925 ( .A1(n455), .A2(n1090), .B1(n274), .B2(n1092), .C1(
        n2120), .C2(n1091), .ZN(register_file_inst1_n2499) );
  INVD1BWP12T U926 ( .I(ALU_MISC_OUT_result[5]), .ZN(n275) );
  TPOAI21D0BWP12T U927 ( .A1(n275), .A2(n1104), .B(n1988), .ZN(
        register_file_inst1_spin[5]) );
  INVD1BWP12T U928 ( .I(ALU_MISC_OUT_result[7]), .ZN(n270) );
  INVD1BWP12T U929 ( .I(register_file_inst1_r11_7_), .ZN(n1516) );
  OAI222D0BWP12T U930 ( .A1(n2113), .A2(n1020), .B1(n270), .B2(n1019), .C1(
        n1021), .C2(n1516), .ZN(register_file_inst1_n2272) );
  INVD1BWP12T U931 ( .I(register_file_inst1_r7_3_), .ZN(n1754) );
  INVD1BWP12T U932 ( .I(ALU_MISC_OUT_result[3]), .ZN(n273) );
  OAI222D0BWP12T U933 ( .A1(n1754), .A2(n1051), .B1(n273), .B2(n1049), .C1(
        n2103), .C2(n1050), .ZN(register_file_inst1_n2396) );
  INVD1BWP12T U934 ( .I(register_file_inst1_tmp1_3_), .ZN(n1767) );
  OAI222D0BWP12T U935 ( .A1(n2103), .A2(n1026), .B1(n273), .B2(n2168), .C1(
        n1027), .C2(n1767), .ZN(register_file_inst1_n2140) );
  INVD1BWP12T U936 ( .I(register_file_inst1_r4_6_), .ZN(n1467) );
  OAI222D0BWP12T U937 ( .A1(n1467), .A2(n1090), .B1(n271), .B2(n1092), .C1(
        n2110), .C2(n1091), .ZN(register_file_inst1_n2495) );
  INVD1BWP12T U938 ( .I(register_file_inst1_r11_6_), .ZN(n1477) );
  OAI222D0BWP12T U939 ( .A1(n2110), .A2(n964), .B1(n271), .B2(n1019), .C1(
        n1021), .C2(n1477), .ZN(register_file_inst1_n2271) );
  CKND0BWP12T U940 ( .I(register_file_inst1_r8_10_), .ZN(n258) );
  OAI222D0BWP12T U941 ( .A1(n258), .A2(n1075), .B1(n274), .B2(n1078), .C1(
        n2120), .C2(n1077), .ZN(register_file_inst1_n2371) );
  CKND0BWP12T U942 ( .I(register_file_inst1_r8_9_), .ZN(n259) );
  INVD1BWP12T U943 ( .I(ALU_MISC_OUT_result[9]), .ZN(n272) );
  OAI222D0BWP12T U944 ( .A1(n259), .A2(n1075), .B1(n272), .B2(n1078), .C1(
        n2117), .C2(n1077), .ZN(register_file_inst1_n2370) );
  INVD1BWP12T U945 ( .I(register_file_inst1_r4_5_), .ZN(n1712) );
  OAI222D0BWP12T U946 ( .A1(n1712), .A2(n1090), .B1(n275), .B2(n1092), .C1(
        n2107), .C2(n1091), .ZN(register_file_inst1_n2494) );
  INVD1BWP12T U947 ( .I(register_file_inst1_r3_9_), .ZN(n1385) );
  OAI222D0BWP12T U948 ( .A1(n2117), .A2(n1066), .B1(n272), .B2(n1067), .C1(
        n1064), .C2(n1385), .ZN(register_file_inst1_n2530) );
  TPOAI21D0BWP12T U949 ( .A1(n274), .A2(n1104), .B(n2014), .ZN(
        register_file_inst1_spin[10]) );
  INVD1BWP12T U950 ( .I(register_file_inst1_r4_9_), .ZN(n1396) );
  OAI222D0BWP12T U951 ( .A1(n1396), .A2(n1090), .B1(n272), .B2(n1092), .C1(
        n2117), .C2(n1091), .ZN(register_file_inst1_n2498) );
  INVD1BWP12T U952 ( .I(register_file_inst1_r12_10_), .ZN(n444) );
  OAI222D0BWP12T U953 ( .A1(n444), .A2(n1071), .B1(n274), .B2(n1074), .C1(
        n2120), .C2(n1073), .ZN(register_file_inst1_n2243) );
  TPOAI21D0BWP12T U954 ( .A1(n270), .A2(n1104), .B(n2023), .ZN(
        register_file_inst1_spin[7]) );
  INVD1BWP12T U955 ( .I(register_file_inst1_r8_7_), .ZN(n1490) );
  OAI222D0BWP12T U956 ( .A1(n1490), .A2(n1075), .B1(n270), .B2(n1078), .C1(
        n2113), .C2(n1077), .ZN(register_file_inst1_n2368) );
  INVD1BWP12T U957 ( .I(register_file_inst1_r11_5_), .ZN(n1713) );
  OAI222D0BWP12T U958 ( .A1(n2107), .A2(n1020), .B1(n275), .B2(n1019), .C1(
        n1021), .C2(n1713), .ZN(register_file_inst1_n2270) );
  INVD1BWP12T U959 ( .I(register_file_inst1_r4_3_), .ZN(n1763) );
  OAI222D0BWP12T U960 ( .A1(n1763), .A2(n1090), .B1(n273), .B2(n1092), .C1(
        n2103), .C2(n1091), .ZN(register_file_inst1_n2492) );
  INVD1BWP12T U961 ( .I(register_file_inst1_r0_10_), .ZN(n445) );
  OAI222D0BWP12T U962 ( .A1(n445), .A2(n1086), .B1(n274), .B2(n1089), .C1(
        n2120), .C2(n1088), .ZN(register_file_inst1_n2627) );
  INVD1BWP12T U963 ( .I(register_file_inst1_r8_6_), .ZN(n260) );
  OAI222D0BWP12T U964 ( .A1(n260), .A2(n1075), .B1(n271), .B2(n1078), .C1(
        n2110), .C2(n1077), .ZN(register_file_inst1_n2367) );
  INVD1BWP12T U965 ( .I(register_file_inst1_r11_10_), .ZN(n1407) );
  OAI222D0BWP12T U966 ( .A1(n2120), .A2(n964), .B1(n274), .B2(n1019), .C1(
        n1021), .C2(n1407), .ZN(register_file_inst1_n2275) );
  INVD1BWP12T U967 ( .I(register_file_inst1_r0_9_), .ZN(n1384) );
  OAI222D0BWP12T U968 ( .A1(n1384), .A2(n1086), .B1(n272), .B2(n1089), .C1(
        n2117), .C2(n1088), .ZN(register_file_inst1_n2626) );
  TPOAI21D0BWP12T U969 ( .A1(n272), .A2(n1104), .B(n2017), .ZN(
        register_file_inst1_spin[9]) );
  INVD1BWP12T U970 ( .I(register_file_inst1_tmp1_5_), .ZN(n1716) );
  OAI222D0BWP12T U971 ( .A1(n2107), .A2(n1026), .B1(n275), .B2(n2168), .C1(
        n1027), .C2(n1716), .ZN(register_file_inst1_n2142) );
  INVD1BWP12T U972 ( .I(register_file_inst1_r6_5_), .ZN(n1715) );
  OAI222D0BWP12T U973 ( .A1(n1715), .A2(n1045), .B1(n275), .B2(n1043), .C1(
        n2107), .C2(n1044), .ZN(register_file_inst1_n2430) );
  CKND0BWP12T U974 ( .I(register_file_inst1_r8_5_), .ZN(n261) );
  OAI222D0BWP12T U975 ( .A1(n261), .A2(n1075), .B1(n275), .B2(n1078), .C1(
        n2107), .C2(n1077), .ZN(register_file_inst1_n2366) );
  INVD1BWP12T U976 ( .I(register_file_inst1_r4_7_), .ZN(n1515) );
  OAI222D0BWP12T U977 ( .A1(n1515), .A2(n1090), .B1(n270), .B2(n1092), .C1(
        n2113), .C2(n1091), .ZN(register_file_inst1_n2496) );
  CKND0BWP12T U978 ( .I(register_file_inst1_r2_10_), .ZN(n262) );
  OAI222D0BWP12T U979 ( .A1(n2120), .A2(n1062), .B1(n274), .B2(n1063), .C1(
        n1060), .C2(n262), .ZN(register_file_inst1_n2563) );
  INVD1BWP12T U980 ( .I(register_file_inst1_r0_7_), .ZN(n1503) );
  OAI222D0BWP12T U981 ( .A1(n1503), .A2(n1086), .B1(n270), .B2(n1089), .C1(
        n2113), .C2(n1088), .ZN(register_file_inst1_n2624) );
  INVD1BWP12T U982 ( .I(register_file_inst1_r11_9_), .ZN(n1397) );
  OAI222D0BWP12T U983 ( .A1(n2117), .A2(n1020), .B1(n272), .B2(n1019), .C1(
        n1021), .C2(n1397), .ZN(register_file_inst1_n2274) );
  INVD1BWP12T U984 ( .I(register_file_inst1_r8_3_), .ZN(n1723) );
  OAI222D0BWP12T U985 ( .A1(n1723), .A2(n1075), .B1(n273), .B2(n1078), .C1(
        n2103), .C2(n1077), .ZN(register_file_inst1_n2364) );
  INVD1BWP12T U986 ( .I(register_file_inst1_lr_10_), .ZN(n447) );
  OAI222D0BWP12T U987 ( .A1(n447), .A2(n1082), .B1(n274), .B2(n1085), .C1(
        n2120), .C2(n1084), .ZN(register_file_inst1_n2211) );
  INVD1BWP12T U988 ( .I(register_file_inst1_lr_9_), .ZN(n1386) );
  OAI222D0BWP12T U989 ( .A1(n1386), .A2(n1082), .B1(n272), .B2(n1085), .C1(
        n2117), .C2(n1084), .ZN(register_file_inst1_n2210) );
  INVD1BWP12T U990 ( .I(register_file_inst1_r0_6_), .ZN(n1457) );
  OAI222D0BWP12T U991 ( .A1(n1457), .A2(n1086), .B1(n271), .B2(n1089), .C1(
        n2110), .C2(n1088), .ZN(register_file_inst1_n2623) );
  INVD1BWP12T U992 ( .I(register_file_inst1_r0_5_), .ZN(n1700) );
  OAI222D0BWP12T U993 ( .A1(n1700), .A2(n1086), .B1(n275), .B2(n1089), .C1(
        n2107), .C2(n1088), .ZN(register_file_inst1_n2622) );
  INVD1BWP12T U994 ( .I(register_file_inst1_r3_3_), .ZN(n1752) );
  OAI222D0BWP12T U995 ( .A1(n2103), .A2(n1066), .B1(n273), .B2(n1067), .C1(
        n1064), .C2(n1752), .ZN(register_file_inst1_n2524) );
  TPOAI21D0BWP12T U996 ( .A1(n273), .A2(n1104), .B(n2032), .ZN(
        register_file_inst1_spin[3]) );
  INVD1BWP12T U997 ( .I(register_file_inst1_r11_3_), .ZN(n1764) );
  OAI222D0BWP12T U998 ( .A1(n2103), .A2(n964), .B1(n273), .B2(n1019), .C1(
        n1021), .C2(n1764), .ZN(register_file_inst1_n2268) );
  INVD1BWP12T U999 ( .I(register_file_inst1_tmp1_6_), .ZN(n1470) );
  OAI222D0BWP12T U1000 ( .A1(n2110), .A2(n1026), .B1(n271), .B2(n2168), .C1(
        n1027), .C2(n1470), .ZN(register_file_inst1_n2143) );
  INVD1BWP12T U1001 ( .I(register_file_inst1_r3_5_), .ZN(n1701) );
  OAI222D0BWP12T U1002 ( .A1(n2107), .A2(n1066), .B1(n275), .B2(n1067), .C1(
        n1064), .C2(n1701), .ZN(register_file_inst1_n2526) );
  INVD1BWP12T U1003 ( .I(register_file_inst1_lr_7_), .ZN(n1505) );
  OAI222D0BWP12T U1004 ( .A1(n1505), .A2(n1082), .B1(n270), .B2(n1085), .C1(
        n2113), .C2(n1084), .ZN(register_file_inst1_n2208) );
  INVD1BWP12T U1005 ( .I(register_file_inst1_r3_6_), .ZN(n1458) );
  OAI222D0BWP12T U1006 ( .A1(n2110), .A2(n1066), .B1(n271), .B2(n1067), .C1(
        n1064), .C2(n1458), .ZN(register_file_inst1_n2527) );
  INVD1BWP12T U1007 ( .I(register_file_inst1_r0_3_), .ZN(n1751) );
  OAI222D0BWP12T U1008 ( .A1(n1751), .A2(n1086), .B1(n273), .B2(n1089), .C1(
        n2103), .C2(n1088), .ZN(register_file_inst1_n2620) );
  INVD1BWP12T U1009 ( .I(register_file_inst1_tmp1_7_), .ZN(n1519) );
  OAI222D0BWP12T U1010 ( .A1(n2113), .A2(n1026), .B1(n270), .B2(n2168), .C1(
        n1027), .C2(n1519), .ZN(register_file_inst1_n2144) );
  INVD1BWP12T U1011 ( .I(register_file_inst1_r3_7_), .ZN(n1504) );
  OAI222D0BWP12T U1012 ( .A1(n2113), .A2(n1066), .B1(n270), .B2(n1067), .C1(
        n1064), .C2(n1504), .ZN(register_file_inst1_n2528) );
  INVD1BWP12T U1013 ( .I(register_file_inst1_r10_3_), .ZN(n1762) );
  OAI222D0BWP12T U1014 ( .A1(n2103), .A2(n1069), .B1(n273), .B2(n1070), .C1(
        n1068), .C2(n1762), .ZN(register_file_inst1_n2300) );
  INVD1BWP12T U1015 ( .I(register_file_inst1_r3_10_), .ZN(n446) );
  OAI222D0BWP12T U1016 ( .A1(n2120), .A2(n1066), .B1(n274), .B2(n1067), .C1(
        n1064), .C2(n446), .ZN(register_file_inst1_n2531) );
  INVD1BWP12T U1017 ( .I(register_file_inst1_r10_5_), .ZN(n1711) );
  OAI222D0BWP12T U1018 ( .A1(n2107), .A2(n1069), .B1(n275), .B2(n1070), .C1(
        n1068), .C2(n1711), .ZN(register_file_inst1_n2302) );
  INVD1BWP12T U1019 ( .I(register_file_inst1_lr_6_), .ZN(n1459) );
  OAI222D0BWP12T U1020 ( .A1(n1459), .A2(n1082), .B1(n271), .B2(n1085), .C1(
        n2110), .C2(n1084), .ZN(register_file_inst1_n2207) );
  INVD1BWP12T U1021 ( .I(register_file_inst1_lr_5_), .ZN(n1702) );
  OAI222D0BWP12T U1022 ( .A1(n1702), .A2(n1082), .B1(n275), .B2(n1085), .C1(
        n2107), .C2(n1084), .ZN(register_file_inst1_n2206) );
  INVD1BWP12T U1023 ( .I(register_file_inst1_r10_6_), .ZN(n1466) );
  OAI222D0BWP12T U1024 ( .A1(n2110), .A2(n1069), .B1(n271), .B2(n1070), .C1(
        n1068), .C2(n1466), .ZN(register_file_inst1_n2303) );
  INVD1BWP12T U1025 ( .I(register_file_inst1_lr_3_), .ZN(n1753) );
  OAI222D0BWP12T U1026 ( .A1(n1753), .A2(n1082), .B1(n273), .B2(n1085), .C1(
        n2103), .C2(n1084), .ZN(register_file_inst1_n2204) );
  INVD1BWP12T U1027 ( .I(register_file_inst1_r10_7_), .ZN(n1514) );
  OAI222D0BWP12T U1028 ( .A1(n2113), .A2(n1069), .B1(n270), .B2(n1070), .C1(
        n1068), .C2(n1514), .ZN(register_file_inst1_n2304) );
  INVD1BWP12T U1029 ( .I(register_file_inst1_tmp1_9_), .ZN(n1400) );
  OAI222D0BWP12T U1030 ( .A1(n2117), .A2(n1026), .B1(n272), .B2(n2168), .C1(
        n1027), .C2(n1400), .ZN(register_file_inst1_n2146) );
  INVD1BWP12T U1031 ( .I(register_file_inst1_r10_9_), .ZN(n1395) );
  OAI222D0BWP12T U1032 ( .A1(n2117), .A2(n1069), .B1(n272), .B2(n1070), .C1(
        n1068), .C2(n1395), .ZN(register_file_inst1_n2306) );
  INVD1BWP12T U1033 ( .I(register_file_inst1_r10_10_), .ZN(n454) );
  OAI222D0BWP12T U1034 ( .A1(n2120), .A2(n1069), .B1(n274), .B2(n1070), .C1(
        n1068), .C2(n454), .ZN(register_file_inst1_n2307) );
  INVD1BWP12T U1035 ( .I(register_file_inst1_r9_10_), .ZN(n1409) );
  OAI222D0BWP12T U1036 ( .A1(n1409), .A2(n1079), .B1(n274), .B2(n1081), .C1(
        n2120), .C2(n1080), .ZN(register_file_inst1_n2339) );
  INVD1BWP12T U1037 ( .I(register_file_inst1_tmp1_10_), .ZN(n458) );
  OAI222D0BWP12T U1038 ( .A1(n2120), .A2(n1026), .B1(n274), .B2(n2168), .C1(
        n1027), .C2(n458), .ZN(register_file_inst1_n2147) );
  INVD1BWP12T U1039 ( .I(register_file_inst1_r9_9_), .ZN(n1372) );
  OAI222D0BWP12T U1040 ( .A1(n1372), .A2(n1079), .B1(n272), .B2(n1081), .C1(
        n2117), .C2(n1080), .ZN(register_file_inst1_n2338) );
  CKND0BWP12T U1041 ( .I(register_file_inst1_r9_7_), .ZN(n263) );
  OAI222D0BWP12T U1042 ( .A1(n263), .A2(n1079), .B1(n270), .B2(n1081), .C1(
        n2113), .C2(n1080), .ZN(register_file_inst1_n2336) );
  INVD1BWP12T U1043 ( .I(register_file_inst1_r9_6_), .ZN(n1479) );
  OAI222D0BWP12T U1044 ( .A1(n1479), .A2(n1079), .B1(n271), .B2(n1081), .C1(
        n2110), .C2(n1080), .ZN(register_file_inst1_n2335) );
  INVD1BWP12T U1045 ( .I(register_file_inst1_r1_10_), .ZN(n1408) );
  OAI222D0BWP12T U1046 ( .A1(n1408), .A2(n1093), .B1(n274), .B2(n1095), .C1(
        n2120), .C2(n1094), .ZN(register_file_inst1_n2595) );
  INVD1BWP12T U1047 ( .I(register_file_inst1_r9_5_), .ZN(n1656) );
  OAI222D0BWP12T U1048 ( .A1(n1656), .A2(n1079), .B1(n275), .B2(n1081), .C1(
        n2107), .C2(n1080), .ZN(register_file_inst1_n2334) );
  CKND0BWP12T U1049 ( .I(register_file_inst1_r2_3_), .ZN(n264) );
  OAI222D0BWP12T U1050 ( .A1(n2103), .A2(n1062), .B1(n273), .B2(n1063), .C1(
        n1060), .C2(n264), .ZN(register_file_inst1_n2556) );
  INVD1BWP12T U1051 ( .I(register_file_inst1_r1_9_), .ZN(n1388) );
  OAI222D0BWP12T U1052 ( .A1(n1388), .A2(n1093), .B1(n272), .B2(n1095), .C1(
        n2117), .C2(n1094), .ZN(register_file_inst1_n2594) );
  INVD1BWP12T U1053 ( .I(register_file_inst1_r1_7_), .ZN(n1507) );
  OAI222D0BWP12T U1054 ( .A1(n1507), .A2(n1093), .B1(n270), .B2(n1095), .C1(
        n2113), .C2(n1094), .ZN(register_file_inst1_n2592) );
  INVD1BWP12T U1055 ( .I(register_file_inst1_r1_6_), .ZN(n1478) );
  OAI222D0BWP12T U1056 ( .A1(n1478), .A2(n1093), .B1(n271), .B2(n1095), .C1(
        n2110), .C2(n1094), .ZN(register_file_inst1_n2591) );
  CKND0BWP12T U1057 ( .I(register_file_inst1_r2_5_), .ZN(n265) );
  OAI222D0BWP12T U1058 ( .A1(n2107), .A2(n1062), .B1(n275), .B2(n1063), .C1(
        n1060), .C2(n265), .ZN(register_file_inst1_n2558) );
  INVD1BWP12T U1059 ( .I(register_file_inst1_r1_5_), .ZN(n1704) );
  OAI222D0BWP12T U1060 ( .A1(n1704), .A2(n1093), .B1(n275), .B2(n1095), .C1(
        n2107), .C2(n1094), .ZN(register_file_inst1_n2590) );
  CKND0BWP12T U1061 ( .I(register_file_inst1_r9_3_), .ZN(n266) );
  OAI222D0BWP12T U1062 ( .A1(n266), .A2(n1079), .B1(n273), .B2(n1081), .C1(
        n2103), .C2(n1080), .ZN(register_file_inst1_n2332) );
  INVD1BWP12T U1063 ( .I(register_file_inst1_r1_3_), .ZN(n1755) );
  OAI222D0BWP12T U1064 ( .A1(n1755), .A2(n1093), .B1(n273), .B2(n1095), .C1(
        n2103), .C2(n1094), .ZN(register_file_inst1_n2588) );
  INVD1BWP12T U1065 ( .I(register_file_inst1_r2_6_), .ZN(n267) );
  OAI222D0BWP12T U1066 ( .A1(n2110), .A2(n1062), .B1(n271), .B2(n1063), .C1(
        n1060), .C2(n267), .ZN(register_file_inst1_n2559) );
  CKND0BWP12T U1067 ( .I(register_file_inst1_r2_7_), .ZN(n268) );
  OAI222D0BWP12T U1068 ( .A1(n2113), .A2(n1062), .B1(n270), .B2(n1063), .C1(
        n1060), .C2(n268), .ZN(register_file_inst1_n2560) );
  CKND0BWP12T U1069 ( .I(register_file_inst1_r2_9_), .ZN(n269) );
  OAI222D0BWP12T U1070 ( .A1(n2117), .A2(n1062), .B1(n272), .B2(n1063), .C1(
        n1060), .C2(n269), .ZN(register_file_inst1_n2562) );
  INVD1BWP12T U1071 ( .I(register_file_inst1_r12_9_), .ZN(n1383) );
  OAI222D0BWP12T U1072 ( .A1(n1383), .A2(n1071), .B1(n272), .B2(n1074), .C1(
        n2117), .C2(n1073), .ZN(register_file_inst1_n2242) );
  INVD1BWP12T U1073 ( .I(register_file_inst1_r12_6_), .ZN(n1456) );
  OAI222D0BWP12T U1074 ( .A1(n1456), .A2(n1071), .B1(n271), .B2(n1074), .C1(
        n2110), .C2(n1073), .ZN(register_file_inst1_n2239) );
  INVD1BWP12T U1075 ( .I(register_file_inst1_r12_7_), .ZN(n1502) );
  OAI222D0BWP12T U1076 ( .A1(n1502), .A2(n1071), .B1(n270), .B2(n1074), .C1(
        n2113), .C2(n1073), .ZN(register_file_inst1_n2240) );
  INVD1BWP12T U1077 ( .I(register_file_inst1_r6_7_), .ZN(n1518) );
  OAI222D0BWP12T U1078 ( .A1(n1518), .A2(n1045), .B1(n270), .B2(n1043), .C1(
        n2113), .C2(n1044), .ZN(register_file_inst1_n2432) );
  INVD1BWP12T U1079 ( .I(register_file_inst1_r6_9_), .ZN(n1399) );
  OAI222D0BWP12T U1080 ( .A1(n1399), .A2(n1045), .B1(n272), .B2(n1043), .C1(
        n2117), .C2(n1044), .ZN(register_file_inst1_n2434) );
  INVD1BWP12T U1081 ( .I(register_file_inst1_r5_3_), .ZN(n1765) );
  OAI222D0BWP12T U1082 ( .A1(n1765), .A2(n1096), .B1(n273), .B2(n1098), .C1(
        n2103), .C2(n1097), .ZN(register_file_inst1_n2460) );
  INVD1BWP12T U1083 ( .I(register_file_inst1_r7_9_), .ZN(n1387) );
  OAI222D0BWP12T U1084 ( .A1(n1387), .A2(n1051), .B1(n272), .B2(n1049), .C1(
        n2117), .C2(n1050), .ZN(register_file_inst1_n2402) );
  INVD1BWP12T U1085 ( .I(register_file_inst1_r6_10_), .ZN(n457) );
  OAI222D0BWP12T U1086 ( .A1(n457), .A2(n1045), .B1(n274), .B2(n1043), .C1(
        n2120), .C2(n1044), .ZN(register_file_inst1_n2435) );
  INVD1BWP12T U1087 ( .I(register_file_inst1_r7_7_), .ZN(n1506) );
  OAI222D0BWP12T U1088 ( .A1(n1506), .A2(n1051), .B1(n270), .B2(n1049), .C1(
        n2113), .C2(n1050), .ZN(register_file_inst1_n2400) );
  INVD1BWP12T U1089 ( .I(register_file_inst1_r5_7_), .ZN(n1517) );
  OAI222D0BWP12T U1090 ( .A1(n1517), .A2(n1096), .B1(n270), .B2(n1098), .C1(
        n2113), .C2(n1097), .ZN(register_file_inst1_n2464) );
  INVD1BWP12T U1091 ( .I(register_file_inst1_r7_6_), .ZN(n1480) );
  OAI222D0BWP12T U1092 ( .A1(n1480), .A2(n1051), .B1(n271), .B2(n1049), .C1(
        n2110), .C2(n1050), .ZN(register_file_inst1_n2399) );
  INVD1BWP12T U1093 ( .I(register_file_inst1_r6_6_), .ZN(n1469) );
  OAI222D0BWP12T U1094 ( .A1(n1469), .A2(n1045), .B1(n271), .B2(n1043), .C1(
        n2110), .C2(n1044), .ZN(register_file_inst1_n2431) );
  OAI222D0BWP12T U1095 ( .A1(n1703), .A2(n1051), .B1(n275), .B2(n1049), .C1(
        n2107), .C2(n1050), .ZN(register_file_inst1_n2398) );
  INVD1BWP12T U1096 ( .I(register_file_inst1_r5_6_), .ZN(n1468) );
  OAI222D0BWP12T U1097 ( .A1(n1468), .A2(n1096), .B1(n271), .B2(n1098), .C1(
        n2110), .C2(n1097), .ZN(register_file_inst1_n2463) );
  INVD1BWP12T U1098 ( .I(register_file_inst1_r12_3_), .ZN(n1750) );
  OAI222D0BWP12T U1099 ( .A1(n1750), .A2(n1071), .B1(n273), .B2(n1074), .C1(
        n2103), .C2(n1073), .ZN(register_file_inst1_n2236) );
  INVD1BWP12T U1100 ( .I(register_file_inst1_r12_5_), .ZN(n1699) );
  OAI222D0BWP12T U1101 ( .A1(n1699), .A2(n1071), .B1(n275), .B2(n1074), .C1(
        n2107), .C2(n1073), .ZN(register_file_inst1_n2238) );
  INVD1BWP12T U1102 ( .I(register_file_inst1_r5_9_), .ZN(n1398) );
  OAI222D0BWP12T U1103 ( .A1(n1398), .A2(n1096), .B1(n272), .B2(n1098), .C1(
        n2117), .C2(n1097), .ZN(register_file_inst1_n2466) );
  INVD1BWP12T U1104 ( .I(register_file_inst1_r7_10_), .ZN(n1410) );
  OAI222D0BWP12T U1105 ( .A1(n1410), .A2(n1051), .B1(n274), .B2(n1049), .C1(
        n2120), .C2(n1050), .ZN(register_file_inst1_n2403) );
  INVD1BWP12T U1106 ( .I(register_file_inst1_r6_3_), .ZN(n1766) );
  OAI222D0BWP12T U1107 ( .A1(n1766), .A2(n1045), .B1(n273), .B2(n1043), .C1(
        n2103), .C2(n1044), .ZN(register_file_inst1_n2428) );
  INVD1BWP12T U1108 ( .I(register_file_inst1_r5_10_), .ZN(n456) );
  OAI222D0BWP12T U1109 ( .A1(n456), .A2(n1096), .B1(n274), .B2(n1098), .C1(
        n2120), .C2(n1097), .ZN(register_file_inst1_n2467) );
  INVD1BWP12T U1110 ( .I(register_file_inst1_r5_5_), .ZN(n1714) );
  OAI222D0BWP12T U1111 ( .A1(n1714), .A2(n1096), .B1(n275), .B2(n1098), .C1(
        n2107), .C2(n1097), .ZN(register_file_inst1_n2462) );
  INVD1BWP12T U1112 ( .I(register_file_inst1_r4_0_), .ZN(n1855) );
  INVD1BWP12T U1113 ( .I(ALU_MISC_OUT_result[0]), .ZN(n279) );
  OAI222D0BWP12T U1114 ( .A1(n1855), .A2(n1090), .B1(n279), .B2(n1092), .C1(
        n2085), .C2(n1091), .ZN(register_file_inst1_n2489) );
  INVD1BWP12T U1115 ( .I(register_file_inst1_r9_0_), .ZN(n1876) );
  OAI222D0BWP12T U1116 ( .A1(n1876), .A2(n1079), .B1(n279), .B2(n1081), .C1(
        n2085), .C2(n1080), .ZN(register_file_inst1_n2329) );
  INVD1BWP12T U1117 ( .I(register_file_inst1_r12_8_), .ZN(n1356) );
  INVD1BWP12T U1118 ( .I(ALU_MISC_OUT_result[8]), .ZN(n280) );
  OAI222D0BWP12T U1119 ( .A1(n1356), .A2(n1071), .B1(n280), .B2(n1074), .C1(
        n2115), .C2(n1073), .ZN(register_file_inst1_n2241) );
  INVD1BWP12T U1120 ( .I(register_file_inst1_r11_8_), .ZN(n1346) );
  OAI222D0BWP12T U1121 ( .A1(n2115), .A2(n964), .B1(n280), .B2(n1019), .C1(
        n1021), .C2(n1346), .ZN(register_file_inst1_n2273) );
  INVD1BWP12T U1122 ( .I(register_file_inst1_r7_0_), .ZN(n1878) );
  OAI222D0BWP12T U1123 ( .A1(n1878), .A2(n1051), .B1(n279), .B2(n1049), .C1(
        n2085), .C2(n1050), .ZN(register_file_inst1_n2393) );
  INVD1BWP12T U1124 ( .I(register_file_inst1_r3_8_), .ZN(n1357) );
  OAI222D0BWP12T U1125 ( .A1(n2115), .A2(n1066), .B1(n280), .B2(n1067), .C1(
        n1064), .C2(n1357), .ZN(register_file_inst1_n2529) );
  INVD1BWP12T U1126 ( .I(register_file_inst1_r12_0_), .ZN(n1851) );
  OAI222D0BWP12T U1127 ( .A1(n1851), .A2(n1071), .B1(n279), .B2(n1074), .C1(
        n2085), .C2(n1073), .ZN(register_file_inst1_n2233) );
  CKND0BWP12T U1128 ( .I(register_file_inst1_r2_8_), .ZN(n276) );
  OAI222D0BWP12T U1129 ( .A1(n2115), .A2(n1062), .B1(n280), .B2(n1063), .C1(
        n1060), .C2(n276), .ZN(register_file_inst1_n2561) );
  CKND0BWP12T U1130 ( .I(register_file_inst1_r9_8_), .ZN(n277) );
  OAI222D0BWP12T U1131 ( .A1(n277), .A2(n1079), .B1(n280), .B2(n1081), .C1(
        n2115), .C2(n1080), .ZN(register_file_inst1_n2337) );
  INVD1BWP12T U1132 ( .I(register_file_inst1_r0_8_), .ZN(n1337) );
  OAI222D0BWP12T U1133 ( .A1(n1337), .A2(n1086), .B1(n280), .B2(n1089), .C1(
        n2115), .C2(n1088), .ZN(register_file_inst1_n2625) );
  INVD1BWP12T U1134 ( .I(register_file_inst1_r7_8_), .ZN(n1338) );
  OAI222D0BWP12T U1135 ( .A1(n1338), .A2(n1051), .B1(n280), .B2(n1049), .C1(
        n2115), .C2(n1050), .ZN(register_file_inst1_n2401) );
  INVD1BWP12T U1136 ( .I(register_file_inst1_r6_0_), .ZN(n1862) );
  OAI222D0BWP12T U1137 ( .A1(n1862), .A2(n1045), .B1(n279), .B2(n1043), .C1(
        n2085), .C2(n1044), .ZN(register_file_inst1_n2425) );
  CKND0BWP12T U1138 ( .I(register_file_inst1_r2_0_), .ZN(n278) );
  OAI222D0BWP12T U1139 ( .A1(n2085), .A2(n1062), .B1(n279), .B2(n1063), .C1(
        n1060), .C2(n278), .ZN(register_file_inst1_n2553) );
  INVD1BWP12T U1140 ( .I(register_file_inst1_lr_8_), .ZN(n1359) );
  OAI222D0BWP12T U1141 ( .A1(n1359), .A2(n1082), .B1(n280), .B2(n1085), .C1(
        n2115), .C2(n1084), .ZN(register_file_inst1_n2209) );
  INVD1BWP12T U1142 ( .I(register_file_inst1_r1_8_), .ZN(n1339) );
  OAI222D0BWP12T U1143 ( .A1(n1339), .A2(n1093), .B1(n280), .B2(n1095), .C1(
        n2115), .C2(n1094), .ZN(register_file_inst1_n2593) );
  INVD1BWP12T U1144 ( .I(register_file_inst1_lr_0_), .ZN(n1857) );
  OAI222D0BWP12T U1145 ( .A1(n1857), .A2(n1082), .B1(n279), .B2(n1085), .C1(
        n2085), .C2(n1084), .ZN(register_file_inst1_n2201) );
  INVD1BWP12T U1146 ( .I(register_file_inst1_r11_0_), .ZN(n1872) );
  OAI222D0BWP12T U1147 ( .A1(n2085), .A2(n964), .B1(n279), .B2(n1019), .C1(
        n1021), .C2(n1872), .ZN(register_file_inst1_n2265) );
  INVD1BWP12T U1148 ( .I(register_file_inst1_r8_0_), .ZN(n1849) );
  OAI222D0BWP12T U1149 ( .A1(n1849), .A2(n1075), .B1(n279), .B2(n1078), .C1(
        n2085), .C2(n1077), .ZN(register_file_inst1_n2361) );
  INVD1BWP12T U1150 ( .I(register_file_inst1_r1_0_), .ZN(n1874) );
  OAI222D0BWP12T U1151 ( .A1(n1874), .A2(n1093), .B1(n279), .B2(n1095), .C1(
        n2085), .C2(n1094), .ZN(register_file_inst1_n2585) );
  INVD1BWP12T U1152 ( .I(register_file_inst1_r0_0_), .ZN(n1880) );
  OAI222D0BWP12T U1153 ( .A1(n1880), .A2(n1086), .B1(n279), .B2(n1089), .C1(
        n2085), .C2(n1088), .ZN(register_file_inst1_n2617) );
  INVD1BWP12T U1154 ( .I(register_file_inst1_r5_0_), .ZN(n1691) );
  OAI222D0BWP12T U1155 ( .A1(n1691), .A2(n1096), .B1(n279), .B2(n1098), .C1(
        n2085), .C2(n1097), .ZN(register_file_inst1_n2457) );
  INVD1BWP12T U1156 ( .I(STACK_RF_next_sp[0]), .ZN(n1684) );
  OAI222D0BWP12T U1157 ( .A1(n1684), .A2(n1099), .B1(n279), .B2(n1104), .C1(
        n2085), .C2(n1102), .ZN(register_file_inst1_spin[0]) );
  INVD1BWP12T U1158 ( .I(register_file_inst1_tmp1_0_), .ZN(n1881) );
  OAI222D0BWP12T U1159 ( .A1(n2085), .A2(n1026), .B1(n279), .B2(n2168), .C1(
        n1027), .C2(n1881), .ZN(register_file_inst1_n2136) );
  INVD1BWP12T U1160 ( .I(register_file_inst1_r3_0_), .ZN(n1853) );
  OAI222D0BWP12T U1161 ( .A1(n2085), .A2(n1066), .B1(n279), .B2(n1067), .C1(
        n1064), .C2(n1853), .ZN(register_file_inst1_n2521) );
  INVD1BWP12T U1162 ( .I(register_file_inst1_r8_8_), .ZN(n1355) );
  OAI222D0BWP12T U1163 ( .A1(n1355), .A2(n1075), .B1(n280), .B2(n1078), .C1(
        n2115), .C2(n1077), .ZN(register_file_inst1_n2369) );
  INVD1BWP12T U1164 ( .I(register_file_inst1_r10_0_), .ZN(n1860) );
  OAI222D0BWP12T U1165 ( .A1(n2085), .A2(n1069), .B1(n279), .B2(n1070), .C1(
        n1068), .C2(n1860), .ZN(register_file_inst1_n2297) );
  INVD1BWP12T U1166 ( .I(register_file_inst1_r4_8_), .ZN(n1358) );
  OAI222D0BWP12T U1167 ( .A1(n1358), .A2(n1090), .B1(n280), .B2(n1092), .C1(
        n2115), .C2(n1091), .ZN(register_file_inst1_n2497) );
  INVD1BWP12T U1168 ( .I(register_file_inst1_r6_8_), .ZN(n1361) );
  OAI222D0BWP12T U1169 ( .A1(n1361), .A2(n1045), .B1(n280), .B2(n1043), .C1(
        n2115), .C2(n1044), .ZN(register_file_inst1_n2433) );
  INVD1BWP12T U1170 ( .I(register_file_inst1_r5_8_), .ZN(n1347) );
  OAI222D0BWP12T U1171 ( .A1(n1347), .A2(n1096), .B1(n280), .B2(n1098), .C1(
        n2115), .C2(n1097), .ZN(register_file_inst1_n2465) );
  INVD1BWP12T U1172 ( .I(register_file_inst1_tmp1_8_), .ZN(n1348) );
  OAI222D0BWP12T U1173 ( .A1(n2115), .A2(n1026), .B1(n280), .B2(n2168), .C1(
        n1027), .C2(n1348), .ZN(register_file_inst1_n2145) );
  TPOAI21D0BWP12T U1174 ( .A1(n280), .A2(n1104), .B(n2020), .ZN(
        register_file_inst1_spin[8]) );
  INVD1BWP12T U1175 ( .I(register_file_inst1_r10_8_), .ZN(n1360) );
  OAI222D0BWP12T U1176 ( .A1(n2115), .A2(n1069), .B1(n280), .B2(n1070), .C1(
        n1068), .C2(n1360), .ZN(register_file_inst1_n2305) );
  INVD1BWP12T U1177 ( .I(ALU_MISC_OUT_result[1]), .ZN(n283) );
  INVD1BWP12T U1178 ( .I(register_file_inst1_r10_1_), .ZN(n1785) );
  OAI222D0BWP12T U1179 ( .A1(n2098), .A2(n1069), .B1(n283), .B2(n1070), .C1(
        n1068), .C2(n1785), .ZN(register_file_inst1_n2298) );
  INVD1BWP12T U1180 ( .I(register_file_inst1_r9_1_), .ZN(n1833) );
  OAI222D0BWP12T U1181 ( .A1(n1833), .A2(n1079), .B1(n283), .B2(n1081), .C1(
        n2098), .C2(n1080), .ZN(register_file_inst1_n2330) );
  INVD1BWP12T U1182 ( .I(register_file_inst1_r0_1_), .ZN(n1776) );
  OAI222D0BWP12T U1183 ( .A1(n1776), .A2(n1086), .B1(n283), .B2(n1089), .C1(
        n2098), .C2(n1088), .ZN(register_file_inst1_n2618) );
  INVD1BWP12T U1184 ( .I(register_file_inst1_r6_1_), .ZN(n1788) );
  OAI222D0BWP12T U1185 ( .A1(n1788), .A2(n1045), .B1(n283), .B2(n1043), .C1(
        n2098), .C2(n1044), .ZN(register_file_inst1_n2426) );
  INVD1BWP12T U1186 ( .I(register_file_inst1_r12_1_), .ZN(n1775) );
  OAI222D0BWP12T U1187 ( .A1(n1775), .A2(n1071), .B1(n283), .B2(n1074), .C1(
        n2098), .C2(n1073), .ZN(register_file_inst1_n2234) );
  INVD1BWP12T U1188 ( .I(register_file_inst1_r4_1_), .ZN(n1786) );
  OAI222D0BWP12T U1189 ( .A1(n1786), .A2(n1090), .B1(n283), .B2(n1092), .C1(
        n2098), .C2(n1091), .ZN(register_file_inst1_n2490) );
  INVD1BWP12T U1190 ( .I(register_file_inst1_r3_1_), .ZN(n1777) );
  OAI222D0BWP12T U1191 ( .A1(n2098), .A2(n1066), .B1(n283), .B2(n1067), .C1(
        n1064), .C2(n1777), .ZN(register_file_inst1_n2522) );
  INVD1BWP12T U1192 ( .I(register_file_inst1_tmp1_1_), .ZN(n1789) );
  OAI222D0BWP12T U1193 ( .A1(n2098), .A2(n1026), .B1(n283), .B2(n2168), .C1(
        n1027), .C2(n1789), .ZN(register_file_inst1_n2138) );
  INVD1BWP12T U1194 ( .I(register_file_inst1_r7_1_), .ZN(n1834) );
  OAI222D0BWP12T U1195 ( .A1(n1834), .A2(n1051), .B1(n283), .B2(n1049), .C1(
        n2098), .C2(n1050), .ZN(register_file_inst1_n2394) );
  TPOAI21D0BWP12T U1196 ( .A1(n283), .A2(n1104), .B(n2036), .ZN(
        register_file_inst1_spin[1]) );
  CKND0BWP12T U1197 ( .I(register_file_inst1_r2_1_), .ZN(n281) );
  OAI222D0BWP12T U1198 ( .A1(n2098), .A2(n1062), .B1(n283), .B2(n1063), .C1(
        n1060), .C2(n281), .ZN(register_file_inst1_n2554) );
  INVD1BWP12T U1199 ( .I(register_file_inst1_r5_1_), .ZN(n1787) );
  OAI222D0BWP12T U1200 ( .A1(n1787), .A2(n1096), .B1(n283), .B2(n1098), .C1(
        n2098), .C2(n1097), .ZN(register_file_inst1_n2458) );
  INVD1BWP12T U1201 ( .I(register_file_inst1_lr_1_), .ZN(n1778) );
  OAI222D0BWP12T U1202 ( .A1(n1778), .A2(n1082), .B1(n283), .B2(n1085), .C1(
        n2098), .C2(n1084), .ZN(register_file_inst1_n2202) );
  CKND0BWP12T U1203 ( .I(register_file_inst1_r8_1_), .ZN(n282) );
  OAI222D0BWP12T U1204 ( .A1(n282), .A2(n1075), .B1(n283), .B2(n1078), .C1(
        n2098), .C2(n1077), .ZN(register_file_inst1_n2362) );
  INVD1BWP12T U1205 ( .I(register_file_inst1_r1_1_), .ZN(n1832) );
  OAI222D0BWP12T U1206 ( .A1(n1832), .A2(n1093), .B1(n283), .B2(n1095), .C1(
        n2098), .C2(n1094), .ZN(register_file_inst1_n2586) );
  INVD1BWP12T U1207 ( .I(register_file_inst1_r11_1_), .ZN(n1831) );
  OAI222D0BWP12T U1208 ( .A1(n2098), .A2(n1020), .B1(n283), .B2(n1019), .C1(
        n1021), .C2(n1831), .ZN(register_file_inst1_n2266) );
  NR2D1BWP12T U1209 ( .A1(n2310), .A2(n289), .ZN(n838) );
  AOI22D0BWP12T U1210 ( .A1(register_file_inst1_r6_1_), .A2(n839), .B1(
        register_file_inst1_r4_1_), .B2(n838), .ZN(n288) );
  ND2D1BWP12T U1211 ( .A1(n2313), .A2(n2312), .ZN(n284) );
  NR2D1BWP12T U1212 ( .A1(n284), .A2(n2307), .ZN(n840) );
  AOI22D0BWP12T U1213 ( .A1(register_file_inst1_r7_1_), .A2(n841), .B1(
        register_file_inst1_r2_1_), .B2(n840), .ZN(n287) );
  NR2D1BWP12T U1214 ( .A1(n284), .A2(n2309), .ZN(n842) );
  AOI22D0BWP12T U1215 ( .A1(register_file_inst1_r0_1_), .A2(n843), .B1(
        register_file_inst1_r3_1_), .B2(n842), .ZN(n286) );
  AOI22D0BWP12T U1216 ( .A1(register_file_inst1_r1_1_), .A2(n845), .B1(
        register_file_inst1_r5_1_), .B2(n844), .ZN(n285) );
  ND4D1BWP12T U1217 ( .A1(n288), .A2(n287), .A3(n286), .A4(n285), .ZN(n294) );
  AOI22D0BWP12T U1218 ( .A1(register_file_inst1_r8_1_), .A2(n1948), .B1(
        STACK_RF_next_sp[1]), .B2(n1927), .ZN(n292) );
  NR2D1BWP12T U1219 ( .A1(n2309), .A2(n2314), .ZN(n851) );
  INVD1BWP12T U1220 ( .I(n851), .ZN(n744) );
  AOI22D0BWP12T U1221 ( .A1(register_file_inst1_r10_1_), .A2(n852), .B1(
        register_file_inst1_r11_1_), .B2(n851), .ZN(n291) );
  NR2XD0BWP12T U1222 ( .A1(n289), .A2(n2308), .ZN(n398) );
  AOI22D0BWP12T U1223 ( .A1(register_file_inst1_r9_1_), .A2(n850), .B1(
        register_file_inst1_r12_1_), .B2(n398), .ZN(n290) );
  ND4D1BWP12T U1224 ( .A1(n2037), .A2(n292), .A3(n291), .A4(n290), .ZN(n293)
         );
  AO21D1BWP12T U1225 ( .A1(n2306), .A2(n294), .B(n293), .Z(
        RF_MEMCTRL_data_reg[1]) );
  AOI22D0BWP12T U1226 ( .A1(register_file_inst1_r6_0_), .A2(n839), .B1(
        register_file_inst1_r4_0_), .B2(n838), .ZN(n298) );
  AOI22D0BWP12T U1227 ( .A1(register_file_inst1_r7_0_), .A2(n841), .B1(
        register_file_inst1_r2_0_), .B2(n840), .ZN(n297) );
  AOI22D0BWP12T U1228 ( .A1(register_file_inst1_r0_0_), .A2(n843), .B1(
        register_file_inst1_r3_0_), .B2(n842), .ZN(n296) );
  AOI22D0BWP12T U1229 ( .A1(register_file_inst1_r1_0_), .A2(n845), .B1(
        register_file_inst1_r5_0_), .B2(n844), .ZN(n295) );
  ND4D1BWP12T U1230 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(n303) );
  AOI22D0BWP12T U1231 ( .A1(STACK_RF_next_sp[0]), .A2(n1927), .B1(
        register_file_inst1_r8_0_), .B2(n1948), .ZN(n301) );
  AOI22D0BWP12T U1232 ( .A1(register_file_inst1_r10_0_), .A2(n852), .B1(
        register_file_inst1_r11_0_), .B2(n851), .ZN(n300) );
  AOI22D0BWP12T U1233 ( .A1(register_file_inst1_r9_0_), .A2(n850), .B1(
        register_file_inst1_r12_0_), .B2(n398), .ZN(n299) );
  ND4D1BWP12T U1234 ( .A1(n2038), .A2(n301), .A3(n300), .A4(n299), .ZN(n302)
         );
  AO21D1BWP12T U1235 ( .A1(n2306), .A2(n303), .B(n302), .Z(
        RF_MEMCTRL_data_reg[0]) );
  AOI22D0BWP12T U1236 ( .A1(register_file_inst1_r6_2_), .A2(n839), .B1(
        register_file_inst1_r4_2_), .B2(n838), .ZN(n307) );
  AOI22D0BWP12T U1237 ( .A1(register_file_inst1_r7_2_), .A2(n841), .B1(
        register_file_inst1_r2_2_), .B2(n840), .ZN(n306) );
  AOI22D0BWP12T U1238 ( .A1(register_file_inst1_r0_2_), .A2(n843), .B1(
        register_file_inst1_r3_2_), .B2(n842), .ZN(n305) );
  AOI22D0BWP12T U1239 ( .A1(register_file_inst1_r1_2_), .A2(n845), .B1(
        register_file_inst1_r5_2_), .B2(n844), .ZN(n304) );
  ND4D1BWP12T U1240 ( .A1(n307), .A2(n306), .A3(n305), .A4(n304), .ZN(n312) );
  AOI22D0BWP12T U1241 ( .A1(register_file_inst1_r8_2_), .A2(n1948), .B1(
        STACK_RF_next_sp[2]), .B2(n1927), .ZN(n310) );
  AOI22D0BWP12T U1242 ( .A1(register_file_inst1_r10_2_), .A2(n852), .B1(
        register_file_inst1_r11_2_), .B2(n851), .ZN(n309) );
  AOI22D0BWP12T U1243 ( .A1(register_file_inst1_r9_2_), .A2(n850), .B1(
        register_file_inst1_r12_2_), .B2(n398), .ZN(n308) );
  ND4D1BWP12T U1244 ( .A1(n1992), .A2(n310), .A3(n309), .A4(n308), .ZN(n311)
         );
  AO21D1BWP12T U1245 ( .A1(n2306), .A2(n312), .B(n311), .Z(
        RF_MEMCTRL_data_reg[2]) );
  AOI22D0BWP12T U1246 ( .A1(register_file_inst1_r6_3_), .A2(n839), .B1(
        register_file_inst1_r4_3_), .B2(n838), .ZN(n316) );
  AOI22D0BWP12T U1247 ( .A1(register_file_inst1_r7_3_), .A2(n841), .B1(
        register_file_inst1_r2_3_), .B2(n840), .ZN(n315) );
  AOI22D0BWP12T U1248 ( .A1(register_file_inst1_r0_3_), .A2(n843), .B1(
        register_file_inst1_r3_3_), .B2(n842), .ZN(n314) );
  AOI22D0BWP12T U1249 ( .A1(register_file_inst1_r1_3_), .A2(n845), .B1(
        register_file_inst1_r5_3_), .B2(n844), .ZN(n313) );
  ND4D1BWP12T U1250 ( .A1(n316), .A2(n315), .A3(n314), .A4(n313), .ZN(n321) );
  AOI22D0BWP12T U1251 ( .A1(register_file_inst1_r8_3_), .A2(n1948), .B1(
        STACK_RF_next_sp[3]), .B2(n1927), .ZN(n319) );
  AOI22D0BWP12T U1252 ( .A1(register_file_inst1_r10_3_), .A2(n852), .B1(
        register_file_inst1_r11_3_), .B2(n851), .ZN(n318) );
  AOI22D0BWP12T U1253 ( .A1(register_file_inst1_r9_3_), .A2(n850), .B1(
        register_file_inst1_r12_3_), .B2(n398), .ZN(n317) );
  ND4D1BWP12T U1254 ( .A1(n2033), .A2(n319), .A3(n318), .A4(n317), .ZN(n320)
         );
  AO21D1BWP12T U1255 ( .A1(n2306), .A2(n321), .B(n320), .Z(
        RF_MEMCTRL_data_reg[3]) );
  AOI22D0BWP12T U1256 ( .A1(register_file_inst1_r6_6_), .A2(n839), .B1(
        register_file_inst1_r4_6_), .B2(n838), .ZN(n325) );
  AOI22D1BWP12T U1257 ( .A1(register_file_inst1_r7_6_), .A2(n841), .B1(
        register_file_inst1_r2_6_), .B2(n840), .ZN(n324) );
  AOI22D1BWP12T U1258 ( .A1(register_file_inst1_r0_6_), .A2(n843), .B1(
        register_file_inst1_r3_6_), .B2(n842), .ZN(n323) );
  AOI22D0BWP12T U1259 ( .A1(register_file_inst1_r1_6_), .A2(n845), .B1(
        register_file_inst1_r5_6_), .B2(n844), .ZN(n322) );
  ND4D1BWP12T U1260 ( .A1(n325), .A2(n324), .A3(n323), .A4(n322), .ZN(n330) );
  AOI22D1BWP12T U1261 ( .A1(register_file_inst1_r8_6_), .A2(n1948), .B1(
        STACK_RF_next_sp[6]), .B2(n1927), .ZN(n328) );
  AOI22D1BWP12T U1262 ( .A1(register_file_inst1_r10_6_), .A2(n852), .B1(
        register_file_inst1_r11_6_), .B2(n851), .ZN(n327) );
  AOI22D0BWP12T U1263 ( .A1(register_file_inst1_r9_6_), .A2(n850), .B1(
        register_file_inst1_r12_6_), .B2(n398), .ZN(n326) );
  ND4D1BWP12T U1264 ( .A1(n2027), .A2(n328), .A3(n327), .A4(n326), .ZN(n329)
         );
  AO21D1BWP12T U1265 ( .A1(n2306), .A2(n330), .B(n329), .Z(
        RF_MEMCTRL_data_reg[6]) );
  AOI22D0BWP12T U1266 ( .A1(register_file_inst1_r6_7_), .A2(n839), .B1(
        register_file_inst1_r4_7_), .B2(n838), .ZN(n334) );
  AOI22D0BWP12T U1267 ( .A1(register_file_inst1_r7_7_), .A2(n841), .B1(
        register_file_inst1_r2_7_), .B2(n840), .ZN(n333) );
  AOI22D0BWP12T U1268 ( .A1(register_file_inst1_r0_7_), .A2(n843), .B1(
        register_file_inst1_r3_7_), .B2(n842), .ZN(n332) );
  AOI22D0BWP12T U1269 ( .A1(register_file_inst1_r1_7_), .A2(n845), .B1(
        register_file_inst1_r5_7_), .B2(n844), .ZN(n331) );
  ND4D1BWP12T U1270 ( .A1(n334), .A2(n333), .A3(n332), .A4(n331), .ZN(n339) );
  AOI22D0BWP12T U1271 ( .A1(register_file_inst1_r8_7_), .A2(n1948), .B1(
        STACK_RF_next_sp[7]), .B2(n1927), .ZN(n337) );
  AOI22D1BWP12T U1272 ( .A1(register_file_inst1_r10_7_), .A2(n852), .B1(
        register_file_inst1_r11_7_), .B2(n851), .ZN(n336) );
  AOI22D0BWP12T U1273 ( .A1(register_file_inst1_r9_7_), .A2(n850), .B1(
        register_file_inst1_r12_7_), .B2(n398), .ZN(n335) );
  ND4D1BWP12T U1274 ( .A1(n2024), .A2(n337), .A3(n336), .A4(n335), .ZN(n338)
         );
  AO21D1BWP12T U1275 ( .A1(n2306), .A2(n339), .B(n338), .Z(
        RF_MEMCTRL_data_reg[7]) );
  AOI22D0BWP12T U1276 ( .A1(register_file_inst1_r6_4_), .A2(n839), .B1(
        register_file_inst1_r4_4_), .B2(n838), .ZN(n343) );
  AOI22D0BWP12T U1277 ( .A1(register_file_inst1_r7_4_), .A2(n841), .B1(
        register_file_inst1_r2_4_), .B2(n840), .ZN(n342) );
  AOI22D0BWP12T U1278 ( .A1(register_file_inst1_r0_4_), .A2(n843), .B1(
        register_file_inst1_r3_4_), .B2(n842), .ZN(n341) );
  AOI22D0BWP12T U1279 ( .A1(register_file_inst1_r1_4_), .A2(n845), .B1(
        register_file_inst1_r5_4_), .B2(n844), .ZN(n340) );
  ND4D1BWP12T U1280 ( .A1(n343), .A2(n342), .A3(n341), .A4(n340), .ZN(n348) );
  AOI22D0BWP12T U1281 ( .A1(register_file_inst1_r8_4_), .A2(n1948), .B1(
        STACK_RF_next_sp[4]), .B2(n1927), .ZN(n346) );
  AOI22D0BWP12T U1282 ( .A1(register_file_inst1_r10_4_), .A2(n852), .B1(
        register_file_inst1_r11_4_), .B2(n851), .ZN(n345) );
  AOI22D0BWP12T U1283 ( .A1(register_file_inst1_r9_4_), .A2(n850), .B1(
        register_file_inst1_r12_4_), .B2(n398), .ZN(n344) );
  ND4D1BWP12T U1284 ( .A1(n2030), .A2(n346), .A3(n345), .A4(n344), .ZN(n347)
         );
  AO21D1BWP12T U1285 ( .A1(n2306), .A2(n348), .B(n347), .Z(
        RF_MEMCTRL_data_reg[4]) );
  AOI22D0BWP12T U1286 ( .A1(register_file_inst1_r6_5_), .A2(n839), .B1(
        register_file_inst1_r4_5_), .B2(n838), .ZN(n352) );
  AOI22D0BWP12T U1287 ( .A1(register_file_inst1_r7_5_), .A2(n841), .B1(
        register_file_inst1_r2_5_), .B2(n840), .ZN(n351) );
  AOI22D0BWP12T U1288 ( .A1(register_file_inst1_r0_5_), .A2(n843), .B1(
        register_file_inst1_r3_5_), .B2(n842), .ZN(n350) );
  AOI22D0BWP12T U1289 ( .A1(register_file_inst1_r1_5_), .A2(n845), .B1(
        register_file_inst1_r5_5_), .B2(n844), .ZN(n349) );
  ND4D1BWP12T U1290 ( .A1(n352), .A2(n351), .A3(n350), .A4(n349), .ZN(n357) );
  AOI22D1BWP12T U1291 ( .A1(register_file_inst1_r8_5_), .A2(n1948), .B1(
        STACK_RF_next_sp[5]), .B2(n1927), .ZN(n355) );
  AOI22D1BWP12T U1292 ( .A1(register_file_inst1_r10_5_), .A2(n852), .B1(
        register_file_inst1_r11_5_), .B2(n851), .ZN(n354) );
  AOI22D0BWP12T U1293 ( .A1(register_file_inst1_r9_5_), .A2(n850), .B1(
        register_file_inst1_r12_5_), .B2(n398), .ZN(n353) );
  ND4D1BWP12T U1294 ( .A1(n1989), .A2(n355), .A3(n354), .A4(n353), .ZN(n356)
         );
  AO21D1BWP12T U1295 ( .A1(n2306), .A2(n357), .B(n356), .Z(
        RF_MEMCTRL_data_reg[5]) );
  TPNR2D0BWP12T U1296 ( .A1(n2105), .A2(n1102), .ZN(n2028) );
  TPNR2D0BWP12T U1297 ( .A1(n2113), .A2(n1102), .ZN(n2022) );
  TPNR2D0BWP12T U1298 ( .A1(n2107), .A2(n1102), .ZN(n1987) );
  TPNR2D0BWP12T U1299 ( .A1(n2110), .A2(n1102), .ZN(n2025) );
  TPNR2D0BWP12T U1300 ( .A1(n2098), .A2(n1102), .ZN(n2034) );
  TPNR2D0BWP12T U1301 ( .A1(n2101), .A2(n1102), .ZN(n1990) );
  TPNR2D0BWP12T U1302 ( .A1(n2103), .A2(n1102), .ZN(n2031) );
  AOI22D0BWP12T U1303 ( .A1(register_file_inst1_r6_10_), .A2(n839), .B1(
        register_file_inst1_r4_10_), .B2(n838), .ZN(n361) );
  AOI22D0BWP12T U1304 ( .A1(register_file_inst1_r7_10_), .A2(n841), .B1(
        register_file_inst1_r2_10_), .B2(n840), .ZN(n360) );
  AOI22D0BWP12T U1305 ( .A1(register_file_inst1_r0_10_), .A2(n843), .B1(
        register_file_inst1_r3_10_), .B2(n842), .ZN(n359) );
  AOI22D0BWP12T U1306 ( .A1(register_file_inst1_r1_10_), .A2(n845), .B1(
        register_file_inst1_r5_10_), .B2(n844), .ZN(n358) );
  ND4D1BWP12T U1307 ( .A1(n361), .A2(n360), .A3(n359), .A4(n358), .ZN(n366) );
  AOI22D0BWP12T U1308 ( .A1(register_file_inst1_lr_10_), .A2(n1947), .B1(
        register_file_inst1_r8_10_), .B2(n1948), .ZN(n364) );
  AOI22D0BWP12T U1309 ( .A1(register_file_inst1_r10_10_), .A2(n852), .B1(
        register_file_inst1_r11_10_), .B2(n851), .ZN(n363) );
  AOI22D0BWP12T U1310 ( .A1(register_file_inst1_r9_10_), .A2(n850), .B1(
        register_file_inst1_r12_10_), .B2(n398), .ZN(n362) );
  ND4D1BWP12T U1311 ( .A1(n364), .A2(n2015), .A3(n363), .A4(n362), .ZN(n365)
         );
  AO21D1BWP12T U1312 ( .A1(n2306), .A2(n366), .B(n365), .Z(
        RF_MEMCTRL_data_reg[10]) );
  AOI22D0BWP12T U1313 ( .A1(register_file_inst1_r6_14_), .A2(n839), .B1(
        register_file_inst1_r4_14_), .B2(n838), .ZN(n370) );
  AOI22D0BWP12T U1314 ( .A1(register_file_inst1_r7_14_), .A2(n841), .B1(
        register_file_inst1_r2_14_), .B2(n840), .ZN(n369) );
  AOI22D0BWP12T U1315 ( .A1(register_file_inst1_r0_14_), .A2(n843), .B1(
        register_file_inst1_r3_14_), .B2(n842), .ZN(n368) );
  AOI22D0BWP12T U1316 ( .A1(register_file_inst1_r1_14_), .A2(n845), .B1(
        register_file_inst1_r5_14_), .B2(n844), .ZN(n367) );
  ND4D1BWP12T U1317 ( .A1(n370), .A2(n369), .A3(n368), .A4(n367), .ZN(n375) );
  AOI22D0BWP12T U1318 ( .A1(STACK_RF_next_sp[14]), .A2(n1927), .B1(
        register_file_inst1_r8_14_), .B2(n1948), .ZN(n373) );
  AOI22D0BWP12T U1319 ( .A1(register_file_inst1_r10_14_), .A2(n852), .B1(
        register_file_inst1_r11_14_), .B2(n851), .ZN(n372) );
  AOI22D0BWP12T U1320 ( .A1(register_file_inst1_r9_14_), .A2(n850), .B1(
        register_file_inst1_r12_14_), .B2(n398), .ZN(n371) );
  ND4D1BWP12T U1321 ( .A1(n1985), .A2(n373), .A3(n372), .A4(n371), .ZN(n374)
         );
  AO21D1BWP12T U1322 ( .A1(n2306), .A2(n375), .B(n374), .Z(
        RF_MEMCTRL_data_reg[14]) );
  AOI22D0BWP12T U1323 ( .A1(register_file_inst1_r6_12_), .A2(n839), .B1(
        register_file_inst1_r4_12_), .B2(n838), .ZN(n379) );
  AOI22D0BWP12T U1324 ( .A1(register_file_inst1_r7_12_), .A2(n841), .B1(
        register_file_inst1_r2_12_), .B2(n840), .ZN(n378) );
  AOI22D0BWP12T U1325 ( .A1(register_file_inst1_r0_12_), .A2(n843), .B1(
        register_file_inst1_r3_12_), .B2(n842), .ZN(n377) );
  AOI22D0BWP12T U1326 ( .A1(register_file_inst1_r1_12_), .A2(n845), .B1(
        register_file_inst1_r5_12_), .B2(n844), .ZN(n376) );
  ND4D1BWP12T U1327 ( .A1(n379), .A2(n378), .A3(n377), .A4(n376), .ZN(n384) );
  AOI22D0BWP12T U1328 ( .A1(register_file_inst1_lr_12_), .A2(n1947), .B1(
        register_file_inst1_r8_12_), .B2(n1948), .ZN(n382) );
  AOI22D0BWP12T U1329 ( .A1(register_file_inst1_r10_12_), .A2(n852), .B1(
        register_file_inst1_r11_12_), .B2(n851), .ZN(n381) );
  AOI22D0BWP12T U1330 ( .A1(register_file_inst1_r9_12_), .A2(n850), .B1(
        register_file_inst1_r12_12_), .B2(n398), .ZN(n380) );
  ND4D1BWP12T U1331 ( .A1(n382), .A2(n2009), .A3(n381), .A4(n380), .ZN(n383)
         );
  AO21D1BWP12T U1332 ( .A1(n2306), .A2(n384), .B(n383), .Z(
        RF_MEMCTRL_data_reg[12]) );
  AOI22D0BWP12T U1333 ( .A1(register_file_inst1_r6_11_), .A2(n839), .B1(
        register_file_inst1_r4_11_), .B2(n838), .ZN(n388) );
  AOI22D0BWP12T U1334 ( .A1(register_file_inst1_r7_11_), .A2(n841), .B1(
        register_file_inst1_r2_11_), .B2(n840), .ZN(n387) );
  AOI22D0BWP12T U1335 ( .A1(register_file_inst1_r0_11_), .A2(n843), .B1(
        register_file_inst1_r3_11_), .B2(n842), .ZN(n386) );
  AOI22D0BWP12T U1336 ( .A1(register_file_inst1_r1_11_), .A2(n845), .B1(
        register_file_inst1_r5_11_), .B2(n844), .ZN(n385) );
  ND4D1BWP12T U1337 ( .A1(n388), .A2(n387), .A3(n386), .A4(n385), .ZN(n393) );
  AOI22D0BWP12T U1338 ( .A1(register_file_inst1_lr_11_), .A2(n1947), .B1(
        register_file_inst1_r10_11_), .B2(n852), .ZN(n391) );
  AOI22D0BWP12T U1339 ( .A1(register_file_inst1_r11_11_), .A2(n851), .B1(
        STACK_RF_next_sp[11]), .B2(n1927), .ZN(n390) );
  AOI22D0BWP12T U1340 ( .A1(register_file_inst1_r9_11_), .A2(n850), .B1(
        register_file_inst1_r12_11_), .B2(n398), .ZN(n389) );
  ND4D1BWP12T U1341 ( .A1(n391), .A2(n2012), .A3(n390), .A4(n389), .ZN(n392)
         );
  AO21D1BWP12T U1342 ( .A1(n2306), .A2(n393), .B(n392), .Z(
        RF_MEMCTRL_data_reg[11]) );
  AOI22D0BWP12T U1343 ( .A1(register_file_inst1_r6_15_), .A2(n839), .B1(
        register_file_inst1_r4_15_), .B2(n838), .ZN(n397) );
  AOI22D0BWP12T U1344 ( .A1(register_file_inst1_r7_15_), .A2(n841), .B1(
        register_file_inst1_r2_15_), .B2(n840), .ZN(n396) );
  AOI22D0BWP12T U1345 ( .A1(register_file_inst1_r0_15_), .A2(n843), .B1(
        register_file_inst1_r3_15_), .B2(n842), .ZN(n395) );
  AOI22D0BWP12T U1346 ( .A1(register_file_inst1_r1_15_), .A2(n845), .B1(
        register_file_inst1_r5_15_), .B2(n844), .ZN(n394) );
  ND4D1BWP12T U1347 ( .A1(n397), .A2(n396), .A3(n395), .A4(n394), .ZN(n403) );
  AOI22D0BWP12T U1348 ( .A1(register_file_inst1_lr_15_), .A2(n1947), .B1(
        STACK_RF_next_sp[15]), .B2(n1927), .ZN(n401) );
  AOI22D0BWP12T U1349 ( .A1(register_file_inst1_r10_15_), .A2(n852), .B1(
        register_file_inst1_r11_15_), .B2(n851), .ZN(n400) );
  AOI22D0BWP12T U1350 ( .A1(register_file_inst1_r9_15_), .A2(n850), .B1(
        register_file_inst1_r12_15_), .B2(n398), .ZN(n399) );
  ND4D1BWP12T U1351 ( .A1(n401), .A2(n2006), .A3(n400), .A4(n399), .ZN(n402)
         );
  AO21D1BWP12T U1352 ( .A1(n2306), .A2(n403), .B(n402), .Z(
        RF_MEMCTRL_data_reg[15]) );
  AOI22D0BWP12T U1353 ( .A1(register_file_inst1_r6_13_), .A2(n839), .B1(
        register_file_inst1_r4_13_), .B2(n838), .ZN(n407) );
  AOI22D0BWP12T U1354 ( .A1(register_file_inst1_r7_13_), .A2(n841), .B1(
        register_file_inst1_r2_13_), .B2(n840), .ZN(n406) );
  AOI22D0BWP12T U1355 ( .A1(register_file_inst1_r0_13_), .A2(n843), .B1(
        register_file_inst1_r3_13_), .B2(n842), .ZN(n405) );
  AOI22D0BWP12T U1356 ( .A1(register_file_inst1_r1_13_), .A2(n845), .B1(
        register_file_inst1_r5_13_), .B2(n844), .ZN(n404) );
  ND4D1BWP12T U1357 ( .A1(n407), .A2(n406), .A3(n405), .A4(n404), .ZN(n412) );
  AOI22D0BWP12T U1358 ( .A1(STACK_RF_next_sp[13]), .A2(n1927), .B1(
        register_file_inst1_r8_13_), .B2(n1948), .ZN(n410) );
  AOI22D0BWP12T U1359 ( .A1(register_file_inst1_r10_13_), .A2(n852), .B1(
        register_file_inst1_r11_13_), .B2(n851), .ZN(n409) );
  AOI22D0BWP12T U1360 ( .A1(register_file_inst1_r9_13_), .A2(n850), .B1(
        register_file_inst1_r12_13_), .B2(n398), .ZN(n408) );
  ND4D1BWP12T U1361 ( .A1(n1986), .A2(n410), .A3(n409), .A4(n408), .ZN(n411)
         );
  AO21D1BWP12T U1362 ( .A1(n2306), .A2(n412), .B(n411), .Z(
        RF_MEMCTRL_data_reg[13]) );
  AOI22D0BWP12T U1363 ( .A1(register_file_inst1_r6_9_), .A2(n839), .B1(
        register_file_inst1_r4_9_), .B2(n838), .ZN(n416) );
  AOI22D0BWP12T U1364 ( .A1(register_file_inst1_r7_9_), .A2(n841), .B1(
        register_file_inst1_r2_9_), .B2(n840), .ZN(n415) );
  AOI22D0BWP12T U1365 ( .A1(register_file_inst1_r0_9_), .A2(n843), .B1(
        register_file_inst1_r3_9_), .B2(n842), .ZN(n414) );
  AOI22D0BWP12T U1366 ( .A1(register_file_inst1_r1_9_), .A2(n845), .B1(
        register_file_inst1_r5_9_), .B2(n844), .ZN(n413) );
  ND4D1BWP12T U1367 ( .A1(n416), .A2(n415), .A3(n414), .A4(n413), .ZN(n421) );
  AOI22D0BWP12T U1368 ( .A1(register_file_inst1_lr_9_), .A2(n1947), .B1(
        register_file_inst1_r8_9_), .B2(n1948), .ZN(n419) );
  AOI22D1BWP12T U1369 ( .A1(register_file_inst1_r10_9_), .A2(n852), .B1(
        register_file_inst1_r11_9_), .B2(n851), .ZN(n418) );
  AOI22D0BWP12T U1370 ( .A1(register_file_inst1_r9_9_), .A2(n850), .B1(
        register_file_inst1_r12_9_), .B2(n398), .ZN(n417) );
  ND4D1BWP12T U1371 ( .A1(n419), .A2(n2018), .A3(n418), .A4(n417), .ZN(n420)
         );
  AO21D1BWP12T U1372 ( .A1(n2306), .A2(n421), .B(n420), .Z(
        RF_MEMCTRL_data_reg[9]) );
  AOI22D0BWP12T U1373 ( .A1(register_file_inst1_r6_8_), .A2(n839), .B1(
        register_file_inst1_r4_8_), .B2(n838), .ZN(n425) );
  AOI22D0BWP12T U1374 ( .A1(register_file_inst1_r7_8_), .A2(n841), .B1(
        register_file_inst1_r2_8_), .B2(n840), .ZN(n424) );
  AOI22D0BWP12T U1375 ( .A1(register_file_inst1_r0_8_), .A2(n843), .B1(
        register_file_inst1_r3_8_), .B2(n842), .ZN(n423) );
  AOI22D0BWP12T U1376 ( .A1(register_file_inst1_r1_8_), .A2(n845), .B1(
        register_file_inst1_r5_8_), .B2(n844), .ZN(n422) );
  ND4D1BWP12T U1377 ( .A1(n425), .A2(n424), .A3(n423), .A4(n422), .ZN(n430) );
  AOI22D0BWP12T U1378 ( .A1(register_file_inst1_lr_8_), .A2(n1947), .B1(
        register_file_inst1_r8_8_), .B2(n1948), .ZN(n428) );
  AOI22D0BWP12T U1379 ( .A1(register_file_inst1_r10_8_), .A2(n852), .B1(
        register_file_inst1_r11_8_), .B2(n851), .ZN(n427) );
  AOI22D0BWP12T U1380 ( .A1(register_file_inst1_r9_8_), .A2(n850), .B1(
        register_file_inst1_r12_8_), .B2(n398), .ZN(n426) );
  ND4D1BWP12T U1381 ( .A1(n428), .A2(n2021), .A3(n427), .A4(n426), .ZN(n429)
         );
  AO21D1BWP12T U1382 ( .A1(n2306), .A2(n430), .B(n429), .Z(
        RF_MEMCTRL_data_reg[8]) );
  OAI22D1BWP12T U1383 ( .A1(n431), .A2(n1873), .B1(n1553), .B2(n1871), .ZN(
        n442) );
  OAI22D1BWP12T U1384 ( .A1(n433), .A2(n1877), .B1(n432), .B2(n1875), .ZN(n441) );
  AOI22D1BWP12T U1385 ( .A1(register_file_inst1_tmp1_25_), .A2(n1835), .B1(
        register_file_inst1_r0_25_), .B2(n1633), .ZN(n435) );
  AOI22D1BWP12T U1386 ( .A1(register_file_inst1_r5_25_), .A2(n1868), .B1(
        STACK_RF_next_sp[25]), .B2(n1867), .ZN(n434) );
  ND3D1BWP12T U1387 ( .A1(n435), .A2(n434), .A3(n2156), .ZN(n440) );
  AOI22D1BWP12T U1388 ( .A1(register_file_inst1_r12_25_), .A2(n1659), .B1(
        register_file_inst1_r8_25_), .B2(n1838), .ZN(n438) );
  AOI22D1BWP12T U1389 ( .A1(register_file_inst1_r4_25_), .A2(n1595), .B1(
        register_file_inst1_r3_25_), .B2(n1839), .ZN(n437) );
  AOI22D1BWP12T U1390 ( .A1(register_file_inst1_r6_25_), .A2(n1596), .B1(
        register_file_inst1_r10_25_), .B2(n1840), .ZN(n436) );
  ND4D1BWP12T U1391 ( .A1(n438), .A2(n437), .A3(n2157), .A4(n436), .ZN(n439)
         );
  OR4D1BWP12T U1392 ( .A1(n442), .A2(n441), .A3(n440), .A4(n439), .Z(
        RF_ALU_operand_b[25]) );
  CKND2D1BWP12T U1393 ( .A1(n501), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[7]), .ZN(n2270) );
  TPND2D0BWP12T U1394 ( .A1(n501), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[8]), .ZN(n2266) );
  CKND2D1BWP12T U1395 ( .A1(n501), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[6]), .ZN(n2271) );
  TPND2D0BWP12T U1396 ( .A1(n501), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[9]), .ZN(n2264) );
  TPND2D0BWP12T U1397 ( .A1(n501), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[10]), .ZN(n2262) );
  TPND2D0BWP12T U1398 ( .A1(n501), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[11]), .ZN(n2260) );
  TPND2D0BWP12T U1399 ( .A1(n501), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[12]), .ZN(n2258) );
  TPND2D0BWP12T U1400 ( .A1(n501), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[13]), .ZN(n2256) );
  TPND2D0BWP12T U1401 ( .A1(n501), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[14]), .ZN(n2254) );
  INVD1BWP12T U1402 ( .I(STACK_RF_next_sp[10]), .ZN(n443) );
  OAI22D1BWP12T U1403 ( .A1(n444), .A2(n1798), .B1(n443), .B2(n1796), .ZN(n451) );
  OAI22D1BWP12T U1404 ( .A1(n2202), .A2(n1802), .B1(n445), .B2(n1800), .ZN(
        n450) );
  OAI22D1BWP12T U1405 ( .A1(n447), .A2(n1805), .B1(n446), .B2(n1803), .ZN(n449) );
  OAI22D1BWP12T U1406 ( .A1(n1408), .A2(n1809), .B1(n1410), .B2(n1807), .ZN(
        n448) );
  NR4D0BWP12T U1407 ( .A1(n451), .A2(n450), .A3(n449), .A4(n448), .ZN(n464) );
  CKND2D1BWP12T U1408 ( .A1(register_file_inst1_r9_10_), .A2(n1911), .ZN(n453)
         );
  CKND2D1BWP12T U1409 ( .A1(register_file_inst1_r8_10_), .A2(n1910), .ZN(n452)
         );
  ND3D1BWP12T U1410 ( .A1(n2203), .A2(n453), .A3(n452), .ZN(n462) );
  OAI22D1BWP12T U1411 ( .A1(n455), .A2(n1903), .B1(n454), .B2(n1901), .ZN(n461) );
  OAI22D1BWP12T U1412 ( .A1(n456), .A2(n1907), .B1(n1407), .B2(n1905), .ZN(
        n460) );
  OAI22D1BWP12T U1413 ( .A1(n458), .A2(n1823), .B1(n457), .B2(n1821), .ZN(n459) );
  NR4D0BWP12T U1414 ( .A1(n462), .A2(n461), .A3(n460), .A4(n459), .ZN(n463) );
  CKND2D1BWP12T U1415 ( .A1(n464), .A2(n463), .ZN(RF_ALU_STACK_operand_a[10])
         );
  OAI22D1BWP12T U1416 ( .A1(n465), .A2(n1873), .B1(n582), .B2(n1871), .ZN(n476) );
  OAI22D1BWP12T U1417 ( .A1(n467), .A2(n1877), .B1(n466), .B2(n1875), .ZN(n475) );
  AOI22D1BWP12T U1418 ( .A1(register_file_inst1_tmp1_26_), .A2(n1835), .B1(
        register_file_inst1_r0_26_), .B2(n1633), .ZN(n469) );
  AOI22D1BWP12T U1419 ( .A1(register_file_inst1_r5_26_), .A2(n1868), .B1(
        STACK_RF_next_sp[26]), .B2(n1867), .ZN(n468) );
  ND3D1BWP12T U1420 ( .A1(n469), .A2(n468), .A3(n2158), .ZN(n474) );
  AOI22D1BWP12T U1421 ( .A1(register_file_inst1_r12_26_), .A2(n1659), .B1(
        register_file_inst1_r8_26_), .B2(n1838), .ZN(n472) );
  AOI22D1BWP12T U1422 ( .A1(register_file_inst1_r4_26_), .A2(n1595), .B1(
        register_file_inst1_r3_26_), .B2(n1839), .ZN(n471) );
  AOI22D1BWP12T U1423 ( .A1(register_file_inst1_r6_26_), .A2(n1596), .B1(
        register_file_inst1_r10_26_), .B2(n1840), .ZN(n470) );
  ND4D1BWP12T U1424 ( .A1(n472), .A2(n471), .A3(n2159), .A4(n470), .ZN(n473)
         );
  OR4D1BWP12T U1425 ( .A1(n476), .A2(n475), .A3(n474), .A4(n473), .Z(
        RF_ALU_operand_b[26]) );
  INVD1BWP12T U1426 ( .I(register_file_inst1_r1_28_), .ZN(n1005) );
  INVD1BWP12T U1427 ( .I(register_file_inst1_r11_28_), .ZN(n1579) );
  OAI22D1BWP12T U1428 ( .A1(n1005), .A2(n1873), .B1(n1579), .B2(n1871), .ZN(
        n485) );
  INVD1BWP12T U1429 ( .I(register_file_inst1_r7_28_), .ZN(n1006) );
  INVD1BWP12T U1430 ( .I(register_file_inst1_r9_28_), .ZN(n1013) );
  OAI22D1BWP12T U1431 ( .A1(n1006), .A2(n1877), .B1(n1013), .B2(n1875), .ZN(
        n484) );
  AOI22D1BWP12T U1432 ( .A1(register_file_inst1_tmp1_28_), .A2(n1835), .B1(
        register_file_inst1_r0_28_), .B2(n1633), .ZN(n478) );
  AOI22D1BWP12T U1433 ( .A1(register_file_inst1_r5_28_), .A2(n1868), .B1(
        STACK_RF_next_sp[28]), .B2(n1867), .ZN(n477) );
  ND3D1BWP12T U1434 ( .A1(n478), .A2(n477), .A3(n2162), .ZN(n483) );
  AOI22D1BWP12T U1435 ( .A1(register_file_inst1_r12_28_), .A2(n1659), .B1(
        register_file_inst1_r8_28_), .B2(n1838), .ZN(n481) );
  AOI22D1BWP12T U1436 ( .A1(register_file_inst1_r4_28_), .A2(n1595), .B1(
        register_file_inst1_r3_28_), .B2(n1839), .ZN(n480) );
  AOI22D1BWP12T U1437 ( .A1(register_file_inst1_r6_28_), .A2(n1596), .B1(
        register_file_inst1_r10_28_), .B2(n1840), .ZN(n479) );
  ND4D1BWP12T U1438 ( .A1(n481), .A2(n480), .A3(n2163), .A4(n479), .ZN(n482)
         );
  OR4D1BWP12T U1439 ( .A1(n485), .A2(n484), .A3(n483), .A4(n482), .Z(
        RF_ALU_operand_b[28]) );
  OAI22D1BWP12T U1440 ( .A1(n486), .A2(n1873), .B1(n1566), .B2(n1871), .ZN(
        n497) );
  OAI22D1BWP12T U1441 ( .A1(n488), .A2(n1877), .B1(n487), .B2(n1875), .ZN(n496) );
  AOI22D1BWP12T U1442 ( .A1(register_file_inst1_tmp1_27_), .A2(n1835), .B1(
        register_file_inst1_r0_27_), .B2(n1633), .ZN(n490) );
  AOI22D1BWP12T U1443 ( .A1(register_file_inst1_r5_27_), .A2(n1868), .B1(
        STACK_RF_next_sp[27]), .B2(n1867), .ZN(n489) );
  ND3D1BWP12T U1444 ( .A1(n490), .A2(n489), .A3(n2160), .ZN(n495) );
  AOI22D1BWP12T U1445 ( .A1(register_file_inst1_r12_27_), .A2(n1659), .B1(
        register_file_inst1_r8_27_), .B2(n1838), .ZN(n493) );
  AOI22D1BWP12T U1446 ( .A1(register_file_inst1_r4_27_), .A2(n1595), .B1(
        register_file_inst1_r3_27_), .B2(n1839), .ZN(n492) );
  AOI22D1BWP12T U1447 ( .A1(register_file_inst1_r6_27_), .A2(n1596), .B1(
        register_file_inst1_r10_27_), .B2(n1840), .ZN(n491) );
  ND4D1BWP12T U1448 ( .A1(n493), .A2(n492), .A3(n2161), .A4(n491), .ZN(n494)
         );
  OR4D1BWP12T U1449 ( .A1(n497), .A2(n496), .A3(n495), .A4(n494), .Z(
        RF_ALU_operand_b[27]) );
  CKND2D0BWP12T U1450 ( .A1(n772), .A2(MEMCTRL_load_in), .ZN(n1957) );
  INR3XD0BWP12T U1451 ( .A1(n498), .B1(n2288), .B2(n501), .ZN(n2040) );
  BUFFD1BWP12T U1452 ( .I(n2285), .Z(n1949) );
  BUFFD1BWP12T U1453 ( .I(n2286), .Z(n1950) );
  CKND0BWP12T U1454 ( .I(n1104), .ZN(n1936) );
  CKND0BWP12T U1455 ( .I(n1081), .ZN(n1935) );
  CKND0BWP12T U1456 ( .I(n1078), .ZN(n1933) );
  CKND0BWP12T U1457 ( .I(n1074), .ZN(n1934) );
  INR2D0BWP12T U1458 ( .A1(memory_interface_inst1_fsm_state_2_), .B1(
        memory_interface_inst1_fsm_state_1_), .ZN(n615) );
  NR2D0BWP12T U1459 ( .A1(n615), .A2(memory_interface_inst1_fsm_state_0_), 
        .ZN(n2249) );
  AOI21D0BWP12T U1460 ( .A1(memory_interface_inst1_fsm_state_2_), .A2(
        memory_interface_inst1_fsm_state_1_), .B(n499), .ZN(n2248) );
  OAI21D0BWP12T U1461 ( .A1(n2279), .A2(n2278), .B(n514), .ZN(n2280) );
  CKND0BWP12T U1462 ( .I(n2275), .ZN(n1967) );
  CKND0BWP12T U1463 ( .I(n2183), .ZN(n2174) );
  AOI21D1BWP12T U1464 ( .A1(MEM_MEMCTRL_from_mem_data[7]), .A2(n501), .B(n500), 
        .ZN(n1101) );
  DCCKND8BWP12T U1465 ( .I(ALU_MISC_OUT_result[30]), .ZN(n1054) );
  AOI21D1BWP12T U1466 ( .A1(n501), .A2(MEM_MEMCTRL_from_mem_data[6]), .B(n500), 
        .ZN(n1055) );
  MUX2ND0BWP12T U1467 ( .I0(n1054), .I1(n1055), .S(n514), .ZN(n1110) );
  INVD3BWP12T U1468 ( .I(ALU_MISC_OUT_result[29]), .ZN(n1030) );
  AOI21D1BWP12T U1469 ( .A1(n501), .A2(MEM_MEMCTRL_from_mem_data[5]), .B(n500), 
        .ZN(n1031) );
  INVD2BWP12T U1470 ( .I(ALU_MISC_OUT_result[28]), .ZN(n1011) );
  AOI21D1BWP12T U1471 ( .A1(n501), .A2(MEM_MEMCTRL_from_mem_data[4]), .B(n500), 
        .ZN(n1012) );
  MUX2NXD0BWP12T U1472 ( .I0(n1011), .I1(n1012), .S(n514), .ZN(n1106) );
  MUX2NXD0BWP12T U1473 ( .I0(n505), .I1(n504), .S(n514), .ZN(n1057) );
  MUX2NXD0BWP12T U1474 ( .I0(n509), .I1(n508), .S(n514), .ZN(n1033) );
  MUX2D1BWP12T U1475 ( .I0(n511), .I1(n510), .S(n514), .Z(n1018) );
  MUX2NXD0BWP12T U1476 ( .I0(n988), .I1(n989), .S(n514), .ZN(n1014) );
  MUX2D1BWP12T U1477 ( .I0(n513), .I1(n512), .S(n514), .Z(n1002) );
  MUX2NXD0BWP12T U1478 ( .I0(n516), .I1(n515), .S(n514), .ZN(n998) );
  NR2XD1BWP12T U1479 ( .A1(n14), .A2(n517), .ZN(n999) );
  TPND2D1BWP12T U1480 ( .A1(n998), .A2(n999), .ZN(n1001) );
  NR2XD1BWP12T U1481 ( .A1(n1002), .A2(n1001), .ZN(n1015) );
  TPNR2D3BWP12T U1482 ( .A1(n1018), .A2(n1017), .ZN(n1034) );
  TPND2D2BWP12T U1483 ( .A1(n1033), .A2(n1034), .ZN(n1036) );
  TPNR2D3BWP12T U1484 ( .A1(n11), .A2(n1036), .ZN(n1058) );
  TPND2D2BWP12T U1485 ( .A1(n1057), .A2(n1058), .ZN(n1105) );
  TPNR2D3BWP12T U1486 ( .A1(n12), .A2(n1105), .ZN(n1107) );
  TPND2D2BWP12T U1487 ( .A1(n1106), .A2(n1107), .ZN(n1109) );
  TPNR2D2BWP12T U1488 ( .A1(n13), .A2(n1109), .ZN(n1111) );
  ND2D1BWP12T U1489 ( .A1(n1110), .A2(n1111), .ZN(n518) );
  XOR2XD1BWP12T U1490 ( .A1(n519), .A2(n518), .Z(n520) );
  IOA21D2BWP12T U1491 ( .A1(n520), .A2(n2287), .B(n2281), .ZN(
        register_file_inst1_n2200) );
  OAI22D1BWP12T U1492 ( .A1(n522), .A2(n1903), .B1(n521), .B2(n1901), .ZN(n532) );
  OAI22D1BWP12T U1493 ( .A1(n523), .A2(n1907), .B1(n533), .B2(n1905), .ZN(n531) );
  AOI22D1BWP12T U1494 ( .A1(register_file_inst1_tmp1_20_), .A2(n2244), .B1(
        register_file_inst1_r6_20_), .B2(n1909), .ZN(n525) );
  AOI22D1BWP12T U1495 ( .A1(register_file_inst1_r9_20_), .A2(n1911), .B1(
        register_file_inst1_r8_20_), .B2(n1910), .ZN(n524) );
  ND3D1BWP12T U1496 ( .A1(n525), .A2(n524), .A3(n2222), .ZN(n530) );
  AOI22D1BWP12T U1497 ( .A1(register_file_inst1_r12_20_), .A2(n1915), .B1(
        STACK_RF_next_sp[20]), .B2(n1914), .ZN(n528) );
  AOI22D1BWP12T U1498 ( .A1(register_file_inst1_lr_20_), .A2(n1917), .B1(
        register_file_inst1_r3_20_), .B2(n1916), .ZN(n527) );
  AOI22D1BWP12T U1499 ( .A1(register_file_inst1_r1_20_), .A2(n1919), .B1(
        register_file_inst1_r7_20_), .B2(n1918), .ZN(n526) );
  ND4D1BWP12T U1500 ( .A1(n528), .A2(n2223), .A3(n527), .A4(n526), .ZN(n529)
         );
  OR4D2BWP12T U1501 ( .A1(n532), .A2(n531), .A3(n530), .A4(n529), .Z(
        RF_ALU_STACK_operand_a[20]) );
  OAI22D1BWP12T U1502 ( .A1(n534), .A2(n1873), .B1(n533), .B2(n1871), .ZN(n545) );
  OAI22D1BWP12T U1503 ( .A1(n536), .A2(n1877), .B1(n535), .B2(n1875), .ZN(n544) );
  AOI22D1BWP12T U1504 ( .A1(register_file_inst1_tmp1_20_), .A2(n1835), .B1(
        register_file_inst1_r0_20_), .B2(n1633), .ZN(n538) );
  AOI22D1BWP12T U1505 ( .A1(register_file_inst1_r5_20_), .A2(n1868), .B1(
        STACK_RF_next_sp[20]), .B2(n1867), .ZN(n537) );
  ND3D1BWP12T U1506 ( .A1(n538), .A2(n537), .A3(n2146), .ZN(n543) );
  AOI22D1BWP12T U1507 ( .A1(register_file_inst1_r12_20_), .A2(n1659), .B1(
        register_file_inst1_r8_20_), .B2(n1838), .ZN(n541) );
  AOI22D1BWP12T U1508 ( .A1(register_file_inst1_r4_20_), .A2(n1595), .B1(
        register_file_inst1_r3_20_), .B2(n1839), .ZN(n540) );
  AOI22D1BWP12T U1509 ( .A1(register_file_inst1_r6_20_), .A2(n1596), .B1(
        register_file_inst1_r10_20_), .B2(n1840), .ZN(n539) );
  ND4D1BWP12T U1510 ( .A1(n541), .A2(n540), .A3(n2147), .A4(n539), .ZN(n542)
         );
  OAI22D1BWP12T U1511 ( .A1(n546), .A2(n1873), .B1(n1906), .B2(n1871), .ZN(
        n557) );
  OAI22D1BWP12T U1512 ( .A1(n548), .A2(n1877), .B1(n547), .B2(n1875), .ZN(n556) );
  AOI22D1BWP12T U1513 ( .A1(register_file_inst1_tmp1_21_), .A2(n1835), .B1(
        register_file_inst1_r0_21_), .B2(n1633), .ZN(n550) );
  AOI22D1BWP12T U1514 ( .A1(register_file_inst1_r5_21_), .A2(n1868), .B1(
        STACK_RF_next_sp[21]), .B2(n1867), .ZN(n549) );
  ND3D1BWP12T U1515 ( .A1(n550), .A2(n549), .A3(n2148), .ZN(n555) );
  AOI22D1BWP12T U1516 ( .A1(register_file_inst1_r12_21_), .A2(n1659), .B1(
        register_file_inst1_r8_21_), .B2(n1838), .ZN(n553) );
  AOI22D1BWP12T U1517 ( .A1(register_file_inst1_r4_21_), .A2(n1595), .B1(
        register_file_inst1_r3_21_), .B2(n1839), .ZN(n552) );
  AOI22D1BWP12T U1518 ( .A1(register_file_inst1_r6_21_), .A2(n1596), .B1(
        register_file_inst1_r10_21_), .B2(n1840), .ZN(n551) );
  ND4D1BWP12T U1519 ( .A1(n553), .A2(n552), .A3(n2149), .A4(n551), .ZN(n554)
         );
  INVD1BWP12T U1520 ( .I(register_file_inst1_r1_22_), .ZN(n979) );
  OAI22D1BWP12T U1521 ( .A1(n979), .A2(n1873), .B1(n593), .B2(n1871), .ZN(n566) );
  INVD1BWP12T U1522 ( .I(register_file_inst1_r7_22_), .ZN(n605) );
  INVD1BWP12T U1523 ( .I(register_file_inst1_r9_22_), .ZN(n990) );
  OAI22D1BWP12T U1524 ( .A1(n605), .A2(n1877), .B1(n990), .B2(n1875), .ZN(n565) );
  AOI22D1BWP12T U1525 ( .A1(register_file_inst1_tmp1_22_), .A2(n1835), .B1(
        register_file_inst1_r0_22_), .B2(n1633), .ZN(n559) );
  AOI22D1BWP12T U1526 ( .A1(register_file_inst1_r5_22_), .A2(n1868), .B1(
        STACK_RF_next_sp[22]), .B2(n1867), .ZN(n558) );
  ND3D1BWP12T U1527 ( .A1(n559), .A2(n558), .A3(n2150), .ZN(n564) );
  AOI22D1BWP12T U1528 ( .A1(register_file_inst1_r12_22_), .A2(n1659), .B1(
        register_file_inst1_r8_22_), .B2(n1838), .ZN(n562) );
  AOI22D1BWP12T U1529 ( .A1(register_file_inst1_r4_22_), .A2(n1595), .B1(
        register_file_inst1_r3_22_), .B2(n1839), .ZN(n561) );
  AOI22D1BWP12T U1530 ( .A1(register_file_inst1_r6_22_), .A2(n1596), .B1(
        register_file_inst1_r10_22_), .B2(n1840), .ZN(n560) );
  ND4D1BWP12T U1531 ( .A1(n562), .A2(n561), .A3(n2151), .A4(n560), .ZN(n563)
         );
  OAI22D1BWP12T U1532 ( .A1(n568), .A2(n1903), .B1(n567), .B2(n1901), .ZN(n579) );
  OAI22D1BWP12T U1533 ( .A1(n570), .A2(n1907), .B1(n569), .B2(n1905), .ZN(n578) );
  AOI22D1BWP12T U1534 ( .A1(register_file_inst1_tmp1_24_), .A2(n2244), .B1(
        register_file_inst1_r6_24_), .B2(n1909), .ZN(n572) );
  AOI22D1BWP12T U1535 ( .A1(register_file_inst1_r9_24_), .A2(n1911), .B1(
        register_file_inst1_r8_24_), .B2(n1910), .ZN(n571) );
  ND3D1BWP12T U1536 ( .A1(n572), .A2(n571), .A3(n2230), .ZN(n577) );
  AOI22D1BWP12T U1537 ( .A1(register_file_inst1_r12_24_), .A2(n1915), .B1(
        STACK_RF_next_sp[24]), .B2(n1914), .ZN(n575) );
  AOI22D1BWP12T U1538 ( .A1(register_file_inst1_lr_24_), .A2(n1917), .B1(
        register_file_inst1_r3_24_), .B2(n1916), .ZN(n574) );
  AOI22D1BWP12T U1539 ( .A1(register_file_inst1_r1_24_), .A2(n1919), .B1(
        register_file_inst1_r7_24_), .B2(n1918), .ZN(n573) );
  ND4D1BWP12T U1540 ( .A1(n575), .A2(n2231), .A3(n574), .A4(n573), .ZN(n576)
         );
  OAI22D1BWP12T U1541 ( .A1(n581), .A2(n1903), .B1(n580), .B2(n1901), .ZN(n592) );
  OAI22D1BWP12T U1542 ( .A1(n583), .A2(n1907), .B1(n582), .B2(n1905), .ZN(n591) );
  AOI22D1BWP12T U1543 ( .A1(register_file_inst1_tmp1_26_), .A2(n2244), .B1(
        register_file_inst1_r6_26_), .B2(n1909), .ZN(n585) );
  AOI22D1BWP12T U1544 ( .A1(register_file_inst1_r8_26_), .A2(n1910), .B1(
        register_file_inst1_r9_26_), .B2(n1911), .ZN(n584) );
  ND3D1BWP12T U1545 ( .A1(n585), .A2(n584), .A3(n2234), .ZN(n590) );
  AOI22D1BWP12T U1546 ( .A1(register_file_inst1_r12_26_), .A2(n1915), .B1(
        STACK_RF_next_sp[26]), .B2(n1914), .ZN(n588) );
  AOI22D1BWP12T U1547 ( .A1(register_file_inst1_lr_26_), .A2(n1917), .B1(
        register_file_inst1_r3_26_), .B2(n1916), .ZN(n587) );
  AOI22D1BWP12T U1548 ( .A1(register_file_inst1_r1_26_), .A2(n1919), .B1(
        register_file_inst1_r7_26_), .B2(n1918), .ZN(n586) );
  ND4D1BWP12T U1549 ( .A1(n588), .A2(n2235), .A3(n587), .A4(n586), .ZN(n589)
         );
  INVD1BWP12T U1550 ( .I(register_file_inst1_r4_22_), .ZN(n981) );
  INVD1BWP12T U1551 ( .I(register_file_inst1_r10_22_), .ZN(n984) );
  OAI22D1BWP12T U1552 ( .A1(n981), .A2(n1903), .B1(n984), .B2(n1901), .ZN(n602) );
  INVD1BWP12T U1553 ( .I(register_file_inst1_r5_22_), .ZN(n977) );
  OAI22D1BWP12T U1554 ( .A1(n977), .A2(n1907), .B1(n593), .B2(n1905), .ZN(n601) );
  AOI22D1BWP12T U1555 ( .A1(register_file_inst1_tmp1_22_), .A2(n2244), .B1(
        register_file_inst1_r6_22_), .B2(n1909), .ZN(n595) );
  AOI22D1BWP12T U1556 ( .A1(register_file_inst1_r9_22_), .A2(n1911), .B1(
        register_file_inst1_r8_22_), .B2(n1910), .ZN(n594) );
  ND3D1BWP12T U1557 ( .A1(n595), .A2(n594), .A3(n2226), .ZN(n600) );
  AOI22D1BWP12T U1558 ( .A1(register_file_inst1_r12_22_), .A2(n1915), .B1(
        STACK_RF_next_sp[22]), .B2(n1914), .ZN(n598) );
  AOI22D1BWP12T U1559 ( .A1(register_file_inst1_lr_22_), .A2(n1917), .B1(
        register_file_inst1_r3_22_), .B2(n1916), .ZN(n597) );
  AOI22D1BWP12T U1560 ( .A1(register_file_inst1_r1_22_), .A2(n1919), .B1(
        register_file_inst1_r7_22_), .B2(n1918), .ZN(n596) );
  ND4D1BWP12T U1561 ( .A1(n598), .A2(n2227), .A3(n597), .A4(n596), .ZN(n599)
         );
  INVD1BWP12T U1562 ( .I(register_file_inst1_r6_16_), .ZN(n1197) );
  OAI222D1BWP12T U1563 ( .A1(n1197), .A2(n1045), .B1(n1044), .B2(n967), .C1(
        n1043), .C2(n966), .ZN(register_file_inst1_n2441) );
  INVD1BWP12T U1564 ( .I(register_file_inst1_r1_16_), .ZN(n1206) );
  OAI222D1BWP12T U1565 ( .A1(n1206), .A2(n1093), .B1(n1094), .B2(n967), .C1(
        n1095), .C2(n966), .ZN(register_file_inst1_n2601) );
  INVD1BWP12T U1566 ( .I(register_file_inst1_r5_16_), .ZN(n1196) );
  OAI222D1BWP12T U1567 ( .A1(n1196), .A2(n1096), .B1(n1097), .B2(n967), .C1(
        n1098), .C2(n966), .ZN(register_file_inst1_n2473) );
  INVD1BWP12T U1568 ( .I(register_file_inst1_r7_16_), .ZN(n1208) );
  OAI222D1BWP12T U1569 ( .A1(n1208), .A2(n1051), .B1(n1050), .B2(n967), .C1(
        n1049), .C2(n966), .ZN(register_file_inst1_n2409) );
  INVD1BWP12T U1570 ( .I(register_file_inst1_lr_16_), .ZN(n1187) );
  OAI222D1BWP12T U1571 ( .A1(n1187), .A2(n1082), .B1(n1084), .B2(n967), .C1(
        n1085), .C2(n966), .ZN(register_file_inst1_n2217) );
  INVD1BWP12T U1572 ( .I(register_file_inst1_r0_19_), .ZN(n1528) );
  OAI222D1BWP12T U1573 ( .A1(n1528), .A2(n1086), .B1(n1088), .B2(n971), .C1(
        n1089), .C2(n970), .ZN(register_file_inst1_n2636) );
  INVD1BWP12T U1574 ( .I(register_file_inst1_r4_19_), .ZN(n1540) );
  OAI222D1BWP12T U1575 ( .A1(n1540), .A2(n1090), .B1(n1091), .B2(n971), .C1(
        n1092), .C2(n970), .ZN(register_file_inst1_n2508) );
  OAI222D1BWP12T U1576 ( .A1(n1532), .A2(n1093), .B1(n1094), .B2(n971), .C1(
        n1095), .C2(n970), .ZN(register_file_inst1_n2604) );
  OAI222D1BWP12T U1577 ( .A1(n1531), .A2(n1051), .B1(n1050), .B2(n971), .C1(
        n1049), .C2(n970), .ZN(register_file_inst1_n2412) );
  INVD1BWP12T U1578 ( .I(register_file_inst1_r6_19_), .ZN(n1543) );
  OAI222D1BWP12T U1579 ( .A1(n1543), .A2(n1045), .B1(n1044), .B2(n971), .C1(
        n1043), .C2(n970), .ZN(register_file_inst1_n2444) );
  INVD1BWP12T U1580 ( .I(register_file_inst1_r5_19_), .ZN(n1542) );
  OAI222D1BWP12T U1581 ( .A1(n1542), .A2(n1096), .B1(n1097), .B2(n971), .C1(
        n1098), .C2(n970), .ZN(register_file_inst1_n2476) );
  INVD1BWP12T U1582 ( .I(register_file_inst1_r3_19_), .ZN(n1529) );
  OAI222D1BWP12T U1583 ( .A1(n1529), .A2(n1064), .B1(n1066), .B2(n971), .C1(
        n1067), .C2(n970), .ZN(register_file_inst1_n2540) );
  CKND0BWP12T U1584 ( .I(register_file_inst1_r2_19_), .ZN(n603) );
  OAI222D1BWP12T U1585 ( .A1(n603), .A2(n1060), .B1(n1062), .B2(n971), .C1(
        n1063), .C2(n970), .ZN(register_file_inst1_n2572) );
  INVD1BWP12T U1586 ( .I(register_file_inst1_r10_19_), .ZN(n1539) );
  OAI222D1BWP12T U1587 ( .A1(n1539), .A2(n1068), .B1(n1069), .B2(n971), .C1(
        n1070), .C2(n970), .ZN(register_file_inst1_n2316) );
  CKND0BWP12T U1588 ( .I(register_file_inst1_r6_22_), .ZN(n604) );
  OAI222D1BWP12T U1589 ( .A1(n604), .A2(n1045), .B1(n1044), .B2(n989), .C1(
        n1043), .C2(n988), .ZN(register_file_inst1_n2447) );
  OAI222D1BWP12T U1590 ( .A1(n605), .A2(n1051), .B1(n1050), .B2(n989), .C1(
        n1049), .C2(n988), .ZN(register_file_inst1_n2415) );
  CKND0BWP12T U1591 ( .I(register_file_inst1_tmp1_28_), .ZN(n606) );
  OAI222D1BWP12T U1592 ( .A1(n606), .A2(n1027), .B1(n1026), .B2(n1012), .C1(
        n2168), .C2(n1011), .ZN(register_file_inst1_n2165) );
  CKND0BWP12T U1593 ( .I(register_file_inst1_r2_28_), .ZN(n607) );
  OAI222D1BWP12T U1594 ( .A1(n607), .A2(n1060), .B1(n1062), .B2(n1012), .C1(
        n1063), .C2(n1011), .ZN(register_file_inst1_n2581) );
  CKND0BWP12T U1595 ( .I(register_file_inst1_r3_28_), .ZN(n608) );
  OAI222D1BWP12T U1596 ( .A1(n608), .A2(n1064), .B1(n1066), .B2(n1012), .C1(
        n1067), .C2(n1011), .ZN(register_file_inst1_n2549) );
  INVD1BWP12T U1597 ( .I(register_file_inst1_r10_28_), .ZN(n1577) );
  OAI222D1BWP12T U1598 ( .A1(n1577), .A2(n1068), .B1(n1069), .B2(n1012), .C1(
        n1070), .C2(n1011), .ZN(register_file_inst1_n2325) );
  OAI222D1BWP12T U1599 ( .A1(n1579), .A2(n1021), .B1(n964), .B2(n1012), .C1(
        n1019), .C2(n1011), .ZN(register_file_inst1_n2293) );
  CKND0BWP12T U1600 ( .I(register_file_inst1_r2_29_), .ZN(n609) );
  OAI222D1BWP12T U1601 ( .A1(n609), .A2(n1060), .B1(n1062), .B2(n1031), .C1(
        n1063), .C2(n1030), .ZN(register_file_inst1_n2582) );
  INVD1BWP12T U1602 ( .I(register_file_inst1_r10_29_), .ZN(n1604) );
  OAI222D1BWP12T U1603 ( .A1(n1604), .A2(n1068), .B1(n1069), .B2(n1031), .C1(
        n1070), .C2(n1030), .ZN(register_file_inst1_n2326) );
  CKND0BWP12T U1604 ( .I(register_file_inst1_r3_29_), .ZN(n610) );
  OAI222D1BWP12T U1605 ( .A1(n610), .A2(n1064), .B1(n1066), .B2(n1031), .C1(
        n1067), .C2(n1030), .ZN(register_file_inst1_n2550) );
  OAI222D1BWP12T U1606 ( .A1(n1617), .A2(n1021), .B1(n1020), .B2(n1055), .C1(
        n1019), .C2(n1054), .ZN(register_file_inst1_n2295) );
  CKND0BWP12T U1607 ( .I(register_file_inst1_tmp1_30_), .ZN(n611) );
  OAI222D1BWP12T U1608 ( .A1(n611), .A2(n1027), .B1(n1026), .B2(n1055), .C1(
        n2168), .C2(n1054), .ZN(register_file_inst1_n2167) );
  INVD1BWP12T U1609 ( .I(register_file_inst1_r11_31_), .ZN(n1645) );
  OAI222D1BWP12T U1610 ( .A1(n1019), .A2(n1103), .B1(n964), .B2(n1101), .C1(
        n1645), .C2(n1021), .ZN(register_file_inst1_n2296) );
  CKND0BWP12T U1611 ( .I(register_file_inst1_r6_31_), .ZN(n612) );
  OAI222D1BWP12T U1612 ( .A1(n1043), .A2(n1103), .B1(n1044), .B2(n1101), .C1(
        n612), .C2(n1045), .ZN(register_file_inst1_n2456) );
  INVD1BWP12T U1613 ( .I(register_file_inst1_r7_31_), .ZN(n1632) );
  OAI222D1BWP12T U1614 ( .A1(n1049), .A2(n1103), .B1(n1050), .B2(n1101), .C1(
        n1632), .C2(n1051), .ZN(register_file_inst1_n2424) );
  CKND0BWP12T U1615 ( .I(register_file_inst1_tmp1_31_), .ZN(n613) );
  OAI222D1BWP12T U1616 ( .A1(n2168), .A2(n1103), .B1(n1026), .B2(n1101), .C1(
        n613), .C2(n1027), .ZN(register_file_inst1_n2168) );
  NR2D1BWP12T U1617 ( .A1(n2322), .A2(n2320), .ZN(n1939) );
  ND2D1BWP12T U1618 ( .A1(n615), .A2(n614), .ZN(n934) );
  CKND0BWP12T U1619 ( .I(memory_interface_inst1_fsm_state_2_), .ZN(n616) );
  OAI21D0BWP12T U1620 ( .A1(n617), .A2(n616), .B(n2247), .ZN(n634) );
  ND2D1BWP12T U1621 ( .A1(n934), .A2(n634), .ZN(n2039) );
  NR2D1BWP12T U1622 ( .A1(n2323), .A2(n2321), .ZN(n1940) );
  NR2D1BWP12T U1623 ( .A1(n2088), .A2(n2094), .ZN(n1944) );
  INVD1BWP12T U1624 ( .I(n1944), .ZN(n1858) );
  INVD1BWP12T U1625 ( .I(n975), .ZN(n2035) );
  CKND1BWP12T U1626 ( .I(n934), .ZN(n860) );
  NR2D1BWP12T U1627 ( .A1(n860), .A2(n618), .ZN(n2045) );
  CKND2D0BWP12T U1628 ( .A1(n2251), .A2(n2041), .ZN(n633) );
  NR2D1BWP12T U1629 ( .A1(n633), .A2(n2044), .ZN(n636) );
  INVD1BWP12T U1630 ( .I(n636), .ZN(n619) );
  OAI21D1BWP12T U1631 ( .A1(n2332), .A2(n619), .B(n2045), .ZN(
        MEMCTRL_MEM_to_mem_write_enable) );
  INVD1BWP12T U1632 ( .I(n633), .ZN(n620) );
  AOI31D1BWP12T U1633 ( .A1(n2042), .A2(n634), .A3(n621), .B(n620), .ZN(n753)
         );
  AOI22D0BWP12T U1634 ( .A1(n772), .A2(RF_MEMCTRL_data_reg[6]), .B1(n753), 
        .B2(memory_interface_inst1_delay_data_in32[6]), .ZN(n632) );
  AOI22D0BWP12T U1635 ( .A1(register_file_inst1_r6_22_), .A2(n839), .B1(
        register_file_inst1_r4_22_), .B2(n838), .ZN(n625) );
  AOI22D0BWP12T U1636 ( .A1(register_file_inst1_r7_22_), .A2(n841), .B1(
        register_file_inst1_r2_22_), .B2(n840), .ZN(n624) );
  AOI22D0BWP12T U1637 ( .A1(register_file_inst1_r0_22_), .A2(n843), .B1(
        register_file_inst1_r3_22_), .B2(n842), .ZN(n623) );
  AOI22D0BWP12T U1638 ( .A1(register_file_inst1_r1_22_), .A2(n845), .B1(
        register_file_inst1_r5_22_), .B2(n844), .ZN(n622) );
  ND4D1BWP12T U1639 ( .A1(n625), .A2(n624), .A3(n623), .A4(n622), .ZN(n630) );
  AOI22D0BWP12T U1640 ( .A1(register_file_inst1_lr_22_), .A2(n1947), .B1(
        register_file_inst1_r10_22_), .B2(n852), .ZN(n628) );
  AOI22D0BWP12T U1641 ( .A1(STACK_RF_next_sp[22]), .A2(n1927), .B1(
        register_file_inst1_r11_22_), .B2(n851), .ZN(n627) );
  AOI22D0BWP12T U1642 ( .A1(register_file_inst1_r9_22_), .A2(n850), .B1(
        register_file_inst1_r12_22_), .B2(n398), .ZN(n626) );
  ND4D1BWP12T U1643 ( .A1(n628), .A2(n2000), .A3(n627), .A4(n626), .ZN(n629)
         );
  AO21D1BWP12T U1644 ( .A1(n2306), .A2(n630), .B(n629), .Z(
        RF_MEMCTRL_data_reg[22]) );
  AOI22D1BWP12T U1645 ( .A1(n860), .A2(
        memory_interface_inst1_delay_data_in32[22]), .B1(n763), .B2(
        RF_MEMCTRL_data_reg[22]), .ZN(n631) );
  ND2D1BWP12T U1646 ( .A1(n632), .A2(n631), .ZN(MEMCTRL_MEM_to_mem_data[14])
         );
  INVD1BWP12T U1647 ( .I(MEMCTRL_load_in), .ZN(n635) );
  AOI22D1BWP12T U1648 ( .A1(n636), .A2(n635), .B1(n634), .B2(n633), .ZN(
        MEMCTRL_MEM_to_mem_read_enable) );
  AOI22D1BWP12T U1649 ( .A1(n2297), .A2(
        memory_interface_inst1_delay_addr_single[4]), .B1(
        MEMCTRL_IN_address[4]), .B2(n2043), .ZN(n638) );
  AN2XD0BWP12T U1650 ( .A1(memory_interface_inst1_delay_addr_for_adder_1_), 
        .A2(memory_interface_inst1_delay_addr_for_adder_0_), .Z(n768) );
  ND2D1BWP12T U1651 ( .A1(n768), .A2(
        memory_interface_inst1_delay_addr_for_adder_2_), .ZN(n766) );
  INVD1BWP12T U1652 ( .I(memory_interface_inst1_delay_addr_for_adder_3_), .ZN(
        n711) );
  NR2D1BWP12T U1653 ( .A1(n766), .A2(n711), .ZN(n710) );
  NR2D1BWP12T U1654 ( .A1(n2297), .A2(n2043), .ZN(n767) );
  ND2D1BWP12T U1655 ( .A1(n710), .A2(
        memory_interface_inst1_delay_addr_for_adder_4_), .ZN(n700) );
  OAI211D1BWP12T U1656 ( .A1(n710), .A2(
        memory_interface_inst1_delay_addr_for_adder_4_), .B(n767), .C(n700), 
        .ZN(n637) );
  ND2D1BWP12T U1657 ( .A1(n638), .A2(n637), .ZN(MEMCTRL_MEM_to_mem_address[4])
         );
  INR2D1BWP12T U1658 ( .A1(n753), .B1(n2297), .ZN(n771) );
  AOI22D1BWP12T U1659 ( .A1(n2297), .A2(MEM_MEMCTRL_from_mem_data[2]), .B1(
        n771), .B2(memory_interface_inst1_delay_data_in32[10]), .ZN(n640) );
  AOI22D0BWP12T U1660 ( .A1(n860), .A2(
        memory_interface_inst1_delay_data_in32[26]), .B1(n772), .B2(
        RF_MEMCTRL_data_reg[10]), .ZN(n639) );
  ND2D1BWP12T U1661 ( .A1(n640), .A2(n639), .ZN(MEMCTRL_MEM_to_mem_data[2]) );
  NR2D1BWP12T U1662 ( .A1(memory_interface_inst1_delay_addr_for_adder_0_), 
        .A2(memory_interface_inst1_delay_addr_for_adder_1_), .ZN(n642) );
  INVD1BWP12T U1663 ( .I(n767), .ZN(n728) );
  AOI22D1BWP12T U1664 ( .A1(n2297), .A2(
        memory_interface_inst1_delay_addr_single[1]), .B1(
        MEMCTRL_IN_address[1]), .B2(n2043), .ZN(n641) );
  OAI31D1BWP12T U1665 ( .A1(n768), .A2(n642), .A3(n728), .B(n641), .ZN(
        MEMCTRL_MEM_to_mem_address[1]) );
  AOI22D0BWP12T U1666 ( .A1(n772), .A2(RF_MEMCTRL_data_reg[3]), .B1(n753), 
        .B2(memory_interface_inst1_delay_data_in32[3]), .ZN(n653) );
  AOI22D0BWP12T U1667 ( .A1(register_file_inst1_r6_19_), .A2(n839), .B1(
        register_file_inst1_r4_19_), .B2(n838), .ZN(n646) );
  AOI22D0BWP12T U1668 ( .A1(register_file_inst1_r7_19_), .A2(n841), .B1(
        register_file_inst1_r2_19_), .B2(n840), .ZN(n645) );
  AOI22D0BWP12T U1669 ( .A1(register_file_inst1_r0_19_), .A2(n843), .B1(
        register_file_inst1_r3_19_), .B2(n842), .ZN(n644) );
  AOI22D0BWP12T U1670 ( .A1(register_file_inst1_r1_19_), .A2(n845), .B1(
        register_file_inst1_r5_19_), .B2(n844), .ZN(n643) );
  ND4D1BWP12T U1671 ( .A1(n646), .A2(n645), .A3(n644), .A4(n643), .ZN(n651) );
  AOI22D0BWP12T U1672 ( .A1(register_file_inst1_lr_19_), .A2(n1947), .B1(
        register_file_inst1_r10_19_), .B2(n852), .ZN(n649) );
  AOI22D0BWP12T U1673 ( .A1(STACK_RF_next_sp[19]), .A2(n1927), .B1(
        register_file_inst1_r11_19_), .B2(n851), .ZN(n648) );
  AOI22D0BWP12T U1674 ( .A1(register_file_inst1_r9_19_), .A2(n850), .B1(
        register_file_inst1_r12_19_), .B2(n398), .ZN(n647) );
  ND4D1BWP12T U1675 ( .A1(n649), .A2(n2002), .A3(n648), .A4(n647), .ZN(n650)
         );
  AO21D1BWP12T U1676 ( .A1(n2306), .A2(n651), .B(n650), .Z(
        RF_MEMCTRL_data_reg[19]) );
  AOI22D1BWP12T U1677 ( .A1(n860), .A2(
        memory_interface_inst1_delay_data_in32[19]), .B1(n763), .B2(
        RF_MEMCTRL_data_reg[19]), .ZN(n652) );
  ND2D1BWP12T U1678 ( .A1(n653), .A2(n652), .ZN(MEMCTRL_MEM_to_mem_data[11])
         );
  AOI22D0BWP12T U1679 ( .A1(n772), .A2(RF_MEMCTRL_data_reg[2]), .B1(n753), 
        .B2(memory_interface_inst1_delay_data_in32[2]), .ZN(n664) );
  AOI22D0BWP12T U1680 ( .A1(register_file_inst1_r6_18_), .A2(n839), .B1(
        register_file_inst1_r4_18_), .B2(n838), .ZN(n657) );
  AOI22D0BWP12T U1681 ( .A1(register_file_inst1_r7_18_), .A2(n841), .B1(
        register_file_inst1_r2_18_), .B2(n840), .ZN(n656) );
  AOI22D0BWP12T U1682 ( .A1(register_file_inst1_r0_18_), .A2(n843), .B1(
        register_file_inst1_r3_18_), .B2(n842), .ZN(n655) );
  AOI22D0BWP12T U1683 ( .A1(register_file_inst1_r1_18_), .A2(n845), .B1(
        register_file_inst1_r5_18_), .B2(n844), .ZN(n654) );
  ND4D1BWP12T U1684 ( .A1(n657), .A2(n656), .A3(n655), .A4(n654), .ZN(n662) );
  OAI22D0BWP12T U1685 ( .A1(n745), .A2(n1113), .B1(n1135), .B2(n744), .ZN(n660) );
  AOI22D0BWP12T U1686 ( .A1(register_file_inst1_r8_18_), .A2(n1948), .B1(
        register_file_inst1_r10_18_), .B2(n852), .ZN(n659) );
  AOI22D0BWP12T U1687 ( .A1(register_file_inst1_r9_18_), .A2(n850), .B1(
        register_file_inst1_r12_18_), .B2(n398), .ZN(n658) );
  IND4D1BWP12T U1688 ( .A1(n660), .B1(n2003), .B2(n659), .B3(n658), .ZN(n661)
         );
  AO21D1BWP12T U1689 ( .A1(n2306), .A2(n662), .B(n661), .Z(
        RF_MEMCTRL_data_reg[18]) );
  AOI22D1BWP12T U1690 ( .A1(n860), .A2(
        memory_interface_inst1_delay_data_in32[18]), .B1(n763), .B2(
        RF_MEMCTRL_data_reg[18]), .ZN(n663) );
  ND2D1BWP12T U1691 ( .A1(n664), .A2(n663), .ZN(MEMCTRL_MEM_to_mem_data[10])
         );
  INVD1BWP12T U1692 ( .I(memory_interface_inst1_delay_addr_for_adder_0_), .ZN(
        n665) );
  AO222D1BWP12T U1693 ( .A1(n2043), .A2(MEMCTRL_IN_address[0]), .B1(n665), 
        .B2(n767), .C1(n2297), .C2(memory_interface_inst1_delay_addr_single[0]), .Z(MEMCTRL_MEM_to_mem_address[0]) );
  AOI22D0BWP12T U1694 ( .A1(n772), .A2(RF_MEMCTRL_data_reg[4]), .B1(n753), 
        .B2(memory_interface_inst1_delay_data_in32[4]), .ZN(n676) );
  AOI22D0BWP12T U1695 ( .A1(register_file_inst1_r6_20_), .A2(n839), .B1(
        register_file_inst1_r4_20_), .B2(n838), .ZN(n669) );
  AOI22D0BWP12T U1696 ( .A1(register_file_inst1_r7_20_), .A2(n841), .B1(
        register_file_inst1_r2_20_), .B2(n840), .ZN(n668) );
  AOI22D0BWP12T U1697 ( .A1(register_file_inst1_r0_20_), .A2(n843), .B1(
        register_file_inst1_r3_20_), .B2(n842), .ZN(n667) );
  AOI22D0BWP12T U1698 ( .A1(register_file_inst1_r1_20_), .A2(n845), .B1(
        register_file_inst1_r5_20_), .B2(n844), .ZN(n666) );
  ND4D1BWP12T U1699 ( .A1(n669), .A2(n668), .A3(n667), .A4(n666), .ZN(n674) );
  AOI22D0BWP12T U1700 ( .A1(STACK_RF_next_sp[20]), .A2(n1927), .B1(
        register_file_inst1_r8_20_), .B2(n1948), .ZN(n672) );
  AOI22D0BWP12T U1701 ( .A1(register_file_inst1_r10_20_), .A2(n852), .B1(
        register_file_inst1_r11_20_), .B2(n851), .ZN(n671) );
  AOI22D0BWP12T U1702 ( .A1(register_file_inst1_r9_20_), .A2(n850), .B1(
        register_file_inst1_r12_20_), .B2(n398), .ZN(n670) );
  ND4D1BWP12T U1703 ( .A1(n1984), .A2(n672), .A3(n671), .A4(n670), .ZN(n673)
         );
  AO21D1BWP12T U1704 ( .A1(n2306), .A2(n674), .B(n673), .Z(
        RF_MEMCTRL_data_reg[20]) );
  AOI22D1BWP12T U1705 ( .A1(n860), .A2(
        memory_interface_inst1_delay_data_in32[20]), .B1(n763), .B2(
        RF_MEMCTRL_data_reg[20]), .ZN(n675) );
  ND2D1BWP12T U1706 ( .A1(n676), .A2(n675), .ZN(MEMCTRL_MEM_to_mem_data[12])
         );
  AOI22D0BWP12T U1707 ( .A1(n772), .A2(RF_MEMCTRL_data_reg[7]), .B1(n753), 
        .B2(memory_interface_inst1_delay_data_in32[7]), .ZN(n687) );
  AOI22D0BWP12T U1708 ( .A1(register_file_inst1_r6_23_), .A2(n839), .B1(
        register_file_inst1_r4_23_), .B2(n838), .ZN(n680) );
  AOI22D0BWP12T U1709 ( .A1(register_file_inst1_r7_23_), .A2(n841), .B1(
        register_file_inst1_r2_23_), .B2(n840), .ZN(n679) );
  AOI22D0BWP12T U1710 ( .A1(register_file_inst1_r0_23_), .A2(n843), .B1(
        register_file_inst1_r3_23_), .B2(n842), .ZN(n678) );
  AOI22D0BWP12T U1711 ( .A1(register_file_inst1_r1_23_), .A2(n845), .B1(
        register_file_inst1_r5_23_), .B2(n844), .ZN(n677) );
  ND4D1BWP12T U1712 ( .A1(n680), .A2(n679), .A3(n678), .A4(n677), .ZN(n685) );
  AOI22D0BWP12T U1713 ( .A1(STACK_RF_next_sp[23]), .A2(n1927), .B1(
        register_file_inst1_r9_23_), .B2(n850), .ZN(n683) );
  AOI22D0BWP12T U1714 ( .A1(register_file_inst1_r8_23_), .A2(n1948), .B1(
        register_file_inst1_r11_23_), .B2(n851), .ZN(n682) );
  AOI22D0BWP12T U1715 ( .A1(register_file_inst1_r12_23_), .A2(n398), .B1(
        register_file_inst1_r10_23_), .B2(n852), .ZN(n681) );
  ND4D1BWP12T U1716 ( .A1(n683), .A2(n1999), .A3(n682), .A4(n681), .ZN(n684)
         );
  AO21D1BWP12T U1717 ( .A1(n2306), .A2(n685), .B(n684), .Z(
        RF_MEMCTRL_data_reg[23]) );
  AOI22D1BWP12T U1718 ( .A1(n860), .A2(
        memory_interface_inst1_delay_data_in32[23]), .B1(n763), .B2(
        RF_MEMCTRL_data_reg[23]), .ZN(n686) );
  ND2D1BWP12T U1719 ( .A1(n687), .A2(n686), .ZN(MEMCTRL_MEM_to_mem_data[15])
         );
  AOI22D0BWP12T U1720 ( .A1(n772), .A2(RF_MEMCTRL_data_reg[5]), .B1(n753), 
        .B2(memory_interface_inst1_delay_data_in32[5]), .ZN(n698) );
  AOI22D0BWP12T U1721 ( .A1(register_file_inst1_r6_21_), .A2(n839), .B1(
        register_file_inst1_r4_21_), .B2(n838), .ZN(n691) );
  AOI22D0BWP12T U1722 ( .A1(register_file_inst1_r7_21_), .A2(n841), .B1(
        register_file_inst1_r2_21_), .B2(n840), .ZN(n690) );
  AOI22D0BWP12T U1723 ( .A1(register_file_inst1_r0_21_), .A2(n843), .B1(
        register_file_inst1_r3_21_), .B2(n842), .ZN(n689) );
  AOI22D0BWP12T U1724 ( .A1(register_file_inst1_r1_21_), .A2(n845), .B1(
        register_file_inst1_r5_21_), .B2(n844), .ZN(n688) );
  ND4D1BWP12T U1725 ( .A1(n691), .A2(n690), .A3(n689), .A4(n688), .ZN(n696) );
  AOI22D0BWP12T U1726 ( .A1(STACK_RF_next_sp[21]), .A2(n1927), .B1(
        register_file_inst1_r10_21_), .B2(n852), .ZN(n694) );
  AOI22D0BWP12T U1727 ( .A1(register_file_inst1_r8_21_), .A2(n1948), .B1(
        register_file_inst1_r11_21_), .B2(n851), .ZN(n693) );
  AOI22D0BWP12T U1728 ( .A1(register_file_inst1_r9_21_), .A2(n850), .B1(
        register_file_inst1_r12_21_), .B2(n398), .ZN(n692) );
  ND4D1BWP12T U1729 ( .A1(n694), .A2(n2001), .A3(n693), .A4(n692), .ZN(n695)
         );
  AO21D1BWP12T U1730 ( .A1(n2306), .A2(n696), .B(n695), .Z(
        RF_MEMCTRL_data_reg[21]) );
  AOI22D1BWP12T U1731 ( .A1(n860), .A2(
        memory_interface_inst1_delay_data_in32[21]), .B1(n763), .B2(
        RF_MEMCTRL_data_reg[21]), .ZN(n697) );
  ND2D1BWP12T U1732 ( .A1(n698), .A2(n697), .ZN(MEMCTRL_MEM_to_mem_data[13])
         );
  AOI22D1BWP12T U1733 ( .A1(n2297), .A2(
        memory_interface_inst1_delay_addr_single[5]), .B1(
        MEMCTRL_IN_address[5]), .B2(n2043), .ZN(n702) );
  INVD1BWP12T U1734 ( .I(memory_interface_inst1_delay_addr_for_adder_5_), .ZN(
        n699) );
  NR2D1BWP12T U1735 ( .A1(n700), .A2(n699), .ZN(n723) );
  AO211D1BWP12T U1736 ( .A1(n700), .A2(n699), .B(n723), .C(n728), .Z(n701) );
  ND2D1BWP12T U1737 ( .A1(n702), .A2(n701), .ZN(MEMCTRL_MEM_to_mem_address[5])
         );
  AOI22D1BWP12T U1738 ( .A1(n2297), .A2(
        memory_interface_inst1_delay_addr_single[10]), .B1(
        MEMCTRL_IN_address[10]), .B2(n2043), .ZN(n704) );
  ND2D1BWP12T U1739 ( .A1(n723), .A2(
        memory_interface_inst1_delay_addr_for_adder_6_), .ZN(n731) );
  INVD1BWP12T U1740 ( .I(memory_interface_inst1_delay_addr_for_adder_7_), .ZN(
        n730) );
  NR2D1BWP12T U1741 ( .A1(n731), .A2(n730), .ZN(n729) );
  ND2D1BWP12T U1742 ( .A1(n729), .A2(
        memory_interface_inst1_delay_addr_for_adder_8_), .ZN(n720) );
  INVD1BWP12T U1743 ( .I(memory_interface_inst1_delay_addr_for_adder_9_), .ZN(
        n715) );
  NR2D1BWP12T U1744 ( .A1(n720), .A2(n715), .ZN(n714) );
  ND2D1BWP12T U1745 ( .A1(n714), .A2(
        memory_interface_inst1_delay_addr_for_adder_10_), .ZN(n707) );
  OAI211D1BWP12T U1746 ( .A1(n714), .A2(
        memory_interface_inst1_delay_addr_for_adder_10_), .B(n767), .C(n707), 
        .ZN(n703) );
  ND2D1BWP12T U1747 ( .A1(n704), .A2(n703), .ZN(MEMCTRL_MEM_to_mem_address[10]) );
  AOI22D1BWP12T U1748 ( .A1(n2297), .A2(MEM_MEMCTRL_from_mem_data[0]), .B1(
        n771), .B2(memory_interface_inst1_delay_data_in32[8]), .ZN(n706) );
  AOI22D0BWP12T U1749 ( .A1(n860), .A2(
        memory_interface_inst1_delay_data_in32[24]), .B1(n772), .B2(
        RF_MEMCTRL_data_reg[8]), .ZN(n705) );
  ND2D1BWP12T U1750 ( .A1(n706), .A2(n705), .ZN(MEMCTRL_MEM_to_mem_data[0]) );
  MAOI22D0BWP12T U1751 ( .A1(memory_interface_inst1_delay_addr_for_adder_11_), 
        .A2(n707), .B1(memory_interface_inst1_delay_addr_for_adder_11_), .B2(
        n707), .ZN(n709) );
  AOI22D1BWP12T U1752 ( .A1(n2297), .A2(
        memory_interface_inst1_delay_addr_single[11]), .B1(
        MEMCTRL_IN_address[11]), .B2(n2043), .ZN(n708) );
  OAI21D1BWP12T U1753 ( .A1(n728), .A2(n709), .B(n708), .ZN(
        MEMCTRL_MEM_to_mem_address[11]) );
  AOI22D1BWP12T U1754 ( .A1(n2297), .A2(
        memory_interface_inst1_delay_addr_single[3]), .B1(
        MEMCTRL_IN_address[3]), .B2(n2043), .ZN(n713) );
  AO211D1BWP12T U1755 ( .A1(n766), .A2(n711), .B(n710), .C(n728), .Z(n712) );
  ND2D1BWP12T U1756 ( .A1(n713), .A2(n712), .ZN(MEMCTRL_MEM_to_mem_address[3])
         );
  AOI22D1BWP12T U1757 ( .A1(n2297), .A2(
        memory_interface_inst1_delay_addr_single[9]), .B1(
        MEMCTRL_IN_address[9]), .B2(n2043), .ZN(n717) );
  AO211D1BWP12T U1758 ( .A1(n720), .A2(n715), .B(n714), .C(n728), .Z(n716) );
  ND2D1BWP12T U1759 ( .A1(n717), .A2(n716), .ZN(MEMCTRL_MEM_to_mem_address[9])
         );
  AOI22D1BWP12T U1760 ( .A1(n2297), .A2(MEM_MEMCTRL_from_mem_data[1]), .B1(
        n771), .B2(memory_interface_inst1_delay_data_in32[9]), .ZN(n719) );
  AOI22D0BWP12T U1761 ( .A1(n860), .A2(
        memory_interface_inst1_delay_data_in32[25]), .B1(n772), .B2(
        RF_MEMCTRL_data_reg[9]), .ZN(n718) );
  ND2D1BWP12T U1762 ( .A1(n719), .A2(n718), .ZN(MEMCTRL_MEM_to_mem_data[1]) );
  AOI22D1BWP12T U1763 ( .A1(n2297), .A2(
        memory_interface_inst1_delay_addr_single[8]), .B1(
        MEMCTRL_IN_address[8]), .B2(n2043), .ZN(n722) );
  OAI211D1BWP12T U1764 ( .A1(n729), .A2(
        memory_interface_inst1_delay_addr_for_adder_8_), .B(n767), .C(n720), 
        .ZN(n721) );
  ND2D1BWP12T U1765 ( .A1(n722), .A2(n721), .ZN(MEMCTRL_MEM_to_mem_address[8])
         );
  AOI22D1BWP12T U1766 ( .A1(n2297), .A2(
        memory_interface_inst1_delay_addr_single[6]), .B1(
        MEMCTRL_IN_address[6]), .B2(n2043), .ZN(n725) );
  OAI211D1BWP12T U1767 ( .A1(n723), .A2(
        memory_interface_inst1_delay_addr_for_adder_6_), .B(n767), .C(n731), 
        .ZN(n724) );
  ND2D1BWP12T U1768 ( .A1(n725), .A2(n724), .ZN(MEMCTRL_MEM_to_mem_address[6])
         );
  AOI22D1BWP12T U1769 ( .A1(n2297), .A2(MEM_MEMCTRL_from_mem_data[5]), .B1(
        n771), .B2(memory_interface_inst1_delay_data_in32[13]), .ZN(n727) );
  AOI22D0BWP12T U1770 ( .A1(n860), .A2(
        memory_interface_inst1_delay_data_in32[29]), .B1(n772), .B2(
        RF_MEMCTRL_data_reg[13]), .ZN(n726) );
  ND2D1BWP12T U1771 ( .A1(n727), .A2(n726), .ZN(MEMCTRL_MEM_to_mem_data[5]) );
  AOI22D1BWP12T U1772 ( .A1(n2297), .A2(
        memory_interface_inst1_delay_addr_single[7]), .B1(
        MEMCTRL_IN_address[7]), .B2(n2043), .ZN(n733) );
  AO211D1BWP12T U1773 ( .A1(n731), .A2(n730), .B(n729), .C(n728), .Z(n732) );
  ND2D1BWP12T U1774 ( .A1(n733), .A2(n732), .ZN(MEMCTRL_MEM_to_mem_address[7])
         );
  AOI22D1BWP12T U1775 ( .A1(n2297), .A2(MEM_MEMCTRL_from_mem_data[3]), .B1(
        n771), .B2(memory_interface_inst1_delay_data_in32[11]), .ZN(n735) );
  AOI22D0BWP12T U1776 ( .A1(n860), .A2(
        memory_interface_inst1_delay_data_in32[27]), .B1(n772), .B2(
        RF_MEMCTRL_data_reg[11]), .ZN(n734) );
  ND2D1BWP12T U1777 ( .A1(n735), .A2(n734), .ZN(MEMCTRL_MEM_to_mem_data[3]) );
  AOI22D1BWP12T U1778 ( .A1(n2297), .A2(MEM_MEMCTRL_from_mem_data[7]), .B1(
        n771), .B2(memory_interface_inst1_delay_data_in32[15]), .ZN(n737) );
  AOI22D0BWP12T U1779 ( .A1(n860), .A2(
        memory_interface_inst1_delay_data_in32[31]), .B1(n772), .B2(
        RF_MEMCTRL_data_reg[15]), .ZN(n736) );
  ND2D1BWP12T U1780 ( .A1(n737), .A2(n736), .ZN(MEMCTRL_MEM_to_mem_data[7]) );
  AOI22D1BWP12T U1781 ( .A1(n2297), .A2(MEM_MEMCTRL_from_mem_data[4]), .B1(
        n771), .B2(memory_interface_inst1_delay_data_in32[12]), .ZN(n739) );
  AOI22D0BWP12T U1782 ( .A1(n860), .A2(
        memory_interface_inst1_delay_data_in32[28]), .B1(n772), .B2(
        RF_MEMCTRL_data_reg[12]), .ZN(n738) );
  ND2D1BWP12T U1783 ( .A1(n739), .A2(n738), .ZN(MEMCTRL_MEM_to_mem_data[4]) );
  AOI22D0BWP12T U1784 ( .A1(n772), .A2(RF_MEMCTRL_data_reg[0]), .B1(n753), 
        .B2(memory_interface_inst1_delay_data_in32[0]), .ZN(n752) );
  AOI22D0BWP12T U1785 ( .A1(register_file_inst1_r6_16_), .A2(n839), .B1(
        register_file_inst1_r4_16_), .B2(n838), .ZN(n743) );
  AOI22D0BWP12T U1786 ( .A1(register_file_inst1_r7_16_), .A2(n841), .B1(
        register_file_inst1_r2_16_), .B2(n840), .ZN(n742) );
  AOI22D0BWP12T U1787 ( .A1(register_file_inst1_r0_16_), .A2(n843), .B1(
        register_file_inst1_r3_16_), .B2(n842), .ZN(n741) );
  AOI22D0BWP12T U1788 ( .A1(register_file_inst1_r1_16_), .A2(n845), .B1(
        register_file_inst1_r5_16_), .B2(n844), .ZN(n740) );
  ND4D1BWP12T U1789 ( .A1(n743), .A2(n742), .A3(n741), .A4(n740), .ZN(n750) );
  INVD1BWP12T U1790 ( .I(STACK_RF_next_sp[16]), .ZN(n1183) );
  INVD1BWP12T U1791 ( .I(register_file_inst1_r11_16_), .ZN(n1205) );
  OAI22D0BWP12T U1792 ( .A1(n745), .A2(n1183), .B1(n1205), .B2(n744), .ZN(n748) );
  AOI22D0BWP12T U1793 ( .A1(register_file_inst1_r8_16_), .A2(n1948), .B1(
        register_file_inst1_r10_16_), .B2(n852), .ZN(n747) );
  AOI22D0BWP12T U1794 ( .A1(register_file_inst1_r9_16_), .A2(n850), .B1(
        register_file_inst1_r12_16_), .B2(n398), .ZN(n746) );
  IND4D1BWP12T U1795 ( .A1(n748), .B1(n2005), .B2(n747), .B3(n746), .ZN(n749)
         );
  AO21D1BWP12T U1796 ( .A1(n2306), .A2(n750), .B(n749), .Z(
        RF_MEMCTRL_data_reg[16]) );
  AOI22D1BWP12T U1797 ( .A1(n860), .A2(
        memory_interface_inst1_delay_data_in32[16]), .B1(n763), .B2(
        RF_MEMCTRL_data_reg[16]), .ZN(n751) );
  ND2D1BWP12T U1798 ( .A1(n752), .A2(n751), .ZN(MEMCTRL_MEM_to_mem_data[8]) );
  AOI22D0BWP12T U1799 ( .A1(n772), .A2(RF_MEMCTRL_data_reg[1]), .B1(n753), 
        .B2(memory_interface_inst1_delay_data_in32[1]), .ZN(n765) );
  AOI22D0BWP12T U1800 ( .A1(register_file_inst1_r6_17_), .A2(n839), .B1(
        register_file_inst1_r4_17_), .B2(n838), .ZN(n757) );
  AOI22D0BWP12T U1801 ( .A1(register_file_inst1_r7_17_), .A2(n841), .B1(
        register_file_inst1_r2_17_), .B2(n840), .ZN(n756) );
  AOI22D0BWP12T U1802 ( .A1(register_file_inst1_r0_17_), .A2(n843), .B1(
        register_file_inst1_r3_17_), .B2(n842), .ZN(n755) );
  AOI22D0BWP12T U1803 ( .A1(register_file_inst1_r1_17_), .A2(n845), .B1(
        register_file_inst1_r5_17_), .B2(n844), .ZN(n754) );
  ND4D1BWP12T U1804 ( .A1(n757), .A2(n756), .A3(n755), .A4(n754), .ZN(n762) );
  AOI22D0BWP12T U1805 ( .A1(STACK_RF_next_sp[17]), .A2(n1927), .B1(
        register_file_inst1_r10_17_), .B2(n852), .ZN(n760) );
  AOI22D0BWP12T U1806 ( .A1(register_file_inst1_r8_17_), .A2(n1948), .B1(
        register_file_inst1_r11_17_), .B2(n851), .ZN(n759) );
  AOI22D0BWP12T U1807 ( .A1(register_file_inst1_r9_17_), .A2(n850), .B1(
        register_file_inst1_r12_17_), .B2(n398), .ZN(n758) );
  ND4D1BWP12T U1808 ( .A1(n760), .A2(n2004), .A3(n759), .A4(n758), .ZN(n761)
         );
  AO21D1BWP12T U1809 ( .A1(n2306), .A2(n762), .B(n761), .Z(
        RF_MEMCTRL_data_reg[17]) );
  AOI22D1BWP12T U1810 ( .A1(n860), .A2(
        memory_interface_inst1_delay_data_in32[17]), .B1(n763), .B2(
        RF_MEMCTRL_data_reg[17]), .ZN(n764) );
  ND2D1BWP12T U1811 ( .A1(n765), .A2(n764), .ZN(MEMCTRL_MEM_to_mem_data[9]) );
  AOI22D1BWP12T U1812 ( .A1(n2297), .A2(
        memory_interface_inst1_delay_addr_single[2]), .B1(
        MEMCTRL_IN_address[2]), .B2(n2043), .ZN(n770) );
  OAI211D1BWP12T U1813 ( .A1(n768), .A2(
        memory_interface_inst1_delay_addr_for_adder_2_), .B(n767), .C(n766), 
        .ZN(n769) );
  ND2D1BWP12T U1814 ( .A1(n770), .A2(n769), .ZN(MEMCTRL_MEM_to_mem_address[2])
         );
  AOI22D1BWP12T U1815 ( .A1(n2297), .A2(MEM_MEMCTRL_from_mem_data[6]), .B1(
        n771), .B2(memory_interface_inst1_delay_data_in32[14]), .ZN(n774) );
  AOI22D0BWP12T U1816 ( .A1(n860), .A2(
        memory_interface_inst1_delay_data_in32[30]), .B1(n772), .B2(
        RF_MEMCTRL_data_reg[14]), .ZN(n773) );
  ND2D1BWP12T U1817 ( .A1(n774), .A2(n773), .ZN(MEMCTRL_MEM_to_mem_data[6]) );
  AOI22D0BWP12T U1818 ( .A1(register_file_inst1_r6_25_), .A2(n839), .B1(
        register_file_inst1_r4_25_), .B2(n838), .ZN(n778) );
  AOI22D0BWP12T U1819 ( .A1(register_file_inst1_r7_25_), .A2(n841), .B1(
        register_file_inst1_r2_25_), .B2(n840), .ZN(n777) );
  AOI22D0BWP12T U1820 ( .A1(register_file_inst1_r0_25_), .A2(n843), .B1(
        register_file_inst1_r3_25_), .B2(n842), .ZN(n776) );
  AOI22D0BWP12T U1821 ( .A1(register_file_inst1_r1_25_), .A2(n845), .B1(
        register_file_inst1_r5_25_), .B2(n844), .ZN(n775) );
  ND4D1BWP12T U1822 ( .A1(n778), .A2(n777), .A3(n776), .A4(n775), .ZN(n783) );
  AOI22D0BWP12T U1823 ( .A1(STACK_RF_next_sp[25]), .A2(n1927), .B1(
        register_file_inst1_r9_25_), .B2(n850), .ZN(n781) );
  AOI22D0BWP12T U1824 ( .A1(register_file_inst1_r8_25_), .A2(n1948), .B1(
        register_file_inst1_r11_25_), .B2(n851), .ZN(n780) );
  AOI22D0BWP12T U1825 ( .A1(register_file_inst1_r12_25_), .A2(n398), .B1(
        register_file_inst1_r10_25_), .B2(n852), .ZN(n779) );
  ND4D1BWP12T U1826 ( .A1(n781), .A2(n1998), .A3(n780), .A4(n779), .ZN(n782)
         );
  AO21D1BWP12T U1827 ( .A1(n2306), .A2(n783), .B(n782), .Z(
        RF_MEMCTRL_data_reg[25]) );
  AOI22D0BWP12T U1828 ( .A1(register_file_inst1_r6_27_), .A2(n839), .B1(
        register_file_inst1_r4_27_), .B2(n838), .ZN(n787) );
  AOI22D0BWP12T U1829 ( .A1(register_file_inst1_r7_27_), .A2(n841), .B1(
        register_file_inst1_r2_27_), .B2(n840), .ZN(n786) );
  AOI22D0BWP12T U1830 ( .A1(register_file_inst1_r0_27_), .A2(n843), .B1(
        register_file_inst1_r3_27_), .B2(n842), .ZN(n785) );
  AOI22D0BWP12T U1831 ( .A1(register_file_inst1_r1_27_), .A2(n845), .B1(
        register_file_inst1_r5_27_), .B2(n844), .ZN(n784) );
  ND4D1BWP12T U1832 ( .A1(n787), .A2(n786), .A3(n785), .A4(n784), .ZN(n792) );
  AOI22D0BWP12T U1833 ( .A1(register_file_inst1_r8_27_), .A2(n1948), .B1(
        STACK_RF_next_sp[27]), .B2(n1927), .ZN(n790) );
  AOI22D0BWP12T U1834 ( .A1(register_file_inst1_r10_27_), .A2(n852), .B1(
        register_file_inst1_r11_27_), .B2(n851), .ZN(n789) );
  AOI22D0BWP12T U1835 ( .A1(register_file_inst1_r9_27_), .A2(n850), .B1(
        register_file_inst1_r12_27_), .B2(n398), .ZN(n788) );
  ND4D1BWP12T U1836 ( .A1(n790), .A2(n1996), .A3(n789), .A4(n788), .ZN(n791)
         );
  AO21D1BWP12T U1837 ( .A1(n2306), .A2(n792), .B(n791), .Z(
        RF_MEMCTRL_data_reg[27]) );
  AOI22D0BWP12T U1838 ( .A1(register_file_inst1_r6_31_), .A2(n839), .B1(
        register_file_inst1_r4_31_), .B2(n838), .ZN(n796) );
  AOI22D0BWP12T U1839 ( .A1(register_file_inst1_r7_31_), .A2(n841), .B1(
        register_file_inst1_r2_31_), .B2(n840), .ZN(n795) );
  AOI22D0BWP12T U1840 ( .A1(register_file_inst1_r0_31_), .A2(n843), .B1(
        register_file_inst1_r3_31_), .B2(n842), .ZN(n794) );
  AOI22D0BWP12T U1841 ( .A1(register_file_inst1_r1_31_), .A2(n845), .B1(
        register_file_inst1_r5_31_), .B2(n844), .ZN(n793) );
  ND4D1BWP12T U1842 ( .A1(n796), .A2(n795), .A3(n794), .A4(n793), .ZN(n801) );
  AOI22D0BWP12T U1843 ( .A1(STACK_RF_next_sp[31]), .A2(n1927), .B1(
        register_file_inst1_r9_31_), .B2(n850), .ZN(n799) );
  AOI22D0BWP12T U1844 ( .A1(register_file_inst1_r8_31_), .A2(n1948), .B1(
        register_file_inst1_r11_31_), .B2(n851), .ZN(n798) );
  AOI22D0BWP12T U1845 ( .A1(register_file_inst1_r12_31_), .A2(n398), .B1(
        register_file_inst1_r10_31_), .B2(n852), .ZN(n797) );
  ND4D1BWP12T U1846 ( .A1(n799), .A2(n1993), .A3(n798), .A4(n797), .ZN(n800)
         );
  AO21D1BWP12T U1847 ( .A1(n2306), .A2(n801), .B(n800), .Z(
        RF_MEMCTRL_data_reg[31]) );
  AOI22D0BWP12T U1848 ( .A1(register_file_inst1_r6_29_), .A2(n839), .B1(
        register_file_inst1_r4_29_), .B2(n838), .ZN(n805) );
  AOI22D0BWP12T U1849 ( .A1(register_file_inst1_r7_29_), .A2(n841), .B1(
        register_file_inst1_r2_29_), .B2(n840), .ZN(n804) );
  AOI22D0BWP12T U1850 ( .A1(register_file_inst1_r0_29_), .A2(n843), .B1(
        register_file_inst1_r3_29_), .B2(n842), .ZN(n803) );
  AOI22D0BWP12T U1851 ( .A1(register_file_inst1_r1_29_), .A2(n845), .B1(
        register_file_inst1_r5_29_), .B2(n844), .ZN(n802) );
  ND4D1BWP12T U1852 ( .A1(n805), .A2(n804), .A3(n803), .A4(n802), .ZN(n810) );
  AOI22D0BWP12T U1853 ( .A1(STACK_RF_next_sp[29]), .A2(n1927), .B1(
        register_file_inst1_r10_29_), .B2(n852), .ZN(n808) );
  AOI22D0BWP12T U1854 ( .A1(register_file_inst1_r8_29_), .A2(n1948), .B1(
        register_file_inst1_r11_29_), .B2(n851), .ZN(n807) );
  AOI22D0BWP12T U1855 ( .A1(register_file_inst1_r9_29_), .A2(n850), .B1(
        register_file_inst1_r12_29_), .B2(n398), .ZN(n806) );
  ND4D1BWP12T U1856 ( .A1(n808), .A2(n1994), .A3(n807), .A4(n806), .ZN(n809)
         );
  AO21D1BWP12T U1857 ( .A1(n2306), .A2(n810), .B(n809), .Z(
        RF_MEMCTRL_data_reg[29]) );
  AOI22D0BWP12T U1858 ( .A1(register_file_inst1_r6_24_), .A2(n839), .B1(
        register_file_inst1_r4_24_), .B2(n838), .ZN(n814) );
  AOI22D0BWP12T U1859 ( .A1(register_file_inst1_r7_24_), .A2(n841), .B1(
        register_file_inst1_r2_24_), .B2(n840), .ZN(n813) );
  AOI22D0BWP12T U1860 ( .A1(register_file_inst1_r0_24_), .A2(n843), .B1(
        register_file_inst1_r3_24_), .B2(n842), .ZN(n812) );
  AOI22D0BWP12T U1861 ( .A1(register_file_inst1_r1_24_), .A2(n845), .B1(
        register_file_inst1_r5_24_), .B2(n844), .ZN(n811) );
  ND4D1BWP12T U1862 ( .A1(n814), .A2(n813), .A3(n812), .A4(n811), .ZN(n819) );
  AOI22D0BWP12T U1863 ( .A1(STACK_RF_next_sp[24]), .A2(n1927), .B1(
        register_file_inst1_r8_24_), .B2(n1948), .ZN(n817) );
  AOI22D0BWP12T U1864 ( .A1(register_file_inst1_r10_24_), .A2(n852), .B1(
        register_file_inst1_r11_24_), .B2(n851), .ZN(n816) );
  AOI22D0BWP12T U1865 ( .A1(register_file_inst1_r9_24_), .A2(n850), .B1(
        register_file_inst1_r12_24_), .B2(n398), .ZN(n815) );
  ND4D1BWP12T U1866 ( .A1(n1983), .A2(n817), .A3(n816), .A4(n815), .ZN(n818)
         );
  AO21D1BWP12T U1867 ( .A1(n2306), .A2(n819), .B(n818), .Z(
        RF_MEMCTRL_data_reg[24]) );
  AOI22D0BWP12T U1868 ( .A1(register_file_inst1_r6_30_), .A2(n839), .B1(
        register_file_inst1_r4_30_), .B2(n838), .ZN(n823) );
  AOI22D0BWP12T U1869 ( .A1(register_file_inst1_r7_30_), .A2(n841), .B1(
        register_file_inst1_r2_30_), .B2(n840), .ZN(n822) );
  AOI22D0BWP12T U1870 ( .A1(register_file_inst1_r0_30_), .A2(n843), .B1(
        register_file_inst1_r3_30_), .B2(n842), .ZN(n821) );
  AOI22D0BWP12T U1871 ( .A1(register_file_inst1_r1_30_), .A2(n845), .B1(
        register_file_inst1_r5_30_), .B2(n844), .ZN(n820) );
  ND4D1BWP12T U1872 ( .A1(n823), .A2(n822), .A3(n821), .A4(n820), .ZN(n828) );
  AOI22D0BWP12T U1873 ( .A1(STACK_RF_next_sp[30]), .A2(n1927), .B1(
        register_file_inst1_r8_30_), .B2(n1948), .ZN(n826) );
  AOI22D0BWP12T U1874 ( .A1(register_file_inst1_r10_30_), .A2(n852), .B1(
        register_file_inst1_r11_30_), .B2(n851), .ZN(n825) );
  AOI22D0BWP12T U1875 ( .A1(register_file_inst1_r9_30_), .A2(n850), .B1(
        register_file_inst1_r12_30_), .B2(n398), .ZN(n824) );
  ND4D1BWP12T U1876 ( .A1(n1982), .A2(n826), .A3(n825), .A4(n824), .ZN(n827)
         );
  AO21D1BWP12T U1877 ( .A1(n2306), .A2(n828), .B(n827), .Z(
        RF_MEMCTRL_data_reg[30]) );
  AOI22D0BWP12T U1878 ( .A1(register_file_inst1_r6_26_), .A2(n839), .B1(
        register_file_inst1_r4_26_), .B2(n838), .ZN(n832) );
  AOI22D0BWP12T U1879 ( .A1(register_file_inst1_r7_26_), .A2(n841), .B1(
        register_file_inst1_r2_26_), .B2(n840), .ZN(n831) );
  AOI22D0BWP12T U1880 ( .A1(register_file_inst1_r0_26_), .A2(n843), .B1(
        register_file_inst1_r3_26_), .B2(n842), .ZN(n830) );
  AOI22D0BWP12T U1881 ( .A1(register_file_inst1_r1_26_), .A2(n845), .B1(
        register_file_inst1_r5_26_), .B2(n844), .ZN(n829) );
  ND4D1BWP12T U1882 ( .A1(n832), .A2(n831), .A3(n830), .A4(n829), .ZN(n837) );
  AOI22D0BWP12T U1883 ( .A1(register_file_inst1_lr_26_), .A2(n1947), .B1(
        register_file_inst1_r9_26_), .B2(n850), .ZN(n835) );
  AOI22D0BWP12T U1884 ( .A1(STACK_RF_next_sp[26]), .A2(n1927), .B1(
        register_file_inst1_r11_26_), .B2(n851), .ZN(n834) );
  AOI22D0BWP12T U1885 ( .A1(register_file_inst1_r12_26_), .A2(n398), .B1(
        register_file_inst1_r10_26_), .B2(n852), .ZN(n833) );
  ND4D1BWP12T U1886 ( .A1(n835), .A2(n1997), .A3(n834), .A4(n833), .ZN(n836)
         );
  AO21D1BWP12T U1887 ( .A1(n2306), .A2(n837), .B(n836), .Z(
        RF_MEMCTRL_data_reg[26]) );
  AOI22D0BWP12T U1888 ( .A1(register_file_inst1_r6_28_), .A2(n839), .B1(
        register_file_inst1_r4_28_), .B2(n838), .ZN(n849) );
  AOI22D0BWP12T U1889 ( .A1(register_file_inst1_r7_28_), .A2(n841), .B1(
        register_file_inst1_r2_28_), .B2(n840), .ZN(n848) );
  AOI22D0BWP12T U1890 ( .A1(register_file_inst1_r0_28_), .A2(n843), .B1(
        register_file_inst1_r3_28_), .B2(n842), .ZN(n847) );
  AOI22D0BWP12T U1891 ( .A1(register_file_inst1_r1_28_), .A2(n845), .B1(
        register_file_inst1_r5_28_), .B2(n844), .ZN(n846) );
  ND4D1BWP12T U1892 ( .A1(n849), .A2(n848), .A3(n847), .A4(n846), .ZN(n857) );
  AOI22D0BWP12T U1893 ( .A1(register_file_inst1_lr_28_), .A2(n1947), .B1(
        register_file_inst1_r9_28_), .B2(n850), .ZN(n855) );
  AOI22D0BWP12T U1894 ( .A1(STACK_RF_next_sp[28]), .A2(n1927), .B1(
        register_file_inst1_r11_28_), .B2(n851), .ZN(n854) );
  AOI22D0BWP12T U1895 ( .A1(register_file_inst1_r12_28_), .A2(n398), .B1(
        register_file_inst1_r10_28_), .B2(n852), .ZN(n853) );
  ND4D1BWP12T U1896 ( .A1(n855), .A2(n1995), .A3(n854), .A4(n853), .ZN(n856)
         );
  AO21D1BWP12T U1897 ( .A1(n2306), .A2(n857), .B(n856), .Z(
        RF_MEMCTRL_data_reg[28]) );
  INVD1BWP12T U1898 ( .I(n1956), .ZN(n861) );
  CKND2D1BWP12T U1899 ( .A1(n858), .A2(memory_interface_inst1_fsm_state_0_), 
        .ZN(n933) );
  NR2D0BWP12T U1900 ( .A1(n933), .A2(memory_interface_inst1_fsm_state_3_), 
        .ZN(n859) );
  AOI211D1BWP12T U1901 ( .A1(n862), .A2(n861), .B(n860), .C(n859), .ZN(n1954)
         );
  ND2D1BWP12T U1902 ( .A1(n862), .A2(n2333), .ZN(n1955) );
  OA21D1BWP12T U1903 ( .A1(n1957), .A2(n1956), .B(n1955), .Z(n1958) );
  NR2D1BWP12T U1904 ( .A1(n2120), .A2(n1102), .ZN(n2013) );
  NR2D1BWP12T U1905 ( .A1(n2126), .A2(n1102), .ZN(n2007) );
  NR2D1BWP12T U1906 ( .A1(n2123), .A2(n1102), .ZN(n2010) );
  NR2D1BWP12T U1907 ( .A1(n2117), .A2(n1102), .ZN(n2016) );
  NR2D1BWP12T U1908 ( .A1(n2115), .A2(n1102), .ZN(n2019) );
  INVD1BWP12T U1909 ( .I(n2280), .ZN(n2284) );
  OAI211D1BWP12T U1910 ( .A1(n2284), .A2(register_file_inst1_pc_write_in_1_), 
        .B(n2283), .C(n2282), .ZN(register_file_inst1_n2170) );
  ND2D1BWP12T U1911 ( .A1(n2324), .A2(n2325), .ZN(n867) );
  NR2D1BWP12T U1912 ( .A1(n2318), .A2(n867), .ZN(n943) );
  NR2D1BWP12T U1913 ( .A1(n2322), .A2(n2319), .ZN(n942) );
  AOI22D0BWP12T U1914 ( .A1(register_file_inst1_r0_2_), .A2(n943), .B1(
        register_file_inst1_r9_2_), .B2(n942), .ZN(n866) );
  NR2D1BWP12T U1915 ( .A1(n2317), .A2(n2320), .ZN(n945) );
  NR2D1BWP12T U1916 ( .A1(n2323), .A2(n2317), .ZN(n944) );
  AOI22D0BWP12T U1917 ( .A1(register_file_inst1_r6_2_), .A2(n945), .B1(
        register_file_inst1_lr_2_), .B2(n944), .ZN(n865) );
  NR2D1BWP12T U1918 ( .A1(n2323), .A2(n2318), .ZN(n947) );
  NR2D1BWP12T U1919 ( .A1(n2323), .A2(n2322), .ZN(n946) );
  AOI22D0BWP12T U1920 ( .A1(register_file_inst1_r12_2_), .A2(n947), .B1(
        STACK_RF_next_sp[2]), .B2(n946), .ZN(n864) );
  NR2D1BWP12T U1921 ( .A1(n2322), .A2(n867), .ZN(n949) );
  NR2D1BWP12T U1922 ( .A1(n867), .A2(n2321), .ZN(n948) );
  AOI22D0BWP12T U1923 ( .A1(register_file_inst1_r1_2_), .A2(n949), .B1(
        register_file_inst1_r3_2_), .B2(n948), .ZN(n863) );
  ND4D1BWP12T U1924 ( .A1(n866), .A2(n865), .A3(n864), .A4(n863), .ZN(n2047)
         );
  NR2D1BWP12T U1925 ( .A1(n2318), .A2(n2319), .ZN(n955) );
  NR2D1BWP12T U1926 ( .A1(n867), .A2(n2317), .ZN(n954) );
  AOI22D0BWP12T U1927 ( .A1(register_file_inst1_r8_2_), .A2(n955), .B1(
        register_file_inst1_r2_2_), .B2(n954), .ZN(n870) );
  NR2D1BWP12T U1928 ( .A1(n2321), .A2(n2320), .ZN(n957) );
  NR2D1BWP12T U1929 ( .A1(n2318), .A2(n2320), .ZN(n956) );
  AOI22D0BWP12T U1930 ( .A1(register_file_inst1_r7_2_), .A2(n957), .B1(
        register_file_inst1_r4_2_), .B2(n956), .ZN(n869) );
  NR2D1BWP12T U1931 ( .A1(n2319), .A2(n2317), .ZN(n958) );
  NR2D1BWP12T U1932 ( .A1(n2321), .A2(n2319), .ZN(n959) );
  AOI22D0BWP12T U1933 ( .A1(register_file_inst1_r10_2_), .A2(n958), .B1(
        register_file_inst1_r11_2_), .B2(n959), .ZN(n868) );
  ND4D1BWP12T U1934 ( .A1(n870), .A2(n869), .A3(n868), .A4(n2046), .ZN(n2048)
         );
  AOI22D0BWP12T U1935 ( .A1(register_file_inst1_r0_3_), .A2(n943), .B1(
        register_file_inst1_r9_3_), .B2(n942), .ZN(n874) );
  AOI22D0BWP12T U1936 ( .A1(register_file_inst1_r6_3_), .A2(n945), .B1(
        register_file_inst1_lr_3_), .B2(n944), .ZN(n873) );
  AOI22D0BWP12T U1937 ( .A1(register_file_inst1_r12_3_), .A2(n947), .B1(
        STACK_RF_next_sp[3]), .B2(n946), .ZN(n872) );
  AOI22D0BWP12T U1938 ( .A1(register_file_inst1_r1_3_), .A2(n949), .B1(
        register_file_inst1_r3_3_), .B2(n948), .ZN(n871) );
  ND4D1BWP12T U1939 ( .A1(n874), .A2(n873), .A3(n872), .A4(n871), .ZN(n2050)
         );
  AOI22D0BWP12T U1940 ( .A1(register_file_inst1_r8_3_), .A2(n955), .B1(
        register_file_inst1_r2_3_), .B2(n954), .ZN(n877) );
  AOI22D0BWP12T U1941 ( .A1(register_file_inst1_r7_3_), .A2(n957), .B1(
        register_file_inst1_r4_3_), .B2(n956), .ZN(n876) );
  AOI22D0BWP12T U1942 ( .A1(register_file_inst1_r10_3_), .A2(n958), .B1(
        register_file_inst1_r11_3_), .B2(n959), .ZN(n875) );
  ND4D1BWP12T U1943 ( .A1(n877), .A2(n876), .A3(n875), .A4(n2049), .ZN(n2051)
         );
  AOI22D0BWP12T U1944 ( .A1(register_file_inst1_r0_4_), .A2(n943), .B1(
        register_file_inst1_r9_4_), .B2(n942), .ZN(n881) );
  AOI22D0BWP12T U1945 ( .A1(register_file_inst1_r6_4_), .A2(n945), .B1(
        register_file_inst1_lr_4_), .B2(n944), .ZN(n880) );
  AOI22D0BWP12T U1946 ( .A1(register_file_inst1_r12_4_), .A2(n947), .B1(
        STACK_RF_next_sp[4]), .B2(n946), .ZN(n879) );
  AOI22D0BWP12T U1947 ( .A1(register_file_inst1_r1_4_), .A2(n949), .B1(
        register_file_inst1_r3_4_), .B2(n948), .ZN(n878) );
  ND4D1BWP12T U1948 ( .A1(n881), .A2(n880), .A3(n879), .A4(n878), .ZN(n2053)
         );
  AOI22D0BWP12T U1949 ( .A1(register_file_inst1_r8_4_), .A2(n955), .B1(
        register_file_inst1_r2_4_), .B2(n954), .ZN(n884) );
  AOI22D0BWP12T U1950 ( .A1(register_file_inst1_r7_4_), .A2(n957), .B1(
        register_file_inst1_r4_4_), .B2(n956), .ZN(n883) );
  AOI22D0BWP12T U1951 ( .A1(register_file_inst1_r10_4_), .A2(n958), .B1(
        register_file_inst1_r11_4_), .B2(n959), .ZN(n882) );
  ND4D1BWP12T U1952 ( .A1(n884), .A2(n883), .A3(n882), .A4(n2052), .ZN(n2054)
         );
  AOI22D0BWP12T U1953 ( .A1(register_file_inst1_r0_5_), .A2(n943), .B1(
        register_file_inst1_r9_5_), .B2(n942), .ZN(n890) );
  AOI22D0BWP12T U1954 ( .A1(register_file_inst1_r6_5_), .A2(n945), .B1(
        register_file_inst1_lr_5_), .B2(n944), .ZN(n889) );
  AOI22D0BWP12T U1955 ( .A1(register_file_inst1_r12_5_), .A2(n947), .B1(
        STACK_RF_next_sp[5]), .B2(n946), .ZN(n888) );
  AOI22D0BWP12T U1956 ( .A1(register_file_inst1_r1_5_), .A2(n949), .B1(
        register_file_inst1_r3_5_), .B2(n948), .ZN(n887) );
  ND4D1BWP12T U1957 ( .A1(n890), .A2(n889), .A3(n888), .A4(n887), .ZN(n2056)
         );
  AOI22D0BWP12T U1958 ( .A1(register_file_inst1_r8_5_), .A2(n955), .B1(
        register_file_inst1_r2_5_), .B2(n954), .ZN(n893) );
  AOI22D0BWP12T U1959 ( .A1(register_file_inst1_r7_5_), .A2(n957), .B1(
        register_file_inst1_r4_5_), .B2(n956), .ZN(n892) );
  AOI22D0BWP12T U1960 ( .A1(register_file_inst1_r10_5_), .A2(n958), .B1(
        register_file_inst1_r11_5_), .B2(n959), .ZN(n891) );
  ND4D1BWP12T U1961 ( .A1(n893), .A2(n892), .A3(n891), .A4(n2055), .ZN(n2057)
         );
  INVD1BWP12T U1962 ( .I(register_file_inst1_pc_write_in_3_), .ZN(n895) );
  XNR2D1BWP12T U1963 ( .A1(n895), .A2(n894), .ZN(
        register_file_inst1_pc_write_in_plus_two[3]) );
  AOI22D1BWP12T U1964 ( .A1(register_file_inst1_r0_6_), .A2(n943), .B1(
        register_file_inst1_r9_6_), .B2(n942), .ZN(n899) );
  AOI22D1BWP12T U1965 ( .A1(register_file_inst1_r6_6_), .A2(n945), .B1(
        register_file_inst1_lr_6_), .B2(n944), .ZN(n898) );
  AOI22D1BWP12T U1966 ( .A1(register_file_inst1_r12_6_), .A2(n947), .B1(
        STACK_RF_next_sp[6]), .B2(n946), .ZN(n897) );
  AOI22D1BWP12T U1967 ( .A1(register_file_inst1_r1_6_), .A2(n949), .B1(
        register_file_inst1_r3_6_), .B2(n948), .ZN(n896) );
  ND4D1BWP12T U1968 ( .A1(n899), .A2(n898), .A3(n897), .A4(n896), .ZN(n2059)
         );
  AOI22D1BWP12T U1969 ( .A1(register_file_inst1_r8_6_), .A2(n955), .B1(
        register_file_inst1_r2_6_), .B2(n954), .ZN(n902) );
  AOI22D0BWP12T U1970 ( .A1(register_file_inst1_r7_6_), .A2(n957), .B1(
        register_file_inst1_r4_6_), .B2(n956), .ZN(n901) );
  AOI22D1BWP12T U1971 ( .A1(register_file_inst1_r10_6_), .A2(n958), .B1(
        register_file_inst1_r11_6_), .B2(n959), .ZN(n900) );
  ND4D1BWP12T U1972 ( .A1(n902), .A2(n901), .A3(n900), .A4(n2058), .ZN(n2060)
         );
  AOI22D0BWP12T U1973 ( .A1(register_file_inst1_r0_7_), .A2(n943), .B1(
        register_file_inst1_r9_7_), .B2(n942), .ZN(n906) );
  AOI22D0BWP12T U1974 ( .A1(register_file_inst1_r6_7_), .A2(n945), .B1(
        register_file_inst1_lr_7_), .B2(n944), .ZN(n905) );
  AOI22D0BWP12T U1975 ( .A1(register_file_inst1_r12_7_), .A2(n947), .B1(
        STACK_RF_next_sp[7]), .B2(n946), .ZN(n904) );
  AOI22D0BWP12T U1976 ( .A1(register_file_inst1_r1_7_), .A2(n949), .B1(
        register_file_inst1_r3_7_), .B2(n948), .ZN(n903) );
  ND4D1BWP12T U1977 ( .A1(n906), .A2(n905), .A3(n904), .A4(n903), .ZN(n2062)
         );
  AOI22D0BWP12T U1978 ( .A1(register_file_inst1_r8_7_), .A2(n955), .B1(
        register_file_inst1_r2_7_), .B2(n954), .ZN(n909) );
  AOI22D0BWP12T U1979 ( .A1(register_file_inst1_r7_7_), .A2(n957), .B1(
        register_file_inst1_r4_7_), .B2(n956), .ZN(n908) );
  AOI22D0BWP12T U1980 ( .A1(register_file_inst1_r10_7_), .A2(n958), .B1(
        register_file_inst1_r11_7_), .B2(n959), .ZN(n907) );
  ND4D1BWP12T U1981 ( .A1(n909), .A2(n908), .A3(n907), .A4(n2061), .ZN(n2063)
         );
  AOI22D0BWP12T U1982 ( .A1(register_file_inst1_r0_10_), .A2(n943), .B1(
        register_file_inst1_r9_10_), .B2(n942), .ZN(n913) );
  AOI22D0BWP12T U1983 ( .A1(register_file_inst1_r6_10_), .A2(n945), .B1(
        register_file_inst1_lr_10_), .B2(n944), .ZN(n912) );
  AOI22D0BWP12T U1984 ( .A1(register_file_inst1_r12_10_), .A2(n947), .B1(
        STACK_RF_next_sp[10]), .B2(n946), .ZN(n911) );
  AOI22D0BWP12T U1985 ( .A1(register_file_inst1_r1_10_), .A2(n949), .B1(
        register_file_inst1_r3_10_), .B2(n948), .ZN(n910) );
  ND4D1BWP12T U1986 ( .A1(n913), .A2(n912), .A3(n911), .A4(n910), .ZN(n2071)
         );
  AOI22D0BWP12T U1987 ( .A1(register_file_inst1_r8_10_), .A2(n955), .B1(
        register_file_inst1_r2_10_), .B2(n954), .ZN(n916) );
  AOI22D0BWP12T U1988 ( .A1(register_file_inst1_r7_10_), .A2(n957), .B1(
        register_file_inst1_r4_10_), .B2(n956), .ZN(n915) );
  AOI22D0BWP12T U1989 ( .A1(register_file_inst1_r10_10_), .A2(n958), .B1(
        register_file_inst1_r11_10_), .B2(n959), .ZN(n914) );
  ND4D1BWP12T U1990 ( .A1(n916), .A2(n915), .A3(n914), .A4(n2070), .ZN(n2072)
         );
  INVD1BWP12T U1991 ( .I(register_file_inst1_pc_write_in_5_), .ZN(n918) );
  XNR2D1BWP12T U1992 ( .A1(n918), .A2(n917), .ZN(
        register_file_inst1_pc_write_in_plus_two[5]) );
  AOI22D0BWP12T U1993 ( .A1(register_file_inst1_r0_8_), .A2(n943), .B1(
        register_file_inst1_r9_8_), .B2(n942), .ZN(n922) );
  AOI22D0BWP12T U1994 ( .A1(register_file_inst1_r6_8_), .A2(n945), .B1(
        register_file_inst1_lr_8_), .B2(n944), .ZN(n921) );
  AOI22D0BWP12T U1995 ( .A1(register_file_inst1_r12_8_), .A2(n947), .B1(
        STACK_RF_next_sp[8]), .B2(n946), .ZN(n920) );
  AOI22D0BWP12T U1996 ( .A1(register_file_inst1_r1_8_), .A2(n949), .B1(
        register_file_inst1_r3_8_), .B2(n948), .ZN(n919) );
  ND4D1BWP12T U1997 ( .A1(n922), .A2(n921), .A3(n920), .A4(n919), .ZN(n2065)
         );
  AOI22D0BWP12T U1998 ( .A1(register_file_inst1_r8_8_), .A2(n955), .B1(
        register_file_inst1_r2_8_), .B2(n954), .ZN(n925) );
  AOI22D0BWP12T U1999 ( .A1(register_file_inst1_r7_8_), .A2(n957), .B1(
        register_file_inst1_r4_8_), .B2(n956), .ZN(n924) );
  AOI22D0BWP12T U2000 ( .A1(register_file_inst1_r10_8_), .A2(n958), .B1(
        register_file_inst1_r11_8_), .B2(n959), .ZN(n923) );
  ND4D1BWP12T U2001 ( .A1(n925), .A2(n924), .A3(n923), .A4(n2064), .ZN(n2066)
         );
  AOI22D0BWP12T U2002 ( .A1(register_file_inst1_r0_9_), .A2(n943), .B1(
        register_file_inst1_r9_9_), .B2(n942), .ZN(n929) );
  AOI22D0BWP12T U2003 ( .A1(register_file_inst1_r6_9_), .A2(n945), .B1(
        register_file_inst1_lr_9_), .B2(n944), .ZN(n928) );
  AOI22D0BWP12T U2004 ( .A1(register_file_inst1_r12_9_), .A2(n947), .B1(
        STACK_RF_next_sp[9]), .B2(n946), .ZN(n927) );
  AOI22D0BWP12T U2005 ( .A1(register_file_inst1_r1_9_), .A2(n949), .B1(
        register_file_inst1_r3_9_), .B2(n948), .ZN(n926) );
  ND4D1BWP12T U2006 ( .A1(n929), .A2(n928), .A3(n927), .A4(n926), .ZN(n2068)
         );
  AOI22D0BWP12T U2007 ( .A1(register_file_inst1_r8_9_), .A2(n955), .B1(
        register_file_inst1_r2_9_), .B2(n954), .ZN(n932) );
  AOI22D0BWP12T U2008 ( .A1(register_file_inst1_r7_9_), .A2(n957), .B1(
        register_file_inst1_r4_9_), .B2(n956), .ZN(n931) );
  AOI22D0BWP12T U2009 ( .A1(register_file_inst1_r10_9_), .A2(n958), .B1(
        register_file_inst1_r11_9_), .B2(n959), .ZN(n930) );
  ND4D1BWP12T U2010 ( .A1(n932), .A2(n931), .A3(n930), .A4(n2067), .ZN(n2069)
         );
  ND2D1BWP12T U2011 ( .A1(n934), .A2(n933), .ZN(n1961) );
  AOI22D0BWP12T U2012 ( .A1(register_file_inst1_r0_12_), .A2(n943), .B1(
        register_file_inst1_r9_12_), .B2(n942), .ZN(n938) );
  AOI22D0BWP12T U2013 ( .A1(register_file_inst1_r6_12_), .A2(n945), .B1(
        register_file_inst1_lr_12_), .B2(n944), .ZN(n937) );
  AOI22D0BWP12T U2014 ( .A1(register_file_inst1_r12_12_), .A2(n947), .B1(
        STACK_RF_next_sp[12]), .B2(n946), .ZN(n936) );
  AOI22D0BWP12T U2015 ( .A1(register_file_inst1_r1_12_), .A2(n949), .B1(
        register_file_inst1_r3_12_), .B2(n948), .ZN(n935) );
  ND4D1BWP12T U2016 ( .A1(n938), .A2(n937), .A3(n936), .A4(n935), .ZN(n2077)
         );
  AOI22D0BWP12T U2017 ( .A1(register_file_inst1_r8_12_), .A2(n955), .B1(
        register_file_inst1_r2_12_), .B2(n954), .ZN(n941) );
  AOI22D0BWP12T U2018 ( .A1(register_file_inst1_r7_12_), .A2(n957), .B1(
        register_file_inst1_r4_12_), .B2(n956), .ZN(n940) );
  AOI22D0BWP12T U2019 ( .A1(register_file_inst1_r10_12_), .A2(n958), .B1(
        register_file_inst1_r11_12_), .B2(n959), .ZN(n939) );
  ND4D1BWP12T U2020 ( .A1(n941), .A2(n940), .A3(n939), .A4(n2076), .ZN(n2078)
         );
  AOI22D0BWP12T U2021 ( .A1(register_file_inst1_r0_11_), .A2(n943), .B1(
        register_file_inst1_r9_11_), .B2(n942), .ZN(n953) );
  AOI22D0BWP12T U2022 ( .A1(register_file_inst1_r6_11_), .A2(n945), .B1(
        register_file_inst1_lr_11_), .B2(n944), .ZN(n952) );
  AOI22D0BWP12T U2023 ( .A1(register_file_inst1_r12_11_), .A2(n947), .B1(
        STACK_RF_next_sp[11]), .B2(n946), .ZN(n951) );
  AOI22D0BWP12T U2024 ( .A1(register_file_inst1_r1_11_), .A2(n949), .B1(
        register_file_inst1_r3_11_), .B2(n948), .ZN(n950) );
  ND4D1BWP12T U2025 ( .A1(n953), .A2(n952), .A3(n951), .A4(n950), .ZN(n2074)
         );
  AOI22D0BWP12T U2026 ( .A1(register_file_inst1_r8_11_), .A2(n955), .B1(
        register_file_inst1_r2_11_), .B2(n954), .ZN(n962) );
  AOI22D0BWP12T U2027 ( .A1(register_file_inst1_r7_11_), .A2(n957), .B1(
        register_file_inst1_r4_11_), .B2(n956), .ZN(n961) );
  AOI22D0BWP12T U2028 ( .A1(register_file_inst1_r11_11_), .A2(n959), .B1(
        register_file_inst1_r10_11_), .B2(n958), .ZN(n960) );
  ND4D1BWP12T U2029 ( .A1(n962), .A2(n961), .A3(n960), .A4(n2073), .ZN(n2075)
         );
  OAI222D1BWP12T U2030 ( .A1(n1183), .A2(n1037), .B1(n1102), .B2(n967), .C1(
        n1104), .C2(n966), .ZN(register_file_inst1_spin[16]) );
  CKND0BWP12T U2031 ( .I(register_file_inst1_r2_16_), .ZN(n963) );
  OAI222D1BWP12T U2032 ( .A1(n963), .A2(n1060), .B1(n1062), .B2(n967), .C1(
        n1063), .C2(n966), .ZN(register_file_inst1_n2569) );
  INVD1BWP12T U2033 ( .I(register_file_inst1_r10_16_), .ZN(n1194) );
  OAI222D1BWP12T U2034 ( .A1(n1194), .A2(n1068), .B1(n1069), .B2(n967), .C1(
        n1070), .C2(n966), .ZN(register_file_inst1_n2313) );
  INVD1BWP12T U2035 ( .I(register_file_inst1_r3_16_), .ZN(n1186) );
  OAI222D1BWP12T U2036 ( .A1(n1186), .A2(n1064), .B1(n1066), .B2(n967), .C1(
        n1067), .C2(n966), .ZN(register_file_inst1_n2537) );
  OAI222D1BWP12T U2037 ( .A1(n1205), .A2(n1021), .B1(n964), .B2(n967), .C1(
        n1019), .C2(n966), .ZN(register_file_inst1_n2281) );
  INVD1BWP12T U2038 ( .I(register_file_inst1_r12_16_), .ZN(n1184) );
  OAI222D1BWP12T U2039 ( .A1(n1184), .A2(n1071), .B1(n1073), .B2(n967), .C1(
        n1074), .C2(n966), .ZN(register_file_inst1_n2249) );
  CKND0BWP12T U2040 ( .I(register_file_inst1_r8_16_), .ZN(n965) );
  OAI222D1BWP12T U2041 ( .A1(n965), .A2(n1075), .B1(n1077), .B2(n967), .C1(
        n1078), .C2(n966), .ZN(register_file_inst1_n2377) );
  INVD1BWP12T U2042 ( .I(register_file_inst1_r9_16_), .ZN(n1207) );
  OAI222D1BWP12T U2043 ( .A1(n1207), .A2(n1079), .B1(n1080), .B2(n967), .C1(
        n1081), .C2(n966), .ZN(register_file_inst1_n2345) );
  INVD1BWP12T U2044 ( .I(register_file_inst1_r0_16_), .ZN(n1185) );
  OAI222D1BWP12T U2045 ( .A1(n1185), .A2(n1086), .B1(n1088), .B2(n967), .C1(
        n1089), .C2(n966), .ZN(register_file_inst1_n2633) );
  INVD1BWP12T U2046 ( .I(register_file_inst1_r4_16_), .ZN(n1195) );
  OAI222D1BWP12T U2047 ( .A1(n1195), .A2(n1090), .B1(n1091), .B2(n967), .C1(
        n1092), .C2(n966), .ZN(register_file_inst1_n2505) );
  INVD1BWP12T U2048 ( .I(register_file_inst1_tmp1_16_), .ZN(n1198) );
  OAI222D1BWP12T U2049 ( .A1(n1198), .A2(n1027), .B1(n1026), .B2(n967), .C1(
        n2168), .C2(n966), .ZN(register_file_inst1_n2153) );
  INVD1BWP12T U2050 ( .I(STACK_RF_next_sp[19]), .ZN(n1526) );
  OAI222D1BWP12T U2051 ( .A1(n1526), .A2(n1037), .B1(n1102), .B2(n971), .C1(
        n1104), .C2(n970), .ZN(register_file_inst1_spin[19]) );
  OAI222D1BWP12T U2052 ( .A1(n1541), .A2(n1021), .B1(n1020), .B2(n971), .C1(
        n1019), .C2(n970), .ZN(register_file_inst1_n2284) );
  CKND0BWP12T U2053 ( .I(register_file_inst1_r8_19_), .ZN(n968) );
  OAI222D1BWP12T U2054 ( .A1(n968), .A2(n1075), .B1(n1077), .B2(n971), .C1(
        n1078), .C2(n970), .ZN(register_file_inst1_n2380) );
  INVD1BWP12T U2055 ( .I(register_file_inst1_r12_19_), .ZN(n1527) );
  OAI222D1BWP12T U2056 ( .A1(n1527), .A2(n1071), .B1(n1073), .B2(n971), .C1(
        n1074), .C2(n970), .ZN(register_file_inst1_n2252) );
  OAI222D1BWP12T U2057 ( .A1(n969), .A2(n1079), .B1(n1080), .B2(n971), .C1(
        n1081), .C2(n970), .ZN(register_file_inst1_n2348) );
  INVD1BWP12T U2058 ( .I(register_file_inst1_tmp1_19_), .ZN(n1544) );
  OAI222D1BWP12T U2059 ( .A1(n1544), .A2(n1027), .B1(n1026), .B2(n971), .C1(
        n2168), .C2(n970), .ZN(register_file_inst1_n2156) );
  NR2D1BWP12T U2060 ( .A1(n17), .A2(n972), .ZN(n973) );
  XNR2D1BWP12T U2061 ( .A1(n1931), .A2(n973), .ZN(
        register_file_inst1_pc_write_in_plus_two[9]) );
  XNR2D1BWP12T U2062 ( .A1(n17), .A2(n974), .ZN(
        register_file_inst1_pc_write_in_plus_two[8]) );
  CKND0BWP12T U2063 ( .I(STACK_RF_next_sp[22]), .ZN(n976) );
  OAI222D1BWP12T U2064 ( .A1(n976), .A2(n975), .B1(n1102), .B2(n989), .C1(
        n1104), .C2(n988), .ZN(register_file_inst1_spin[22]) );
  OAI222D1BWP12T U2065 ( .A1(n977), .A2(n1096), .B1(n1097), .B2(n989), .C1(
        n1098), .C2(n988), .ZN(register_file_inst1_n2479) );
  CKND0BWP12T U2066 ( .I(register_file_inst1_r0_22_), .ZN(n978) );
  OAI222D1BWP12T U2067 ( .A1(n978), .A2(n1086), .B1(n1088), .B2(n989), .C1(
        n1089), .C2(n988), .ZN(register_file_inst1_n2639) );
  OAI222D1BWP12T U2068 ( .A1(n979), .A2(n1093), .B1(n1094), .B2(n989), .C1(
        n1095), .C2(n988), .ZN(register_file_inst1_n2607) );
  CKND0BWP12T U2069 ( .I(register_file_inst1_tmp1_22_), .ZN(n980) );
  OAI222D1BWP12T U2070 ( .A1(n980), .A2(n1027), .B1(n1026), .B2(n989), .C1(
        n2168), .C2(n988), .ZN(register_file_inst1_n2159) );
  OAI222D1BWP12T U2071 ( .A1(n981), .A2(n1090), .B1(n1091), .B2(n989), .C1(
        n1092), .C2(n988), .ZN(register_file_inst1_n2511) );
  CKND0BWP12T U2072 ( .I(register_file_inst1_lr_22_), .ZN(n982) );
  OAI222D1BWP12T U2073 ( .A1(n982), .A2(n1082), .B1(n1084), .B2(n989), .C1(
        n1085), .C2(n988), .ZN(register_file_inst1_n2223) );
  CKND0BWP12T U2074 ( .I(register_file_inst1_r2_22_), .ZN(n983) );
  OAI222D1BWP12T U2075 ( .A1(n983), .A2(n1060), .B1(n1062), .B2(n989), .C1(
        n1063), .C2(n988), .ZN(register_file_inst1_n2575) );
  OAI222D1BWP12T U2076 ( .A1(n984), .A2(n1068), .B1(n1069), .B2(n989), .C1(
        n1070), .C2(n988), .ZN(register_file_inst1_n2319) );
  CKND0BWP12T U2077 ( .I(register_file_inst1_r3_22_), .ZN(n985) );
  OAI222D1BWP12T U2078 ( .A1(n985), .A2(n1064), .B1(n1066), .B2(n989), .C1(
        n1067), .C2(n988), .ZN(register_file_inst1_n2543) );
  CKND0BWP12T U2079 ( .I(register_file_inst1_r12_22_), .ZN(n986) );
  OAI222D1BWP12T U2080 ( .A1(n986), .A2(n1071), .B1(n1073), .B2(n989), .C1(
        n1074), .C2(n988), .ZN(register_file_inst1_n2255) );
  CKND0BWP12T U2081 ( .I(register_file_inst1_r8_22_), .ZN(n987) );
  OAI222D1BWP12T U2082 ( .A1(n987), .A2(n1075), .B1(n1077), .B2(n989), .C1(
        n1078), .C2(n988), .ZN(register_file_inst1_n2383) );
  OAI222D1BWP12T U2083 ( .A1(n990), .A2(n1079), .B1(n1080), .B2(n989), .C1(
        n1081), .C2(n988), .ZN(register_file_inst1_n2351) );
  INVD1BWP12T U2084 ( .I(register_file_inst1_pc_write_in_14_), .ZN(n992) );
  XNR2D1BWP12T U2085 ( .A1(n992), .A2(n991), .ZN(
        register_file_inst1_pc_write_in_plus_two[14]) );
  INVD1BWP12T U2086 ( .I(register_file_inst1_pc_write_in_12_), .ZN(n994) );
  XNR2D1BWP12T U2087 ( .A1(n994), .A2(n993), .ZN(
        register_file_inst1_pc_write_in_plus_two[12]) );
  INVD1BWP12T U2088 ( .I(n995), .ZN(n997) );
  XNR2D1BWP12T U2089 ( .A1(n997), .A2(n996), .ZN(
        register_file_inst1_pc_write_in_plus_two[18]) );
  INVD1BWP12T U2090 ( .I(n998), .ZN(n1000) );
  XNR2D1BWP12T U2091 ( .A1(n1000), .A2(n999), .ZN(
        register_file_inst1_pc_write_in_plus_two[20]) );
  XOR2D1BWP12T U2092 ( .A1(n1002), .A2(n1001), .Z(
        register_file_inst1_pc_write_in_plus_two[21]) );
  CKND0BWP12T U2093 ( .I(register_file_inst1_r6_28_), .ZN(n1003) );
  OAI222D1BWP12T U2094 ( .A1(n1003), .A2(n1045), .B1(n1044), .B2(n1012), .C1(
        n1043), .C2(n1011), .ZN(register_file_inst1_n2453) );
  CKND0BWP12T U2095 ( .I(register_file_inst1_lr_28_), .ZN(n1004) );
  OAI222D1BWP12T U2096 ( .A1(n1004), .A2(n1082), .B1(n1084), .B2(n1012), .C1(
        n1085), .C2(n1011), .ZN(register_file_inst1_n2229) );
  INVD1BWP12T U2097 ( .I(register_file_inst1_r4_28_), .ZN(n1578) );
  OAI222D1BWP12T U2098 ( .A1(n1578), .A2(n1090), .B1(n1091), .B2(n1012), .C1(
        n1092), .C2(n1011), .ZN(register_file_inst1_n2517) );
  OAI222D1BWP12T U2099 ( .A1(n1005), .A2(n1093), .B1(n1094), .B2(n1012), .C1(
        n1095), .C2(n1011), .ZN(register_file_inst1_n2613) );
  INVD1BWP12T U2100 ( .I(register_file_inst1_r5_28_), .ZN(n1580) );
  OAI222D1BWP12T U2101 ( .A1(n1580), .A2(n1096), .B1(n1097), .B2(n1012), .C1(
        n1098), .C2(n1011), .ZN(register_file_inst1_n2485) );
  OAI222D1BWP12T U2102 ( .A1(n1006), .A2(n1051), .B1(n1050), .B2(n1012), .C1(
        n1049), .C2(n1011), .ZN(register_file_inst1_n2421) );
  CKND0BWP12T U2103 ( .I(register_file_inst1_r0_28_), .ZN(n1007) );
  OAI222D1BWP12T U2104 ( .A1(n1007), .A2(n1086), .B1(n1088), .B2(n1012), .C1(
        n1089), .C2(n1011), .ZN(register_file_inst1_n2645) );
  CKND0BWP12T U2105 ( .I(STACK_RF_next_sp[28]), .ZN(n1008) );
  OAI222D1BWP12T U2106 ( .A1(n1008), .A2(n1037), .B1(n1102), .B2(n1012), .C1(
        n1104), .C2(n1011), .ZN(register_file_inst1_spin[28]) );
  CKND0BWP12T U2107 ( .I(register_file_inst1_r8_28_), .ZN(n1009) );
  OAI222D1BWP12T U2108 ( .A1(n1009), .A2(n1075), .B1(n1077), .B2(n1012), .C1(
        n1078), .C2(n1011), .ZN(register_file_inst1_n2389) );
  CKND0BWP12T U2109 ( .I(register_file_inst1_r12_28_), .ZN(n1010) );
  OAI222D1BWP12T U2110 ( .A1(n1010), .A2(n1071), .B1(n1073), .B2(n1012), .C1(
        n1074), .C2(n1011), .ZN(register_file_inst1_n2261) );
  OAI222D1BWP12T U2111 ( .A1(n1013), .A2(n1079), .B1(n1080), .B2(n1012), .C1(
        n1081), .C2(n1011), .ZN(register_file_inst1_n2357) );
  INVD0BWP12T U2112 ( .I(n1014), .ZN(n1016) );
  XOR2D1BWP12T U2113 ( .A1(n1018), .A2(n1017), .Z(
        register_file_inst1_pc_write_in_plus_two[23]) );
  INVD1BWP12T U2114 ( .I(register_file_inst1_r11_29_), .ZN(n1606) );
  OAI222D1BWP12T U2115 ( .A1(n1606), .A2(n1021), .B1(n1020), .B2(n1031), .C1(
        n1019), .C2(n1030), .ZN(register_file_inst1_n2294) );
  INVD1BWP12T U2116 ( .I(register_file_inst1_r7_29_), .ZN(n1592) );
  OAI222D1BWP12T U2117 ( .A1(n1592), .A2(n1051), .B1(n1050), .B2(n1031), .C1(
        n1049), .C2(n1030), .ZN(register_file_inst1_n2422) );
  CKND0BWP12T U2118 ( .I(register_file_inst1_lr_29_), .ZN(n1022) );
  OAI222D1BWP12T U2119 ( .A1(n1022), .A2(n1082), .B1(n1084), .B2(n1031), .C1(
        n1085), .C2(n1030), .ZN(register_file_inst1_n2230) );
  INVD1BWP12T U2120 ( .I(register_file_inst1_r4_29_), .ZN(n1605) );
  OAI222D1BWP12T U2121 ( .A1(n1605), .A2(n1090), .B1(n1091), .B2(n1031), .C1(
        n1092), .C2(n1030), .ZN(register_file_inst1_n2518) );
  CKND0BWP12T U2122 ( .I(register_file_inst1_r6_29_), .ZN(n1023) );
  OAI222D1BWP12T U2123 ( .A1(n1023), .A2(n1045), .B1(n1044), .B2(n1031), .C1(
        n1043), .C2(n1030), .ZN(register_file_inst1_n2454) );
  CKND0BWP12T U2124 ( .I(STACK_RF_next_sp[29]), .ZN(n1024) );
  OAI222D1BWP12T U2125 ( .A1(n1024), .A2(n1099), .B1(n1102), .B2(n1031), .C1(
        n1104), .C2(n1030), .ZN(register_file_inst1_spin[29]) );
  INVD1BWP12T U2126 ( .I(register_file_inst1_r1_29_), .ZN(n1590) );
  OAI222D1BWP12T U2127 ( .A1(n1590), .A2(n1093), .B1(n1094), .B2(n1031), .C1(
        n1095), .C2(n1030), .ZN(register_file_inst1_n2614) );
  CKND0BWP12T U2128 ( .I(register_file_inst1_r0_29_), .ZN(n1025) );
  OAI222D1BWP12T U2129 ( .A1(n1025), .A2(n1086), .B1(n1088), .B2(n1031), .C1(
        n1089), .C2(n1030), .ZN(register_file_inst1_n2646) );
  INVD1BWP12T U2130 ( .I(register_file_inst1_r5_29_), .ZN(n1607) );
  OAI222D1BWP12T U2131 ( .A1(n1607), .A2(n1096), .B1(n1097), .B2(n1031), .C1(
        n1098), .C2(n1030), .ZN(register_file_inst1_n2486) );
  CKND0BWP12T U2132 ( .I(register_file_inst1_tmp1_29_), .ZN(n1028) );
  OAI222D1BWP12T U2133 ( .A1(n1028), .A2(n1027), .B1(n1026), .B2(n1031), .C1(
        n2168), .C2(n1030), .ZN(register_file_inst1_n2166) );
  INVD1BWP12T U2134 ( .I(register_file_inst1_r9_29_), .ZN(n1591) );
  OAI222D1BWP12T U2135 ( .A1(n1591), .A2(n1079), .B1(n1080), .B2(n1031), .C1(
        n1081), .C2(n1030), .ZN(register_file_inst1_n2358) );
  CKND0BWP12T U2136 ( .I(register_file_inst1_r8_29_), .ZN(n1029) );
  OAI222D1BWP12T U2137 ( .A1(n1029), .A2(n1075), .B1(n1077), .B2(n1031), .C1(
        n1078), .C2(n1030), .ZN(register_file_inst1_n2390) );
  CKND0BWP12T U2138 ( .I(register_file_inst1_r12_29_), .ZN(n1032) );
  OAI222D1BWP12T U2139 ( .A1(n1032), .A2(n1071), .B1(n1073), .B2(n1031), .C1(
        n1074), .C2(n1030), .ZN(register_file_inst1_n2262) );
  INVD1BWP12T U2140 ( .I(n1033), .ZN(n1035) );
  XNR2D1BWP12T U2141 ( .A1(n1035), .A2(n1034), .ZN(
        register_file_inst1_pc_write_in_plus_two[24]) );
  XOR2D1BWP12T U2142 ( .A1(n11), .A2(n1036), .Z(
        register_file_inst1_pc_write_in_plus_two[25]) );
  CKND0BWP12T U2143 ( .I(STACK_RF_next_sp[30]), .ZN(n1038) );
  OAI222D1BWP12T U2144 ( .A1(n1038), .A2(n1037), .B1(n1102), .B2(n1055), .C1(
        n1104), .C2(n1054), .ZN(register_file_inst1_spin[30]) );
  CKND0BWP12T U2145 ( .I(register_file_inst1_r2_30_), .ZN(n1039) );
  OAI222D1BWP12T U2146 ( .A1(n1039), .A2(n1060), .B1(n1062), .B2(n1055), .C1(
        n1063), .C2(n1054), .ZN(register_file_inst1_n2583) );
  CKND0BWP12T U2147 ( .I(register_file_inst1_r3_30_), .ZN(n1040) );
  OAI222D1BWP12T U2148 ( .A1(n1040), .A2(n1064), .B1(n1066), .B2(n1055), .C1(
        n1067), .C2(n1054), .ZN(register_file_inst1_n2551) );
  OAI222D1BWP12T U2149 ( .A1(n1041), .A2(n1068), .B1(n1069), .B2(n1055), .C1(
        n1070), .C2(n1054), .ZN(register_file_inst1_n2327) );
  INVD1BWP12T U2150 ( .I(register_file_inst1_r1_30_), .ZN(n1618) );
  OAI222D1BWP12T U2151 ( .A1(n1618), .A2(n1093), .B1(n1094), .B2(n1055), .C1(
        n1095), .C2(n1054), .ZN(register_file_inst1_n2615) );
  OAI222D1BWP12T U2152 ( .A1(n1042), .A2(n1096), .B1(n1097), .B2(n1055), .C1(
        n1098), .C2(n1054), .ZN(register_file_inst1_n2487) );
  CKND0BWP12T U2153 ( .I(register_file_inst1_r6_30_), .ZN(n1046) );
  OAI222D1BWP12T U2154 ( .A1(n1046), .A2(n1045), .B1(n1044), .B2(n1055), .C1(
        n1043), .C2(n1054), .ZN(register_file_inst1_n2455) );
  CKND0BWP12T U2155 ( .I(register_file_inst1_r0_30_), .ZN(n1047) );
  OAI222D1BWP12T U2156 ( .A1(n1047), .A2(n1086), .B1(n1088), .B2(n1055), .C1(
        n1089), .C2(n1054), .ZN(register_file_inst1_n2647) );
  OAI222D1BWP12T U2157 ( .A1(n1048), .A2(n1090), .B1(n1091), .B2(n1055), .C1(
        n1092), .C2(n1054), .ZN(register_file_inst1_n2519) );
  INVD1BWP12T U2158 ( .I(register_file_inst1_r7_30_), .ZN(n1620) );
  OAI222D1BWP12T U2159 ( .A1(n1620), .A2(n1051), .B1(n1050), .B2(n1055), .C1(
        n1049), .C2(n1054), .ZN(register_file_inst1_n2423) );
  CKND0BWP12T U2160 ( .I(register_file_inst1_lr_30_), .ZN(n1052) );
  OAI222D1BWP12T U2161 ( .A1(n1052), .A2(n1082), .B1(n1084), .B2(n1055), .C1(
        n1085), .C2(n1054), .ZN(register_file_inst1_n2231) );
  CKND0BWP12T U2162 ( .I(register_file_inst1_r12_30_), .ZN(n1053) );
  OAI222D1BWP12T U2163 ( .A1(n1053), .A2(n1071), .B1(n1073), .B2(n1055), .C1(
        n1074), .C2(n1054), .ZN(register_file_inst1_n2263) );
  INVD1BWP12T U2164 ( .I(register_file_inst1_r9_30_), .ZN(n1619) );
  OAI222D1BWP12T U2165 ( .A1(n1619), .A2(n1079), .B1(n1080), .B2(n1055), .C1(
        n1081), .C2(n1054), .ZN(register_file_inst1_n2359) );
  CKND0BWP12T U2166 ( .I(register_file_inst1_r8_30_), .ZN(n1056) );
  OAI222D1BWP12T U2167 ( .A1(n1056), .A2(n1075), .B1(n1077), .B2(n1055), .C1(
        n1078), .C2(n1054), .ZN(register_file_inst1_n2391) );
  INVD1BWP12T U2168 ( .I(n1057), .ZN(n1059) );
  XNR2D1BWP12T U2169 ( .A1(n1059), .A2(n1058), .ZN(
        register_file_inst1_pc_write_in_plus_two[26]) );
  INVD1BWP12T U2170 ( .I(ALU_OUT_z), .ZN(n2292) );
  CKND0BWP12T U2171 ( .I(register_file_inst1_r2_31_), .ZN(n1061) );
  OAI222D1BWP12T U2172 ( .A1(n1063), .A2(n1103), .B1(n1062), .B2(n1101), .C1(
        n1061), .C2(n1060), .ZN(register_file_inst1_n2584) );
  CKND0BWP12T U2173 ( .I(register_file_inst1_r3_31_), .ZN(n1065) );
  OAI222D1BWP12T U2174 ( .A1(n1067), .A2(n1103), .B1(n1066), .B2(n1101), .C1(
        n1065), .C2(n1064), .ZN(register_file_inst1_n2552) );
  INVD1BWP12T U2175 ( .I(register_file_inst1_r10_31_), .ZN(n1643) );
  OAI222D1BWP12T U2176 ( .A1(n1070), .A2(n1103), .B1(n1069), .B2(n1101), .C1(
        n1643), .C2(n1068), .ZN(register_file_inst1_n2328) );
  CKND0BWP12T U2177 ( .I(register_file_inst1_r12_31_), .ZN(n1072) );
  OAI222D1BWP12T U2178 ( .A1(n1074), .A2(n1103), .B1(n1073), .B2(n1101), .C1(
        n1072), .C2(n1071), .ZN(register_file_inst1_n2264) );
  CKND0BWP12T U2179 ( .I(register_file_inst1_r8_31_), .ZN(n1076) );
  OAI222D1BWP12T U2180 ( .A1(n1078), .A2(n1103), .B1(n1077), .B2(n1101), .C1(
        n1076), .C2(n1075), .ZN(register_file_inst1_n2392) );
  INVD1BWP12T U2181 ( .I(register_file_inst1_r9_31_), .ZN(n1631) );
  OAI222D1BWP12T U2182 ( .A1(n1081), .A2(n1103), .B1(n1080), .B2(n1101), .C1(
        n1631), .C2(n1079), .ZN(register_file_inst1_n2360) );
  CKND0BWP12T U2183 ( .I(register_file_inst1_lr_31_), .ZN(n1083) );
  OAI222D1BWP12T U2184 ( .A1(n1085), .A2(n1103), .B1(n1084), .B2(n1101), .C1(
        n1083), .C2(n1082), .ZN(register_file_inst1_n2232) );
  CKND0BWP12T U2185 ( .I(register_file_inst1_r0_31_), .ZN(n1087) );
  OAI222D1BWP12T U2186 ( .A1(n1089), .A2(n1103), .B1(n1088), .B2(n1101), .C1(
        n1087), .C2(n1086), .ZN(register_file_inst1_n2648) );
  INVD1BWP12T U2187 ( .I(register_file_inst1_r4_31_), .ZN(n1644) );
  OAI222D1BWP12T U2188 ( .A1(n1092), .A2(n1103), .B1(n1091), .B2(n1101), .C1(
        n1644), .C2(n1090), .ZN(register_file_inst1_n2520) );
  INVD1BWP12T U2189 ( .I(register_file_inst1_r1_31_), .ZN(n1630) );
  OAI222D1BWP12T U2190 ( .A1(n1095), .A2(n1103), .B1(n1094), .B2(n1101), .C1(
        n1630), .C2(n1093), .ZN(register_file_inst1_n2616) );
  INVD1BWP12T U2191 ( .I(register_file_inst1_r5_31_), .ZN(n1646) );
  OAI222D1BWP12T U2192 ( .A1(n1098), .A2(n1103), .B1(n1097), .B2(n1101), .C1(
        n1646), .C2(n1096), .ZN(register_file_inst1_n2488) );
  CKND0BWP12T U2193 ( .I(STACK_RF_next_sp[31]), .ZN(n1100) );
  OAI222D1BWP12T U2194 ( .A1(n1104), .A2(n1103), .B1(n1102), .B2(n1101), .C1(
        n1100), .C2(n1099), .ZN(register_file_inst1_spin[31]) );
  XOR2D1BWP12T U2195 ( .A1(n12), .A2(n1105), .Z(
        register_file_inst1_pc_write_in_plus_two[27]) );
  INVD1BWP12T U2196 ( .I(n1106), .ZN(n1108) );
  XNR2D1BWP12T U2197 ( .A1(n1108), .A2(n1107), .ZN(
        register_file_inst1_pc_write_in_plus_two[28]) );
  INVD1BWP12T U2198 ( .I(ALU_OUT_v), .ZN(n2296) );
  XOR2D1BWP12T U2199 ( .A1(n13), .A2(n1109), .Z(
        register_file_inst1_pc_write_in_plus_two[29]) );
  INVD1BWP12T U2200 ( .I(n1110), .ZN(n1112) );
  XNR2D1BWP12T U2201 ( .A1(n1112), .A2(n1111), .ZN(
        register_file_inst1_pc_write_in_plus_two[30]) );
  OAI22D1BWP12T U2202 ( .A1(n1114), .A2(n1798), .B1(n1113), .B2(n1796), .ZN(
        n1121) );
  OAI22D1BWP12T U2203 ( .A1(n2218), .A2(n1802), .B1(n1115), .B2(n1800), .ZN(
        n1120) );
  OAI22D1BWP12T U2204 ( .A1(n1117), .A2(n1805), .B1(n1116), .B2(n1803), .ZN(
        n1119) );
  OAI22D1BWP12T U2205 ( .A1(n1136), .A2(n1809), .B1(n1138), .B2(n1807), .ZN(
        n1118) );
  NR4D0BWP12T U2206 ( .A1(n1121), .A2(n1120), .A3(n1119), .A4(n1118), .ZN(
        n1134) );
  CKND2D1BWP12T U2207 ( .A1(register_file_inst1_r9_18_), .A2(n1911), .ZN(n1123) );
  CKND2D1BWP12T U2208 ( .A1(register_file_inst1_r8_18_), .A2(n1910), .ZN(n1122) );
  ND3D1BWP12T U2209 ( .A1(n2219), .A2(n1123), .A3(n1122), .ZN(n1132) );
  OAI22D1BWP12T U2210 ( .A1(n1125), .A2(n1903), .B1(n1124), .B2(n1901), .ZN(
        n1131) );
  OAI22D1BWP12T U2211 ( .A1(n1126), .A2(n1907), .B1(n1135), .B2(n1905), .ZN(
        n1130) );
  OAI22D1BWP12T U2212 ( .A1(n1128), .A2(n1823), .B1(n1127), .B2(n1821), .ZN(
        n1129) );
  NR4D0BWP12T U2213 ( .A1(n1132), .A2(n1131), .A3(n1130), .A4(n1129), .ZN(
        n1133) );
  ND2D1BWP12T U2214 ( .A1(n1134), .A2(n1133), .ZN(RF_ALU_STACK_operand_a[18])
         );
  OAI22D1BWP12T U2215 ( .A1(n1136), .A2(n1873), .B1(n1135), .B2(n1871), .ZN(
        n1147) );
  OAI22D1BWP12T U2216 ( .A1(n1138), .A2(n1877), .B1(n1137), .B2(n1875), .ZN(
        n1146) );
  AOI22D1BWP12T U2217 ( .A1(register_file_inst1_tmp1_18_), .A2(n1835), .B1(
        register_file_inst1_r0_18_), .B2(n1633), .ZN(n1140) );
  AOI22D1BWP12T U2218 ( .A1(register_file_inst1_r5_18_), .A2(n1868), .B1(
        STACK_RF_next_sp[18]), .B2(n1867), .ZN(n1139) );
  ND3D1BWP12T U2219 ( .A1(n1140), .A2(n1139), .A3(n2142), .ZN(n1145) );
  AOI22D1BWP12T U2220 ( .A1(register_file_inst1_r12_18_), .A2(n1659), .B1(
        register_file_inst1_r8_18_), .B2(n1838), .ZN(n1143) );
  AOI22D1BWP12T U2221 ( .A1(register_file_inst1_r4_18_), .A2(n1595), .B1(
        register_file_inst1_r3_18_), .B2(n1839), .ZN(n1142) );
  AOI22D1BWP12T U2222 ( .A1(register_file_inst1_r6_18_), .A2(n1596), .B1(
        register_file_inst1_r10_18_), .B2(n1840), .ZN(n1141) );
  ND4D1BWP12T U2223 ( .A1(n1143), .A2(n1142), .A3(n2143), .A4(n1141), .ZN(
        n1144) );
  OR4XD1BWP12T U2224 ( .A1(n1147), .A2(n1146), .A3(n1145), .A4(n1144), .Z(
        RF_ALU_operand_b[18]) );
  OAI22D1BWP12T U2225 ( .A1(n1164), .A2(n1873), .B1(n1173), .B2(n1871), .ZN(
        n1157) );
  OAI22D1BWP12T U2226 ( .A1(n1163), .A2(n1877), .B1(n1148), .B2(n1875), .ZN(
        n1156) );
  AOI22D1BWP12T U2227 ( .A1(register_file_inst1_tmp1_17_), .A2(n1835), .B1(
        register_file_inst1_r0_17_), .B2(n1633), .ZN(n1150) );
  AOI22D1BWP12T U2228 ( .A1(register_file_inst1_r5_17_), .A2(n1868), .B1(
        STACK_RF_next_sp[17]), .B2(n1867), .ZN(n1149) );
  ND3D1BWP12T U2229 ( .A1(n1150), .A2(n1149), .A3(n2140), .ZN(n1155) );
  AOI22D1BWP12T U2230 ( .A1(register_file_inst1_r12_17_), .A2(n1659), .B1(
        register_file_inst1_r8_17_), .B2(n1838), .ZN(n1153) );
  AOI22D1BWP12T U2231 ( .A1(register_file_inst1_r4_17_), .A2(n1595), .B1(
        register_file_inst1_r3_17_), .B2(n1839), .ZN(n1152) );
  AOI22D1BWP12T U2232 ( .A1(register_file_inst1_r6_17_), .A2(n1596), .B1(
        register_file_inst1_r10_17_), .B2(n1840), .ZN(n1151) );
  ND4D1BWP12T U2233 ( .A1(n1153), .A2(n1152), .A3(n2141), .A4(n1151), .ZN(
        n1154) );
  OR4XD1BWP12T U2234 ( .A1(n1157), .A2(n1156), .A3(n1155), .A4(n1154), .Z(
        RF_ALU_operand_b[17]) );
  OAI22D1BWP12T U2235 ( .A1(n1159), .A2(n1798), .B1(n1158), .B2(n1796), .ZN(
        n1168) );
  OAI22D1BWP12T U2236 ( .A1(n2216), .A2(n1802), .B1(n1160), .B2(n1800), .ZN(
        n1167) );
  OAI22D1BWP12T U2237 ( .A1(n1162), .A2(n1805), .B1(n1161), .B2(n1803), .ZN(
        n1166) );
  OAI22D1BWP12T U2238 ( .A1(n1164), .A2(n1809), .B1(n1163), .B2(n1807), .ZN(
        n1165) );
  NR4D0BWP12T U2239 ( .A1(n1168), .A2(n1167), .A3(n1166), .A4(n1165), .ZN(
        n1182) );
  CKND2D1BWP12T U2240 ( .A1(register_file_inst1_r9_17_), .A2(n1911), .ZN(n1170) );
  ND2D1BWP12T U2241 ( .A1(register_file_inst1_r8_17_), .A2(n1910), .ZN(n1169)
         );
  ND3D1BWP12T U2242 ( .A1(n2217), .A2(n1170), .A3(n1169), .ZN(n1180) );
  OAI22D1BWP12T U2243 ( .A1(n1172), .A2(n1903), .B1(n1171), .B2(n1901), .ZN(
        n1179) );
  OAI22D1BWP12T U2244 ( .A1(n1174), .A2(n1907), .B1(n1173), .B2(n1905), .ZN(
        n1178) );
  OAI22D1BWP12T U2245 ( .A1(n1176), .A2(n1823), .B1(n1175), .B2(n1821), .ZN(
        n1177) );
  NR4D0BWP12T U2246 ( .A1(n1180), .A2(n1179), .A3(n1178), .A4(n1177), .ZN(
        n1181) );
  ND2D1BWP12T U2247 ( .A1(n1182), .A2(n1181), .ZN(RF_ALU_STACK_operand_a[17])
         );
  OAI22D1BWP12T U2248 ( .A1(n1184), .A2(n1798), .B1(n1183), .B2(n1796), .ZN(
        n1191) );
  OAI22D1BWP12T U2249 ( .A1(n2214), .A2(n1802), .B1(n1185), .B2(n1800), .ZN(
        n1190) );
  OAI22D1BWP12T U2250 ( .A1(n1187), .A2(n1805), .B1(n1186), .B2(n1803), .ZN(
        n1189) );
  OAI22D1BWP12T U2251 ( .A1(n1206), .A2(n1809), .B1(n1208), .B2(n1807), .ZN(
        n1188) );
  NR4D0BWP12T U2252 ( .A1(n1191), .A2(n1190), .A3(n1189), .A4(n1188), .ZN(
        n1204) );
  CKND2D1BWP12T U2253 ( .A1(register_file_inst1_r9_16_), .A2(n1911), .ZN(n1193) );
  CKND2D1BWP12T U2254 ( .A1(register_file_inst1_r8_16_), .A2(n1910), .ZN(n1192) );
  ND3D1BWP12T U2255 ( .A1(n2215), .A2(n1193), .A3(n1192), .ZN(n1202) );
  OAI22D1BWP12T U2256 ( .A1(n1195), .A2(n1903), .B1(n1194), .B2(n1901), .ZN(
        n1201) );
  OAI22D1BWP12T U2257 ( .A1(n1196), .A2(n1907), .B1(n1205), .B2(n1905), .ZN(
        n1200) );
  OAI22D1BWP12T U2258 ( .A1(n1198), .A2(n1823), .B1(n1197), .B2(n1821), .ZN(
        n1199) );
  NR4D0BWP12T U2259 ( .A1(n1202), .A2(n1201), .A3(n1200), .A4(n1199), .ZN(
        n1203) );
  ND2D1BWP12T U2260 ( .A1(n1204), .A2(n1203), .ZN(RF_ALU_STACK_operand_a[16])
         );
  OAI22D1BWP12T U2261 ( .A1(n1206), .A2(n1873), .B1(n1205), .B2(n1871), .ZN(
        n1217) );
  OAI22D1BWP12T U2262 ( .A1(n1208), .A2(n1877), .B1(n1207), .B2(n1875), .ZN(
        n1216) );
  AOI22D1BWP12T U2263 ( .A1(register_file_inst1_tmp1_16_), .A2(n1835), .B1(
        register_file_inst1_r0_16_), .B2(n1633), .ZN(n1210) );
  AOI22D1BWP12T U2264 ( .A1(register_file_inst1_r5_16_), .A2(n1868), .B1(
        STACK_RF_next_sp[16]), .B2(n1867), .ZN(n1209) );
  ND3D1BWP12T U2265 ( .A1(n1210), .A2(n1209), .A3(n2138), .ZN(n1215) );
  AOI22D1BWP12T U2266 ( .A1(register_file_inst1_r12_16_), .A2(n1659), .B1(
        register_file_inst1_r8_16_), .B2(n1838), .ZN(n1213) );
  AOI22D1BWP12T U2267 ( .A1(register_file_inst1_r4_16_), .A2(n1595), .B1(
        register_file_inst1_r3_16_), .B2(n1839), .ZN(n1212) );
  AOI22D1BWP12T U2268 ( .A1(register_file_inst1_r6_16_), .A2(n1596), .B1(
        register_file_inst1_r10_16_), .B2(n1840), .ZN(n1211) );
  ND4D1BWP12T U2269 ( .A1(n1213), .A2(n1212), .A3(n2139), .A4(n1211), .ZN(
        n1214) );
  OR4XD1BWP12T U2270 ( .A1(n1217), .A2(n1216), .A3(n1215), .A4(n1214), .Z(
        RF_ALU_operand_b[16]) );
  OAI22D1BWP12T U2271 ( .A1(n1234), .A2(n1873), .B1(n1243), .B2(n1871), .ZN(
        n1227) );
  OAI22D1BWP12T U2272 ( .A1(n1233), .A2(n1877), .B1(n1218), .B2(n1875), .ZN(
        n1226) );
  AOI22D1BWP12T U2273 ( .A1(register_file_inst1_tmp1_15_), .A2(n1835), .B1(
        register_file_inst1_r0_15_), .B2(n1633), .ZN(n1220) );
  AOI22D1BWP12T U2274 ( .A1(register_file_inst1_r5_15_), .A2(n1868), .B1(
        STACK_RF_next_sp[15]), .B2(n1867), .ZN(n1219) );
  ND3D1BWP12T U2275 ( .A1(n1220), .A2(n1219), .A3(n2136), .ZN(n1225) );
  AOI22D1BWP12T U2276 ( .A1(register_file_inst1_r12_15_), .A2(n1659), .B1(
        register_file_inst1_r8_15_), .B2(n1838), .ZN(n1223) );
  AOI22D1BWP12T U2277 ( .A1(register_file_inst1_r4_15_), .A2(n1595), .B1(
        register_file_inst1_r3_15_), .B2(n1839), .ZN(n1222) );
  AOI22D1BWP12T U2278 ( .A1(register_file_inst1_r6_15_), .A2(n1596), .B1(
        register_file_inst1_r10_15_), .B2(n1840), .ZN(n1221) );
  ND4D1BWP12T U2279 ( .A1(n1223), .A2(n1222), .A3(n2137), .A4(n1221), .ZN(
        n1224) );
  OR4XD1BWP12T U2280 ( .A1(n1227), .A2(n1226), .A3(n1225), .A4(n1224), .Z(
        RF_ALU_operand_b[15]) );
  OAI22D1BWP12T U2281 ( .A1(n1229), .A2(n1798), .B1(n1228), .B2(n1796), .ZN(
        n1238) );
  OAI22D1BWP12T U2282 ( .A1(n2212), .A2(n1802), .B1(n1230), .B2(n1800), .ZN(
        n1237) );
  OAI22D1BWP12T U2283 ( .A1(n1232), .A2(n1805), .B1(n1231), .B2(n1803), .ZN(
        n1236) );
  OAI22D1BWP12T U2284 ( .A1(n1234), .A2(n1809), .B1(n1233), .B2(n1807), .ZN(
        n1235) );
  NR4D0BWP12T U2285 ( .A1(n1238), .A2(n1237), .A3(n1236), .A4(n1235), .ZN(
        n1252) );
  CKND2D1BWP12T U2286 ( .A1(register_file_inst1_r9_15_), .A2(n1911), .ZN(n1240) );
  ND2D1BWP12T U2287 ( .A1(register_file_inst1_r8_15_), .A2(n1910), .ZN(n1239)
         );
  ND3D1BWP12T U2288 ( .A1(n2213), .A2(n1240), .A3(n1239), .ZN(n1250) );
  OAI22D1BWP12T U2289 ( .A1(n1242), .A2(n1903), .B1(n1241), .B2(n1901), .ZN(
        n1249) );
  OAI22D1BWP12T U2290 ( .A1(n1244), .A2(n1907), .B1(n1243), .B2(n1905), .ZN(
        n1248) );
  OAI22D1BWP12T U2291 ( .A1(n1246), .A2(n1823), .B1(n1245), .B2(n1821), .ZN(
        n1247) );
  NR4D0BWP12T U2292 ( .A1(n1250), .A2(n1249), .A3(n1248), .A4(n1247), .ZN(
        n1251) );
  ND2D1BWP12T U2293 ( .A1(n1252), .A2(n1251), .ZN(RF_ALU_STACK_operand_a[15])
         );
  OAI22D1BWP12T U2294 ( .A1(n1254), .A2(n1873), .B1(n1253), .B2(n1871), .ZN(
        n1265) );
  OAI22D1BWP12T U2295 ( .A1(n1256), .A2(n1877), .B1(n1255), .B2(n1875), .ZN(
        n1264) );
  AOI22D1BWP12T U2296 ( .A1(register_file_inst1_tmp1_14_), .A2(n1835), .B1(
        register_file_inst1_r0_14_), .B2(n1633), .ZN(n1258) );
  AOI22D1BWP12T U2297 ( .A1(register_file_inst1_r5_14_), .A2(n1868), .B1(
        STACK_RF_next_sp[14]), .B2(n1867), .ZN(n1257) );
  ND3D1BWP12T U2298 ( .A1(n1258), .A2(n1257), .A3(n2133), .ZN(n1263) );
  AOI22D1BWP12T U2299 ( .A1(register_file_inst1_r12_14_), .A2(n1659), .B1(
        register_file_inst1_r8_14_), .B2(n1838), .ZN(n1261) );
  AOI22D1BWP12T U2300 ( .A1(register_file_inst1_r4_14_), .A2(n1595), .B1(
        register_file_inst1_r3_14_), .B2(n1839), .ZN(n1260) );
  AOI22D1BWP12T U2301 ( .A1(register_file_inst1_r6_14_), .A2(n1596), .B1(
        register_file_inst1_r10_14_), .B2(n1840), .ZN(n1259) );
  ND4D1BWP12T U2302 ( .A1(n1261), .A2(n1260), .A3(n2134), .A4(n1259), .ZN(
        n1262) );
  OR4XD1BWP12T U2303 ( .A1(n1265), .A2(n1264), .A3(n1263), .A4(n1262), .Z(
        RF_ALU_operand_b[14]) );
  OAI22D1BWP12T U2304 ( .A1(n1282), .A2(n1873), .B1(n1291), .B2(n1871), .ZN(
        n1275) );
  OAI22D1BWP12T U2305 ( .A1(n1281), .A2(n1877), .B1(n1266), .B2(n1875), .ZN(
        n1274) );
  AOI22D1BWP12T U2306 ( .A1(register_file_inst1_tmp1_13_), .A2(n1835), .B1(
        register_file_inst1_r0_13_), .B2(n1633), .ZN(n1268) );
  AOI22D1BWP12T U2307 ( .A1(register_file_inst1_r5_13_), .A2(n1868), .B1(
        STACK_RF_next_sp[13]), .B2(n1867), .ZN(n1267) );
  ND3D1BWP12T U2308 ( .A1(n1268), .A2(n1267), .A3(n2130), .ZN(n1273) );
  AOI22D1BWP12T U2309 ( .A1(register_file_inst1_r12_13_), .A2(n1659), .B1(
        register_file_inst1_r8_13_), .B2(n1838), .ZN(n1271) );
  AOI22D1BWP12T U2310 ( .A1(register_file_inst1_r4_13_), .A2(n1595), .B1(
        register_file_inst1_r3_13_), .B2(n1839), .ZN(n1270) );
  AOI22D1BWP12T U2311 ( .A1(register_file_inst1_r6_13_), .A2(n1596), .B1(
        register_file_inst1_r10_13_), .B2(n1840), .ZN(n1269) );
  ND4D1BWP12T U2312 ( .A1(n1271), .A2(n1270), .A3(n2131), .A4(n1269), .ZN(
        n1272) );
  OR4XD1BWP12T U2313 ( .A1(n1275), .A2(n1274), .A3(n1273), .A4(n1272), .Z(
        RF_ALU_operand_b[13]) );
  OAI22D1BWP12T U2314 ( .A1(n1277), .A2(n1798), .B1(n1276), .B2(n1796), .ZN(
        n1286) );
  OAI22D1BWP12T U2315 ( .A1(n2208), .A2(n1802), .B1(n1278), .B2(n1800), .ZN(
        n1285) );
  OAI22D1BWP12T U2316 ( .A1(n1280), .A2(n1805), .B1(n1279), .B2(n1803), .ZN(
        n1284) );
  OAI22D1BWP12T U2317 ( .A1(n1282), .A2(n1809), .B1(n1281), .B2(n1807), .ZN(
        n1283) );
  NR4D0BWP12T U2318 ( .A1(n1286), .A2(n1285), .A3(n1284), .A4(n1283), .ZN(
        n1300) );
  CKND2D1BWP12T U2319 ( .A1(register_file_inst1_r9_13_), .A2(n1911), .ZN(n1288) );
  ND2D1BWP12T U2320 ( .A1(register_file_inst1_r8_13_), .A2(n1910), .ZN(n1287)
         );
  ND3D1BWP12T U2321 ( .A1(n2209), .A2(n1288), .A3(n1287), .ZN(n1298) );
  OAI22D1BWP12T U2322 ( .A1(n1290), .A2(n1903), .B1(n1289), .B2(n1901), .ZN(
        n1297) );
  OAI22D1BWP12T U2323 ( .A1(n1292), .A2(n1907), .B1(n1291), .B2(n1905), .ZN(
        n1296) );
  OAI22D1BWP12T U2324 ( .A1(n1294), .A2(n1823), .B1(n1293), .B2(n1821), .ZN(
        n1295) );
  NR4D0BWP12T U2325 ( .A1(n1298), .A2(n1297), .A3(n1296), .A4(n1295), .ZN(
        n1299) );
  ND2D1BWP12T U2326 ( .A1(n1300), .A2(n1299), .ZN(RF_ALU_STACK_operand_a[13])
         );
  INVD1BWP12T U2327 ( .I(STACK_RF_next_sp[12]), .ZN(n1301) );
  OAI22D1BWP12T U2328 ( .A1(n1302), .A2(n1798), .B1(n1301), .B2(n1796), .ZN(
        n1309) );
  OAI22D1BWP12T U2329 ( .A1(n2206), .A2(n1802), .B1(n1303), .B2(n1800), .ZN(
        n1308) );
  OAI22D1BWP12T U2330 ( .A1(n1305), .A2(n1805), .B1(n1304), .B2(n1803), .ZN(
        n1307) );
  OAI22D1BWP12T U2331 ( .A1(n1324), .A2(n1809), .B1(n1326), .B2(n1807), .ZN(
        n1306) );
  NR4D0BWP12T U2332 ( .A1(n1309), .A2(n1308), .A3(n1307), .A4(n1306), .ZN(
        n1322) );
  CKND2D1BWP12T U2333 ( .A1(register_file_inst1_r9_12_), .A2(n1911), .ZN(n1311) );
  CKND2D1BWP12T U2334 ( .A1(register_file_inst1_r8_12_), .A2(n1910), .ZN(n1310) );
  ND3D1BWP12T U2335 ( .A1(n2207), .A2(n1311), .A3(n1310), .ZN(n1320) );
  OAI22D1BWP12T U2336 ( .A1(n1313), .A2(n1903), .B1(n1312), .B2(n1901), .ZN(
        n1319) );
  OAI22D1BWP12T U2337 ( .A1(n1314), .A2(n1907), .B1(n1323), .B2(n1905), .ZN(
        n1318) );
  OAI22D1BWP12T U2338 ( .A1(n1316), .A2(n1823), .B1(n1315), .B2(n1821), .ZN(
        n1317) );
  NR4D0BWP12T U2339 ( .A1(n1320), .A2(n1319), .A3(n1318), .A4(n1317), .ZN(
        n1321) );
  ND2D1BWP12T U2340 ( .A1(n1322), .A2(n1321), .ZN(RF_ALU_STACK_operand_a[12])
         );
  OAI22D1BWP12T U2341 ( .A1(n1324), .A2(n1873), .B1(n1323), .B2(n1871), .ZN(
        n1335) );
  OAI22D1BWP12T U2342 ( .A1(n1326), .A2(n1877), .B1(n1325), .B2(n1875), .ZN(
        n1334) );
  INVD1BWP12T U2343 ( .I(n1633), .ZN(n1879) );
  AOI22D1BWP12T U2344 ( .A1(register_file_inst1_tmp1_12_), .A2(n1835), .B1(
        register_file_inst1_r0_12_), .B2(n1633), .ZN(n1328) );
  AOI22D1BWP12T U2345 ( .A1(register_file_inst1_r5_12_), .A2(n1868), .B1(
        STACK_RF_next_sp[12]), .B2(n1867), .ZN(n1327) );
  ND3D1BWP12T U2346 ( .A1(n1328), .A2(n1327), .A3(n2127), .ZN(n1333) );
  AOI22D1BWP12T U2347 ( .A1(register_file_inst1_r12_12_), .A2(n1659), .B1(
        register_file_inst1_r8_12_), .B2(n1838), .ZN(n1331) );
  AOI22D1BWP12T U2348 ( .A1(register_file_inst1_r4_12_), .A2(n1595), .B1(
        register_file_inst1_r3_12_), .B2(n1839), .ZN(n1330) );
  AOI22D1BWP12T U2349 ( .A1(register_file_inst1_r6_12_), .A2(n1596), .B1(
        register_file_inst1_r10_12_), .B2(n1840), .ZN(n1329) );
  ND4D1BWP12T U2350 ( .A1(n1331), .A2(n1330), .A3(n2128), .A4(n1329), .ZN(
        n1332) );
  OR4XD1BWP12T U2351 ( .A1(n1335), .A2(n1334), .A3(n1333), .A4(n1332), .Z(
        RF_ALU_operand_b[12]) );
  INVD1BWP12T U2352 ( .I(STACK_RF_next_sp[8]), .ZN(n1336) );
  OAI22D1BWP12T U2353 ( .A1(n1356), .A2(n1798), .B1(n1336), .B2(n1796), .ZN(
        n1343) );
  OAI22D1BWP12T U2354 ( .A1(n2198), .A2(n1802), .B1(n1337), .B2(n1800), .ZN(
        n1342) );
  OAI22D1BWP12T U2355 ( .A1(n1359), .A2(n1805), .B1(n1357), .B2(n1803), .ZN(
        n1341) );
  OAI22D1BWP12T U2356 ( .A1(n1339), .A2(n1809), .B1(n1338), .B2(n1807), .ZN(
        n1340) );
  NR4D0BWP12T U2357 ( .A1(n1343), .A2(n1342), .A3(n1341), .A4(n1340), .ZN(
        n1354) );
  CKND2D1BWP12T U2358 ( .A1(register_file_inst1_r9_8_), .A2(n1911), .ZN(n1345)
         );
  CKND2D1BWP12T U2359 ( .A1(register_file_inst1_r8_8_), .A2(n1910), .ZN(n1344)
         );
  ND3D1BWP12T U2360 ( .A1(n2199), .A2(n1345), .A3(n1344), .ZN(n1352) );
  OAI22D1BWP12T U2361 ( .A1(n1358), .A2(n1903), .B1(n1360), .B2(n1901), .ZN(
        n1351) );
  OAI22D1BWP12T U2362 ( .A1(n1347), .A2(n1907), .B1(n1346), .B2(n1905), .ZN(
        n1350) );
  OAI22D1BWP12T U2363 ( .A1(n1348), .A2(n1823), .B1(n1361), .B2(n1821), .ZN(
        n1349) );
  NR4D0BWP12T U2364 ( .A1(n1352), .A2(n1351), .A3(n1350), .A4(n1349), .ZN(
        n1353) );
  ND2D1BWP12T U2365 ( .A1(n1354), .A2(n1353), .ZN(RF_ALU_STACK_operand_a[8])
         );
  INVD1BWP12T U2366 ( .I(n1838), .ZN(n1848) );
  OAI22D1BWP12T U2367 ( .A1(n1356), .A2(n1850), .B1(n1355), .B2(n1848), .ZN(
        n1365) );
  INVD1BWP12T U2368 ( .I(n1839), .ZN(n1852) );
  OAI22D1BWP12T U2369 ( .A1(n1358), .A2(n1854), .B1(n1357), .B2(n1852), .ZN(
        n1364) );
  INVD1BWP12T U2370 ( .I(n1943), .ZN(n1856) );
  OAI22D1BWP12T U2371 ( .A1(n2198), .A2(n1858), .B1(n1359), .B2(n1856), .ZN(
        n1363) );
  INVD1BWP12T U2372 ( .I(n1840), .ZN(n1859) );
  OAI22D1BWP12T U2373 ( .A1(n1361), .A2(n1861), .B1(n1360), .B2(n1859), .ZN(
        n1362) );
  NR4D0BWP12T U2374 ( .A1(n1365), .A2(n1364), .A3(n1363), .A4(n1362), .ZN(
        n1371) );
  AOI22D1BWP12T U2375 ( .A1(register_file_inst1_tmp1_8_), .A2(n1835), .B1(
        register_file_inst1_r0_8_), .B2(n1633), .ZN(n1367) );
  AOI22D1BWP12T U2376 ( .A1(register_file_inst1_r5_8_), .A2(n1868), .B1(
        STACK_RF_next_sp[8]), .B2(n1867), .ZN(n1366) );
  AN3XD1BWP12T U2377 ( .A1(n1367), .A2(n1366), .A3(n2116), .Z(n1370) );
  AOI22D1BWP12T U2378 ( .A1(register_file_inst1_r1_8_), .A2(n1742), .B1(
        register_file_inst1_r11_8_), .B2(n1741), .ZN(n1369) );
  INVD1BWP12T U2379 ( .I(n1877), .ZN(n1744) );
  AOI22D1BWP12T U2380 ( .A1(register_file_inst1_r7_8_), .A2(n1744), .B1(
        register_file_inst1_r9_8_), .B2(n1743), .ZN(n1368) );
  ND4D1BWP12T U2381 ( .A1(n1371), .A2(n1370), .A3(n1369), .A4(n1368), .ZN(
        RF_ALU_operand_b[8]) );
  OAI22D1BWP12T U2382 ( .A1(n1388), .A2(n1873), .B1(n1397), .B2(n1871), .ZN(
        n1381) );
  OAI22D1BWP12T U2383 ( .A1(n1387), .A2(n1877), .B1(n1372), .B2(n1875), .ZN(
        n1380) );
  AOI22D1BWP12T U2384 ( .A1(register_file_inst1_tmp1_9_), .A2(n1835), .B1(
        register_file_inst1_r0_9_), .B2(n1633), .ZN(n1374) );
  AOI22D1BWP12T U2385 ( .A1(register_file_inst1_r5_9_), .A2(n1868), .B1(
        STACK_RF_next_sp[9]), .B2(n1867), .ZN(n1373) );
  ND3D1BWP12T U2386 ( .A1(n1374), .A2(n1373), .A3(n2118), .ZN(n1379) );
  AOI22D1BWP12T U2387 ( .A1(register_file_inst1_r12_9_), .A2(n1659), .B1(
        register_file_inst1_r8_9_), .B2(n1838), .ZN(n1377) );
  AOI22D1BWP12T U2388 ( .A1(register_file_inst1_r4_9_), .A2(n1595), .B1(
        register_file_inst1_r3_9_), .B2(n1839), .ZN(n1376) );
  AOI22D1BWP12T U2389 ( .A1(register_file_inst1_r6_9_), .A2(n1596), .B1(
        register_file_inst1_r10_9_), .B2(n1840), .ZN(n1375) );
  ND4D1BWP12T U2390 ( .A1(n1377), .A2(n1376), .A3(n2119), .A4(n1375), .ZN(
        n1378) );
  OR4XD1BWP12T U2391 ( .A1(n1381), .A2(n1380), .A3(n1379), .A4(n1378), .Z(
        RF_ALU_operand_b[9]) );
  INVD1BWP12T U2392 ( .I(STACK_RF_next_sp[9]), .ZN(n1382) );
  OAI22D1BWP12T U2393 ( .A1(n1383), .A2(n1798), .B1(n1382), .B2(n1796), .ZN(
        n1392) );
  OAI22D1BWP12T U2394 ( .A1(n2200), .A2(n1802), .B1(n1384), .B2(n1800), .ZN(
        n1391) );
  OAI22D1BWP12T U2395 ( .A1(n1386), .A2(n1805), .B1(n1385), .B2(n1803), .ZN(
        n1390) );
  OAI22D1BWP12T U2396 ( .A1(n1388), .A2(n1809), .B1(n1387), .B2(n1807), .ZN(
        n1389) );
  NR4D0BWP12T U2397 ( .A1(n1392), .A2(n1391), .A3(n1390), .A4(n1389), .ZN(
        n1406) );
  CKND2D1BWP12T U2398 ( .A1(register_file_inst1_r9_9_), .A2(n1911), .ZN(n1394)
         );
  ND2D1BWP12T U2399 ( .A1(register_file_inst1_r8_9_), .A2(n1910), .ZN(n1393)
         );
  ND3D1BWP12T U2400 ( .A1(n2201), .A2(n1394), .A3(n1393), .ZN(n1404) );
  OAI22D1BWP12T U2401 ( .A1(n1396), .A2(n1903), .B1(n1395), .B2(n1901), .ZN(
        n1403) );
  OAI22D1BWP12T U2402 ( .A1(n1398), .A2(n1907), .B1(n1397), .B2(n1905), .ZN(
        n1402) );
  OAI22D1BWP12T U2403 ( .A1(n1400), .A2(n1823), .B1(n1399), .B2(n1821), .ZN(
        n1401) );
  NR4D0BWP12T U2404 ( .A1(n1404), .A2(n1403), .A3(n1402), .A4(n1401), .ZN(
        n1405) );
  ND2D1BWP12T U2405 ( .A1(n1406), .A2(n1405), .ZN(RF_ALU_STACK_operand_a[9])
         );
  OAI22D1BWP12T U2406 ( .A1(n1408), .A2(n1873), .B1(n1407), .B2(n1871), .ZN(
        n1419) );
  OAI22D1BWP12T U2407 ( .A1(n1410), .A2(n1877), .B1(n1409), .B2(n1875), .ZN(
        n1418) );
  AOI22D1BWP12T U2408 ( .A1(register_file_inst1_tmp1_10_), .A2(n1835), .B1(
        register_file_inst1_r0_10_), .B2(n1633), .ZN(n1412) );
  AOI22D1BWP12T U2409 ( .A1(register_file_inst1_r5_10_), .A2(n1868), .B1(
        STACK_RF_next_sp[10]), .B2(n1867), .ZN(n1411) );
  ND3D1BWP12T U2410 ( .A1(n1412), .A2(n1411), .A3(n2121), .ZN(n1417) );
  AOI22D1BWP12T U2411 ( .A1(register_file_inst1_r12_10_), .A2(n1659), .B1(
        register_file_inst1_r8_10_), .B2(n1838), .ZN(n1415) );
  AOI22D1BWP12T U2412 ( .A1(register_file_inst1_r4_10_), .A2(n1595), .B1(
        register_file_inst1_r3_10_), .B2(n1839), .ZN(n1414) );
  AOI22D1BWP12T U2413 ( .A1(register_file_inst1_r6_10_), .A2(n1596), .B1(
        register_file_inst1_r10_10_), .B2(n1840), .ZN(n1413) );
  ND4D1BWP12T U2414 ( .A1(n1415), .A2(n1414), .A3(n2122), .A4(n1413), .ZN(
        n1416) );
  OR4XD1BWP12T U2415 ( .A1(n1419), .A2(n1418), .A3(n1417), .A4(n1416), .Z(
        RF_ALU_operand_b[10]) );
  OAI22D1BWP12T U2416 ( .A1(n1436), .A2(n1873), .B1(n1445), .B2(n1871), .ZN(
        n1429) );
  OAI22D1BWP12T U2417 ( .A1(n1435), .A2(n1877), .B1(n1420), .B2(n1875), .ZN(
        n1428) );
  AOI22D1BWP12T U2418 ( .A1(register_file_inst1_tmp1_11_), .A2(n1835), .B1(
        register_file_inst1_r0_11_), .B2(n1633), .ZN(n1422) );
  AOI22D1BWP12T U2419 ( .A1(register_file_inst1_r5_11_), .A2(n1868), .B1(
        STACK_RF_next_sp[11]), .B2(n1867), .ZN(n1421) );
  ND3D1BWP12T U2420 ( .A1(n1422), .A2(n1421), .A3(n2124), .ZN(n1427) );
  AOI22D1BWP12T U2421 ( .A1(register_file_inst1_r12_11_), .A2(n1659), .B1(
        register_file_inst1_r8_11_), .B2(n1838), .ZN(n1425) );
  AOI22D1BWP12T U2422 ( .A1(register_file_inst1_r4_11_), .A2(n1595), .B1(
        register_file_inst1_r3_11_), .B2(n1839), .ZN(n1424) );
  AOI22D1BWP12T U2423 ( .A1(register_file_inst1_r6_11_), .A2(n1596), .B1(
        register_file_inst1_r10_11_), .B2(n1840), .ZN(n1423) );
  ND4D1BWP12T U2424 ( .A1(n1425), .A2(n1424), .A3(n2125), .A4(n1423), .ZN(
        n1426) );
  OR4XD1BWP12T U2425 ( .A1(n1429), .A2(n1428), .A3(n1427), .A4(n1426), .Z(
        RF_ALU_operand_b[11]) );
  INVD1BWP12T U2426 ( .I(STACK_RF_next_sp[11]), .ZN(n1430) );
  OAI22D1BWP12T U2427 ( .A1(n1431), .A2(n1798), .B1(n1430), .B2(n1796), .ZN(
        n1440) );
  OAI22D1BWP12T U2428 ( .A1(n2204), .A2(n1802), .B1(n1432), .B2(n1800), .ZN(
        n1439) );
  OAI22D1BWP12T U2429 ( .A1(n1434), .A2(n1805), .B1(n1433), .B2(n1803), .ZN(
        n1438) );
  OAI22D1BWP12T U2430 ( .A1(n1436), .A2(n1809), .B1(n1435), .B2(n1807), .ZN(
        n1437) );
  NR4D0BWP12T U2431 ( .A1(n1440), .A2(n1439), .A3(n1438), .A4(n1437), .ZN(
        n1454) );
  CKND2D1BWP12T U2432 ( .A1(register_file_inst1_r9_11_), .A2(n1911), .ZN(n1442) );
  ND2D1BWP12T U2433 ( .A1(register_file_inst1_r8_11_), .A2(n1910), .ZN(n1441)
         );
  ND3D1BWP12T U2434 ( .A1(n2205), .A2(n1442), .A3(n1441), .ZN(n1452) );
  OAI22D1BWP12T U2435 ( .A1(n1444), .A2(n1903), .B1(n1443), .B2(n1901), .ZN(
        n1451) );
  OAI22D1BWP12T U2436 ( .A1(n1446), .A2(n1907), .B1(n1445), .B2(n1905), .ZN(
        n1450) );
  OAI22D1BWP12T U2437 ( .A1(n1448), .A2(n1823), .B1(n1447), .B2(n1821), .ZN(
        n1449) );
  NR4D0BWP12T U2438 ( .A1(n1452), .A2(n1451), .A3(n1450), .A4(n1449), .ZN(
        n1453) );
  ND2D1BWP12T U2439 ( .A1(n1454), .A2(n1453), .ZN(RF_ALU_STACK_operand_a[11])
         );
  INVD1BWP12T U2440 ( .I(STACK_RF_next_sp[6]), .ZN(n1455) );
  OAI22D1BWP12T U2441 ( .A1(n1456), .A2(n1798), .B1(n1455), .B2(n1796), .ZN(
        n1463) );
  OAI22D1BWP12T U2442 ( .A1(n2194), .A2(n1802), .B1(n1457), .B2(n1800), .ZN(
        n1462) );
  OAI22D1BWP12T U2443 ( .A1(n1459), .A2(n1805), .B1(n1458), .B2(n1803), .ZN(
        n1461) );
  OAI22D1BWP12T U2444 ( .A1(n1478), .A2(n1809), .B1(n1480), .B2(n1807), .ZN(
        n1460) );
  NR4D0BWP12T U2445 ( .A1(n1463), .A2(n1462), .A3(n1461), .A4(n1460), .ZN(
        n1476) );
  CKND2D1BWP12T U2446 ( .A1(register_file_inst1_r9_6_), .A2(n1911), .ZN(n1465)
         );
  ND2D1BWP12T U2447 ( .A1(register_file_inst1_r8_6_), .A2(n1910), .ZN(n1464)
         );
  ND3D1BWP12T U2448 ( .A1(n2195), .A2(n1465), .A3(n1464), .ZN(n1474) );
  OAI22D1BWP12T U2449 ( .A1(n1467), .A2(n1903), .B1(n1466), .B2(n1901), .ZN(
        n1473) );
  OAI22D1BWP12T U2450 ( .A1(n1468), .A2(n1907), .B1(n1477), .B2(n1905), .ZN(
        n1472) );
  OAI22D1BWP12T U2451 ( .A1(n1470), .A2(n1823), .B1(n1469), .B2(n1821), .ZN(
        n1471) );
  NR4D0BWP12T U2452 ( .A1(n1474), .A2(n1473), .A3(n1472), .A4(n1471), .ZN(
        n1475) );
  ND2D1BWP12T U2453 ( .A1(n1476), .A2(n1475), .ZN(RF_ALU_STACK_operand_a[6])
         );
  OAI22D1BWP12T U2454 ( .A1(n1478), .A2(n1873), .B1(n1477), .B2(n1871), .ZN(
        n1489) );
  OAI22D1BWP12T U2455 ( .A1(n1480), .A2(n1877), .B1(n1479), .B2(n1875), .ZN(
        n1488) );
  AOI22D1BWP12T U2456 ( .A1(register_file_inst1_tmp1_6_), .A2(n1835), .B1(
        register_file_inst1_r0_6_), .B2(n1633), .ZN(n1482) );
  AOI22D1BWP12T U2457 ( .A1(register_file_inst1_r5_6_), .A2(n1868), .B1(
        STACK_RF_next_sp[6]), .B2(n1867), .ZN(n1481) );
  ND3D1BWP12T U2458 ( .A1(n1482), .A2(n1481), .A3(n2111), .ZN(n1487) );
  AOI22D1BWP12T U2459 ( .A1(register_file_inst1_r12_6_), .A2(n1659), .B1(
        register_file_inst1_r8_6_), .B2(n1838), .ZN(n1485) );
  AOI22D1BWP12T U2460 ( .A1(register_file_inst1_r4_6_), .A2(n1595), .B1(
        register_file_inst1_r3_6_), .B2(n1839), .ZN(n1484) );
  AOI22D1BWP12T U2461 ( .A1(register_file_inst1_r6_6_), .A2(n1596), .B1(
        register_file_inst1_r10_6_), .B2(n1840), .ZN(n1483) );
  ND4D1BWP12T U2462 ( .A1(n1485), .A2(n1484), .A3(n2112), .A4(n1483), .ZN(
        n1486) );
  OAI22D1BWP12T U2463 ( .A1(n1502), .A2(n1850), .B1(n1490), .B2(n1848), .ZN(
        n1494) );
  OAI22D1BWP12T U2464 ( .A1(n1515), .A2(n1854), .B1(n1504), .B2(n1852), .ZN(
        n1493) );
  OAI22D1BWP12T U2465 ( .A1(n2196), .A2(n1858), .B1(n1505), .B2(n1856), .ZN(
        n1492) );
  OAI22D1BWP12T U2466 ( .A1(n1518), .A2(n1861), .B1(n1514), .B2(n1859), .ZN(
        n1491) );
  NR4D0BWP12T U2467 ( .A1(n1494), .A2(n1493), .A3(n1492), .A4(n1491), .ZN(
        n1500) );
  AOI22D1BWP12T U2468 ( .A1(register_file_inst1_tmp1_7_), .A2(n1835), .B1(
        register_file_inst1_r0_7_), .B2(n1633), .ZN(n1496) );
  AOI22D1BWP12T U2469 ( .A1(register_file_inst1_r5_7_), .A2(n1868), .B1(
        STACK_RF_next_sp[7]), .B2(n1867), .ZN(n1495) );
  AN3XD1BWP12T U2470 ( .A1(n1496), .A2(n1495), .A3(n2114), .Z(n1499) );
  AOI22D1BWP12T U2471 ( .A1(register_file_inst1_r1_7_), .A2(n1742), .B1(
        register_file_inst1_r11_7_), .B2(n1741), .ZN(n1498) );
  AOI22D1BWP12T U2472 ( .A1(register_file_inst1_r7_7_), .A2(n1744), .B1(
        register_file_inst1_r9_7_), .B2(n1743), .ZN(n1497) );
  ND4D1BWP12T U2473 ( .A1(n1500), .A2(n1499), .A3(n1498), .A4(n1497), .ZN(
        RF_ALU_operand_b[7]) );
  INVD1BWP12T U2474 ( .I(STACK_RF_next_sp[7]), .ZN(n1501) );
  OAI22D1BWP12T U2475 ( .A1(n1502), .A2(n1798), .B1(n1501), .B2(n1796), .ZN(
        n1511) );
  OAI22D1BWP12T U2476 ( .A1(n2196), .A2(n1802), .B1(n1503), .B2(n1800), .ZN(
        n1510) );
  OAI22D1BWP12T U2477 ( .A1(n1505), .A2(n1805), .B1(n1504), .B2(n1803), .ZN(
        n1509) );
  OAI22D1BWP12T U2478 ( .A1(n1507), .A2(n1809), .B1(n1506), .B2(n1807), .ZN(
        n1508) );
  NR4D0BWP12T U2479 ( .A1(n1511), .A2(n1510), .A3(n1509), .A4(n1508), .ZN(
        n1525) );
  CKND2D1BWP12T U2480 ( .A1(register_file_inst1_r9_7_), .A2(n1911), .ZN(n1513)
         );
  CKND2D1BWP12T U2481 ( .A1(register_file_inst1_r8_7_), .A2(n1910), .ZN(n1512)
         );
  ND3D1BWP12T U2482 ( .A1(n2197), .A2(n1513), .A3(n1512), .ZN(n1523) );
  OAI22D1BWP12T U2483 ( .A1(n1515), .A2(n1903), .B1(n1514), .B2(n1901), .ZN(
        n1522) );
  OAI22D1BWP12T U2484 ( .A1(n1517), .A2(n1907), .B1(n1516), .B2(n1905), .ZN(
        n1521) );
  OAI22D1BWP12T U2485 ( .A1(n1519), .A2(n1823), .B1(n1518), .B2(n1821), .ZN(
        n1520) );
  NR4D0BWP12T U2486 ( .A1(n1523), .A2(n1522), .A3(n1521), .A4(n1520), .ZN(
        n1524) );
  ND2D1BWP12T U2487 ( .A1(n1525), .A2(n1524), .ZN(RF_ALU_STACK_operand_a[7])
         );
  OAI22D1BWP12T U2488 ( .A1(n1527), .A2(n1798), .B1(n1526), .B2(n1796), .ZN(
        n1536) );
  OAI22D1BWP12T U2489 ( .A1(n2220), .A2(n1802), .B1(n1528), .B2(n1800), .ZN(
        n1535) );
  OAI22D1BWP12T U2490 ( .A1(n1530), .A2(n1805), .B1(n1529), .B2(n1803), .ZN(
        n1534) );
  OAI22D1BWP12T U2491 ( .A1(n1532), .A2(n1809), .B1(n1531), .B2(n1807), .ZN(
        n1533) );
  NR4D0BWP12T U2492 ( .A1(n1536), .A2(n1535), .A3(n1534), .A4(n1533), .ZN(
        n1550) );
  CKND2D1BWP12T U2493 ( .A1(register_file_inst1_r9_19_), .A2(n1911), .ZN(n1538) );
  ND2D1BWP12T U2494 ( .A1(register_file_inst1_r8_19_), .A2(n1910), .ZN(n1537)
         );
  ND3D1BWP12T U2495 ( .A1(n2221), .A2(n1538), .A3(n1537), .ZN(n1548) );
  OAI22D1BWP12T U2496 ( .A1(n1540), .A2(n1903), .B1(n1539), .B2(n1901), .ZN(
        n1547) );
  OAI22D1BWP12T U2497 ( .A1(n1542), .A2(n1907), .B1(n1541), .B2(n1905), .ZN(
        n1546) );
  OAI22D1BWP12T U2498 ( .A1(n1544), .A2(n1823), .B1(n1543), .B2(n1821), .ZN(
        n1545) );
  NR4D0BWP12T U2499 ( .A1(n1548), .A2(n1547), .A3(n1546), .A4(n1545), .ZN(
        n1549) );
  ND2D1BWP12T U2500 ( .A1(n1550), .A2(n1549), .ZN(RF_ALU_STACK_operand_a[19])
         );
  OAI22D1BWP12T U2501 ( .A1(n1552), .A2(n1903), .B1(n1551), .B2(n1901), .ZN(
        n1563) );
  OAI22D1BWP12T U2502 ( .A1(n1554), .A2(n1907), .B1(n1553), .B2(n1905), .ZN(
        n1562) );
  AOI22D1BWP12T U2503 ( .A1(register_file_inst1_tmp1_25_), .A2(n2244), .B1(
        register_file_inst1_r6_25_), .B2(n1909), .ZN(n1556) );
  AOI22D1BWP12T U2504 ( .A1(register_file_inst1_r8_25_), .A2(n1910), .B1(
        register_file_inst1_r9_25_), .B2(n1911), .ZN(n1555) );
  ND3D1BWP12T U2505 ( .A1(n1556), .A2(n1555), .A3(n2232), .ZN(n1561) );
  AOI22D1BWP12T U2506 ( .A1(register_file_inst1_r12_25_), .A2(n1915), .B1(
        STACK_RF_next_sp[25]), .B2(n1914), .ZN(n1559) );
  AOI22D1BWP12T U2507 ( .A1(register_file_inst1_lr_25_), .A2(n1917), .B1(
        register_file_inst1_r3_25_), .B2(n1916), .ZN(n1558) );
  AOI22D1BWP12T U2508 ( .A1(register_file_inst1_r1_25_), .A2(n1919), .B1(
        register_file_inst1_r7_25_), .B2(n1918), .ZN(n1557) );
  ND4D1BWP12T U2509 ( .A1(n1559), .A2(n2233), .A3(n1558), .A4(n1557), .ZN(
        n1560) );
  OR4XD1BWP12T U2510 ( .A1(n1563), .A2(n1562), .A3(n1561), .A4(n1560), .Z(
        RF_ALU_STACK_operand_a[25]) );
  OAI22D1BWP12T U2511 ( .A1(n1565), .A2(n1903), .B1(n1564), .B2(n1901), .ZN(
        n1576) );
  OAI22D1BWP12T U2512 ( .A1(n1567), .A2(n1907), .B1(n1566), .B2(n1905), .ZN(
        n1575) );
  AOI22D1BWP12T U2513 ( .A1(register_file_inst1_tmp1_27_), .A2(n2244), .B1(
        register_file_inst1_r6_27_), .B2(n1909), .ZN(n1569) );
  AOI22D1BWP12T U2514 ( .A1(register_file_inst1_r9_27_), .A2(n1911), .B1(
        register_file_inst1_r8_27_), .B2(n1910), .ZN(n1568) );
  ND3D1BWP12T U2515 ( .A1(n1569), .A2(n1568), .A3(n2236), .ZN(n1574) );
  AOI22D1BWP12T U2516 ( .A1(register_file_inst1_r12_27_), .A2(n1915), .B1(
        STACK_RF_next_sp[27]), .B2(n1914), .ZN(n1572) );
  AOI22D1BWP12T U2517 ( .A1(register_file_inst1_lr_27_), .A2(n1917), .B1(
        register_file_inst1_r3_27_), .B2(n1916), .ZN(n1571) );
  AOI22D1BWP12T U2518 ( .A1(register_file_inst1_r1_27_), .A2(n1919), .B1(
        register_file_inst1_r7_27_), .B2(n1918), .ZN(n1570) );
  ND4D1BWP12T U2519 ( .A1(n1572), .A2(n2237), .A3(n1571), .A4(n1570), .ZN(
        n1573) );
  OR4XD1BWP12T U2520 ( .A1(n1576), .A2(n1575), .A3(n1574), .A4(n1573), .Z(
        RF_ALU_STACK_operand_a[27]) );
  OAI22D1BWP12T U2521 ( .A1(n1578), .A2(n1903), .B1(n1577), .B2(n1901), .ZN(
        n1589) );
  OAI22D1BWP12T U2522 ( .A1(n1580), .A2(n1907), .B1(n1579), .B2(n1905), .ZN(
        n1588) );
  AOI22D1BWP12T U2523 ( .A1(register_file_inst1_tmp1_28_), .A2(n2244), .B1(
        register_file_inst1_r6_28_), .B2(n1909), .ZN(n1582) );
  AOI22D1BWP12T U2524 ( .A1(register_file_inst1_r8_28_), .A2(n1910), .B1(
        register_file_inst1_r9_28_), .B2(n1911), .ZN(n1581) );
  ND3D1BWP12T U2525 ( .A1(n1582), .A2(n1581), .A3(n2238), .ZN(n1587) );
  AOI22D1BWP12T U2526 ( .A1(register_file_inst1_r12_28_), .A2(n1915), .B1(
        STACK_RF_next_sp[28]), .B2(n1914), .ZN(n1585) );
  AOI22D1BWP12T U2527 ( .A1(register_file_inst1_lr_28_), .A2(n1917), .B1(
        register_file_inst1_r3_28_), .B2(n1916), .ZN(n1584) );
  AOI22D1BWP12T U2528 ( .A1(register_file_inst1_r1_28_), .A2(n1919), .B1(
        register_file_inst1_r7_28_), .B2(n1918), .ZN(n1583) );
  ND4D1BWP12T U2529 ( .A1(n1585), .A2(n2239), .A3(n1584), .A4(n1583), .ZN(
        n1586) );
  OR4XD1BWP12T U2530 ( .A1(n1589), .A2(n1588), .A3(n1587), .A4(n1586), .Z(
        RF_ALU_STACK_operand_a[28]) );
  OAI22D1BWP12T U2531 ( .A1(n1590), .A2(n1873), .B1(n1606), .B2(n1871), .ZN(
        n1603) );
  OAI22D1BWP12T U2532 ( .A1(n1592), .A2(n1877), .B1(n1591), .B2(n1875), .ZN(
        n1602) );
  AOI22D1BWP12T U2533 ( .A1(register_file_inst1_tmp1_29_), .A2(n1835), .B1(
        register_file_inst1_r0_29_), .B2(n1633), .ZN(n1594) );
  AOI22D1BWP12T U2534 ( .A1(register_file_inst1_r5_29_), .A2(n1868), .B1(
        STACK_RF_next_sp[29]), .B2(n1867), .ZN(n1593) );
  ND3D1BWP12T U2535 ( .A1(n1594), .A2(n1593), .A3(n2164), .ZN(n1601) );
  AOI22D1BWP12T U2536 ( .A1(register_file_inst1_r12_29_), .A2(n1659), .B1(
        register_file_inst1_r8_29_), .B2(n1838), .ZN(n1599) );
  AOI22D1BWP12T U2537 ( .A1(register_file_inst1_r4_29_), .A2(n1595), .B1(
        register_file_inst1_r3_29_), .B2(n1839), .ZN(n1598) );
  AOI22D1BWP12T U2538 ( .A1(register_file_inst1_r6_29_), .A2(n1596), .B1(
        register_file_inst1_r10_29_), .B2(n1840), .ZN(n1597) );
  ND4D1BWP12T U2539 ( .A1(n1599), .A2(n1598), .A3(n2165), .A4(n1597), .ZN(
        n1600) );
  OR4XD1BWP12T U2540 ( .A1(n1603), .A2(n1602), .A3(n1601), .A4(n1600), .Z(
        RF_ALU_operand_b[29]) );
  OAI22D1BWP12T U2541 ( .A1(n1605), .A2(n1903), .B1(n1604), .B2(n1901), .ZN(
        n1616) );
  OAI22D1BWP12T U2542 ( .A1(n1607), .A2(n1907), .B1(n1606), .B2(n1905), .ZN(
        n1615) );
  AOI22D1BWP12T U2543 ( .A1(register_file_inst1_tmp1_29_), .A2(n2244), .B1(
        register_file_inst1_r6_29_), .B2(n1909), .ZN(n1609) );
  AOI22D1BWP12T U2544 ( .A1(register_file_inst1_r9_29_), .A2(n1911), .B1(
        register_file_inst1_r8_29_), .B2(n1910), .ZN(n1608) );
  ND3D1BWP12T U2545 ( .A1(n1609), .A2(n1608), .A3(n2240), .ZN(n1614) );
  AOI22D1BWP12T U2546 ( .A1(register_file_inst1_r12_29_), .A2(n1915), .B1(
        STACK_RF_next_sp[29]), .B2(n1914), .ZN(n1612) );
  AOI22D1BWP12T U2547 ( .A1(register_file_inst1_lr_29_), .A2(n1917), .B1(
        register_file_inst1_r3_29_), .B2(n1916), .ZN(n1611) );
  AOI22D1BWP12T U2548 ( .A1(register_file_inst1_r1_29_), .A2(n1919), .B1(
        register_file_inst1_r7_29_), .B2(n1918), .ZN(n1610) );
  ND4D1BWP12T U2549 ( .A1(n1612), .A2(n2241), .A3(n1611), .A4(n1610), .ZN(
        n1613) );
  OR4XD1BWP12T U2550 ( .A1(n1616), .A2(n1615), .A3(n1614), .A4(n1613), .Z(
        RF_ALU_STACK_operand_a[29]) );
  OAI22D1BWP12T U2551 ( .A1(n1618), .A2(n1873), .B1(n1617), .B2(n1871), .ZN(
        n1629) );
  OAI22D1BWP12T U2552 ( .A1(n1620), .A2(n1877), .B1(n1619), .B2(n1875), .ZN(
        n1628) );
  AOI22D1BWP12T U2553 ( .A1(register_file_inst1_tmp1_30_), .A2(n1835), .B1(
        register_file_inst1_r0_30_), .B2(n1633), .ZN(n1622) );
  AOI22D1BWP12T U2554 ( .A1(register_file_inst1_r5_30_), .A2(n1868), .B1(
        STACK_RF_next_sp[30]), .B2(n1867), .ZN(n1621) );
  ND3D1BWP12T U2555 ( .A1(n1622), .A2(n1621), .A3(n2166), .ZN(n1627) );
  AOI22D1BWP12T U2556 ( .A1(register_file_inst1_r12_30_), .A2(n1659), .B1(
        register_file_inst1_r8_30_), .B2(n1838), .ZN(n1625) );
  AOI22D1BWP12T U2557 ( .A1(register_file_inst1_r4_30_), .A2(n1595), .B1(
        register_file_inst1_r3_30_), .B2(n1839), .ZN(n1624) );
  AOI22D1BWP12T U2558 ( .A1(register_file_inst1_r6_30_), .A2(n1596), .B1(
        register_file_inst1_r10_30_), .B2(n1840), .ZN(n1623) );
  ND4D1BWP12T U2559 ( .A1(n1625), .A2(n1624), .A3(n2167), .A4(n1623), .ZN(
        n1626) );
  OR4XD1BWP12T U2560 ( .A1(n1629), .A2(n1628), .A3(n1627), .A4(n1626), .Z(
        RF_ALU_operand_b[30]) );
  OAI22D1BWP12T U2561 ( .A1(n1630), .A2(n1873), .B1(n1645), .B2(n1871), .ZN(
        n1642) );
  OAI22D1BWP12T U2562 ( .A1(n1632), .A2(n1877), .B1(n1631), .B2(n1875), .ZN(
        n1641) );
  AOI22D1BWP12T U2563 ( .A1(register_file_inst1_tmp1_31_), .A2(n1835), .B1(
        register_file_inst1_r0_31_), .B2(n1633), .ZN(n1635) );
  AOI22D1BWP12T U2564 ( .A1(register_file_inst1_r5_31_), .A2(n1868), .B1(
        STACK_RF_next_sp[31]), .B2(n1867), .ZN(n1634) );
  ND3D1BWP12T U2565 ( .A1(n1635), .A2(n1634), .A3(n2169), .ZN(n1640) );
  AOI22D1BWP12T U2566 ( .A1(register_file_inst1_r12_31_), .A2(n1659), .B1(
        register_file_inst1_r8_31_), .B2(n1838), .ZN(n1638) );
  AOI22D1BWP12T U2567 ( .A1(register_file_inst1_r4_31_), .A2(n1595), .B1(
        register_file_inst1_r3_31_), .B2(n1839), .ZN(n1637) );
  AOI22D1BWP12T U2568 ( .A1(register_file_inst1_r6_31_), .A2(n1596), .B1(
        register_file_inst1_r10_31_), .B2(n1840), .ZN(n1636) );
  ND4D1BWP12T U2569 ( .A1(n1638), .A2(n1637), .A3(n2170), .A4(n1636), .ZN(
        n1639) );
  OR4XD1BWP12T U2570 ( .A1(n1642), .A2(n1641), .A3(n1640), .A4(n1639), .Z(
        RF_ALU_operand_b[31]) );
  OAI22D1BWP12T U2571 ( .A1(n1644), .A2(n1903), .B1(n1643), .B2(n1901), .ZN(
        n1655) );
  OAI22D1BWP12T U2572 ( .A1(n1646), .A2(n1907), .B1(n1645), .B2(n1905), .ZN(
        n1654) );
  AOI22D1BWP12T U2573 ( .A1(register_file_inst1_tmp1_31_), .A2(n2244), .B1(
        register_file_inst1_r6_31_), .B2(n1909), .ZN(n1648) );
  AOI22D1BWP12T U2574 ( .A1(register_file_inst1_r8_31_), .A2(n1910), .B1(
        register_file_inst1_r9_31_), .B2(n1911), .ZN(n1647) );
  ND3D1BWP12T U2575 ( .A1(n1648), .A2(n1647), .A3(n2245), .ZN(n1653) );
  AOI22D1BWP12T U2576 ( .A1(register_file_inst1_r12_31_), .A2(n1915), .B1(
        STACK_RF_next_sp[31]), .B2(n1914), .ZN(n1651) );
  AOI22D1BWP12T U2577 ( .A1(register_file_inst1_lr_31_), .A2(n1917), .B1(
        register_file_inst1_r3_31_), .B2(n1916), .ZN(n1650) );
  AOI22D1BWP12T U2578 ( .A1(register_file_inst1_r1_31_), .A2(n1919), .B1(
        register_file_inst1_r7_31_), .B2(n1918), .ZN(n1649) );
  ND4D1BWP12T U2579 ( .A1(n1651), .A2(n2246), .A3(n1650), .A4(n1649), .ZN(
        n1652) );
  OR4XD1BWP12T U2580 ( .A1(n1655), .A2(n1654), .A3(n1653), .A4(n1652), .Z(
        RF_ALU_STACK_operand_a[31]) );
  OAI22D1BWP12T U2581 ( .A1(n1704), .A2(n1873), .B1(n1713), .B2(n1871), .ZN(
        n1666) );
  OAI22D1BWP12T U2582 ( .A1(n1703), .A2(n1877), .B1(n1656), .B2(n1875), .ZN(
        n1665) );
  AOI22D1BWP12T U2583 ( .A1(register_file_inst1_tmp1_5_), .A2(n1835), .B1(
        register_file_inst1_r0_5_), .B2(n1633), .ZN(n1658) );
  AOI22D1BWP12T U2584 ( .A1(register_file_inst1_r5_5_), .A2(n1868), .B1(
        STACK_RF_next_sp[5]), .B2(n1867), .ZN(n1657) );
  ND3D1BWP12T U2585 ( .A1(n1658), .A2(n1657), .A3(n2108), .ZN(n1664) );
  AOI22D1BWP12T U2586 ( .A1(register_file_inst1_r12_5_), .A2(n1659), .B1(
        register_file_inst1_r8_5_), .B2(n1838), .ZN(n1662) );
  AOI22D1BWP12T U2587 ( .A1(register_file_inst1_r4_5_), .A2(n1595), .B1(
        register_file_inst1_r3_5_), .B2(n1839), .ZN(n1661) );
  AOI22D1BWP12T U2588 ( .A1(register_file_inst1_r6_5_), .A2(n1596), .B1(
        register_file_inst1_r10_5_), .B2(n1840), .ZN(n1660) );
  ND4D1BWP12T U2589 ( .A1(n1662), .A2(n1661), .A3(n2109), .A4(n1660), .ZN(
        n1663) );
  OR4XD1BWP12T U2590 ( .A1(n1666), .A2(n1665), .A3(n1664), .A4(n1663), .Z(
        RF_ALU_operand_b[5]) );
  OAI22D1BWP12T U2591 ( .A1(n1668), .A2(n1850), .B1(n1667), .B2(n1848), .ZN(
        n1677) );
  OAI22D1BWP12T U2592 ( .A1(n1670), .A2(n1854), .B1(n1669), .B2(n1852), .ZN(
        n1676) );
  OAI22D1BWP12T U2593 ( .A1(n2190), .A2(n1858), .B1(n1671), .B2(n1856), .ZN(
        n1675) );
  OAI22D1BWP12T U2594 ( .A1(n1673), .A2(n1861), .B1(n1672), .B2(n1859), .ZN(
        n1674) );
  AOI22D1BWP12T U2595 ( .A1(register_file_inst1_tmp1_4_), .A2(n1835), .B1(
        register_file_inst1_r0_4_), .B2(n1633), .ZN(n1679) );
  AOI22D1BWP12T U2596 ( .A1(register_file_inst1_r5_4_), .A2(n1868), .B1(
        STACK_RF_next_sp[4]), .B2(n1867), .ZN(n1678) );
  AN3XD1BWP12T U2597 ( .A1(n1679), .A2(n1678), .A3(n2106), .Z(n1682) );
  AOI22D1BWP12T U2598 ( .A1(register_file_inst1_r1_4_), .A2(n1742), .B1(
        register_file_inst1_r11_4_), .B2(n1741), .ZN(n1681) );
  AOI22D1BWP12T U2599 ( .A1(register_file_inst1_r7_4_), .A2(n1744), .B1(
        register_file_inst1_r9_4_), .B2(n1743), .ZN(n1680) );
  ND4D1BWP12T U2600 ( .A1(n1683), .A2(n1682), .A3(n1681), .A4(n1680), .ZN(
        RF_ALU_operand_b[4]) );
  OAI22D1BWP12T U2601 ( .A1(n1851), .A2(n1798), .B1(n1684), .B2(n1796), .ZN(
        n1688) );
  OAI22D1BWP12T U2602 ( .A1(n2172), .A2(n1802), .B1(n1880), .B2(n1800), .ZN(
        n1687) );
  OAI22D1BWP12T U2603 ( .A1(n1857), .A2(n1805), .B1(n1853), .B2(n1803), .ZN(
        n1686) );
  OAI22D1BWP12T U2604 ( .A1(n1874), .A2(n1809), .B1(n1878), .B2(n1807), .ZN(
        n1685) );
  NR4D0BWP12T U2605 ( .A1(n1688), .A2(n1687), .A3(n1686), .A4(n1685), .ZN(
        n1697) );
  CKND2D1BWP12T U2606 ( .A1(register_file_inst1_r9_0_), .A2(n1911), .ZN(n1690)
         );
  CKND2D1BWP12T U2607 ( .A1(register_file_inst1_r8_0_), .A2(n1910), .ZN(n1689)
         );
  ND3D1BWP12T U2608 ( .A1(n2177), .A2(n1690), .A3(n1689), .ZN(n1695) );
  OAI22D1BWP12T U2609 ( .A1(n1855), .A2(n1903), .B1(n1860), .B2(n1901), .ZN(
        n1694) );
  OAI22D1BWP12T U2610 ( .A1(n1691), .A2(n1907), .B1(n1872), .B2(n1905), .ZN(
        n1693) );
  OAI22D1BWP12T U2611 ( .A1(n1881), .A2(n1823), .B1(n1862), .B2(n1821), .ZN(
        n1692) );
  NR4D0BWP12T U2612 ( .A1(n1695), .A2(n1694), .A3(n1693), .A4(n1692), .ZN(
        n1696) );
  ND2D1BWP12T U2613 ( .A1(n1697), .A2(n1696), .ZN(RF_ALU_STACK_operand_a[0])
         );
  INVD1BWP12T U2614 ( .I(STACK_RF_next_sp[5]), .ZN(n1698) );
  OAI22D1BWP12T U2615 ( .A1(n1699), .A2(n1798), .B1(n1698), .B2(n1796), .ZN(
        n1708) );
  OAI22D1BWP12T U2616 ( .A1(n2192), .A2(n1802), .B1(n1700), .B2(n1800), .ZN(
        n1707) );
  OAI22D1BWP12T U2617 ( .A1(n1702), .A2(n1805), .B1(n1701), .B2(n1803), .ZN(
        n1706) );
  OAI22D1BWP12T U2618 ( .A1(n1704), .A2(n1809), .B1(n1703), .B2(n1807), .ZN(
        n1705) );
  NR4D0BWP12T U2619 ( .A1(n1708), .A2(n1707), .A3(n1706), .A4(n1705), .ZN(
        n1722) );
  CKND2D1BWP12T U2620 ( .A1(register_file_inst1_r9_5_), .A2(n1911), .ZN(n1710)
         );
  ND2D1BWP12T U2621 ( .A1(register_file_inst1_r8_5_), .A2(n1910), .ZN(n1709)
         );
  ND3D1BWP12T U2622 ( .A1(n2193), .A2(n1710), .A3(n1709), .ZN(n1720) );
  OAI22D1BWP12T U2623 ( .A1(n1712), .A2(n1903), .B1(n1711), .B2(n1901), .ZN(
        n1719) );
  OAI22D1BWP12T U2624 ( .A1(n1714), .A2(n1907), .B1(n1713), .B2(n1905), .ZN(
        n1718) );
  OAI22D1BWP12T U2625 ( .A1(n1716), .A2(n1823), .B1(n1715), .B2(n1821), .ZN(
        n1717) );
  NR4D0BWP12T U2626 ( .A1(n1720), .A2(n1719), .A3(n1718), .A4(n1717), .ZN(
        n1721) );
  ND2D1BWP12T U2627 ( .A1(n1722), .A2(n1721), .ZN(RF_ALU_STACK_operand_a[5])
         );
  OAI22D1BWP12T U2628 ( .A1(n1750), .A2(n1850), .B1(n1723), .B2(n1848), .ZN(
        n1727) );
  OAI22D1BWP12T U2629 ( .A1(n1763), .A2(n1854), .B1(n1752), .B2(n1852), .ZN(
        n1726) );
  OAI22D1BWP12T U2630 ( .A1(n2188), .A2(n1858), .B1(n1753), .B2(n1856), .ZN(
        n1725) );
  OAI22D1BWP12T U2631 ( .A1(n1766), .A2(n1861), .B1(n1762), .B2(n1859), .ZN(
        n1724) );
  NR4D0BWP12T U2632 ( .A1(n1727), .A2(n1726), .A3(n1725), .A4(n1724), .ZN(
        n1733) );
  AOI22D1BWP12T U2633 ( .A1(register_file_inst1_tmp1_3_), .A2(n1835), .B1(
        register_file_inst1_r0_3_), .B2(n1633), .ZN(n1729) );
  AOI22D1BWP12T U2634 ( .A1(register_file_inst1_r5_3_), .A2(n1868), .B1(
        STACK_RF_next_sp[3]), .B2(n1867), .ZN(n1728) );
  AN3XD1BWP12T U2635 ( .A1(n1729), .A2(n1728), .A3(n2104), .Z(n1732) );
  AOI22D1BWP12T U2636 ( .A1(register_file_inst1_r1_3_), .A2(n1742), .B1(
        register_file_inst1_r11_3_), .B2(n1741), .ZN(n1731) );
  AOI22D1BWP12T U2637 ( .A1(register_file_inst1_r7_3_), .A2(n1744), .B1(
        register_file_inst1_r9_3_), .B2(n1743), .ZN(n1730) );
  ND4D1BWP12T U2638 ( .A1(n1733), .A2(n1732), .A3(n1731), .A4(n1730), .ZN(
        RF_ALU_operand_b[3]) );
  OAI22D1BWP12T U2639 ( .A1(n1799), .A2(n1850), .B1(n1734), .B2(n1848), .ZN(
        n1738) );
  OAI22D1BWP12T U2640 ( .A1(n1818), .A2(n1854), .B1(n1804), .B2(n1852), .ZN(
        n1737) );
  OAI22D1BWP12T U2641 ( .A1(n2186), .A2(n1858), .B1(n1806), .B2(n1856), .ZN(
        n1736) );
  NR4D0BWP12T U2642 ( .A1(n1738), .A2(n1737), .A3(n1736), .A4(n1735), .ZN(
        n1748) );
  AOI22D1BWP12T U2643 ( .A1(register_file_inst1_tmp1_2_), .A2(n1835), .B1(
        register_file_inst1_r0_2_), .B2(n1633), .ZN(n1740) );
  AOI22D1BWP12T U2644 ( .A1(register_file_inst1_r5_2_), .A2(n1868), .B1(
        STACK_RF_next_sp[2]), .B2(n1867), .ZN(n1739) );
  AN3XD1BWP12T U2645 ( .A1(n1740), .A2(n1739), .A3(n2102), .Z(n1747) );
  AOI22D1BWP12T U2646 ( .A1(register_file_inst1_r1_2_), .A2(n1742), .B1(
        register_file_inst1_r11_2_), .B2(n1741), .ZN(n1746) );
  AOI22D1BWP12T U2647 ( .A1(register_file_inst1_r7_2_), .A2(n1744), .B1(
        register_file_inst1_r9_2_), .B2(n1743), .ZN(n1745) );
  ND4D1BWP12T U2648 ( .A1(n1748), .A2(n1747), .A3(n1746), .A4(n1745), .ZN(
        RF_ALU_operand_b[2]) );
  INVD1BWP12T U2649 ( .I(STACK_RF_next_sp[3]), .ZN(n1749) );
  OAI22D1BWP12T U2650 ( .A1(n1750), .A2(n1798), .B1(n1749), .B2(n1796), .ZN(
        n1759) );
  OAI22D1BWP12T U2651 ( .A1(n2188), .A2(n1802), .B1(n1751), .B2(n1800), .ZN(
        n1758) );
  OAI22D1BWP12T U2652 ( .A1(n1753), .A2(n1805), .B1(n1752), .B2(n1803), .ZN(
        n1757) );
  OAI22D1BWP12T U2653 ( .A1(n1755), .A2(n1809), .B1(n1754), .B2(n1807), .ZN(
        n1756) );
  NR4D0BWP12T U2654 ( .A1(n1759), .A2(n1758), .A3(n1757), .A4(n1756), .ZN(
        n1773) );
  CKND2D1BWP12T U2655 ( .A1(register_file_inst1_r9_3_), .A2(n1911), .ZN(n1761)
         );
  CKND2D1BWP12T U2656 ( .A1(register_file_inst1_r8_3_), .A2(n1910), .ZN(n1760)
         );
  ND3D1BWP12T U2657 ( .A1(n2189), .A2(n1761), .A3(n1760), .ZN(n1771) );
  OAI22D1BWP12T U2658 ( .A1(n1763), .A2(n1903), .B1(n1762), .B2(n1901), .ZN(
        n1770) );
  OAI22D1BWP12T U2659 ( .A1(n1765), .A2(n1907), .B1(n1764), .B2(n1905), .ZN(
        n1769) );
  OAI22D1BWP12T U2660 ( .A1(n1767), .A2(n1823), .B1(n1766), .B2(n1821), .ZN(
        n1768) );
  NR4D0BWP12T U2661 ( .A1(n1771), .A2(n1770), .A3(n1769), .A4(n1768), .ZN(
        n1772) );
  ND2D1BWP12T U2662 ( .A1(n1773), .A2(n1772), .ZN(RF_ALU_STACK_operand_a[3])
         );
  INVD1BWP12T U2663 ( .I(STACK_RF_next_sp[1]), .ZN(n1774) );
  OAI22D1BWP12T U2664 ( .A1(n1775), .A2(n1798), .B1(n1774), .B2(n1796), .ZN(
        n1782) );
  OAI22D1BWP12T U2665 ( .A1(n2184), .A2(n1802), .B1(n1776), .B2(n1800), .ZN(
        n1781) );
  OAI22D1BWP12T U2666 ( .A1(n1778), .A2(n1805), .B1(n1777), .B2(n1803), .ZN(
        n1780) );
  OAI22D1BWP12T U2667 ( .A1(n1832), .A2(n1809), .B1(n1834), .B2(n1807), .ZN(
        n1779) );
  NR4D0BWP12T U2668 ( .A1(n1782), .A2(n1781), .A3(n1780), .A4(n1779), .ZN(
        n1795) );
  CKND2D1BWP12T U2669 ( .A1(register_file_inst1_r9_1_), .A2(n1911), .ZN(n1784)
         );
  CKND2D1BWP12T U2670 ( .A1(register_file_inst1_r8_1_), .A2(n1910), .ZN(n1783)
         );
  ND3D1BWP12T U2671 ( .A1(n2185), .A2(n1784), .A3(n1783), .ZN(n1793) );
  OAI22D1BWP12T U2672 ( .A1(n1786), .A2(n1903), .B1(n1785), .B2(n1901), .ZN(
        n1792) );
  OAI22D1BWP12T U2673 ( .A1(n1787), .A2(n1907), .B1(n1831), .B2(n1905), .ZN(
        n1791) );
  OAI22D1BWP12T U2674 ( .A1(n1789), .A2(n1823), .B1(n1788), .B2(n1821), .ZN(
        n1790) );
  NR4D0BWP12T U2675 ( .A1(n1793), .A2(n1792), .A3(n1791), .A4(n1790), .ZN(
        n1794) );
  ND2D1BWP12T U2676 ( .A1(n1795), .A2(n1794), .ZN(RF_ALU_STACK_operand_a[1])
         );
  INVD1BWP12T U2677 ( .I(STACK_RF_next_sp[2]), .ZN(n1797) );
  OAI22D1BWP12T U2678 ( .A1(n1799), .A2(n1798), .B1(n1797), .B2(n1796), .ZN(
        n1814) );
  OAI22D1BWP12T U2679 ( .A1(n2186), .A2(n1802), .B1(n1801), .B2(n1800), .ZN(
        n1813) );
  OAI22D1BWP12T U2680 ( .A1(n1806), .A2(n1805), .B1(n1804), .B2(n1803), .ZN(
        n1812) );
  OAI22D1BWP12T U2681 ( .A1(n1810), .A2(n1809), .B1(n1808), .B2(n1807), .ZN(
        n1811) );
  NR4D0BWP12T U2682 ( .A1(n1814), .A2(n1813), .A3(n1812), .A4(n1811), .ZN(
        n1830) );
  CKND2D1BWP12T U2683 ( .A1(register_file_inst1_r9_2_), .A2(n1911), .ZN(n1816)
         );
  CKND2D1BWP12T U2684 ( .A1(register_file_inst1_r8_2_), .A2(n1910), .ZN(n1815)
         );
  ND3D1BWP12T U2685 ( .A1(n2187), .A2(n1816), .A3(n1815), .ZN(n1828) );
  OAI22D1BWP12T U2686 ( .A1(n1818), .A2(n1903), .B1(n1817), .B2(n1901), .ZN(
        n1827) );
  OAI22D1BWP12T U2687 ( .A1(n1820), .A2(n1907), .B1(n1819), .B2(n1905), .ZN(
        n1826) );
  OAI22D1BWP12T U2688 ( .A1(n1824), .A2(n1823), .B1(n1822), .B2(n1821), .ZN(
        n1825) );
  NR4D0BWP12T U2689 ( .A1(n1828), .A2(n1827), .A3(n1826), .A4(n1825), .ZN(
        n1829) );
  ND2D1BWP12T U2690 ( .A1(n1830), .A2(n1829), .ZN(RF_ALU_STACK_operand_a[2])
         );
  OAI22D1BWP12T U2691 ( .A1(n1832), .A2(n1873), .B1(n1831), .B2(n1871), .ZN(
        n1847) );
  OAI22D1BWP12T U2692 ( .A1(n1834), .A2(n1877), .B1(n1833), .B2(n1875), .ZN(
        n1846) );
  AOI22D1BWP12T U2693 ( .A1(register_file_inst1_tmp1_1_), .A2(n1835), .B1(
        register_file_inst1_r0_1_), .B2(n1633), .ZN(n1837) );
  AOI22D1BWP12T U2694 ( .A1(register_file_inst1_r5_1_), .A2(n1868), .B1(
        STACK_RF_next_sp[1]), .B2(n1867), .ZN(n1836) );
  ND3D1BWP12T U2695 ( .A1(n1837), .A2(n1836), .A3(n2099), .ZN(n1845) );
  AOI22D1BWP12T U2696 ( .A1(register_file_inst1_r12_1_), .A2(n1659), .B1(
        register_file_inst1_r8_1_), .B2(n1838), .ZN(n1843) );
  AOI22D1BWP12T U2697 ( .A1(register_file_inst1_r4_1_), .A2(n1595), .B1(
        register_file_inst1_r3_1_), .B2(n1839), .ZN(n1842) );
  AOI22D1BWP12T U2698 ( .A1(register_file_inst1_r6_1_), .A2(n1596), .B1(
        register_file_inst1_r10_1_), .B2(n1840), .ZN(n1841) );
  ND4D1BWP12T U2699 ( .A1(n1843), .A2(n1842), .A3(n2100), .A4(n1841), .ZN(
        n1844) );
  OR4XD1BWP12T U2700 ( .A1(n1847), .A2(n1846), .A3(n1845), .A4(n1844), .Z(
        RF_ALU_operand_b[1]) );
  OAI22D1BWP12T U2701 ( .A1(n1851), .A2(n1850), .B1(n1849), .B2(n1848), .ZN(
        n1866) );
  OAI22D1BWP12T U2702 ( .A1(n1855), .A2(n1854), .B1(n1853), .B2(n1852), .ZN(
        n1865) );
  OAI22D1BWP12T U2703 ( .A1(n2172), .A2(n1858), .B1(n1857), .B2(n1856), .ZN(
        n1864) );
  OAI22D1BWP12T U2704 ( .A1(n1862), .A2(n1861), .B1(n1860), .B2(n1859), .ZN(
        n1863) );
  NR4D0BWP12T U2705 ( .A1(n1866), .A2(n1865), .A3(n1864), .A4(n1863), .ZN(
        n1887) );
  ND2D1BWP12T U2706 ( .A1(STACK_RF_next_sp[0]), .A2(n1867), .ZN(n1870) );
  CKND2D1BWP12T U2707 ( .A1(register_file_inst1_r5_0_), .A2(n1868), .ZN(n1869)
         );
  ND3D1BWP12T U2708 ( .A1(n2091), .A2(n1870), .A3(n1869), .ZN(n1885) );
  OAI22D1BWP12T U2709 ( .A1(n1874), .A2(n1873), .B1(n1872), .B2(n1871), .ZN(
        n1884) );
  OAI22D1BWP12T U2710 ( .A1(n1878), .A2(n1877), .B1(n1876), .B2(n1875), .ZN(
        n1883) );
  OAI22D1BWP12T U2711 ( .A1(n1881), .A2(n1928), .B1(n1880), .B2(n1879), .ZN(
        n1882) );
  NR4D0BWP12T U2712 ( .A1(n1885), .A2(n1884), .A3(n1883), .A4(n1882), .ZN(
        n1886) );
  ND2D1BWP12T U2713 ( .A1(n1887), .A2(n1886), .ZN(RF_ALU_operand_b[0]) );
  OAI22D1BWP12T U2714 ( .A1(n1889), .A2(n1903), .B1(n1888), .B2(n1901), .ZN(
        n1900) );
  OAI22D1BWP12T U2715 ( .A1(n1891), .A2(n1907), .B1(n1890), .B2(n1905), .ZN(
        n1899) );
  AOI22D1BWP12T U2716 ( .A1(register_file_inst1_tmp1_23_), .A2(n2244), .B1(
        register_file_inst1_r6_23_), .B2(n1909), .ZN(n1893) );
  AOI22D1BWP12T U2717 ( .A1(register_file_inst1_r8_23_), .A2(n1910), .B1(
        register_file_inst1_r9_23_), .B2(n1911), .ZN(n1892) );
  ND3D1BWP12T U2718 ( .A1(n1893), .A2(n1892), .A3(n2228), .ZN(n1898) );
  AOI22D1BWP12T U2719 ( .A1(register_file_inst1_r12_23_), .A2(n1915), .B1(
        STACK_RF_next_sp[23]), .B2(n1914), .ZN(n1896) );
  AOI22D1BWP12T U2720 ( .A1(register_file_inst1_lr_23_), .A2(n1917), .B1(
        register_file_inst1_r3_23_), .B2(n1916), .ZN(n1895) );
  AOI22D1BWP12T U2721 ( .A1(register_file_inst1_r1_23_), .A2(n1919), .B1(
        register_file_inst1_r7_23_), .B2(n1918), .ZN(n1894) );
  ND4D1BWP12T U2722 ( .A1(n1896), .A2(n2229), .A3(n1895), .A4(n1894), .ZN(
        n1897) );
  OR4XD1BWP12T U2723 ( .A1(n1900), .A2(n1899), .A3(n1898), .A4(n1897), .Z(
        RF_ALU_STACK_operand_a[23]) );
  OAI22D1BWP12T U2724 ( .A1(n1904), .A2(n1903), .B1(n1902), .B2(n1901), .ZN(
        n1926) );
  OAI22D1BWP12T U2725 ( .A1(n1908), .A2(n1907), .B1(n1906), .B2(n1905), .ZN(
        n1925) );
  AOI22D1BWP12T U2726 ( .A1(register_file_inst1_tmp1_21_), .A2(n2244), .B1(
        register_file_inst1_r6_21_), .B2(n1909), .ZN(n1913) );
  AOI22D1BWP12T U2727 ( .A1(register_file_inst1_r9_21_), .A2(n1911), .B1(
        register_file_inst1_r8_21_), .B2(n1910), .ZN(n1912) );
  ND3D1BWP12T U2728 ( .A1(n1913), .A2(n1912), .A3(n2224), .ZN(n1924) );
  AOI22D1BWP12T U2729 ( .A1(register_file_inst1_r12_21_), .A2(n1915), .B1(
        STACK_RF_next_sp[21]), .B2(n1914), .ZN(n1922) );
  AOI22D1BWP12T U2730 ( .A1(register_file_inst1_lr_21_), .A2(n1917), .B1(
        register_file_inst1_r3_21_), .B2(n1916), .ZN(n1921) );
  AOI22D1BWP12T U2731 ( .A1(register_file_inst1_r1_21_), .A2(n1919), .B1(
        register_file_inst1_r7_21_), .B2(n1918), .ZN(n1920) );
  ND4D1BWP12T U2732 ( .A1(n1922), .A2(n2225), .A3(n1921), .A4(n1920), .ZN(
        n1923) );
  OR4XD1BWP12T U2733 ( .A1(n1926), .A2(n1925), .A3(n1924), .A4(n1923), .Z(
        RF_ALU_STACK_operand_a[21]) );
  RCAOI211D0BWP12T U2734 ( .A1(n2035), .A2(STACK_RF_next_sp[8]), .B(n2019), 
        .C(reset), .ZN(n2020) );
  RCAOI211D0BWP12T U2735 ( .A1(n2035), .A2(STACK_RF_next_sp[11]), .B(n2010), 
        .C(reset), .ZN(n2011) );
  RCAOI211D0BWP12T U2736 ( .A1(n2035), .A2(STACK_RF_next_sp[12]), .B(n2007), 
        .C(reset), .ZN(n2008) );
  RCAOI211D0BWP12T U2737 ( .A1(n2035), .A2(STACK_RF_next_sp[7]), .B(n2022), 
        .C(reset), .ZN(n2023) );
  AOI21D0BWP12T U2738 ( .A1(n2286), .A2(IF_RF_incremented_pc_out[1]), .B(reset), .ZN(n2283) );
  AOI22D0BWP12T U2739 ( .A1(RF_pc_out[10]), .A2(n1932), .B1(
        STACK_RF_next_sp[10]), .B2(n1927), .ZN(n2015) );
  INVD1BWP12T U2740 ( .I(RF_pc_out[1]), .ZN(n2184) );
  INVD1BWP12T U2741 ( .I(RF_pc_out[4]), .ZN(n2190) );
  MUX2D1BWP12T U2742 ( .I0(MEMCTRL_RF_IF_data_in[15]), .I1(
        ALU_MISC_OUT_result[15]), .S(n2277), .Z(
        register_file_inst1_pc_write_in_15_) );
  MUX2D1BWP12T U2743 ( .I0(MEMCTRL_RF_IF_data_in[11]), .I1(
        ALU_MISC_OUT_result[11]), .S(n2277), .Z(
        register_file_inst1_pc_write_in_11_) );
  MUX2D1BWP12T U2744 ( .I0(MEMCTRL_RF_IF_data_in[13]), .I1(
        ALU_MISC_OUT_result[13]), .S(n2277), .Z(
        register_file_inst1_pc_write_in_13_) );
  MUX2D1BWP12T U2745 ( .I0(MEMCTRL_RF_IF_data_in[7]), .I1(
        ALU_MISC_OUT_result[7]), .S(n2277), .Z(
        register_file_inst1_pc_write_in_7_) );
  MUX2D1BWP12T U2746 ( .I0(MEMCTRL_RF_IF_data_in[5]), .I1(
        ALU_MISC_OUT_result[5]), .S(n2277), .Z(
        register_file_inst1_pc_write_in_5_) );
  MUX2ND1BWP12T U2747 ( .I0(MEMCTRL_RF_IF_data_in[9]), .I1(
        ALU_MISC_OUT_result[9]), .S(n2277), .ZN(n1931) );
  MUX2D1BWP12T U2748 ( .I0(MEMCTRL_RF_IF_data_in[3]), .I1(
        ALU_MISC_OUT_result[3]), .S(n2277), .Z(
        register_file_inst1_pc_write_in_3_) );
  MUX2XD0BWP12T U2749 ( .I0(MEMCTRL_RF_IF_data_in[0]), .I1(
        ALU_MISC_OUT_result[0]), .S(n2277), .Z(
        register_file_inst1_pc_write_in_0_) );
  MUX2D1BWP12T U2750 ( .I0(MEMCTRL_RF_IF_data_in[1]), .I1(
        ALU_MISC_OUT_result[1]), .S(n2277), .Z(
        register_file_inst1_pc_write_in_1_) );
  RCAOI211D0BWP12T U2751 ( .A1(n2035), .A2(STACK_RF_next_sp[9]), .B(n2016), 
        .C(reset), .ZN(n2017) );
  RCAOI211D0BWP12T U2752 ( .A1(n2035), .A2(STACK_RF_next_sp[4]), .B(n2028), 
        .C(reset), .ZN(n2029) );
  RCAOI211D0BWP12T U2753 ( .A1(n2035), .A2(STACK_RF_next_sp[2]), .B(n1990), 
        .C(reset), .ZN(n1991) );
  TPNR2D1BWP12T U2754 ( .A1(reset), .A2(n2284), .ZN(n2287) );
  AOI22D0BWP12T U2755 ( .A1(RF_pc_out[12]), .A2(n1932), .B1(
        STACK_RF_next_sp[12]), .B2(n1927), .ZN(n2009) );
  OR2D1BWP12T U2756 ( .A1(DEC_RF_operand_b[0]), .A2(n2096), .Z(n1928) );
  NR2D1BWP12T U2757 ( .A1(reset), .A2(n1973), .ZN(n1976) );
  INVD1BWP12T U2758 ( .I(RF_pc_out[8]), .ZN(n2198) );
  INVD1BWP12T U2759 ( .I(RF_pc_out[3]), .ZN(n2188) );
  INVD1BWP12T U2760 ( .I(RF_pc_out[7]), .ZN(n2196) );
  INVD1BWP12T U2761 ( .I(RF_pc_out[2]), .ZN(n2186) );
  ND2D1BWP12T U2762 ( .A1(DEC_RF_alu_stack_write_to_reg[1]), .A2(n1964), .ZN(
        n1973) );
  AO222D1BWP12T U2763 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[29]), .B1(n2286), .B2(
        IF_RF_incremented_pc_out[29]), .C1(RF_pc_out[29]), .C2(n1949), .Z(
        register_file_inst1_n2198) );
  AO222D1BWP12T U2764 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[17]), .B1(n2286), .B2(
        IF_RF_incremented_pc_out[17]), .C1(RF_pc_out[17]), .C2(n2285), .Z(
        register_file_inst1_n2186) );
  AOI211D1BWP12T U2765 ( .A1(n2296), .A2(DEC_CPSR_update_flag_v), .B(reset), 
        .C(n2295), .ZN(register_file_inst1_cpsrin[0]) );
  IND2XD1BWP12T U2766 ( .A1(ALU_OUT_n), .B1(DEC_CPSR_update_flag_n), .ZN(n2290) );
  IND2XD1BWP12T U2767 ( .A1(ALU_OUT_c), .B1(DEC_CPSR_update_flag_c), .ZN(n2294) );
  AO222D1BWP12T U2768 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[10]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[10]), .C1(RF_pc_out[10]), .C2(n2285), .Z(
        register_file_inst1_n2179) );
  AO222D1BWP12T U2769 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[9]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[9]), .C1(RF_pc_out[9]), .C2(n2285), .Z(
        register_file_inst1_n2178) );
  AO222D1BWP12T U2770 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[8]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[8]), .C1(RF_pc_out[8]), .C2(n2285), .Z(
        register_file_inst1_n2177) );
  AO222D1BWP12T U2771 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[7]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[7]), .C1(RF_pc_out[7]), .C2(n2285), .Z(
        register_file_inst1_n2176) );
  AO222D1BWP12T U2772 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[6]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[6]), .C1(RF_pc_out[6]), .C2(n2285), .Z(
        register_file_inst1_n2175) );
  AO222D1BWP12T U2773 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[4]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[4]), .C1(RF_pc_out[4]), .C2(n2285), .Z(
        register_file_inst1_n2173) );
  AO222D1BWP12T U2774 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[3]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[3]), .C1(RF_pc_out[3]), .C2(n2285), .Z(
        register_file_inst1_n2172) );
  MUX2NXD0BWP12T U2775 ( .I0(MEMCTRL_RF_IF_data_in[10]), .I1(
        ALU_MISC_OUT_result[10]), .S(n2277), .ZN(n1929) );
  MUX2NXD0BWP12T U2776 ( .I0(MEMCTRL_RF_IF_data_in[6]), .I1(
        ALU_MISC_OUT_result[6]), .S(n2277), .ZN(n1930) );
  AOI211XD0BWP12T U2777 ( .A1(n2035), .A2(STACK_RF_next_sp[5]), .B(n1987), .C(
        reset), .ZN(n1988) );
  AOI211XD0BWP12T U2778 ( .A1(n2035), .A2(STACK_RF_next_sp[6]), .B(n2025), .C(
        reset), .ZN(n2026) );
  RCAOI211D0BWP12T U2779 ( .A1(n2035), .A2(STACK_RF_next_sp[1]), .B(n2034), 
        .C(reset), .ZN(n2036) );
  RCAOI211D0BWP12T U2780 ( .A1(n2035), .A2(STACK_RF_next_sp[3]), .B(n2031), 
        .C(reset), .ZN(n2032) );
  AO211D0BWP12T U2781 ( .A1(memory_interface_inst1_fsm_state_0_), .A2(n2289), 
        .B(n2288), .C(n501), .Z(MEMCTRL_read_finished) );
  NR2XD0BWP12T U2782 ( .A1(n1957), .A2(DEC_MEMCTRL_load_store_width[0]), .ZN(
        n1951) );
  RCAOI22D0BWP12T U2783 ( .A1(RF_pc_out[9]), .A2(n1944), .B1(
        register_file_inst1_lr_9_), .B2(n1943), .ZN(n2119) );
  AOI22D0BWP12T U2784 ( .A1(RF_pc_out[18]), .A2(n1932), .B1(
        register_file_inst1_lr_18_), .B2(n1947), .ZN(n2003) );
  AOI22D0BWP12T U2785 ( .A1(RF_pc_out[5]), .A2(n1932), .B1(
        register_file_inst1_lr_5_), .B2(n1947), .ZN(n1989) );
  AOI22D0BWP12T U2786 ( .A1(RF_pc_out[20]), .A2(n1932), .B1(
        register_file_inst1_lr_20_), .B2(n1947), .ZN(n1984) );
  AOI22D0BWP12T U2787 ( .A1(RF_pc_out[23]), .A2(n1932), .B1(
        register_file_inst1_lr_23_), .B2(n1947), .ZN(n1999) );
  AOI22D0BWP12T U2788 ( .A1(RF_pc_out[16]), .A2(n1932), .B1(
        register_file_inst1_lr_16_), .B2(n1947), .ZN(n2005) );
  AOI22D0BWP12T U2789 ( .A1(RF_pc_out[28]), .A2(n1932), .B1(
        register_file_inst1_r8_28_), .B2(n1948), .ZN(n1995) );
  AOI22D0BWP12T U2790 ( .A1(RF_pc_out[29]), .A2(n1932), .B1(
        register_file_inst1_lr_29_), .B2(n1947), .ZN(n1994) );
  AOI22D0BWP12T U2791 ( .A1(RF_pc_out[30]), .A2(n1932), .B1(
        register_file_inst1_lr_30_), .B2(n1947), .ZN(n1982) );
  AOI22D0BWP12T U2792 ( .A1(RF_pc_out[31]), .A2(n1932), .B1(
        register_file_inst1_lr_31_), .B2(n1947), .ZN(n1993) );
  AOI22D0BWP12T U2793 ( .A1(RF_pc_out[19]), .A2(n1932), .B1(
        register_file_inst1_r8_19_), .B2(n1948), .ZN(n2002) );
  AOI22D0BWP12T U2794 ( .A1(RF_pc_out[24]), .A2(n1932), .B1(
        register_file_inst1_lr_24_), .B2(n1947), .ZN(n1983) );
  AOI22D0BWP12T U2795 ( .A1(RF_pc_out[25]), .A2(n1932), .B1(
        register_file_inst1_lr_25_), .B2(n1947), .ZN(n1998) );
  AOI22D0BWP12T U2796 ( .A1(RF_pc_out[17]), .A2(n1932), .B1(
        register_file_inst1_lr_17_), .B2(n1947), .ZN(n2004) );
  AOI22D0BWP12T U2797 ( .A1(RF_pc_out[26]), .A2(n1932), .B1(
        register_file_inst1_r8_26_), .B2(n1948), .ZN(n1997) );
  AOI22D0BWP12T U2798 ( .A1(RF_pc_out[27]), .A2(n1932), .B1(
        register_file_inst1_lr_27_), .B2(n1947), .ZN(n1996) );
  AOI22D0BWP12T U2799 ( .A1(RF_pc_out[0]), .A2(n1932), .B1(
        register_file_inst1_lr_0_), .B2(n1947), .ZN(n2038) );
  AOI22D0BWP12T U2800 ( .A1(RF_pc_out[11]), .A2(n1932), .B1(
        register_file_inst1_r8_11_), .B2(n1948), .ZN(n2012) );
  AOI22D0BWP12T U2801 ( .A1(RF_pc_out[21]), .A2(n1932), .B1(
        register_file_inst1_lr_21_), .B2(n1947), .ZN(n2001) );
  AOI22D0BWP12T U2802 ( .A1(RF_pc_out[15]), .A2(n1932), .B1(
        register_file_inst1_r8_15_), .B2(n1948), .ZN(n2006) );
  AOI22D0BWP12T U2803 ( .A1(RF_pc_out[14]), .A2(n1932), .B1(
        register_file_inst1_lr_14_), .B2(n1947), .ZN(n1985) );
  AOI22D0BWP12T U2804 ( .A1(RF_pc_out[13]), .A2(n1932), .B1(
        register_file_inst1_lr_13_), .B2(n1947), .ZN(n1986) );
  RCAOI22D0BWP12T U2805 ( .A1(RF_pc_out[22]), .A2(n1937), .B1(
        register_file_inst1_r0_22_), .B2(n1938), .ZN(n2227) );
  AOI22D0BWP12T U2806 ( .A1(RF_pc_out[11]), .A2(n1940), .B1(
        register_file_inst1_r5_11_), .B2(n1939), .ZN(n2073) );
  AOI22D1BWP12T U2807 ( .A1(RF_pc_out[24]), .A2(n1937), .B1(
        register_file_inst1_r0_24_), .B2(n1938), .ZN(n2231) );
  AOI22D0BWP12T U2808 ( .A1(RF_pc_out[10]), .A2(n1940), .B1(
        register_file_inst1_r5_10_), .B2(n1939), .ZN(n2070) );
  AOI22D0BWP12T U2809 ( .A1(RF_pc_out[9]), .A2(n1940), .B1(
        register_file_inst1_r5_9_), .B2(n1939), .ZN(n2067) );
  AOI22D0BWP12T U2810 ( .A1(RF_pc_out[12]), .A2(n1940), .B1(
        register_file_inst1_r5_12_), .B2(n1939), .ZN(n2076) );
  NR2D1BWP12T U2811 ( .A1(RF_OUT_v), .A2(DEC_CPSR_update_flag_v), .ZN(n2295)
         );
  XOR2XD1BWP12T U2812 ( .A1(DEC_MEMCTRL_load_store_width[0]), .A2(n1953), .Z(
        n1956) );
  OR2D1BWP12T U2813 ( .A1(DEC_RF_operand_a[1]), .A2(DEC_RF_operand_a[2]), .Z(
        n2176) );
  AN2XD1BWP12T U2814 ( .A1(DEC_RF_alu_stack_write_to_reg[1]), .A2(
        DEC_RF_alu_stack_write_to_reg[2]), .Z(n2275) );
  OR2D1BWP12T U2815 ( .A1(DEC_RF_operand_b[2]), .A2(DEC_RF_operand_b[1]), .Z(
        n2097) );
  INR2D1BWP12T U2816 ( .A1(DEC_MISC_OUT_memory_address_source_is_reg), .B1(
        IF_memory_load_req), .ZN(n3) );
  ND3D0BWP12T U2817 ( .A1(DEC_RF_memory_write_to_reg[1]), .A2(n2293), .A3(
        n1972), .ZN(n1975) );
  NR3D1BWP12T U2818 ( .A1(DEC_RF_alu_stack_write_to_reg[4]), .A2(
        DEC_RF_alu_stack_write_to_reg[0]), .A3(n2084), .ZN(n1981) );
  NR2D1BWP12T U2819 ( .A1(DEC_RF_alu_stack_write_to_reg[0]), .A2(n1965), .ZN(
        n1968) );
  INVD1BWP12T U2820 ( .I(DEC_RF_memory_write_to_reg[2]), .ZN(n1972) );
  NR2D1BWP12T U2821 ( .A1(DEC_RF_alu_stack_write_to_reg[2]), .A2(n1962), .ZN(
        n1979) );
  IND3D1BWP12T U2822 ( .A1(DEC_RF_alu_stack_write_to_reg[3]), .B1(
        DEC_RF_alu_stack_write_to_reg_enable), .B2(n1959), .ZN(n1965) );
  IND4D1BWP12T U2823 ( .A1(n2084), .B1(DEC_RF_alu_stack_write_to_reg[4]), .B2(
        n2083), .B3(n2082), .ZN(n2168) );
  INVD1BWP12T U2824 ( .I(DEC_RF_alu_stack_write_to_reg[0]), .ZN(n2082) );
  INVD1BWP12T U2825 ( .I(DEC_RF_memory_write_to_reg[1]), .ZN(n1963) );
  AN3XD1BWP12T U2826 ( .A1(DEC_RF_memory_write_to_reg_enable), .A2(
        DEC_RF_memory_write_to_reg[0]), .A3(n2298), .Z(n2301) );
  INVD1BWP12T U2827 ( .I(DEC_RF_memory_write_to_reg[4]), .ZN(n2298) );
  INVD1BWP12T U2828 ( .I(DEC_RF_alu_stack_write_to_reg[1]), .ZN(n1960) );
  INVD1BWP12T U2829 ( .I(DEC_RF_alu_stack_write_to_reg[2]), .ZN(n1964) );
  INR3D0BWP12T U2830 ( .A1(DEC_RF_alu_stack_write_to_reg[0]), .B1(
        DEC_RF_alu_stack_write_to_reg[4]), .B2(n2084), .ZN(n2276) );
  ND2D1BWP12T U2831 ( .A1(DEC_RF_alu_stack_write_to_reg_enable), .A2(
        DEC_RF_alu_stack_write_to_reg[3]), .ZN(n2084) );
  INR2D1BWP12T U2832 ( .A1(DEC_RF_operand_b[3]), .B1(DEC_RF_operand_b[4]), 
        .ZN(n2305) );
  NR2D1BWP12T U2833 ( .A1(DEC_RF_operand_a[0]), .A2(n2182), .ZN(n2244) );
  ND2D1BWP12T U2834 ( .A1(DEC_RF_operand_a[2]), .A2(DEC_RF_operand_a[1]), .ZN(
        n2183) );
  INR2D1BWP12T U2835 ( .A1(DEC_RF_operand_a[3]), .B1(DEC_RF_operand_a[4]), 
        .ZN(n2303) );
  INVD1BWP12T U2836 ( .I(DEC_RF_operand_a[0]), .ZN(n2175) );
  NR2D1BWP12T U2837 ( .A1(DEC_RF_operand_a[3]), .A2(DEC_RF_operand_a[4]), .ZN(
        n2302) );
  NR2D1BWP12T U2838 ( .A1(DEC_MEMCTRL_load_store_width[1]), .A2(
        DEC_MEMCTRL_load_store_width[0]), .ZN(n2044) );
  ND3D1BWP12T U2839 ( .A1(DEC_RF_memory_store_data_reg[3]), .A2(n2306), .A3(
        n2313), .ZN(n2314) );
  ND3D1BWP12T U2840 ( .A1(DEC_RF_memory_store_data_reg[2]), .A2(
        DEC_RF_memory_store_data_reg[3]), .A3(n2306), .ZN(n2308) );
  ND2D1BWP12T U2841 ( .A1(DEC_RF_memory_store_data_reg[0]), .A2(n2316), .ZN(
        n2311) );
  INVD1BWP12T U2842 ( .I(DEC_RF_memory_store_data_reg[2]), .ZN(n2313) );
  ND2D1BWP12T U2843 ( .A1(DEC_RF_memory_store_data_reg[1]), .A2(
        DEC_RF_memory_store_data_reg[0]), .ZN(n2309) );
  INVD1BWP12T U2844 ( .I(DEC_RF_memory_store_data_reg[1]), .ZN(n2316) );
  ND2D1BWP12T U2845 ( .A1(DEC_RF_memory_store_data_reg[1]), .A2(n2315), .ZN(
        n2307) );
  INVD1BWP12T U2846 ( .I(DEC_RF_memory_store_data_reg[0]), .ZN(n2315) );
  ND2D1BWP12T U2847 ( .A1(DEC_RF_memory_store_data_reg[2]), .A2(n2312), .ZN(
        n2310) );
  INVD1BWP12T U2848 ( .I(DEC_RF_memory_store_data_reg[3]), .ZN(n2312) );
  ND2D1BWP12T U2849 ( .A1(DEC_MEMCTRL_load_store_width[0]), .A2(
        DEC_MEMCTRL_load_store_width[1]), .ZN(n2333) );
  INVD1BWP12T U2850 ( .I(DEC_MEMCTRL_CTRL_memory_store_request), .ZN(n2332) );
  INVD1BWP12T U2851 ( .I(DEC_MEMCTRL_load_store_width[1]), .ZN(n1953) );
  ND2D1BWP12T U2852 ( .A1(DEC_RF_memory_store_address_reg[2]), .A2(
        DEC_RF_memory_store_address_reg[3]), .ZN(n2323) );
  ND2D1BWP12T U2853 ( .A1(DEC_RF_memory_store_address_reg[0]), .A2(n2326), 
        .ZN(n2322) );
  ND2D1BWP12T U2854 ( .A1(DEC_RF_memory_store_address_reg[2]), .A2(n2325), 
        .ZN(n2320) );
  ND2D1BWP12T U2855 ( .A1(DEC_RF_memory_store_address_reg[0]), .A2(
        DEC_RF_memory_store_address_reg[1]), .ZN(n2321) );
  INVD1BWP12T U2856 ( .I(DEC_RF_memory_store_address_reg[3]), .ZN(n2325) );
  ND2D1BWP12T U2857 ( .A1(DEC_RF_memory_store_address_reg[3]), .A2(n2324), 
        .ZN(n2319) );
  INVD1BWP12T U2858 ( .I(DEC_RF_memory_store_address_reg[2]), .ZN(n2324) );
  INVD1BWP12T U2859 ( .I(DEC_RF_memory_store_address_reg[1]), .ZN(n2326) );
  ND2D1BWP12T U2860 ( .A1(DEC_RF_memory_write_to_reg[1]), .A2(n1972), .ZN(
        n1974) );
  INVD1BWP12T U2861 ( .I(DEC_RF_memory_write_to_reg[0]), .ZN(n1966) );
  INVD1BWP12T U2862 ( .I(DEC_RF_alu_stack_write_to_reg[4]), .ZN(n1959) );
  ND2D1BWP12T U2863 ( .A1(DEC_RF_memory_write_to_reg[2]), .A2(
        DEC_RF_memory_write_to_reg[1]), .ZN(n2278) );
  INVD1BWP12T U2864 ( .I(DEC_RF_memory_write_to_reg[3]), .ZN(n2299) );
  ND2D1BWP12T U2865 ( .A1(DEC_RF_memory_write_to_reg[2]), .A2(n1963), .ZN(
        n1977) );
  ND2D1BWP12T U2866 ( .A1(DEC_RF_memory_write_to_reg[3]), .A2(n2301), .ZN(
        n2279) );
  OAI21D1BWP12T U2867 ( .A1(n2081), .A2(DEC_ALU_alu_opcode[4]), .B(n2080), 
        .ZN(ALU_IN_c) );
  ND4D1BWP12T U2868 ( .A1(DEC_ALU_alu_opcode[1]), .A2(DEC_ALU_alu_opcode[2]), 
        .A3(DEC_ALU_alu_opcode[4]), .A4(n2079), .ZN(n2080) );
  NR2D1BWP12T U2869 ( .A1(DEC_ALU_alu_opcode[0]), .A2(DEC_ALU_alu_opcode[3]), 
        .ZN(n2079) );
  AOI22D1BWP12T U2870 ( .A1(register_file_inst1_r2_18_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[18]), .ZN(n2219) );
  AOI22D1BWP12T U2871 ( .A1(register_file_inst1_r2_18_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[18]), .ZN(n2142) );
  AOI22D1BWP12T U2872 ( .A1(register_file_inst1_r2_17_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[17]), .ZN(n2140) );
  AOI22D1BWP12T U2873 ( .A1(register_file_inst1_r2_17_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[17]), .ZN(n2217) );
  AOI22D1BWP12T U2874 ( .A1(register_file_inst1_r2_16_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[16]), .ZN(n2215) );
  AOI22D1BWP12T U2875 ( .A1(register_file_inst1_r2_16_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[16]), .ZN(n2138) );
  AOI22D1BWP12T U2876 ( .A1(register_file_inst1_r2_15_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[15]), .ZN(n2136) );
  AOI22D1BWP12T U2877 ( .A1(register_file_inst1_r2_15_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[15]), .ZN(n2213) );
  AOI22D1BWP12T U2878 ( .A1(register_file_inst1_r2_14_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[14]), .ZN(n2211) );
  AOI22D1BWP12T U2879 ( .A1(register_file_inst1_r2_14_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[14]), .ZN(n2133) );
  AOI22D1BWP12T U2880 ( .A1(register_file_inst1_r2_13_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[13]), .ZN(n2130) );
  AOI22D1BWP12T U2881 ( .A1(register_file_inst1_r2_13_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[13]), .ZN(n2209) );
  AOI22D1BWP12T U2882 ( .A1(register_file_inst1_r2_12_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[12]), .ZN(n2207) );
  AOI22D1BWP12T U2883 ( .A1(register_file_inst1_r2_12_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[12]), .ZN(n2127) );
  AOI22D1BWP12T U2884 ( .A1(register_file_inst1_r2_8_), .A2(n1946), .B1(n1945), 
        .B2(DEC_RF_offset_a[8]), .ZN(n2199) );
  AOI22D1BWP12T U2885 ( .A1(register_file_inst1_r2_8_), .A2(n1942), .B1(n1941), 
        .B2(DEC_RF_offset_b[8]), .ZN(n2116) );
  AOI22D1BWP12T U2886 ( .A1(register_file_inst1_r2_9_), .A2(n1942), .B1(n1941), 
        .B2(DEC_RF_offset_b[9]), .ZN(n2118) );
  AOI22D1BWP12T U2887 ( .A1(register_file_inst1_r2_9_), .A2(n1946), .B1(n1945), 
        .B2(DEC_RF_offset_a[9]), .ZN(n2201) );
  AOI22D1BWP12T U2888 ( .A1(register_file_inst1_r2_10_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[10]), .ZN(n2203) );
  AOI22D1BWP12T U2889 ( .A1(register_file_inst1_r2_10_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[10]), .ZN(n2121) );
  AOI22D1BWP12T U2890 ( .A1(register_file_inst1_r2_11_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[11]), .ZN(n2124) );
  AOI22D1BWP12T U2891 ( .A1(register_file_inst1_r2_11_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[11]), .ZN(n2205) );
  AOI22D1BWP12T U2892 ( .A1(register_file_inst1_r2_6_), .A2(n1946), .B1(n1945), 
        .B2(DEC_RF_offset_a[6]), .ZN(n2195) );
  AOI22D1BWP12T U2893 ( .A1(register_file_inst1_r2_6_), .A2(n1942), .B1(n1941), 
        .B2(DEC_RF_offset_b[6]), .ZN(n2111) );
  AOI22D1BWP12T U2894 ( .A1(register_file_inst1_r2_7_), .A2(n1942), .B1(n1941), 
        .B2(DEC_RF_offset_b[7]), .ZN(n2114) );
  AOI22D1BWP12T U2895 ( .A1(register_file_inst1_r2_7_), .A2(n1946), .B1(n1945), 
        .B2(DEC_RF_offset_a[7]), .ZN(n2197) );
  AOI22D1BWP12T U2896 ( .A1(register_file_inst1_r2_19_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[19]), .ZN(n2144) );
  AOI22D1BWP12T U2897 ( .A1(register_file_inst1_r2_19_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[19]), .ZN(n2221) );
  AOI22D1BWP12T U2898 ( .A1(register_file_inst1_r2_20_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[20]), .ZN(n2222) );
  AOI22D1BWP12T U2899 ( .A1(register_file_inst1_r2_20_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[20]), .ZN(n2146) );
  AOI22D1BWP12T U2900 ( .A1(register_file_inst1_r2_21_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[21]), .ZN(n2148) );
  AOI22D1BWP12T U2901 ( .A1(register_file_inst1_r2_22_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[22]), .ZN(n2150) );
  AOI22D1BWP12T U2902 ( .A1(register_file_inst1_r2_23_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[23]), .ZN(n2152) );
  AOI22D1BWP12T U2903 ( .A1(register_file_inst1_r2_24_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[24]), .ZN(n2230) );
  AOI22D1BWP12T U2904 ( .A1(register_file_inst1_r2_24_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[24]), .ZN(n2154) );
  AOI22D1BWP12T U2905 ( .A1(register_file_inst1_r2_25_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[25]), .ZN(n2156) );
  AOI22D1BWP12T U2906 ( .A1(register_file_inst1_r2_25_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[25]), .ZN(n2232) );
  AOI22D1BWP12T U2907 ( .A1(register_file_inst1_r2_26_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[26]), .ZN(n2158) );
  AOI22D1BWP12T U2908 ( .A1(register_file_inst1_r2_26_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[26]), .ZN(n2234) );
  AOI22D1BWP12T U2909 ( .A1(register_file_inst1_r2_27_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[27]), .ZN(n2160) );
  AOI22D1BWP12T U2910 ( .A1(register_file_inst1_r2_27_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[27]), .ZN(n2236) );
  AOI22D1BWP12T U2911 ( .A1(register_file_inst1_r2_28_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[28]), .ZN(n2162) );
  AOI22D1BWP12T U2912 ( .A1(register_file_inst1_r2_28_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[28]), .ZN(n2238) );
  AOI22D1BWP12T U2913 ( .A1(register_file_inst1_r2_29_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[29]), .ZN(n2164) );
  AOI22D1BWP12T U2914 ( .A1(register_file_inst1_r2_29_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[29]), .ZN(n2240) );
  AOI22D1BWP12T U2915 ( .A1(register_file_inst1_r2_30_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[30]), .ZN(n2166) );
  AOI22D1BWP12T U2916 ( .A1(register_file_inst1_r2_30_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[30]), .ZN(n2242) );
  AOI22D1BWP12T U2917 ( .A1(register_file_inst1_r2_31_), .A2(n1942), .B1(n1941), .B2(DEC_RF_offset_b[31]), .ZN(n2169) );
  AOI22D1BWP12T U2918 ( .A1(register_file_inst1_r2_31_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[31]), .ZN(n2245) );
  AOI22D1BWP12T U2919 ( .A1(register_file_inst1_r2_5_), .A2(n1942), .B1(n1941), 
        .B2(DEC_RF_offset_b[5]), .ZN(n2108) );
  AOI22D1BWP12T U2920 ( .A1(register_file_inst1_r2_4_), .A2(n1942), .B1(n1941), 
        .B2(DEC_RF_offset_b[4]), .ZN(n2106) );
  AOI22D1BWP12T U2921 ( .A1(register_file_inst1_r2_0_), .A2(n1946), .B1(n1945), 
        .B2(DEC_RF_offset_a[0]), .ZN(n2177) );
  AOI22D1BWP12T U2922 ( .A1(register_file_inst1_r2_4_), .A2(n1946), .B1(n1945), 
        .B2(DEC_RF_offset_a[4]), .ZN(n2191) );
  AOI22D1BWP12T U2923 ( .A1(register_file_inst1_r2_5_), .A2(n1946), .B1(n1945), 
        .B2(DEC_RF_offset_a[5]), .ZN(n2193) );
  AOI22D1BWP12T U2924 ( .A1(register_file_inst1_r2_3_), .A2(n1942), .B1(n1941), 
        .B2(DEC_RF_offset_b[3]), .ZN(n2104) );
  AOI22D1BWP12T U2925 ( .A1(register_file_inst1_r2_2_), .A2(n1942), .B1(n1941), 
        .B2(DEC_RF_offset_b[2]), .ZN(n2102) );
  AOI22D1BWP12T U2926 ( .A1(register_file_inst1_r2_3_), .A2(n1946), .B1(n1945), 
        .B2(DEC_RF_offset_a[3]), .ZN(n2189) );
  AOI22D1BWP12T U2927 ( .A1(register_file_inst1_r2_1_), .A2(n1946), .B1(n1945), 
        .B2(DEC_RF_offset_a[1]), .ZN(n2185) );
  AOI22D1BWP12T U2928 ( .A1(register_file_inst1_r2_2_), .A2(n1946), .B1(n1945), 
        .B2(DEC_RF_offset_a[2]), .ZN(n2187) );
  AOI22D1BWP12T U2929 ( .A1(register_file_inst1_r2_1_), .A2(n1942), .B1(n1941), 
        .B2(DEC_RF_offset_b[1]), .ZN(n2099) );
  AOI22D1BWP12T U2930 ( .A1(register_file_inst1_r2_0_), .A2(n1942), .B1(n1941), 
        .B2(DEC_RF_offset_b[0]), .ZN(n2091) );
  ND3D1BWP12T U2931 ( .A1(n2095), .A2(DEC_RF_operand_b[4]), .A3(
        DEC_RF_operand_b[3]), .ZN(n2096) );
  INVD1BWP12T U2932 ( .I(DEC_RF_operand_b[2]), .ZN(n2087) );
  NR2D1BWP12T U2933 ( .A1(DEC_RF_operand_b[4]), .A2(DEC_RF_operand_b[3]), .ZN(
        n2304) );
  ND2D1BWP12T U2934 ( .A1(DEC_RF_operand_b[2]), .A2(n2086), .ZN(n2090) );
  INVD1BWP12T U2935 ( .I(DEC_RF_operand_b[1]), .ZN(n2086) );
  INVD1BWP12T U2936 ( .I(DEC_RF_operand_b[0]), .ZN(n2089) );
  AOI22D1BWP12T U2937 ( .A1(register_file_inst1_r2_23_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[23]), .ZN(n2228) );
  AOI22D1BWP12T U2938 ( .A1(register_file_inst1_r2_21_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[21]), .ZN(n2224) );
  AOI22D1BWP12T U2939 ( .A1(register_file_inst1_r2_22_), .A2(n1946), .B1(n1945), .B2(DEC_RF_offset_a[22]), .ZN(n2226) );
  ND3D1BWP12T U2940 ( .A1(n2174), .A2(DEC_RF_operand_a[4]), .A3(
        DEC_RF_operand_a[3]), .ZN(n2182) );
  ND2D1BWP12T U2941 ( .A1(n2303), .A2(DEC_RF_operand_a[0]), .ZN(n2181) );
  ND2D1BWP12T U2942 ( .A1(DEC_RF_operand_a[0]), .A2(n2302), .ZN(n2180) );
  ND2D1BWP12T U2943 ( .A1(DEC_RF_operand_a[1]), .A2(n2173), .ZN(n2179) );
  INVD1BWP12T U2944 ( .I(DEC_RF_operand_a[2]), .ZN(n2173) );
  ND2D1BWP12T U2945 ( .A1(DEC_RF_operand_a[2]), .A2(n2171), .ZN(n2178) );
  INVD1BWP12T U2946 ( .I(DEC_RF_operand_a[1]), .ZN(n2171) );
  IND4D1BWP12T U2947 ( .A1(DEC_RF_memory_write_to_reg[4]), .B1(
        DEC_RF_memory_write_to_reg_enable), .B2(n2299), .B3(n1966), .ZN(n1969)
         );
  INR3D0BWP12T U2948 ( .A1(DEC_RF_memory_write_to_reg_enable), .B1(
        DEC_RF_memory_write_to_reg[0]), .B2(n2299), .ZN(n2300) );
  ND2D1BWP12T U2949 ( .A1(n2305), .A2(DEC_RF_operand_b[0]), .ZN(n2094) );
  ND2D1BWP12T U2950 ( .A1(DEC_RF_operand_b[2]), .A2(DEC_RF_operand_b[1]), .ZN(
        n2088) );
  ND2D1BWP12T U2951 ( .A1(n2304), .A2(DEC_RF_operand_b[0]), .ZN(n2092) );
  ND2D1BWP12T U2952 ( .A1(DEC_RF_operand_b[1]), .A2(n2087), .ZN(n2093) );
  IND2D1BWP12T U2953 ( .A1(DEC_RF_memory_store_address_reg[0]), .B1(
        DEC_RF_memory_store_address_reg[1]), .ZN(n2317) );
  IND2D1BWP12T U2954 ( .A1(DEC_RF_memory_store_address_reg[0]), .B1(n2326), 
        .ZN(n2318) );
  NR2D1BWP12T U2955 ( .A1(IF_memory_load_req), .A2(
        DEC_MISC_OUT_memory_address_source_is_reg), .ZN(n4) );
  AOI22D0BWP12T U2956 ( .A1(RF_pc_out[22]), .A2(n1932), .B1(
        register_file_inst1_r8_22_), .B2(n1948), .ZN(n2000) );
  AOI22D0BWP12T U2957 ( .A1(RF_pc_out[7]), .A2(n1932), .B1(
        register_file_inst1_lr_7_), .B2(n1947), .ZN(n2024) );
  AOI22D1BWP12T U2958 ( .A1(RF_pc_out[6]), .A2(n1932), .B1(
        register_file_inst1_lr_6_), .B2(n1947), .ZN(n2027) );
  AOI22D0BWP12T U2959 ( .A1(RF_pc_out[4]), .A2(n1932), .B1(
        register_file_inst1_lr_4_), .B2(n1947), .ZN(n2030) );
  AOI22D0BWP12T U2960 ( .A1(RF_pc_out[3]), .A2(n1932), .B1(
        register_file_inst1_lr_3_), .B2(n1947), .ZN(n2033) );
  AOI22D0BWP12T U2961 ( .A1(RF_pc_out[2]), .A2(n1932), .B1(
        register_file_inst1_lr_2_), .B2(n1947), .ZN(n1992) );
  OAI21D1BWP12T U2962 ( .A1(n2327), .A2(n501), .B(n2270), .ZN(
        MEMCTRL_RF_IF_data_in[7]) );
  OAI21D1BWP12T U2963 ( .A1(n501), .A2(n2331), .B(n2274), .ZN(
        MEMCTRL_RF_IF_data_in[0]) );
  OAI21D1BWP12T U2964 ( .A1(n501), .A2(n2330), .B(n2273), .ZN(
        MEMCTRL_RF_IF_data_in[4]) );
  OAI21D1BWP12T U2965 ( .A1(n501), .A2(n2329), .B(n2272), .ZN(
        MEMCTRL_RF_IF_data_in[5]) );
  OAI21D1BWP12T U2966 ( .A1(n501), .A2(n2328), .B(n2271), .ZN(
        MEMCTRL_RF_IF_data_in[6]) );
  AOI22D0BWP12T U2967 ( .A1(RF_pc_out[1]), .A2(n1932), .B1(
        register_file_inst1_lr_1_), .B2(n1947), .ZN(n2037) );
  AOI22D1BWP12T U2968 ( .A1(RF_pc_out[12]), .A2(n1944), .B1(
        register_file_inst1_lr_12_), .B2(n1943), .ZN(n2128) );
  AOI22D1BWP12T U2969 ( .A1(RF_pc_out[14]), .A2(n1944), .B1(
        register_file_inst1_lr_14_), .B2(n1943), .ZN(n2134) );
  AOI22D1BWP12T U2970 ( .A1(RF_pc_out[16]), .A2(n1944), .B1(
        register_file_inst1_lr_16_), .B2(n1943), .ZN(n2139) );
  AOI22D1BWP12T U2971 ( .A1(RF_pc_out[18]), .A2(n1944), .B1(
        register_file_inst1_lr_18_), .B2(n1943), .ZN(n2143) );
  AOI22D1BWP12T U2972 ( .A1(RF_pc_out[20]), .A2(n1944), .B1(
        register_file_inst1_lr_20_), .B2(n1943), .ZN(n2147) );
  AOI22D1BWP12T U2973 ( .A1(RF_pc_out[22]), .A2(n1944), .B1(
        register_file_inst1_lr_22_), .B2(n1943), .ZN(n2151) );
  AOI22D1BWP12T U2974 ( .A1(RF_pc_out[24]), .A2(n1944), .B1(
        register_file_inst1_lr_24_), .B2(n1943), .ZN(n2155) );
  AOI22D1BWP12T U2975 ( .A1(RF_pc_out[26]), .A2(n1944), .B1(
        register_file_inst1_lr_26_), .B2(n1943), .ZN(n2159) );
  AOI22D1BWP12T U2976 ( .A1(RF_pc_out[28]), .A2(n1944), .B1(
        register_file_inst1_lr_28_), .B2(n1943), .ZN(n2163) );
  AOI22D1BWP12T U2977 ( .A1(RF_pc_out[29]), .A2(n1944), .B1(
        register_file_inst1_lr_29_), .B2(n1943), .ZN(n2165) );
  AOI22D1BWP12T U2978 ( .A1(RF_pc_out[21]), .A2(n1937), .B1(
        register_file_inst1_r0_21_), .B2(n1938), .ZN(n2225) );
  AOI22D1BWP12T U2979 ( .A1(RF_pc_out[20]), .A2(n1937), .B1(
        register_file_inst1_r0_20_), .B2(n1938), .ZN(n2223) );
  AOI22D1BWP12T U2980 ( .A1(RF_pc_out[23]), .A2(n1937), .B1(
        register_file_inst1_r0_23_), .B2(n1938), .ZN(n2229) );
  AOI22D1BWP12T U2981 ( .A1(RF_pc_out[25]), .A2(n1937), .B1(
        register_file_inst1_r0_25_), .B2(n1938), .ZN(n2233) );
  AOI22D1BWP12T U2982 ( .A1(RF_pc_out[26]), .A2(n1937), .B1(
        register_file_inst1_r0_26_), .B2(n1938), .ZN(n2235) );
  AOI22D1BWP12T U2983 ( .A1(RF_pc_out[27]), .A2(n1937), .B1(
        register_file_inst1_r0_27_), .B2(n1938), .ZN(n2237) );
  AOI22D1BWP12T U2984 ( .A1(RF_pc_out[28]), .A2(n1937), .B1(
        register_file_inst1_r0_28_), .B2(n1938), .ZN(n2239) );
  AOI22D1BWP12T U2985 ( .A1(RF_pc_out[29]), .A2(n1937), .B1(
        register_file_inst1_r0_29_), .B2(n1938), .ZN(n2241) );
  AOI22D1BWP12T U2986 ( .A1(RF_pc_out[30]), .A2(n1937), .B1(
        register_file_inst1_r0_30_), .B2(n1938), .ZN(n2243) );
  AOI22D1BWP12T U2987 ( .A1(RF_pc_out[31]), .A2(n1937), .B1(
        register_file_inst1_r0_31_), .B2(n1938), .ZN(n2246) );
  AOI22D1BWP12T U2988 ( .A1(RF_pc_out[1]), .A2(n1944), .B1(
        register_file_inst1_lr_1_), .B2(n1943), .ZN(n2100) );
  AOI22D1BWP12T U2989 ( .A1(RF_pc_out[5]), .A2(n1944), .B1(
        register_file_inst1_lr_5_), .B2(n1943), .ZN(n2109) );
  AOI22D1BWP12T U2990 ( .A1(RF_pc_out[6]), .A2(n1944), .B1(
        register_file_inst1_lr_6_), .B2(n1943), .ZN(n2112) );
  AOI22D1BWP12T U2991 ( .A1(RF_pc_out[10]), .A2(n1944), .B1(
        register_file_inst1_lr_10_), .B2(n1943), .ZN(n2122) );
  AOI22D1BWP12T U2992 ( .A1(RF_pc_out[11]), .A2(n1944), .B1(
        register_file_inst1_lr_11_), .B2(n1943), .ZN(n2125) );
  AOI22D1BWP12T U2993 ( .A1(RF_pc_out[13]), .A2(n1944), .B1(
        register_file_inst1_lr_13_), .B2(n1943), .ZN(n2131) );
  AOI22D1BWP12T U2994 ( .A1(RF_pc_out[15]), .A2(n1944), .B1(
        register_file_inst1_lr_15_), .B2(n1943), .ZN(n2137) );
  AOI22D1BWP12T U2995 ( .A1(RF_pc_out[17]), .A2(n1944), .B1(
        register_file_inst1_lr_17_), .B2(n1943), .ZN(n2141) );
  AOI22D1BWP12T U2996 ( .A1(RF_pc_out[19]), .A2(n1944), .B1(
        register_file_inst1_lr_19_), .B2(n1943), .ZN(n2145) );
  AOI22D1BWP12T U2997 ( .A1(RF_pc_out[21]), .A2(n1944), .B1(
        register_file_inst1_lr_21_), .B2(n1943), .ZN(n2149) );
  AOI22D1BWP12T U2998 ( .A1(RF_pc_out[23]), .A2(n1944), .B1(
        register_file_inst1_lr_23_), .B2(n1943), .ZN(n2153) );
  AOI22D1BWP12T U2999 ( .A1(RF_pc_out[25]), .A2(n1944), .B1(
        register_file_inst1_lr_25_), .B2(n1943), .ZN(n2157) );
  AOI22D1BWP12T U3000 ( .A1(RF_pc_out[27]), .A2(n1944), .B1(
        register_file_inst1_lr_27_), .B2(n1943), .ZN(n2161) );
  AOI22D1BWP12T U3001 ( .A1(RF_pc_out[30]), .A2(n1944), .B1(
        register_file_inst1_lr_30_), .B2(n1943), .ZN(n2167) );
  AOI22D1BWP12T U3002 ( .A1(RF_pc_out[31]), .A2(n1944), .B1(
        register_file_inst1_lr_31_), .B2(n1943), .ZN(n2170) );
  AOI211D1BWP12T U3003 ( .A1(n2250), .A2(n2249), .B(n2248), .C(n2247), .ZN(
        MEMCTRL_write_finished) );
  AOI22D0BWP12T U3004 ( .A1(RF_pc_out[9]), .A2(n1932), .B1(STACK_RF_next_sp[9]), .B2(n1927), .ZN(n2018) );
  AOI22D0BWP12T U3005 ( .A1(RF_pc_out[8]), .A2(n1932), .B1(STACK_RF_next_sp[8]), .B2(n1927), .ZN(n2021) );
  AOI22D0BWP12T U3006 ( .A1(RF_pc_out[2]), .A2(n1940), .B1(
        register_file_inst1_r5_2_), .B2(n1939), .ZN(n2046) );
  AOI22D0BWP12T U3007 ( .A1(RF_pc_out[3]), .A2(n1940), .B1(
        register_file_inst1_r5_3_), .B2(n1939), .ZN(n2049) );
  AOI22D0BWP12T U3008 ( .A1(RF_pc_out[4]), .A2(n1940), .B1(
        register_file_inst1_r5_4_), .B2(n1939), .ZN(n2052) );
  AOI22D0BWP12T U3009 ( .A1(RF_pc_out[5]), .A2(n1940), .B1(
        register_file_inst1_r5_5_), .B2(n1939), .ZN(n2055) );
  AOI22D0BWP12T U3010 ( .A1(RF_pc_out[6]), .A2(n1940), .B1(
        register_file_inst1_r5_6_), .B2(n1939), .ZN(n2058) );
  AOI22D0BWP12T U3011 ( .A1(RF_pc_out[7]), .A2(n1940), .B1(
        register_file_inst1_r5_7_), .B2(n1939), .ZN(n2061) );
  AOI22D0BWP12T U3012 ( .A1(RF_pc_out[8]), .A2(n1940), .B1(
        register_file_inst1_r5_8_), .B2(n1939), .ZN(n2064) );
  OAI211D1BWP12T U3013 ( .A1(n2269), .A2(n2255), .B(n2267), .C(n2254), .ZN(
        MEMCTRL_RF_IF_data_in[14]) );
  AOI22D1BWP12T U3014 ( .A1(RF_pc_out[31]), .A2(n1949), .B1(n2286), .B2(
        IF_RF_incremented_pc_out[31]), .ZN(n2281) );
  OAI211D1BWP12T U3015 ( .A1(n2269), .A2(n2268), .B(n2267), .C(n2266), .ZN(
        MEMCTRL_RF_IF_data_in[8]) );
  OAI211D1BWP12T U3016 ( .A1(n2269), .A2(n2261), .B(n2267), .C(n2260), .ZN(
        MEMCTRL_RF_IF_data_in[11]) );
  OAI211D1BWP12T U3017 ( .A1(n2269), .A2(n2259), .B(n2267), .C(n2258), .ZN(
        MEMCTRL_RF_IF_data_in[12]) );
  OAI211D1BWP12T U3018 ( .A1(n2269), .A2(n2257), .B(n2267), .C(n2256), .ZN(
        MEMCTRL_RF_IF_data_in[13]) );
  OAI211D1BWP12T U3019 ( .A1(n2269), .A2(n2253), .B(n2267), .C(n2252), .ZN(
        MEMCTRL_RF_IF_data_in[15]) );
  OAI211D1BWP12T U3020 ( .A1(n2269), .A2(n2265), .B(n2267), .C(n2264), .ZN(
        MEMCTRL_RF_IF_data_in[9]) );
  OAI211D1BWP12T U3021 ( .A1(n2269), .A2(n2263), .B(n2267), .C(n2262), .ZN(
        MEMCTRL_RF_IF_data_in[10]) );
  INVD1BWP12T U3022 ( .I(MEMCTRL_RF_IF_data_in[7]), .ZN(n2113) );
  INVD1BWP12T U3023 ( .I(MEMCTRL_RF_IF_data_in[4]), .ZN(n2105) );
  INVD1BWP12T U3024 ( .I(MEMCTRL_RF_IF_data_in[5]), .ZN(n2107) );
  INVD1BWP12T U3025 ( .I(MEMCTRL_RF_IF_data_in[6]), .ZN(n2110) );
  INVD1BWP12T U3026 ( .I(MEMCTRL_RF_IF_data_in[0]), .ZN(n2085) );
  MUX2D1BWP12T U3027 ( .I0(MEM_MEMCTRL_from_mem_data[9]), .I1(
        memory_interface_inst1_delay_first_two_bytes_out[1]), .S(n501), .Z(
        MEMCTRL_RF_IF_data_in[1]) );
  MUX2D1BWP12T U3028 ( .I0(MEM_MEMCTRL_from_mem_data[10]), .I1(
        memory_interface_inst1_delay_first_two_bytes_out[2]), .S(n501), .Z(
        MEMCTRL_RF_IF_data_in[2]) );
  MUX2D1BWP12T U3029 ( .I0(MEM_MEMCTRL_from_mem_data[11]), .I1(
        memory_interface_inst1_delay_first_two_bytes_out[3]), .S(n501), .Z(
        MEMCTRL_RF_IF_data_in[3]) );
  NR2D1BWP12T U3030 ( .A1(MEMCTRL_write_finished), .A2(n1961), .ZN(n2251) );
  INVD1BWP12T U3031 ( .I(MEMCTRL_RF_IF_data_in[1]), .ZN(n2098) );
  INVD1BWP12T U3032 ( .I(MEMCTRL_RF_IF_data_in[2]), .ZN(n2101) );
  INVD1BWP12T U3033 ( .I(MEMCTRL_RF_IF_data_in[3]), .ZN(n2103) );
  AOI211D1BWP12T U3034 ( .A1(n2035), .A2(STACK_RF_next_sp[10]), .B(n2013), .C(
        reset), .ZN(n2014) );
  AO222D1BWP12T U3035 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[28]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[28]), .C1(RF_pc_out[28]), .C2(n1949), .Z(
        register_file_inst1_n2197) );
  AO222D1BWP12T U3036 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[27]), .B1(n2286), .B2(
        IF_RF_incremented_pc_out[27]), .C1(RF_pc_out[27]), .C2(n1949), .Z(
        register_file_inst1_n2196) );
  AO222D1BWP12T U3037 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[26]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[26]), .C1(RF_pc_out[26]), .C2(n1949), .Z(
        register_file_inst1_n2195) );
  AO222D1BWP12T U3038 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[25]), .B1(n2286), .B2(
        IF_RF_incremented_pc_out[25]), .C1(RF_pc_out[25]), .C2(n1949), .Z(
        register_file_inst1_n2194) );
  AO222D1BWP12T U3039 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[24]), .B1(n2286), .B2(
        IF_RF_incremented_pc_out[24]), .C1(RF_pc_out[24]), .C2(n1949), .Z(
        register_file_inst1_n2193) );
  AO222D1BWP12T U3040 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[23]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[23]), .C1(RF_pc_out[23]), .C2(n1949), .Z(
        register_file_inst1_n2192) );
  AO222D1BWP12T U3041 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[21]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[21]), .C1(RF_pc_out[21]), .C2(n1949), .Z(
        register_file_inst1_n2190) );
  AO222D1BWP12T U3042 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[18]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[18]), .C1(RF_pc_out[18]), .C2(n2285), .Z(
        register_file_inst1_n2187) );
  AO222D1BWP12T U3043 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[16]), .B1(n2286), .B2(
        IF_RF_incremented_pc_out[16]), .C1(RF_pc_out[16]), .C2(n2285), .Z(
        register_file_inst1_n2185) );
  AO222D1BWP12T U3044 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[14]), .B1(n2286), .B2(
        IF_RF_incremented_pc_out[14]), .C1(RF_pc_out[14]), .C2(n1949), .Z(
        register_file_inst1_n2183) );
  AO222D1BWP12T U3045 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[5]), .B1(n2286), .B2(
        IF_RF_incremented_pc_out[5]), .C1(RF_pc_out[5]), .C2(n1949), .Z(
        register_file_inst1_n2174) );
  AO222D1BWP12T U3046 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[2]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[2]), .C1(RF_pc_out[2]), .C2(n1949), .Z(
        register_file_inst1_n2171) );
  AO222D1BWP12T U3047 ( .A1(register_file_inst1_pc_write_in_0_), .A2(n2287), 
        .B1(n1950), .B2(IF_RF_incremented_pc_out[0]), .C1(n2285), .C2(
        RF_pc_out[0]), .Z(register_file_inst1_n2169) );
  AO222D1BWP12T U3048 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[20]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[20]), .C1(RF_pc_out[20]), .C2(n1949), .Z(
        register_file_inst1_n2189) );
  AO222D1BWP12T U3049 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[15]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[15]), .C1(RF_pc_out[15]), .C2(n2285), .Z(
        register_file_inst1_n2184) );
  AO222D1BWP12T U3050 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[13]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[13]), .C1(RF_pc_out[13]), .C2(n1949), .Z(
        register_file_inst1_n2182) );
  AO222D1BWP12T U3051 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[12]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[12]), .C1(RF_pc_out[12]), .C2(n2285), .Z(
        register_file_inst1_n2181) );
  AO222D1BWP12T U3052 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[11]), .B1(n1950), .B2(
        IF_RF_incremented_pc_out[11]), .C1(RF_pc_out[11]), .C2(n2285), .Z(
        register_file_inst1_n2180) );
  ND2D1BWP12T U3053 ( .A1(RF_pc_out[1]), .A2(n1949), .ZN(n2282) );
  AO222D1BWP12T U3054 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[22]), .B1(n2286), .B2(
        IF_RF_incremented_pc_out[22]), .C1(RF_pc_out[22]), .C2(n1949), .Z(
        register_file_inst1_n2191) );
  AO222D1BWP12T U3055 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[19]), .B1(n2286), .B2(
        IF_RF_incremented_pc_out[19]), .C1(RF_pc_out[19]), .C2(n1949), .Z(
        register_file_inst1_n2188) );
  AOI211D1BWP12T U3056 ( .A1(n2292), .A2(DEC_CPSR_update_flag_z), .B(reset), 
        .C(n2291), .ZN(register_file_inst1_cpsrin[1]) );
  NR2D1BWP12T U3057 ( .A1(RF_OUT_z), .A2(DEC_CPSR_update_flag_z), .ZN(n2291)
         );
  INVD1BWP12T U3058 ( .I(RF_pc_out[5]), .ZN(n2192) );
  INVD1BWP12T U3059 ( .I(RF_pc_out[6]), .ZN(n2194) );
  INVD1BWP12T U3060 ( .I(RF_pc_out[9]), .ZN(n2200) );
  INVD1BWP12T U3061 ( .I(RF_pc_out[10]), .ZN(n2202) );
  INVD1BWP12T U3062 ( .I(RF_pc_out[11]), .ZN(n2204) );
  INVD1BWP12T U3063 ( .I(RF_pc_out[12]), .ZN(n2206) );
  INVD1BWP12T U3064 ( .I(RF_pc_out[13]), .ZN(n2208) );
  INVD1BWP12T U3065 ( .I(RF_pc_out[14]), .ZN(n2210) );
  INVD1BWP12T U3066 ( .I(RF_pc_out[15]), .ZN(n2212) );
  INVD1BWP12T U3067 ( .I(RF_pc_out[16]), .ZN(n2214) );
  INVD1BWP12T U3068 ( .I(RF_pc_out[17]), .ZN(n2216) );
  INVD1BWP12T U3069 ( .I(RF_pc_out[18]), .ZN(n2218) );
  INVD1BWP12T U3070 ( .I(RF_pc_out[19]), .ZN(n2220) );
  INVD1BWP12T U3071 ( .I(RF_pc_out[0]), .ZN(n2172) );
  AOI21D1BWP12T U3072 ( .A1(n2045), .A2(n1955), .B(reset), .ZN(
        memory_interface_inst1_fsm_N35) );
  NR2D1BWP12T U3073 ( .A1(n1954), .A2(reset), .ZN(
        memory_interface_inst1_fsm_N34) );
  NR2D1BWP12T U3074 ( .A1(n1952), .A2(reset), .ZN(
        memory_interface_inst1_fsm_N33) );
  NR2D1BWP12T U3075 ( .A1(n1958), .A2(reset), .ZN(
        memory_interface_inst1_fsm_N32) );
  INVD1BWP12T U3076 ( .I(RF_OUT_c), .ZN(n2081) );
  NR3D1BWP12T U3077 ( .A1(reset), .A2(IF_RF_incremented_pc_write_enable), .A3(
        n2280), .ZN(n2285) );
  INR3D0BWP12T U3078 ( .A1(IF_RF_incremented_pc_write_enable), .B1(reset), 
        .B2(n2280), .ZN(n2286) );
  NR2D1BWP12T U3079 ( .A1(MEMCTRL_write_finished), .A2(n2039), .ZN(n2297) );
  IND2D1BWP12T U3080 ( .A1(MEMCTRL_write_finished), .B1(n2040), .ZN(n2043) );
  NR2D1BWP12T U3081 ( .A1(reset), .A2(n1936), .ZN(n1978) );
  NR2D1BWP12T U3082 ( .A1(reset), .A2(n1935), .ZN(n1970) );
  NR2D1BWP12T U3083 ( .A1(reset), .A2(n1934), .ZN(n1971) );
  NR2D1BWP12T U3084 ( .A1(reset), .A2(n1933), .ZN(n1980) );
  INVD1BWP12T U3085 ( .I(MEMCTRL_write_finished), .ZN(n2042) );
  NR2D1BWP12T U3086 ( .A1(reset), .A2(n1967), .ZN(n2083) );
  INVD1BWP12T U3087 ( .I(MEMCTRL_read_finished), .ZN(n2041) );
  INVD1BWP12T U3088 ( .I(reset), .ZN(n2293) );
  AO222D1BWP12T U3089 ( .A1(n2287), .A2(
        register_file_inst1_pc_write_in_plus_two[30]), .B1(n2286), .B2(
        IF_RF_incremented_pc_out[30]), .C1(RF_pc_out[30]), .C2(n1949), .Z(
        register_file_inst1_n2199) );
  RCIAO21D0BWP12T U3090 ( .A1(n2048), .A2(n2047), .B(
        DEC_RF_memory_store_address_reg[4]), .ZN(RF_MEMCTRL_address_reg[2]) );
  RCIAO21D0BWP12T U3091 ( .A1(n2051), .A2(n2050), .B(
        DEC_RF_memory_store_address_reg[4]), .ZN(RF_MEMCTRL_address_reg[3]) );
  RCIAO21D0BWP12T U3092 ( .A1(n2054), .A2(n2053), .B(
        DEC_RF_memory_store_address_reg[4]), .ZN(RF_MEMCTRL_address_reg[4]) );
  RCIAO21D0BWP12T U3093 ( .A1(n2057), .A2(n2056), .B(
        DEC_RF_memory_store_address_reg[4]), .ZN(RF_MEMCTRL_address_reg[5]) );
  RCIAO21D0BWP12T U3094 ( .A1(n2060), .A2(n2059), .B(
        DEC_RF_memory_store_address_reg[4]), .ZN(RF_MEMCTRL_address_reg[6]) );
  RCIAO21D0BWP12T U3095 ( .A1(n2063), .A2(n2062), .B(
        DEC_RF_memory_store_address_reg[4]), .ZN(RF_MEMCTRL_address_reg[7]) );
  RCIAO21D0BWP12T U3096 ( .A1(n2066), .A2(n2065), .B(
        DEC_RF_memory_store_address_reg[4]), .ZN(RF_MEMCTRL_address_reg[8]) );
  RCIAO21D0BWP12T U3097 ( .A1(n2069), .A2(n2068), .B(
        DEC_RF_memory_store_address_reg[4]), .ZN(RF_MEMCTRL_address_reg[9]) );
  RCIAO21D0BWP12T U3098 ( .A1(n2072), .A2(n2071), .B(
        DEC_RF_memory_store_address_reg[4]), .ZN(RF_MEMCTRL_address_reg[10])
         );
  RCIAO21D0BWP12T U3099 ( .A1(n2075), .A2(n2074), .B(
        DEC_RF_memory_store_address_reg[4]), .ZN(RF_MEMCTRL_address_reg[11])
         );
  RCIAO21D0BWP12T U3100 ( .A1(n2078), .A2(n2077), .B(
        DEC_RF_memory_store_address_reg[4]), .ZN(RF_MEMCTRL_address_reg[12])
         );
  OA211D1BWP12T U3101 ( .A1(DEC_CPSR_update_flag_n), .A2(RF_OUT_n), .B(n2290), 
        .C(n2293), .Z(register_file_inst1_cpsrin[3]) );
  OA211D1BWP12T U3102 ( .A1(DEC_CPSR_update_flag_c), .A2(RF_OUT_c), .B(n2294), 
        .C(n2293), .Z(register_file_inst1_cpsrin[2]) );
endmodule

