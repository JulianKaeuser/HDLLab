`define R0 4'b0000
`define R1 4'b0001
`define R2 4'b0010
`define R3 4'b0011
`define R4 4'b0100
`define R5 4'b0101
`define R6 4'b0110
`define R7 4'b0111

`define SP 4'b1000
`define PC 4'b1001
`define LR 4'b1010
`define IMM 4'b1111

`timescale 1ns/10ps
module register_file_tb ();

// needed wires
reg [31:0] write_in, immediate_in, next_pc, cpsr_in;
wire [31:0] regA, regB, pc_out, cpsr_out;
reg clk, write_en, pc_en;
reg [3:0] regA_sel, regB_sel, write_dest;

//dut
register_file rf (
.regA_select(regA_sel),
.regB_select(regB_sel),
.write_dest(write_dest),
.write_en(write_en),
.write_in(write_in),
.immediate_in(immediate_in),
.cpsr_in(cpsr_in),
.next_pc(next_pc),
.pc_en(pc_en),
.clk(clk),
.regA_out(regA),
.regB_out(regB),
.pc_out(pc_out),
.cpsr_out(cpsr_out)
);


initial begin
   // 1 bit signals
   clk = 0;
   pc_en = 1;
   write_en = 0;

   // 4 bit signals
   regA_sel = `R0;
   regB_sel = `R0;
   write_dest = `R1;

   // 32 bit signals
   write_in = 31'b0;
   immediate_in = 31'b11;
   cpsr_in = 31'b0;
   next_pc = 31'b0;
end

// some clock action
always begin
#5 clk = !clk;
end

initial begin
   $dumpfile("register_file.vcd");
   $dumpvars;

   $display("\t\ttime,\tclk"); 
   $monitor("%d,\t%b, \t%b, \t%b ",$time, clk, pc_en, write_en, regA_sel, regB_sel, write_dest, ); 
end

initial begin

   #5;
   #100;
   $finish;
end
endmodule

`undef R0
`undef R1
`undef R2
`undef R3
`undef R4
`undef R5
`undef R6
`undef R7

`undef PC
`undef LR
`undef IMM
`undef SP
