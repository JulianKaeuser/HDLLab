
module register_file ( readA_sel, readB_sel, readC_sel, readD_sel, write1_sel, 
        write2_sel, write1_en, write2_en, write1_in, write2_in, immediate1_in, 
        immediate2_in, next_pc_in, next_cpsr_in, next_sp_in, clk, reset, 
        regA_out, regB_out, regC_out, regD_out, pc_out, cpsr_out, sp_out, 
        next_pc_en_BAR );
  input [4:0] readA_sel;
  input [4:0] readB_sel;
  input [4:0] readC_sel;
  input [4:0] readD_sel;
  input [4:0] write1_sel;
  input [4:0] write2_sel;
  input [31:0] write1_in;
  input [31:0] write2_in;
  input [31:0] immediate1_in;
  input [31:0] immediate2_in;
  input [31:0] next_pc_in;
  input [3:0] next_cpsr_in;
  input [31:0] next_sp_in;
  output [31:0] regA_out;
  output [31:0] regB_out;
  output [31:0] regC_out;
  output [31:0] regD_out;
  output [31:0] pc_out;
  output [3:0] cpsr_out;
  output [31:0] sp_out;
  input write1_en, write2_en, clk, reset, next_pc_en_BAR;
  wire   n2136, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008;
  wire   [2010:2041] n;
  wire   [31:0] r0;
  wire   [31:0] r1;
  wire   [31:0] r2;
  wire   [31:0] r3;
  wire   [31:0] r4;
  wire   [31:0] r5;
  wire   [31:0] r6;
  wire   [31:0] r7;
  wire   [31:0] r8;
  wire   [31:0] r9;
  wire   [31:0] r10;
  wire   [31:0] r11;
  wire   [31:0] r12;
  wire   [31:0] lr;
  wire   [31:0] tmp1;
  wire   [31:0] spin;
  wire   [3:0] cpsrin;

  DFQD1BWP12T r0_reg_31_ ( .D(n2648), .CP(clk), .Q(r0[31]) );
  DFQD1BWP12T r0_reg_30_ ( .D(n2647), .CP(clk), .Q(r0[30]) );
  DFQD1BWP12T r0_reg_29_ ( .D(n2646), .CP(clk), .Q(r0[29]) );
  DFQD1BWP12T r0_reg_28_ ( .D(n2645), .CP(clk), .Q(r0[28]) );
  DFQD1BWP12T r0_reg_27_ ( .D(n2644), .CP(clk), .Q(r0[27]) );
  DFQD1BWP12T r0_reg_26_ ( .D(n2643), .CP(clk), .Q(r0[26]) );
  DFQD1BWP12T r0_reg_25_ ( .D(n2642), .CP(clk), .Q(r0[25]) );
  DFQD1BWP12T r0_reg_24_ ( .D(n2641), .CP(clk), .Q(r0[24]) );
  DFQD1BWP12T r0_reg_23_ ( .D(n2640), .CP(clk), .Q(r0[23]) );
  DFQD1BWP12T r0_reg_22_ ( .D(n2639), .CP(clk), .Q(r0[22]) );
  DFQD1BWP12T r0_reg_21_ ( .D(n2638), .CP(clk), .Q(r0[21]) );
  DFQD1BWP12T r0_reg_20_ ( .D(n2637), .CP(clk), .Q(r0[20]) );
  DFQD1BWP12T r0_reg_19_ ( .D(n2636), .CP(clk), .Q(r0[19]) );
  DFQD1BWP12T r0_reg_18_ ( .D(n2635), .CP(clk), .Q(r0[18]) );
  DFQD1BWP12T r0_reg_17_ ( .D(n2634), .CP(clk), .Q(r0[17]) );
  DFQD1BWP12T r0_reg_16_ ( .D(n2633), .CP(clk), .Q(r0[16]) );
  DFQD1BWP12T r0_reg_15_ ( .D(n2632), .CP(clk), .Q(r0[15]) );
  DFQD1BWP12T r0_reg_14_ ( .D(n2631), .CP(clk), .Q(r0[14]) );
  DFQD1BWP12T r0_reg_13_ ( .D(n2630), .CP(clk), .Q(r0[13]) );
  DFQD1BWP12T r0_reg_12_ ( .D(n2629), .CP(clk), .Q(r0[12]) );
  DFQD1BWP12T r0_reg_11_ ( .D(n2628), .CP(clk), .Q(r0[11]) );
  DFQD1BWP12T r0_reg_10_ ( .D(n2627), .CP(clk), .Q(r0[10]) );
  DFQD1BWP12T r0_reg_9_ ( .D(n2626), .CP(clk), .Q(r0[9]) );
  DFQD1BWP12T r0_reg_8_ ( .D(n2625), .CP(clk), .Q(r0[8]) );
  DFQD1BWP12T r0_reg_7_ ( .D(n2624), .CP(clk), .Q(r0[7]) );
  DFQD1BWP12T r0_reg_6_ ( .D(n2623), .CP(clk), .Q(r0[6]) );
  DFQD1BWP12T r0_reg_5_ ( .D(n2622), .CP(clk), .Q(r0[5]) );
  DFQD1BWP12T r0_reg_4_ ( .D(n2621), .CP(clk), .Q(r0[4]) );
  DFQD1BWP12T r0_reg_3_ ( .D(n2620), .CP(clk), .Q(r0[3]) );
  DFQD1BWP12T r0_reg_2_ ( .D(n2619), .CP(clk), .Q(r0[2]) );
  DFQD1BWP12T r0_reg_1_ ( .D(n2618), .CP(clk), .Q(r0[1]) );
  DFQD1BWP12T r0_reg_0_ ( .D(n2617), .CP(clk), .Q(r0[0]) );
  DFQD1BWP12T r1_reg_31_ ( .D(n2616), .CP(clk), .Q(r1[31]) );
  DFQD1BWP12T r1_reg_30_ ( .D(n2615), .CP(clk), .Q(r1[30]) );
  DFQD1BWP12T r1_reg_29_ ( .D(n2614), .CP(clk), .Q(r1[29]) );
  DFQD1BWP12T r1_reg_28_ ( .D(n2613), .CP(clk), .Q(r1[28]) );
  DFQD1BWP12T r1_reg_27_ ( .D(n2612), .CP(clk), .Q(r1[27]) );
  DFQD1BWP12T r1_reg_26_ ( .D(n2611), .CP(clk), .Q(r1[26]) );
  DFQD1BWP12T r1_reg_25_ ( .D(n2610), .CP(clk), .Q(r1[25]) );
  DFQD1BWP12T r1_reg_24_ ( .D(n2609), .CP(clk), .Q(r1[24]) );
  DFQD1BWP12T r1_reg_23_ ( .D(n2608), .CP(clk), .Q(r1[23]) );
  DFQD1BWP12T r1_reg_22_ ( .D(n2607), .CP(clk), .Q(r1[22]) );
  DFQD1BWP12T r1_reg_21_ ( .D(n2606), .CP(clk), .Q(r1[21]) );
  DFQD1BWP12T r1_reg_20_ ( .D(n2605), .CP(clk), .Q(r1[20]) );
  DFQD1BWP12T r1_reg_19_ ( .D(n2604), .CP(clk), .Q(r1[19]) );
  DFQD1BWP12T r1_reg_18_ ( .D(n2603), .CP(clk), .Q(r1[18]) );
  DFQD1BWP12T r1_reg_17_ ( .D(n2602), .CP(clk), .Q(r1[17]) );
  DFQD1BWP12T r1_reg_16_ ( .D(n2601), .CP(clk), .Q(r1[16]) );
  DFQD1BWP12T r1_reg_15_ ( .D(n2600), .CP(clk), .Q(r1[15]) );
  DFQD1BWP12T r1_reg_14_ ( .D(n2599), .CP(clk), .Q(r1[14]) );
  DFQD1BWP12T r1_reg_13_ ( .D(n2598), .CP(clk), .Q(r1[13]) );
  DFQD1BWP12T r1_reg_12_ ( .D(n2597), .CP(clk), .Q(r1[12]) );
  DFQD1BWP12T r1_reg_11_ ( .D(n2596), .CP(clk), .Q(r1[11]) );
  DFQD1BWP12T r1_reg_10_ ( .D(n2595), .CP(clk), .Q(r1[10]) );
  DFQD1BWP12T r1_reg_9_ ( .D(n2594), .CP(clk), .Q(r1[9]) );
  DFQD1BWP12T r1_reg_8_ ( .D(n2593), .CP(clk), .Q(r1[8]) );
  DFQD1BWP12T r1_reg_7_ ( .D(n2592), .CP(clk), .Q(r1[7]) );
  DFQD1BWP12T r1_reg_6_ ( .D(n2591), .CP(clk), .Q(r1[6]) );
  DFQD1BWP12T r1_reg_5_ ( .D(n2590), .CP(clk), .Q(r1[5]) );
  DFQD1BWP12T r1_reg_4_ ( .D(n2589), .CP(clk), .Q(r1[4]) );
  DFQD1BWP12T r1_reg_3_ ( .D(n2588), .CP(clk), .Q(r1[3]) );
  DFQD1BWP12T r1_reg_2_ ( .D(n2587), .CP(clk), .Q(r1[2]) );
  DFQD1BWP12T r1_reg_1_ ( .D(n2586), .CP(clk), .Q(r1[1]) );
  DFQD1BWP12T r1_reg_0_ ( .D(n2585), .CP(clk), .Q(r1[0]) );
  DFQD1BWP12T r2_reg_31_ ( .D(n2584), .CP(clk), .Q(r2[31]) );
  DFQD1BWP12T r2_reg_30_ ( .D(n2583), .CP(clk), .Q(r2[30]) );
  DFQD1BWP12T r2_reg_29_ ( .D(n2582), .CP(clk), .Q(r2[29]) );
  DFQD1BWP12T r2_reg_28_ ( .D(n2581), .CP(clk), .Q(r2[28]) );
  DFQD1BWP12T r2_reg_27_ ( .D(n2580), .CP(clk), .Q(r2[27]) );
  DFQD1BWP12T r2_reg_26_ ( .D(n2579), .CP(clk), .Q(r2[26]) );
  DFQD1BWP12T r2_reg_25_ ( .D(n2578), .CP(clk), .Q(r2[25]) );
  DFQD1BWP12T r2_reg_24_ ( .D(n2577), .CP(clk), .Q(r2[24]) );
  DFQD1BWP12T r2_reg_23_ ( .D(n2576), .CP(clk), .Q(r2[23]) );
  DFQD1BWP12T r2_reg_22_ ( .D(n2575), .CP(clk), .Q(r2[22]) );
  DFQD1BWP12T r2_reg_21_ ( .D(n2574), .CP(clk), .Q(r2[21]) );
  DFQD1BWP12T r2_reg_20_ ( .D(n2573), .CP(clk), .Q(r2[20]) );
  DFQD1BWP12T r2_reg_19_ ( .D(n2572), .CP(clk), .Q(r2[19]) );
  DFQD1BWP12T r2_reg_18_ ( .D(n2571), .CP(clk), .Q(r2[18]) );
  DFQD1BWP12T r2_reg_17_ ( .D(n2570), .CP(clk), .Q(r2[17]) );
  DFQD1BWP12T r2_reg_16_ ( .D(n2569), .CP(clk), .Q(r2[16]) );
  DFQD1BWP12T r2_reg_15_ ( .D(n2568), .CP(clk), .Q(r2[15]) );
  DFQD1BWP12T r2_reg_14_ ( .D(n2567), .CP(clk), .Q(r2[14]) );
  DFQD1BWP12T r2_reg_13_ ( .D(n2566), .CP(clk), .Q(r2[13]) );
  DFQD1BWP12T r2_reg_12_ ( .D(n2565), .CP(clk), .Q(r2[12]) );
  DFQD1BWP12T r2_reg_11_ ( .D(n2564), .CP(clk), .Q(r2[11]) );
  DFQD1BWP12T r2_reg_10_ ( .D(n2563), .CP(clk), .Q(r2[10]) );
  DFQD1BWP12T r2_reg_9_ ( .D(n2562), .CP(clk), .Q(r2[9]) );
  DFQD1BWP12T r2_reg_8_ ( .D(n2561), .CP(clk), .Q(r2[8]) );
  DFQD1BWP12T r2_reg_7_ ( .D(n2560), .CP(clk), .Q(r2[7]) );
  DFQD1BWP12T r2_reg_6_ ( .D(n2559), .CP(clk), .Q(r2[6]) );
  DFQD1BWP12T r2_reg_5_ ( .D(n2558), .CP(clk), .Q(r2[5]) );
  DFQD1BWP12T r2_reg_4_ ( .D(n2557), .CP(clk), .Q(r2[4]) );
  DFQD1BWP12T r2_reg_3_ ( .D(n2556), .CP(clk), .Q(r2[3]) );
  DFQD1BWP12T r2_reg_2_ ( .D(n2555), .CP(clk), .Q(r2[2]) );
  DFQD1BWP12T r2_reg_1_ ( .D(n2554), .CP(clk), .Q(r2[1]) );
  DFQD1BWP12T r2_reg_0_ ( .D(n2553), .CP(clk), .Q(r2[0]) );
  DFQD1BWP12T r3_reg_31_ ( .D(n2552), .CP(clk), .Q(r3[31]) );
  DFQD1BWP12T r3_reg_30_ ( .D(n2551), .CP(clk), .Q(r3[30]) );
  DFQD1BWP12T r3_reg_29_ ( .D(n2550), .CP(clk), .Q(r3[29]) );
  DFQD1BWP12T r3_reg_28_ ( .D(n2549), .CP(clk), .Q(r3[28]) );
  DFQD1BWP12T r3_reg_27_ ( .D(n2548), .CP(clk), .Q(r3[27]) );
  DFQD1BWP12T r3_reg_26_ ( .D(n2547), .CP(clk), .Q(r3[26]) );
  DFQD1BWP12T r3_reg_25_ ( .D(n2546), .CP(clk), .Q(r3[25]) );
  DFQD1BWP12T r3_reg_24_ ( .D(n2545), .CP(clk), .Q(r3[24]) );
  DFQD1BWP12T r3_reg_23_ ( .D(n2544), .CP(clk), .Q(r3[23]) );
  DFQD1BWP12T r3_reg_22_ ( .D(n2543), .CP(clk), .Q(r3[22]) );
  DFQD1BWP12T r3_reg_21_ ( .D(n2542), .CP(clk), .Q(r3[21]) );
  DFQD1BWP12T r3_reg_20_ ( .D(n2541), .CP(clk), .Q(r3[20]) );
  DFQD1BWP12T r3_reg_19_ ( .D(n2540), .CP(clk), .Q(r3[19]) );
  DFQD1BWP12T r3_reg_18_ ( .D(n2539), .CP(clk), .Q(r3[18]) );
  DFQD1BWP12T r3_reg_17_ ( .D(n2538), .CP(clk), .Q(r3[17]) );
  DFQD1BWP12T r3_reg_16_ ( .D(n2537), .CP(clk), .Q(r3[16]) );
  DFQD1BWP12T r3_reg_15_ ( .D(n2536), .CP(clk), .Q(r3[15]) );
  DFQD1BWP12T r3_reg_14_ ( .D(n2535), .CP(clk), .Q(r3[14]) );
  DFQD1BWP12T r3_reg_13_ ( .D(n2534), .CP(clk), .Q(r3[13]) );
  DFQD1BWP12T r3_reg_12_ ( .D(n2533), .CP(clk), .Q(r3[12]) );
  DFQD1BWP12T r3_reg_11_ ( .D(n2532), .CP(clk), .Q(r3[11]) );
  DFQD1BWP12T r3_reg_10_ ( .D(n2531), .CP(clk), .Q(r3[10]) );
  DFQD1BWP12T r3_reg_9_ ( .D(n2530), .CP(clk), .Q(r3[9]) );
  DFQD1BWP12T r3_reg_8_ ( .D(n2529), .CP(clk), .Q(r3[8]) );
  DFQD1BWP12T r3_reg_7_ ( .D(n2528), .CP(clk), .Q(r3[7]) );
  DFQD1BWP12T r3_reg_6_ ( .D(n2527), .CP(clk), .Q(r3[6]) );
  DFQD1BWP12T r3_reg_5_ ( .D(n2526), .CP(clk), .Q(r3[5]) );
  DFQD1BWP12T r3_reg_4_ ( .D(n2525), .CP(clk), .Q(r3[4]) );
  DFQD1BWP12T r3_reg_3_ ( .D(n2524), .CP(clk), .Q(r3[3]) );
  DFQD1BWP12T r3_reg_2_ ( .D(n2523), .CP(clk), .Q(r3[2]) );
  DFQD1BWP12T r3_reg_1_ ( .D(n2522), .CP(clk), .Q(r3[1]) );
  DFQD1BWP12T r3_reg_0_ ( .D(n2521), .CP(clk), .Q(r3[0]) );
  DFQD1BWP12T r4_reg_31_ ( .D(n2520), .CP(clk), .Q(r4[31]) );
  DFQD1BWP12T r4_reg_30_ ( .D(n2519), .CP(clk), .Q(r4[30]) );
  DFQD1BWP12T r4_reg_29_ ( .D(n2518), .CP(clk), .Q(r4[29]) );
  DFQD1BWP12T r4_reg_28_ ( .D(n2517), .CP(clk), .Q(r4[28]) );
  DFQD1BWP12T r4_reg_27_ ( .D(n2516), .CP(clk), .Q(r4[27]) );
  DFQD1BWP12T r4_reg_26_ ( .D(n2515), .CP(clk), .Q(r4[26]) );
  DFQD1BWP12T r4_reg_25_ ( .D(n2514), .CP(clk), .Q(r4[25]) );
  DFQD1BWP12T r4_reg_24_ ( .D(n2513), .CP(clk), .Q(r4[24]) );
  DFQD1BWP12T r4_reg_23_ ( .D(n2512), .CP(clk), .Q(r4[23]) );
  DFQD1BWP12T r4_reg_22_ ( .D(n2511), .CP(clk), .Q(r4[22]) );
  DFQD1BWP12T r4_reg_21_ ( .D(n2510), .CP(clk), .Q(r4[21]) );
  DFQD1BWP12T r4_reg_20_ ( .D(n2509), .CP(clk), .Q(r4[20]) );
  DFQD1BWP12T r4_reg_19_ ( .D(n2508), .CP(clk), .Q(r4[19]) );
  DFQD1BWP12T r4_reg_18_ ( .D(n2507), .CP(clk), .Q(r4[18]) );
  DFQD1BWP12T r4_reg_17_ ( .D(n2506), .CP(clk), .Q(r4[17]) );
  DFQD1BWP12T r4_reg_16_ ( .D(n2505), .CP(clk), .Q(r4[16]) );
  DFQD1BWP12T r4_reg_15_ ( .D(n2504), .CP(clk), .Q(r4[15]) );
  DFQD1BWP12T r4_reg_14_ ( .D(n2503), .CP(clk), .Q(r4[14]) );
  DFQD1BWP12T r4_reg_13_ ( .D(n2502), .CP(clk), .Q(r4[13]) );
  DFQD1BWP12T r4_reg_12_ ( .D(n2501), .CP(clk), .Q(r4[12]) );
  DFQD1BWP12T r4_reg_11_ ( .D(n2500), .CP(clk), .Q(r4[11]) );
  DFQD1BWP12T r4_reg_10_ ( .D(n2499), .CP(clk), .Q(r4[10]) );
  DFQD1BWP12T r4_reg_9_ ( .D(n2498), .CP(clk), .Q(r4[9]) );
  DFQD1BWP12T r4_reg_8_ ( .D(n2497), .CP(clk), .Q(r4[8]) );
  DFQD1BWP12T r4_reg_7_ ( .D(n2496), .CP(clk), .Q(r4[7]) );
  DFQD1BWP12T r4_reg_6_ ( .D(n2495), .CP(clk), .Q(r4[6]) );
  DFQD1BWP12T r4_reg_5_ ( .D(n2494), .CP(clk), .Q(r4[5]) );
  DFQD1BWP12T r4_reg_4_ ( .D(n2493), .CP(clk), .Q(r4[4]) );
  DFQD1BWP12T r4_reg_3_ ( .D(n2492), .CP(clk), .Q(r4[3]) );
  DFQD1BWP12T r4_reg_2_ ( .D(n2491), .CP(clk), .Q(r4[2]) );
  DFQD1BWP12T r4_reg_1_ ( .D(n2490), .CP(clk), .Q(r4[1]) );
  DFQD1BWP12T r4_reg_0_ ( .D(n2489), .CP(clk), .Q(r4[0]) );
  DFQD1BWP12T r5_reg_31_ ( .D(n2488), .CP(clk), .Q(r5[31]) );
  DFQD1BWP12T r5_reg_30_ ( .D(n2487), .CP(clk), .Q(r5[30]) );
  DFQD1BWP12T r5_reg_29_ ( .D(n2486), .CP(clk), .Q(r5[29]) );
  DFQD1BWP12T r5_reg_28_ ( .D(n2485), .CP(clk), .Q(r5[28]) );
  DFQD1BWP12T r5_reg_27_ ( .D(n2484), .CP(clk), .Q(r5[27]) );
  DFQD1BWP12T r5_reg_26_ ( .D(n2483), .CP(clk), .Q(r5[26]) );
  DFQD1BWP12T r5_reg_25_ ( .D(n2482), .CP(clk), .Q(r5[25]) );
  DFQD1BWP12T r5_reg_24_ ( .D(n2481), .CP(clk), .Q(r5[24]) );
  DFQD1BWP12T r5_reg_23_ ( .D(n2480), .CP(clk), .Q(r5[23]) );
  DFQD1BWP12T r5_reg_22_ ( .D(n2479), .CP(clk), .Q(r5[22]) );
  DFQD1BWP12T r5_reg_21_ ( .D(n2478), .CP(clk), .Q(r5[21]) );
  DFQD1BWP12T r5_reg_20_ ( .D(n2477), .CP(clk), .Q(r5[20]) );
  DFQD1BWP12T r5_reg_19_ ( .D(n2476), .CP(clk), .Q(r5[19]) );
  DFQD1BWP12T r5_reg_18_ ( .D(n2475), .CP(clk), .Q(r5[18]) );
  DFQD1BWP12T r5_reg_17_ ( .D(n2474), .CP(clk), .Q(r5[17]) );
  DFQD1BWP12T r5_reg_16_ ( .D(n2473), .CP(clk), .Q(r5[16]) );
  DFQD1BWP12T r5_reg_15_ ( .D(n2472), .CP(clk), .Q(r5[15]) );
  DFQD1BWP12T r5_reg_14_ ( .D(n2471), .CP(clk), .Q(r5[14]) );
  DFQD1BWP12T r5_reg_13_ ( .D(n2470), .CP(clk), .Q(r5[13]) );
  DFQD1BWP12T r5_reg_12_ ( .D(n2469), .CP(clk), .Q(r5[12]) );
  DFQD1BWP12T r5_reg_11_ ( .D(n2468), .CP(clk), .Q(r5[11]) );
  DFQD1BWP12T r5_reg_10_ ( .D(n2467), .CP(clk), .Q(r5[10]) );
  DFQD1BWP12T r5_reg_9_ ( .D(n2466), .CP(clk), .Q(r5[9]) );
  DFQD1BWP12T r5_reg_8_ ( .D(n2465), .CP(clk), .Q(r5[8]) );
  DFQD1BWP12T r5_reg_7_ ( .D(n2464), .CP(clk), .Q(r5[7]) );
  DFQD1BWP12T r5_reg_6_ ( .D(n2463), .CP(clk), .Q(r5[6]) );
  DFQD1BWP12T r5_reg_5_ ( .D(n2462), .CP(clk), .Q(r5[5]) );
  DFQD1BWP12T r5_reg_4_ ( .D(n2461), .CP(clk), .Q(r5[4]) );
  DFQD1BWP12T r5_reg_3_ ( .D(n2460), .CP(clk), .Q(r5[3]) );
  DFQD1BWP12T r5_reg_2_ ( .D(n2459), .CP(clk), .Q(r5[2]) );
  DFQD1BWP12T r5_reg_1_ ( .D(n2458), .CP(clk), .Q(r5[1]) );
  DFQD1BWP12T r5_reg_0_ ( .D(n2457), .CP(clk), .Q(r5[0]) );
  DFQD1BWP12T r6_reg_31_ ( .D(n2456), .CP(clk), .Q(r6[31]) );
  DFQD1BWP12T r6_reg_30_ ( .D(n2455), .CP(clk), .Q(r6[30]) );
  DFQD1BWP12T r6_reg_29_ ( .D(n2454), .CP(clk), .Q(r6[29]) );
  DFQD1BWP12T r6_reg_28_ ( .D(n2453), .CP(clk), .Q(r6[28]) );
  DFQD1BWP12T r6_reg_27_ ( .D(n2452), .CP(clk), .Q(r6[27]) );
  DFQD1BWP12T r6_reg_26_ ( .D(n2451), .CP(clk), .Q(r6[26]) );
  DFQD1BWP12T r6_reg_25_ ( .D(n2450), .CP(clk), .Q(r6[25]) );
  DFQD1BWP12T r6_reg_24_ ( .D(n2449), .CP(clk), .Q(r6[24]) );
  DFQD1BWP12T r6_reg_23_ ( .D(n2448), .CP(clk), .Q(r6[23]) );
  DFQD1BWP12T r6_reg_22_ ( .D(n2447), .CP(clk), .Q(r6[22]) );
  DFQD1BWP12T r6_reg_21_ ( .D(n2446), .CP(clk), .Q(r6[21]) );
  DFQD1BWP12T r6_reg_20_ ( .D(n2445), .CP(clk), .Q(r6[20]) );
  DFQD1BWP12T r6_reg_19_ ( .D(n2444), .CP(clk), .Q(r6[19]) );
  DFQD1BWP12T r6_reg_18_ ( .D(n2443), .CP(clk), .Q(r6[18]) );
  DFQD1BWP12T r6_reg_17_ ( .D(n2442), .CP(clk), .Q(r6[17]) );
  DFQD1BWP12T r6_reg_16_ ( .D(n2441), .CP(clk), .Q(r6[16]) );
  DFQD1BWP12T r6_reg_15_ ( .D(n2440), .CP(clk), .Q(r6[15]) );
  DFQD1BWP12T r6_reg_14_ ( .D(n2439), .CP(clk), .Q(r6[14]) );
  DFQD1BWP12T r6_reg_13_ ( .D(n2438), .CP(clk), .Q(r6[13]) );
  DFQD1BWP12T r6_reg_12_ ( .D(n2437), .CP(clk), .Q(r6[12]) );
  DFQD1BWP12T r6_reg_11_ ( .D(n2436), .CP(clk), .Q(r6[11]) );
  DFQD1BWP12T r6_reg_10_ ( .D(n2435), .CP(clk), .Q(r6[10]) );
  DFQD1BWP12T r6_reg_9_ ( .D(n2434), .CP(clk), .Q(r6[9]) );
  DFQD1BWP12T r6_reg_8_ ( .D(n2433), .CP(clk), .Q(r6[8]) );
  DFQD1BWP12T r6_reg_7_ ( .D(n2432), .CP(clk), .Q(r6[7]) );
  DFQD1BWP12T r6_reg_6_ ( .D(n2431), .CP(clk), .Q(r6[6]) );
  DFQD1BWP12T r6_reg_5_ ( .D(n2430), .CP(clk), .Q(r6[5]) );
  DFQD1BWP12T r6_reg_4_ ( .D(n2429), .CP(clk), .Q(r6[4]) );
  DFQD1BWP12T r6_reg_3_ ( .D(n2428), .CP(clk), .Q(r6[3]) );
  DFQD1BWP12T r6_reg_2_ ( .D(n2427), .CP(clk), .Q(r6[2]) );
  DFQD1BWP12T r6_reg_1_ ( .D(n2426), .CP(clk), .Q(r6[1]) );
  DFQD1BWP12T r6_reg_0_ ( .D(n2425), .CP(clk), .Q(r6[0]) );
  DFQD1BWP12T r7_reg_31_ ( .D(n2424), .CP(clk), .Q(r7[31]) );
  DFQD1BWP12T r7_reg_30_ ( .D(n2423), .CP(clk), .Q(r7[30]) );
  DFQD1BWP12T r7_reg_29_ ( .D(n2422), .CP(clk), .Q(r7[29]) );
  DFQD1BWP12T r7_reg_28_ ( .D(n2421), .CP(clk), .Q(r7[28]) );
  DFQD1BWP12T r7_reg_27_ ( .D(n2420), .CP(clk), .Q(r7[27]) );
  DFQD1BWP12T r7_reg_26_ ( .D(n2419), .CP(clk), .Q(r7[26]) );
  DFQD1BWP12T r7_reg_25_ ( .D(n2418), .CP(clk), .Q(r7[25]) );
  DFQD1BWP12T r7_reg_24_ ( .D(n2417), .CP(clk), .Q(r7[24]) );
  DFQD1BWP12T r7_reg_23_ ( .D(n2416), .CP(clk), .Q(r7[23]) );
  DFQD1BWP12T r7_reg_22_ ( .D(n2415), .CP(clk), .Q(r7[22]) );
  DFQD1BWP12T r7_reg_21_ ( .D(n2414), .CP(clk), .Q(r7[21]) );
  DFQD1BWP12T r7_reg_20_ ( .D(n2413), .CP(clk), .Q(r7[20]) );
  DFQD1BWP12T r7_reg_19_ ( .D(n2412), .CP(clk), .Q(r7[19]) );
  DFQD1BWP12T r7_reg_18_ ( .D(n2411), .CP(clk), .Q(r7[18]) );
  DFQD1BWP12T r7_reg_17_ ( .D(n2410), .CP(clk), .Q(r7[17]) );
  DFQD1BWP12T r7_reg_16_ ( .D(n2409), .CP(clk), .Q(r7[16]) );
  DFQD1BWP12T r7_reg_15_ ( .D(n2408), .CP(clk), .Q(r7[15]) );
  DFQD1BWP12T r7_reg_14_ ( .D(n2407), .CP(clk), .Q(r7[14]) );
  DFQD1BWP12T r7_reg_13_ ( .D(n2406), .CP(clk), .Q(r7[13]) );
  DFQD1BWP12T r7_reg_12_ ( .D(n2405), .CP(clk), .Q(r7[12]) );
  DFQD1BWP12T r7_reg_11_ ( .D(n2404), .CP(clk), .Q(r7[11]) );
  DFQD1BWP12T r7_reg_10_ ( .D(n2403), .CP(clk), .Q(r7[10]) );
  DFQD1BWP12T r7_reg_9_ ( .D(n2402), .CP(clk), .Q(r7[9]) );
  DFQD1BWP12T r7_reg_8_ ( .D(n2401), .CP(clk), .Q(r7[8]) );
  DFQD1BWP12T r7_reg_7_ ( .D(n2400), .CP(clk), .Q(r7[7]) );
  DFQD1BWP12T r7_reg_6_ ( .D(n2399), .CP(clk), .Q(r7[6]) );
  DFQD1BWP12T r7_reg_5_ ( .D(n2398), .CP(clk), .Q(r7[5]) );
  DFQD1BWP12T r7_reg_4_ ( .D(n2397), .CP(clk), .Q(r7[4]) );
  DFQD1BWP12T r7_reg_3_ ( .D(n2396), .CP(clk), .Q(r7[3]) );
  DFQD1BWP12T r7_reg_2_ ( .D(n2395), .CP(clk), .Q(r7[2]) );
  DFQD1BWP12T r7_reg_1_ ( .D(n2394), .CP(clk), .Q(r7[1]) );
  DFQD1BWP12T r7_reg_0_ ( .D(n2393), .CP(clk), .Q(r7[0]) );
  DFQD1BWP12T r8_reg_31_ ( .D(n2392), .CP(clk), .Q(r8[31]) );
  DFQD1BWP12T r8_reg_30_ ( .D(n2391), .CP(clk), .Q(r8[30]) );
  DFQD1BWP12T r8_reg_29_ ( .D(n2390), .CP(clk), .Q(r8[29]) );
  DFQD1BWP12T r8_reg_28_ ( .D(n2389), .CP(clk), .Q(r8[28]) );
  DFQD1BWP12T r8_reg_27_ ( .D(n2388), .CP(clk), .Q(r8[27]) );
  DFQD1BWP12T r8_reg_26_ ( .D(n2387), .CP(clk), .Q(r8[26]) );
  DFQD1BWP12T r8_reg_25_ ( .D(n2386), .CP(clk), .Q(r8[25]) );
  DFQD1BWP12T r8_reg_24_ ( .D(n2385), .CP(clk), .Q(r8[24]) );
  DFQD1BWP12T r8_reg_23_ ( .D(n2384), .CP(clk), .Q(r8[23]) );
  DFQD1BWP12T r8_reg_22_ ( .D(n2383), .CP(clk), .Q(r8[22]) );
  DFQD1BWP12T r8_reg_21_ ( .D(n2382), .CP(clk), .Q(r8[21]) );
  DFQD1BWP12T r8_reg_20_ ( .D(n2381), .CP(clk), .Q(r8[20]) );
  DFQD1BWP12T r8_reg_19_ ( .D(n2380), .CP(clk), .Q(r8[19]) );
  DFQD1BWP12T r8_reg_18_ ( .D(n2379), .CP(clk), .Q(r8[18]) );
  DFQD1BWP12T r8_reg_17_ ( .D(n2378), .CP(clk), .Q(r8[17]) );
  DFQD1BWP12T r8_reg_16_ ( .D(n2377), .CP(clk), .Q(r8[16]) );
  DFQD1BWP12T r8_reg_15_ ( .D(n2376), .CP(clk), .Q(r8[15]) );
  DFQD1BWP12T r8_reg_14_ ( .D(n2375), .CP(clk), .Q(r8[14]) );
  DFQD1BWP12T r8_reg_13_ ( .D(n2374), .CP(clk), .Q(r8[13]) );
  DFQD1BWP12T r8_reg_12_ ( .D(n2373), .CP(clk), .Q(r8[12]) );
  DFQD1BWP12T r8_reg_11_ ( .D(n2372), .CP(clk), .Q(r8[11]) );
  DFQD1BWP12T r8_reg_10_ ( .D(n2371), .CP(clk), .Q(r8[10]) );
  DFQD1BWP12T r8_reg_9_ ( .D(n2370), .CP(clk), .Q(r8[9]) );
  DFQD1BWP12T r8_reg_8_ ( .D(n2369), .CP(clk), .Q(r8[8]) );
  DFQD1BWP12T r8_reg_7_ ( .D(n2368), .CP(clk), .Q(r8[7]) );
  DFQD1BWP12T r8_reg_6_ ( .D(n2367), .CP(clk), .Q(r8[6]) );
  DFQD1BWP12T r8_reg_5_ ( .D(n2366), .CP(clk), .Q(r8[5]) );
  DFQD1BWP12T r8_reg_4_ ( .D(n2365), .CP(clk), .Q(r8[4]) );
  DFQD1BWP12T r8_reg_3_ ( .D(n2364), .CP(clk), .Q(r8[3]) );
  DFQD1BWP12T r8_reg_2_ ( .D(n2363), .CP(clk), .Q(r8[2]) );
  DFQD1BWP12T r8_reg_1_ ( .D(n2362), .CP(clk), .Q(r8[1]) );
  DFQD1BWP12T r8_reg_0_ ( .D(n2361), .CP(clk), .Q(r8[0]) );
  DFQD1BWP12T r9_reg_31_ ( .D(n2360), .CP(clk), .Q(r9[31]) );
  DFQD1BWP12T r9_reg_30_ ( .D(n2359), .CP(clk), .Q(r9[30]) );
  DFQD1BWP12T r9_reg_29_ ( .D(n2358), .CP(clk), .Q(r9[29]) );
  DFQD1BWP12T r9_reg_28_ ( .D(n2357), .CP(clk), .Q(r9[28]) );
  DFQD1BWP12T r9_reg_27_ ( .D(n2356), .CP(clk), .Q(r9[27]) );
  DFQD1BWP12T r9_reg_26_ ( .D(n2355), .CP(clk), .Q(r9[26]) );
  DFQD1BWP12T r9_reg_25_ ( .D(n2354), .CP(clk), .Q(r9[25]) );
  DFQD1BWP12T r9_reg_24_ ( .D(n2353), .CP(clk), .Q(r9[24]) );
  DFQD1BWP12T r9_reg_23_ ( .D(n2352), .CP(clk), .Q(r9[23]) );
  DFQD1BWP12T r9_reg_22_ ( .D(n2351), .CP(clk), .Q(r9[22]) );
  DFQD1BWP12T r9_reg_21_ ( .D(n2350), .CP(clk), .Q(r9[21]) );
  DFQD1BWP12T r9_reg_20_ ( .D(n2349), .CP(clk), .Q(r9[20]) );
  DFQD1BWP12T r9_reg_19_ ( .D(n2348), .CP(clk), .Q(r9[19]) );
  DFQD1BWP12T r9_reg_18_ ( .D(n2347), .CP(clk), .Q(r9[18]) );
  DFQD1BWP12T r9_reg_17_ ( .D(n2346), .CP(clk), .Q(r9[17]) );
  DFQD1BWP12T r9_reg_16_ ( .D(n2345), .CP(clk), .Q(r9[16]) );
  DFQD1BWP12T r9_reg_15_ ( .D(n2344), .CP(clk), .Q(r9[15]) );
  DFQD1BWP12T r9_reg_14_ ( .D(n2343), .CP(clk), .Q(r9[14]) );
  DFQD1BWP12T r9_reg_13_ ( .D(n2342), .CP(clk), .Q(r9[13]) );
  DFQD1BWP12T r9_reg_12_ ( .D(n2341), .CP(clk), .Q(r9[12]) );
  DFQD1BWP12T r9_reg_11_ ( .D(n2340), .CP(clk), .Q(r9[11]) );
  DFQD1BWP12T r9_reg_10_ ( .D(n2339), .CP(clk), .Q(r9[10]) );
  DFQD1BWP12T r9_reg_9_ ( .D(n2338), .CP(clk), .Q(r9[9]) );
  DFQD1BWP12T r9_reg_8_ ( .D(n2337), .CP(clk), .Q(r9[8]) );
  DFQD1BWP12T r9_reg_7_ ( .D(n2336), .CP(clk), .Q(r9[7]) );
  DFQD1BWP12T r9_reg_6_ ( .D(n2335), .CP(clk), .Q(r9[6]) );
  DFQD1BWP12T r9_reg_5_ ( .D(n2334), .CP(clk), .Q(r9[5]) );
  DFQD1BWP12T r9_reg_4_ ( .D(n2333), .CP(clk), .Q(r9[4]) );
  DFQD1BWP12T r9_reg_3_ ( .D(n2332), .CP(clk), .Q(r9[3]) );
  DFQD1BWP12T r9_reg_2_ ( .D(n2331), .CP(clk), .Q(r9[2]) );
  DFQD1BWP12T r9_reg_1_ ( .D(n2330), .CP(clk), .Q(r9[1]) );
  DFQD1BWP12T r9_reg_0_ ( .D(n2329), .CP(clk), .Q(r9[0]) );
  DFQD1BWP12T r10_reg_31_ ( .D(n2328), .CP(clk), .Q(r10[31]) );
  DFQD1BWP12T r10_reg_30_ ( .D(n2327), .CP(clk), .Q(r10[30]) );
  DFQD1BWP12T r10_reg_29_ ( .D(n2326), .CP(clk), .Q(r10[29]) );
  DFQD1BWP12T r10_reg_28_ ( .D(n2325), .CP(clk), .Q(r10[28]) );
  DFQD1BWP12T r10_reg_27_ ( .D(n2324), .CP(clk), .Q(r10[27]) );
  DFQD1BWP12T r10_reg_26_ ( .D(n2323), .CP(clk), .Q(r10[26]) );
  DFQD1BWP12T r10_reg_25_ ( .D(n2322), .CP(clk), .Q(r10[25]) );
  DFQD1BWP12T r10_reg_24_ ( .D(n2321), .CP(clk), .Q(r10[24]) );
  DFQD1BWP12T r10_reg_23_ ( .D(n2320), .CP(clk), .Q(r10[23]) );
  DFQD1BWP12T r10_reg_22_ ( .D(n2319), .CP(clk), .Q(r10[22]) );
  DFQD1BWP12T r10_reg_21_ ( .D(n2318), .CP(clk), .Q(r10[21]) );
  DFQD1BWP12T r10_reg_20_ ( .D(n2317), .CP(clk), .Q(r10[20]) );
  DFQD1BWP12T r10_reg_19_ ( .D(n2316), .CP(clk), .Q(r10[19]) );
  DFQD1BWP12T r10_reg_18_ ( .D(n2315), .CP(clk), .Q(r10[18]) );
  DFQD1BWP12T r10_reg_17_ ( .D(n2314), .CP(clk), .Q(r10[17]) );
  DFQD1BWP12T r10_reg_16_ ( .D(n2313), .CP(clk), .Q(r10[16]) );
  DFQD1BWP12T r10_reg_15_ ( .D(n2312), .CP(clk), .Q(r10[15]) );
  DFQD1BWP12T r10_reg_14_ ( .D(n2311), .CP(clk), .Q(r10[14]) );
  DFQD1BWP12T r10_reg_13_ ( .D(n2310), .CP(clk), .Q(r10[13]) );
  DFQD1BWP12T r10_reg_12_ ( .D(n2309), .CP(clk), .Q(r10[12]) );
  DFQD1BWP12T r10_reg_11_ ( .D(n2308), .CP(clk), .Q(r10[11]) );
  DFQD1BWP12T r10_reg_10_ ( .D(n2307), .CP(clk), .Q(r10[10]) );
  DFQD1BWP12T r10_reg_9_ ( .D(n2306), .CP(clk), .Q(r10[9]) );
  DFQD1BWP12T r10_reg_8_ ( .D(n2305), .CP(clk), .Q(r10[8]) );
  DFQD1BWP12T r10_reg_7_ ( .D(n2304), .CP(clk), .Q(r10[7]) );
  DFQD1BWP12T r10_reg_6_ ( .D(n2303), .CP(clk), .Q(r10[6]) );
  DFQD1BWP12T r10_reg_5_ ( .D(n2302), .CP(clk), .Q(r10[5]) );
  DFQD1BWP12T r10_reg_4_ ( .D(n2301), .CP(clk), .Q(r10[4]) );
  DFQD1BWP12T r10_reg_3_ ( .D(n2300), .CP(clk), .Q(r10[3]) );
  DFQD1BWP12T r10_reg_2_ ( .D(n2299), .CP(clk), .Q(r10[2]) );
  DFQD1BWP12T r10_reg_1_ ( .D(n2298), .CP(clk), .Q(r10[1]) );
  DFQD1BWP12T r10_reg_0_ ( .D(n2297), .CP(clk), .Q(r10[0]) );
  DFQD1BWP12T r11_reg_31_ ( .D(n2296), .CP(clk), .Q(r11[31]) );
  DFQD1BWP12T r11_reg_30_ ( .D(n2295), .CP(clk), .Q(r11[30]) );
  DFQD1BWP12T r11_reg_29_ ( .D(n2294), .CP(clk), .Q(r11[29]) );
  DFQD1BWP12T r11_reg_28_ ( .D(n2293), .CP(clk), .Q(r11[28]) );
  DFQD1BWP12T r11_reg_27_ ( .D(n2292), .CP(clk), .Q(r11[27]) );
  DFQD1BWP12T r11_reg_26_ ( .D(n2291), .CP(clk), .Q(r11[26]) );
  DFQD1BWP12T r11_reg_25_ ( .D(n2290), .CP(clk), .Q(r11[25]) );
  DFQD1BWP12T r11_reg_24_ ( .D(n2289), .CP(clk), .Q(r11[24]) );
  DFQD1BWP12T r11_reg_23_ ( .D(n2288), .CP(clk), .Q(r11[23]) );
  DFQD1BWP12T r11_reg_22_ ( .D(n2287), .CP(clk), .Q(r11[22]) );
  DFQD1BWP12T r11_reg_21_ ( .D(n2286), .CP(clk), .Q(r11[21]) );
  DFQD1BWP12T r11_reg_20_ ( .D(n2285), .CP(clk), .Q(r11[20]) );
  DFQD1BWP12T r11_reg_19_ ( .D(n2284), .CP(clk), .Q(r11[19]) );
  DFQD1BWP12T r11_reg_18_ ( .D(n2283), .CP(clk), .Q(r11[18]) );
  DFQD1BWP12T r11_reg_17_ ( .D(n2282), .CP(clk), .Q(r11[17]) );
  DFQD1BWP12T r11_reg_16_ ( .D(n2281), .CP(clk), .Q(r11[16]) );
  DFQD1BWP12T r11_reg_15_ ( .D(n2280), .CP(clk), .Q(r11[15]) );
  DFQD1BWP12T r11_reg_14_ ( .D(n2279), .CP(clk), .Q(r11[14]) );
  DFQD1BWP12T r11_reg_13_ ( .D(n2278), .CP(clk), .Q(r11[13]) );
  DFQD1BWP12T r11_reg_12_ ( .D(n2277), .CP(clk), .Q(r11[12]) );
  DFQD1BWP12T r11_reg_11_ ( .D(n2276), .CP(clk), .Q(r11[11]) );
  DFQD1BWP12T r11_reg_10_ ( .D(n2275), .CP(clk), .Q(r11[10]) );
  DFQD1BWP12T r11_reg_9_ ( .D(n2274), .CP(clk), .Q(r11[9]) );
  DFQD1BWP12T r11_reg_8_ ( .D(n2273), .CP(clk), .Q(r11[8]) );
  DFQD1BWP12T r11_reg_7_ ( .D(n2272), .CP(clk), .Q(r11[7]) );
  DFQD1BWP12T r11_reg_6_ ( .D(n2271), .CP(clk), .Q(r11[6]) );
  DFQD1BWP12T r11_reg_5_ ( .D(n2270), .CP(clk), .Q(r11[5]) );
  DFQD1BWP12T r11_reg_4_ ( .D(n2269), .CP(clk), .Q(r11[4]) );
  DFQD1BWP12T r11_reg_3_ ( .D(n2268), .CP(clk), .Q(r11[3]) );
  DFQD1BWP12T r11_reg_2_ ( .D(n2267), .CP(clk), .Q(r11[2]) );
  DFQD1BWP12T r11_reg_1_ ( .D(n2266), .CP(clk), .Q(r11[1]) );
  DFQD1BWP12T r11_reg_0_ ( .D(n2265), .CP(clk), .Q(r11[0]) );
  DFQD1BWP12T r12_reg_31_ ( .D(n2264), .CP(clk), .Q(r12[31]) );
  DFQD1BWP12T r12_reg_30_ ( .D(n2263), .CP(clk), .Q(r12[30]) );
  DFQD1BWP12T r12_reg_29_ ( .D(n2262), .CP(clk), .Q(r12[29]) );
  DFQD1BWP12T r12_reg_28_ ( .D(n2261), .CP(clk), .Q(r12[28]) );
  DFQD1BWP12T r12_reg_27_ ( .D(n2260), .CP(clk), .Q(r12[27]) );
  DFQD1BWP12T r12_reg_26_ ( .D(n2259), .CP(clk), .Q(r12[26]) );
  DFQD1BWP12T r12_reg_25_ ( .D(n2258), .CP(clk), .Q(r12[25]) );
  DFQD1BWP12T r12_reg_24_ ( .D(n2257), .CP(clk), .Q(r12[24]) );
  DFQD1BWP12T r12_reg_23_ ( .D(n2256), .CP(clk), .Q(r12[23]) );
  DFQD1BWP12T r12_reg_22_ ( .D(n2255), .CP(clk), .Q(r12[22]) );
  DFQD1BWP12T r12_reg_21_ ( .D(n2254), .CP(clk), .Q(r12[21]) );
  DFQD1BWP12T r12_reg_20_ ( .D(n2253), .CP(clk), .Q(r12[20]) );
  DFQD1BWP12T r12_reg_19_ ( .D(n2252), .CP(clk), .Q(r12[19]) );
  DFQD1BWP12T r12_reg_18_ ( .D(n2251), .CP(clk), .Q(r12[18]) );
  DFQD1BWP12T r12_reg_17_ ( .D(n2250), .CP(clk), .Q(r12[17]) );
  DFQD1BWP12T r12_reg_16_ ( .D(n2249), .CP(clk), .Q(r12[16]) );
  DFQD1BWP12T r12_reg_15_ ( .D(n2248), .CP(clk), .Q(r12[15]) );
  DFQD1BWP12T r12_reg_14_ ( .D(n2247), .CP(clk), .Q(r12[14]) );
  DFQD1BWP12T r12_reg_13_ ( .D(n2246), .CP(clk), .Q(r12[13]) );
  DFQD1BWP12T r12_reg_12_ ( .D(n2245), .CP(clk), .Q(r12[12]) );
  DFQD1BWP12T r12_reg_11_ ( .D(n2244), .CP(clk), .Q(r12[11]) );
  DFQD1BWP12T r12_reg_10_ ( .D(n2243), .CP(clk), .Q(r12[10]) );
  DFQD1BWP12T r12_reg_9_ ( .D(n2242), .CP(clk), .Q(r12[9]) );
  DFQD1BWP12T r12_reg_8_ ( .D(n2241), .CP(clk), .Q(r12[8]) );
  DFQD1BWP12T r12_reg_7_ ( .D(n2240), .CP(clk), .Q(r12[7]) );
  DFQD1BWP12T r12_reg_6_ ( .D(n2239), .CP(clk), .Q(r12[6]) );
  DFQD1BWP12T r12_reg_5_ ( .D(n2238), .CP(clk), .Q(r12[5]) );
  DFQD1BWP12T r12_reg_4_ ( .D(n2237), .CP(clk), .Q(r12[4]) );
  DFQD1BWP12T r12_reg_3_ ( .D(n2236), .CP(clk), .Q(r12[3]) );
  DFQD1BWP12T r12_reg_2_ ( .D(n2235), .CP(clk), .Q(r12[2]) );
  DFQD1BWP12T r12_reg_1_ ( .D(n2234), .CP(clk), .Q(r12[1]) );
  DFQD1BWP12T r12_reg_0_ ( .D(n2233), .CP(clk), .Q(r12[0]) );
  DFQD1BWP12T lr_reg_31_ ( .D(n2232), .CP(clk), .Q(lr[31]) );
  DFQD1BWP12T lr_reg_30_ ( .D(n2231), .CP(clk), .Q(lr[30]) );
  DFQD1BWP12T lr_reg_29_ ( .D(n2230), .CP(clk), .Q(lr[29]) );
  DFQD1BWP12T lr_reg_28_ ( .D(n2229), .CP(clk), .Q(lr[28]) );
  DFQD1BWP12T lr_reg_27_ ( .D(n2228), .CP(clk), .Q(lr[27]) );
  DFQD1BWP12T lr_reg_26_ ( .D(n2227), .CP(clk), .Q(lr[26]) );
  DFQD1BWP12T lr_reg_25_ ( .D(n2226), .CP(clk), .Q(lr[25]) );
  DFQD1BWP12T lr_reg_24_ ( .D(n2225), .CP(clk), .Q(lr[24]) );
  DFQD1BWP12T lr_reg_23_ ( .D(n2224), .CP(clk), .Q(lr[23]) );
  DFQD1BWP12T lr_reg_22_ ( .D(n2223), .CP(clk), .Q(lr[22]) );
  DFQD1BWP12T lr_reg_21_ ( .D(n2222), .CP(clk), .Q(lr[21]) );
  DFQD1BWP12T lr_reg_20_ ( .D(n2221), .CP(clk), .Q(lr[20]) );
  DFQD1BWP12T lr_reg_19_ ( .D(n2220), .CP(clk), .Q(lr[19]) );
  DFQD1BWP12T lr_reg_18_ ( .D(n2219), .CP(clk), .Q(lr[18]) );
  DFQD1BWP12T lr_reg_17_ ( .D(n2218), .CP(clk), .Q(lr[17]) );
  DFQD1BWP12T lr_reg_16_ ( .D(n2217), .CP(clk), .Q(lr[16]) );
  DFQD1BWP12T lr_reg_15_ ( .D(n2216), .CP(clk), .Q(lr[15]) );
  DFQD1BWP12T lr_reg_14_ ( .D(n2215), .CP(clk), .Q(lr[14]) );
  DFQD1BWP12T lr_reg_13_ ( .D(n2214), .CP(clk), .Q(lr[13]) );
  DFQD1BWP12T lr_reg_12_ ( .D(n2213), .CP(clk), .Q(lr[12]) );
  DFQD1BWP12T lr_reg_11_ ( .D(n2212), .CP(clk), .Q(lr[11]) );
  DFQD1BWP12T lr_reg_10_ ( .D(n2211), .CP(clk), .Q(lr[10]) );
  DFQD1BWP12T lr_reg_9_ ( .D(n2210), .CP(clk), .Q(lr[9]) );
  DFQD1BWP12T lr_reg_8_ ( .D(n2209), .CP(clk), .Q(lr[8]) );
  DFQD1BWP12T lr_reg_7_ ( .D(n2208), .CP(clk), .Q(lr[7]) );
  DFQD1BWP12T lr_reg_6_ ( .D(n2207), .CP(clk), .Q(lr[6]) );
  DFQD1BWP12T lr_reg_5_ ( .D(n2206), .CP(clk), .Q(lr[5]) );
  DFQD1BWP12T lr_reg_4_ ( .D(n2205), .CP(clk), .Q(lr[4]) );
  DFQD1BWP12T lr_reg_3_ ( .D(n2204), .CP(clk), .Q(lr[3]) );
  DFQD1BWP12T lr_reg_2_ ( .D(n2203), .CP(clk), .Q(lr[2]) );
  DFQD1BWP12T lr_reg_1_ ( .D(n2202), .CP(clk), .Q(lr[1]) );
  DFQD1BWP12T lr_reg_0_ ( .D(n2201), .CP(clk), .Q(lr[0]) );
  DFQD1BWP12T sp_reg_31_ ( .D(spin[31]), .CP(clk), .Q(n[2010]) );
  DFQD1BWP12T sp_reg_30_ ( .D(spin[30]), .CP(clk), .Q(n[2011]) );
  DFQD1BWP12T sp_reg_29_ ( .D(spin[29]), .CP(clk), .Q(n[2012]) );
  DFQD1BWP12T sp_reg_28_ ( .D(spin[28]), .CP(clk), .Q(n[2013]) );
  DFQD1BWP12T sp_reg_27_ ( .D(spin[27]), .CP(clk), .Q(n[2014]) );
  DFQD1BWP12T sp_reg_26_ ( .D(spin[26]), .CP(clk), .Q(n[2015]) );
  DFQD1BWP12T sp_reg_25_ ( .D(spin[25]), .CP(clk), .Q(n[2016]) );
  DFQD1BWP12T sp_reg_24_ ( .D(spin[24]), .CP(clk), .Q(n[2017]) );
  DFQD1BWP12T sp_reg_23_ ( .D(spin[23]), .CP(clk), .Q(n[2018]) );
  DFQD1BWP12T sp_reg_22_ ( .D(spin[22]), .CP(clk), .Q(n[2019]) );
  DFQD1BWP12T sp_reg_21_ ( .D(spin[21]), .CP(clk), .Q(n[2020]) );
  DFQD1BWP12T sp_reg_20_ ( .D(spin[20]), .CP(clk), .Q(n[2021]) );
  DFQD1BWP12T sp_reg_19_ ( .D(spin[19]), .CP(clk), .Q(n[2022]) );
  DFQD1BWP12T sp_reg_18_ ( .D(spin[18]), .CP(clk), .Q(n[2023]) );
  DFQD1BWP12T sp_reg_17_ ( .D(spin[17]), .CP(clk), .Q(n[2024]) );
  DFQD1BWP12T sp_reg_16_ ( .D(spin[16]), .CP(clk), .Q(n[2025]) );
  DFQD1BWP12T sp_reg_15_ ( .D(spin[15]), .CP(clk), .Q(n[2026]) );
  DFQD1BWP12T sp_reg_14_ ( .D(spin[14]), .CP(clk), .Q(n[2027]) );
  DFQD1BWP12T sp_reg_13_ ( .D(spin[13]), .CP(clk), .Q(n[2028]) );
  DFQD1BWP12T sp_reg_12_ ( .D(spin[12]), .CP(clk), .Q(n[2029]) );
  DFQD1BWP12T sp_reg_11_ ( .D(spin[11]), .CP(clk), .Q(n[2030]) );
  DFQD1BWP12T sp_reg_10_ ( .D(spin[10]), .CP(clk), .Q(n[2031]) );
  DFQD1BWP12T sp_reg_9_ ( .D(spin[9]), .CP(clk), .Q(n[2032]) );
  DFQD1BWP12T sp_reg_8_ ( .D(spin[8]), .CP(clk), .Q(n[2033]) );
  DFQD1BWP12T sp_reg_7_ ( .D(spin[7]), .CP(clk), .Q(n[2034]) );
  DFQD1BWP12T sp_reg_6_ ( .D(spin[6]), .CP(clk), .Q(n[2035]) );
  DFQD1BWP12T sp_reg_5_ ( .D(spin[5]), .CP(clk), .Q(n[2036]) );
  DFQD1BWP12T sp_reg_4_ ( .D(spin[4]), .CP(clk), .Q(n[2037]) );
  DFQD1BWP12T sp_reg_3_ ( .D(spin[3]), .CP(clk), .Q(n[2038]) );
  DFQD1BWP12T sp_reg_2_ ( .D(spin[2]), .CP(clk), .Q(n[2039]) );
  DFQD1BWP12T sp_reg_1_ ( .D(spin[1]), .CP(clk), .Q(n[2040]) );
  DFQD1BWP12T sp_reg_0_ ( .D(spin[0]), .CP(clk), .Q(n[2041]) );
  DFQD1BWP12T pc_reg_31_ ( .D(n2200), .CP(clk), .Q(pc_out[31]) );
  DFQD1BWP12T pc_reg_30_ ( .D(n2199), .CP(clk), .Q(pc_out[30]) );
  DFQD1BWP12T pc_reg_28_ ( .D(n2197), .CP(clk), .Q(pc_out[28]) );
  DFQD1BWP12T pc_reg_27_ ( .D(n2196), .CP(clk), .Q(pc_out[27]) );
  DFQD1BWP12T pc_reg_25_ ( .D(n2194), .CP(clk), .Q(pc_out[25]) );
  DFQD1BWP12T pc_reg_24_ ( .D(n2193), .CP(clk), .Q(pc_out[24]) );
  DFQD1BWP12T pc_reg_23_ ( .D(n2192), .CP(clk), .Q(pc_out[23]) );
  DFQD1BWP12T pc_reg_22_ ( .D(n2191), .CP(clk), .Q(pc_out[22]) );
  DFQD1BWP12T pc_reg_21_ ( .D(n2190), .CP(clk), .Q(pc_out[21]) );
  DFQD1BWP12T pc_reg_20_ ( .D(n2189), .CP(clk), .Q(pc_out[20]) );
  DFQD1BWP12T pc_reg_19_ ( .D(n2188), .CP(clk), .Q(pc_out[19]) );
  DFQD1BWP12T pc_reg_18_ ( .D(n2187), .CP(clk), .Q(pc_out[18]) );
  DFQD1BWP12T pc_reg_17_ ( .D(n2186), .CP(clk), .Q(pc_out[17]) );
  DFQD1BWP12T pc_reg_16_ ( .D(n2185), .CP(clk), .Q(pc_out[16]) );
  DFQD1BWP12T pc_reg_15_ ( .D(n2184), .CP(clk), .Q(pc_out[15]) );
  DFQD1BWP12T pc_reg_14_ ( .D(n2183), .CP(clk), .Q(pc_out[14]) );
  DFQD1BWP12T pc_reg_13_ ( .D(n2182), .CP(clk), .Q(pc_out[13]) );
  DFQD1BWP12T pc_reg_12_ ( .D(n2181), .CP(clk), .Q(pc_out[12]) );
  DFQD1BWP12T pc_reg_11_ ( .D(n2180), .CP(clk), .Q(pc_out[11]) );
  DFQD1BWP12T pc_reg_10_ ( .D(n2179), .CP(clk), .Q(pc_out[10]) );
  DFQD1BWP12T pc_reg_9_ ( .D(n2178), .CP(clk), .Q(pc_out[9]) );
  DFQD1BWP12T pc_reg_8_ ( .D(n2177), .CP(clk), .Q(pc_out[8]) );
  DFQD1BWP12T pc_reg_7_ ( .D(n2176), .CP(clk), .Q(pc_out[7]) );
  DFQD1BWP12T pc_reg_6_ ( .D(n2175), .CP(clk), .Q(pc_out[6]) );
  DFQD1BWP12T pc_reg_5_ ( .D(n2174), .CP(clk), .Q(pc_out[5]) );
  DFQD1BWP12T pc_reg_4_ ( .D(n2173), .CP(clk), .Q(pc_out[4]) );
  DFQD1BWP12T pc_reg_0_ ( .D(n2169), .CP(clk), .Q(pc_out[0]) );
  DFQD1BWP12T cpsr_reg_3_ ( .D(cpsrin[3]), .CP(clk), .Q(cpsr_out[3]) );
  DFQD1BWP12T cpsr_reg_2_ ( .D(cpsrin[2]), .CP(clk), .Q(cpsr_out[2]) );
  DFQD1BWP12T cpsr_reg_1_ ( .D(cpsrin[1]), .CP(clk), .Q(cpsr_out[1]) );
  DFQD1BWP12T cpsr_reg_0_ ( .D(cpsrin[0]), .CP(clk), .Q(cpsr_out[0]) );
  DFQD1BWP12T tmp1_reg_31_ ( .D(n2168), .CP(clk), .Q(tmp1[31]) );
  DFQD1BWP12T tmp1_reg_30_ ( .D(n2167), .CP(clk), .Q(tmp1[30]) );
  DFQD1BWP12T tmp1_reg_29_ ( .D(n2166), .CP(clk), .Q(tmp1[29]) );
  DFQD1BWP12T tmp1_reg_28_ ( .D(n2165), .CP(clk), .Q(tmp1[28]) );
  DFQD1BWP12T tmp1_reg_27_ ( .D(n2164), .CP(clk), .Q(tmp1[27]) );
  DFQD1BWP12T tmp1_reg_26_ ( .D(n2163), .CP(clk), .Q(tmp1[26]) );
  DFQD1BWP12T tmp1_reg_25_ ( .D(n2162), .CP(clk), .Q(tmp1[25]) );
  DFQD1BWP12T tmp1_reg_24_ ( .D(n2161), .CP(clk), .Q(tmp1[24]) );
  DFQD1BWP12T tmp1_reg_23_ ( .D(n2160), .CP(clk), .Q(tmp1[23]) );
  DFQD1BWP12T tmp1_reg_22_ ( .D(n2159), .CP(clk), .Q(tmp1[22]) );
  DFQD1BWP12T tmp1_reg_21_ ( .D(n2158), .CP(clk), .Q(tmp1[21]) );
  DFQD1BWP12T tmp1_reg_20_ ( .D(n2157), .CP(clk), .Q(tmp1[20]) );
  DFQD1BWP12T tmp1_reg_19_ ( .D(n2156), .CP(clk), .Q(tmp1[19]) );
  DFQD1BWP12T tmp1_reg_18_ ( .D(n2155), .CP(clk), .Q(tmp1[18]) );
  DFQD1BWP12T tmp1_reg_17_ ( .D(n2154), .CP(clk), .Q(tmp1[17]) );
  DFQD1BWP12T tmp1_reg_16_ ( .D(n2153), .CP(clk), .Q(tmp1[16]) );
  DFQD1BWP12T tmp1_reg_15_ ( .D(n2152), .CP(clk), .Q(tmp1[15]) );
  DFQD1BWP12T tmp1_reg_14_ ( .D(n2151), .CP(clk), .Q(tmp1[14]) );
  DFQD1BWP12T tmp1_reg_13_ ( .D(n2150), .CP(clk), .Q(tmp1[13]) );
  DFQD1BWP12T tmp1_reg_12_ ( .D(n2149), .CP(clk), .Q(tmp1[12]) );
  DFQD1BWP12T tmp1_reg_11_ ( .D(n2148), .CP(clk), .Q(tmp1[11]) );
  DFQD1BWP12T tmp1_reg_10_ ( .D(n2147), .CP(clk), .Q(tmp1[10]) );
  DFQD1BWP12T tmp1_reg_9_ ( .D(n2146), .CP(clk), .Q(tmp1[9]) );
  DFQD1BWP12T tmp1_reg_8_ ( .D(n2145), .CP(clk), .Q(tmp1[8]) );
  DFQD1BWP12T tmp1_reg_7_ ( .D(n2144), .CP(clk), .Q(tmp1[7]) );
  DFQD1BWP12T tmp1_reg_6_ ( .D(n2143), .CP(clk), .Q(tmp1[6]) );
  DFQD1BWP12T tmp1_reg_5_ ( .D(n2142), .CP(clk), .Q(tmp1[5]) );
  DFQD1BWP12T tmp1_reg_4_ ( .D(n2141), .CP(clk), .Q(tmp1[4]) );
  DFQD1BWP12T tmp1_reg_3_ ( .D(n2140), .CP(clk), .Q(tmp1[3]) );
  DFQD1BWP12T tmp1_reg_2_ ( .D(n2139), .CP(clk), .Q(tmp1[2]) );
  DFQD1BWP12T tmp1_reg_1_ ( .D(n2138), .CP(clk), .Q(tmp1[1]) );
  DFQD1BWP12T tmp1_reg_0_ ( .D(n2136), .CP(clk), .Q(tmp1[0]) );
  DFQD2BWP12T pc_reg_1_ ( .D(n2170), .CP(clk), .Q(pc_out[1]) );
  DFQD1BWP12T pc_reg_3_ ( .D(n2172), .CP(clk), .Q(pc_out[3]) );
  DFQD1BWP12T pc_reg_26_ ( .D(n2195), .CP(clk), .Q(pc_out[26]) );
  DFQD1BWP12T pc_reg_29_ ( .D(n2198), .CP(clk), .Q(pc_out[29]) );
  DFQD2BWP12T pc_reg_2_ ( .D(n2171), .CP(clk), .Q(pc_out[2]) );
  INVD1BWP12T U3 ( .I(n151), .ZN(n152) );
  ND2D1BWP12T U4 ( .A1(n1850), .A2(n1849), .ZN(n1854) );
  AOI22D1BWP12T U5 ( .A1(r11[1]), .A2(n537), .B1(n205), .B2(r0[1]), .ZN(n1849)
         );
  CKND2D2BWP12T U6 ( .A1(n1871), .A2(n1870), .ZN(regB_out[1]) );
  NR4D0BWP12T U7 ( .A1(n1869), .A2(n1868), .A3(n1867), .A4(n1866), .ZN(n1870)
         );
  INVD1BWP12T U8 ( .I(n172), .ZN(n144) );
  INR2D2BWP12T U9 ( .A1(n153), .B1(n152), .ZN(n521) );
  OAI22D1BWP12T U10 ( .A1(n1852), .A2(n1940), .B1(n1851), .B2(n1928), .ZN(
        n1853) );
  MOAI22D0BWP12T U11 ( .A1(n1848), .A2(n1847), .B1(n200), .B2(immediate2_in[1]), .ZN(n1855) );
  CKBD1BWP12T U12 ( .I(write1_in[17]), .Z(n1239) );
  OAI22D1BWP12T U13 ( .A1(n1852), .A2(n1915), .B1(n1851), .B2(n1903), .ZN(
        n1834) );
  OAI22D1BWP12T U14 ( .A1(n1969), .A2(n1690), .B1(n1967), .B2(n1689), .ZN(
        n1700) );
  OAI22D1BWP12T U15 ( .A1(n1719), .A2(n1976), .B1(n1975), .B2(n1729), .ZN(
        n1710) );
  OAI22D1BWP12T U16 ( .A1(n1973), .A2(n1731), .B1(n1971), .B2(n1730), .ZN(
        n1711) );
  AOI22D1BWP12T U17 ( .A1(tmp1[0]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[0]), .ZN(n652) );
  INVD1BWP12T U18 ( .I(n1239), .ZN(n53) );
  ND2D1BWP12T U19 ( .A1(n182), .A2(n181), .ZN(regA_out[13]) );
  NR2D1BWP12T U20 ( .A1(n112), .A2(n111), .ZN(n1315) );
  INVD1BWP12T U21 ( .I(n53), .ZN(n55) );
  INVD1BWP12T U22 ( .I(n1162), .ZN(n1205) );
  INVD1BWP12T U23 ( .I(n1163), .ZN(n1206) );
  INVD1BWP12T U24 ( .I(n1158), .ZN(n1203) );
  INVD1BWP12T U25 ( .I(n1159), .ZN(n1204) );
  INVD1BWP12T U26 ( .I(n1156), .ZN(n1199) );
  INVD1BWP12T U27 ( .I(n1157), .ZN(n1200) );
  INVD1BWP12T U28 ( .I(n1160), .ZN(n1201) );
  INVD1BWP12T U29 ( .I(n1161), .ZN(n1202) );
  ND4D2BWP12T U30 ( .A1(n587), .A2(n586), .A3(n585), .A4(n584), .ZN(
        regA_out[28]) );
  OA211D1BWP12T U31 ( .A1(n236), .A2(n1458), .B(n235), .C(n234), .Z(n244) );
  INR2XD2BWP12T U32 ( .A1(n209), .B1(n203), .ZN(n1994) );
  TPNR2D1BWP12T U33 ( .A1(n218), .A2(n202), .ZN(n536) );
  INVD2BWP12T U34 ( .I(n185), .ZN(n1861) );
  TPNR2D2BWP12T U35 ( .A1(n173), .A2(n170), .ZN(n171) );
  INVD3BWP12T U36 ( .I(n141), .ZN(n1949) );
  INVD2BWP12T U37 ( .I(n1555), .ZN(n1959) );
  INVD1BWP12T U38 ( .I(n1591), .ZN(n1969) );
  XNR2D1BWP12T U39 ( .A1(n1349), .A2(n1346), .ZN(n383) );
  OAI21D1BWP12T U40 ( .A1(n1346), .A2(n1348), .B(n1345), .ZN(n1347) );
  OAI22D1BWP12T U41 ( .A1(n1852), .A2(n1890), .B1(n1851), .B2(n1878), .ZN(n540) );
  OAI22D1BWP12T U42 ( .A1(n1852), .A2(n822), .B1(n1851), .B2(n828), .ZN(n602)
         );
  OAI22D1BWP12T U43 ( .A1(n1865), .A2(n836), .B1(n1864), .B2(n827), .ZN(n607)
         );
  INR2D1BWP12T U44 ( .A1(readA_sel[4]), .B1(n172), .ZN(n151) );
  INR2D0BWP12T U45 ( .A1(n116), .B1(n115), .ZN(n1291) );
  INR2D0BWP12T U46 ( .A1(n133), .B1(n132), .ZN(n1288) );
  AO22D1BWP12T U47 ( .A1(n1328), .A2(write2_in[8]), .B1(n1330), .B2(
        write1_in[8]), .Z(n1231) );
  INR2D0BWP12T U48 ( .A1(n78), .B1(n77), .ZN(n1303) );
  INR2D0BWP12T U49 ( .A1(n57), .B1(n56), .ZN(n1297) );
  AO22D0BWP12T U50 ( .A1(n1328), .A2(write2_in[10]), .B1(n1330), .B2(
        write1_in[10]), .Z(n1236) );
  INR2D0BWP12T U51 ( .A1(n73), .B1(n72), .ZN(n1282) );
  INR3D0BWP12T U52 ( .A1(n128), .B1(n129), .B2(reset), .ZN(n1309) );
  AN2XD2BWP12T U53 ( .A1(readB_sel[2]), .A2(readB_sel[1]), .Z(n214) );
  MAOI22D0BWP12T U54 ( .A1(n1247), .A2(n1246), .B1(n1247), .B2(n1246), .ZN(n1)
         );
  AO222D0BWP12T U55 ( .A1(pc_out[13]), .A2(n1361), .B1(n1), .B2(n1363), .C1(
        next_pc_in[13]), .C2(n1355), .Z(n2182) );
  MAOI22D0BWP12T U56 ( .A1(n1249), .A2(n1248), .B1(n1249), .B2(n1248), .ZN(n2)
         );
  AO222D0BWP12T U57 ( .A1(pc_out[14]), .A2(n1361), .B1(n2), .B2(n1363), .C1(
        next_pc_in[14]), .C2(n1355), .Z(n2183) );
  MAOI22D0BWP12T U58 ( .A1(n1252), .A2(n1251), .B1(n1252), .B2(n1251), .ZN(n3)
         );
  AO222D0BWP12T U59 ( .A1(pc_out[15]), .A2(n1361), .B1(n3), .B2(n1363), .C1(
        next_pc_in[15]), .C2(n1355), .Z(n2184) );
  IND3D0BWP12T U60 ( .A1(write1_sel[0]), .B1(write1_sel[3]), .B2(write1_en), 
        .ZN(n62) );
  AOI22D1BWP12T U61 ( .A1(n1328), .A2(write2_in[11]), .B1(n1330), .B2(
        write1_in[11]), .ZN(n1241) );
  AOI22D0BWP12T U62 ( .A1(n1328), .A2(write2_in[21]), .B1(n1330), .B2(
        write1_in[21]), .ZN(n1271) );
  INR3D0BWP12T U63 ( .A1(n122), .B1(n123), .B2(reset), .ZN(n1273) );
  INR2D0BWP12T U64 ( .A1(n140), .B1(n139), .ZN(n1300) );
  OA211D0BWP12T U65 ( .A1(n1458), .A2(n615), .B(n614), .C(n613), .Z(n4) );
  AN4XD1BWP12T U66 ( .A1(n616), .A2(n617), .A3(n618), .A4(n619), .Z(n5) );
  AOI22D1BWP12T U67 ( .A1(n1561), .A2(lr[30]), .B1(n1560), .B2(r10[30]), .ZN(
        n6) );
  AOI22D1BWP12T U68 ( .A1(n141), .A2(pc_out[30]), .B1(n1559), .B2(r11[30]), 
        .ZN(n7) );
  ND4D1BWP12T U69 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(regA_out[30]) );
  MAOI22D0BWP12T U70 ( .A1(n1262), .A2(n1261), .B1(n1262), .B2(n1261), .ZN(n8)
         );
  AO222D0BWP12T U71 ( .A1(pc_out[18]), .A2(n1361), .B1(n8), .B2(n1363), .C1(
        next_pc_in[18]), .C2(n1355), .Z(n2187) );
  NR2D0BWP12T U72 ( .A1(write1_sel[3]), .A2(n85), .ZN(n67) );
  AO22D1BWP12T U73 ( .A1(n1328), .A2(write2_in[14]), .B1(n1330), .B2(
        write1_in[14]), .Z(n1249) );
  INR2D0BWP12T U74 ( .A1(n71), .B1(n70), .ZN(n1294) );
  AO222D1BWP12T U75 ( .A1(r6[30]), .A2(n1995), .B1(r8[30]), .B2(n187), .C1(
        n[2011]), .C2(n1994), .Z(n9) );
  AOI22D0BWP12T U76 ( .A1(n1992), .A2(r12[30]), .B1(r1[30]), .B2(n183), .ZN(
        n10) );
  AOI22D0BWP12T U77 ( .A1(r3[30]), .A2(n185), .B1(lr[30]), .B2(n1993), .ZN(n11) );
  ND4D1BWP12T U78 ( .A1(n1399), .A2(n1398), .A3(n10), .A4(n11), .ZN(n12) );
  AOI211D1BWP12T U79 ( .A1(n188), .A2(pc_out[30]), .B(n9), .C(n12), .ZN(n13)
         );
  AOI22D0BWP12T U80 ( .A1(r2[30]), .A2(n1989), .B1(r7[30]), .B2(n215), .ZN(n14) );
  AOI22D0BWP12T U81 ( .A1(n1988), .A2(r10[30]), .B1(r5[30]), .B2(n210), .ZN(
        n15) );
  ND4D1BWP12T U82 ( .A1(n13), .A2(n1400), .A3(n14), .A4(n15), .ZN(regB_out[30]) );
  MAOI22D0BWP12T U83 ( .A1(n1266), .A2(n1265), .B1(n1266), .B2(n1265), .ZN(n16) );
  AO222D0BWP12T U84 ( .A1(pc_out[19]), .A2(n1361), .B1(n16), .B2(n1363), .C1(
        next_pc_in[19]), .C2(n1362), .Z(n2188) );
  IND3D0BWP12T U85 ( .A1(n62), .B1(n79), .B2(write1_sel[4]), .ZN(n63) );
  INR3D0BWP12T U86 ( .A1(write1_sel[2]), .B1(write1_sel[1]), .B2(reset), .ZN(
        n109) );
  NR4D0BWP12T U87 ( .A1(n1664), .A2(n1663), .A3(n1662), .A4(n1661), .ZN(n17)
         );
  ND2D1BWP12T U88 ( .A1(n1677), .A2(n17), .ZN(regA_out[11]) );
  AO22D1BWP12T U89 ( .A1(n1328), .A2(write2_in[22]), .B1(n1330), .B2(n1250), 
        .Z(n1318) );
  MAOI22D0BWP12T U90 ( .A1(n1270), .A2(n1269), .B1(n1270), .B2(n1269), .ZN(n18) );
  AO222D0BWP12T U91 ( .A1(pc_out[20]), .A2(n1361), .B1(n18), .B2(n1363), .C1(
        next_pc_in[20]), .C2(n1362), .Z(n2189) );
  OAI22D0BWP12T U92 ( .A1(n1949), .A2(n1733), .B1(n1948), .B2(n1703), .ZN(n19)
         );
  OAI22D0BWP12T U93 ( .A1(n1953), .A2(n1728), .B1(n1952), .B2(n1718), .ZN(n20)
         );
  NR4D0BWP12T U94 ( .A1(n1706), .A2(n1705), .A3(n19), .A4(n20), .ZN(n1714) );
  NR2D0BWP12T U95 ( .A1(n62), .A2(write1_sel[4]), .ZN(n130) );
  AN2D0BWP12T U96 ( .A1(write1_sel[0]), .A2(n67), .Z(n135) );
  INR2D0BWP12T U97 ( .A1(n118), .B1(n117), .ZN(n1276) );
  MAOI22D0BWP12T U98 ( .A1(n108), .A2(n430), .B1(n108), .B2(n430), .ZN(n21) );
  AO222D0BWP12T U99 ( .A1(pc_out[2]), .A2(n1361), .B1(n1363), .B2(n21), .C1(
        next_pc_in[2]), .C2(n1355), .Z(n2171) );
  MAOI22D0BWP12T U100 ( .A1(n1272), .A2(n1271), .B1(n1272), .B2(n1271), .ZN(
        n22) );
  AO222D0BWP12T U101 ( .A1(pc_out[21]), .A2(n1361), .B1(n22), .B2(n1363), .C1(
        next_pc_in[21]), .C2(n1355), .Z(n2190) );
  NR2D0BWP12T U102 ( .A1(write2_sel[0]), .A2(n99), .ZN(n23) );
  ND4D0BWP12T U103 ( .A1(write2_en), .A2(write2_sel[4]), .A3(write2_sel[3]), 
        .A4(n23), .ZN(n64) );
  AO222D1BWP12T U104 ( .A1(n1957), .A2(r4[17]), .B1(n1809), .B2(tmp1[17]), 
        .C1(r12[17]), .C2(n150), .Z(n1529) );
  AOI22D0BWP12T U105 ( .A1(n1361), .A2(pc_out[31]), .B1(n1355), .B2(
        next_pc_in[31]), .ZN(n1337) );
  INR2D1BWP12T U106 ( .A1(n112), .B1(n111), .ZN(n421) );
  MAOI22D0BWP12T U107 ( .A1(n107), .A2(n106), .B1(n107), .B2(n106), .ZN(n24)
         );
  AO222D0BWP12T U108 ( .A1(pc_out[3]), .A2(n1361), .B1(n24), .B2(n1363), .C1(
        next_pc_in[3]), .C2(n1355), .Z(n2172) );
  INR2D0BWP12T U109 ( .A1(next_cpsr_in[2]), .B1(reset), .ZN(cpsrin[2]) );
  MAOI22D0BWP12T U110 ( .A1(n373), .A2(n372), .B1(n373), .B2(n372), .ZN(n25)
         );
  AO222D0BWP12T U111 ( .A1(pc_out[5]), .A2(n1361), .B1(n25), .B2(n1363), .C1(
        next_pc_in[5]), .C2(n1355), .Z(n2174) );
  MAOI22D0BWP12T U112 ( .A1(n1229), .A2(n1228), .B1(n1229), .B2(n1228), .ZN(
        n26) );
  AO222D0BWP12T U113 ( .A1(pc_out[7]), .A2(n1361), .B1(n26), .B2(n1363), .C1(
        next_pc_in[7]), .C2(n1355), .Z(n2176) );
  MAOI22D0BWP12T U114 ( .A1(n1235), .A2(n1234), .B1(n1235), .B2(n1234), .ZN(
        n27) );
  AO222D0BWP12T U115 ( .A1(pc_out[9]), .A2(n1361), .B1(n27), .B2(n1363), .C1(
        next_pc_in[9]), .C2(n1355), .Z(n2178) );
  MAOI22D0BWP12T U116 ( .A1(n1241), .A2(n1240), .B1(n1241), .B2(n1240), .ZN(
        n28) );
  AO222D0BWP12T U117 ( .A1(pc_out[11]), .A2(n1361), .B1(n28), .B2(n1363), .C1(
        next_pc_in[11]), .C2(n1355), .Z(n2180) );
  MAOI22D0BWP12T U118 ( .A1(n1319), .A2(n1318), .B1(n1319), .B2(n1318), .ZN(
        n29) );
  AO222D0BWP12T U119 ( .A1(pc_out[22]), .A2(n1361), .B1(n29), .B2(n1363), .C1(
        next_pc_in[22]), .C2(n1355), .Z(n2191) );
  CKND0BWP12T U120 ( .I(r7[14]), .ZN(n30) );
  OAI22D0BWP12T U121 ( .A1(n1852), .A2(n30), .B1(n1851), .B2(n624), .ZN(n625)
         );
  OAI22D0BWP12T U122 ( .A1(n1948), .A2(n1482), .B1(n1483), .B2(n1949), .ZN(n31) );
  OAI22D0BWP12T U123 ( .A1(n1959), .A2(n1488), .B1(n1961), .B2(n1489), .ZN(n32) );
  NR4D0BWP12T U124 ( .A1(n1491), .A2(n1490), .A3(n31), .A4(n32), .ZN(n1497) );
  AO222D0BWP12T U125 ( .A1(n1957), .A2(r4[20]), .B1(n1486), .B2(tmp1[20]), 
        .C1(r12[20]), .C2(n150), .Z(n496) );
  AN2D0BWP12T U126 ( .A1(write1_sel[2]), .A2(write1_sel[1]), .Z(n93) );
  IND2D0BWP12T U127 ( .A1(n76), .B1(n75), .ZN(n448) );
  OAI22D0BWP12T U128 ( .A1(write1_in[0]), .A2(n1328), .B1(write2_in[0]), .B2(
        n1330), .ZN(n33) );
  AOI22D0BWP12T U129 ( .A1(pc_out[0]), .A2(n1361), .B1(next_pc_in[0]), .B2(
        n1355), .ZN(n34) );
  OAI21D0BWP12T U130 ( .A1(n1334), .A2(n33), .B(n34), .ZN(n2169) );
  MAOI22D0BWP12T U131 ( .A1(n105), .A2(n104), .B1(n105), .B2(n104), .ZN(n35)
         );
  AO222D0BWP12T U132 ( .A1(pc_out[4]), .A2(n1361), .B1(n35), .B2(n1363), .C1(
        next_pc_in[4]), .C2(n1355), .Z(n2173) );
  MAOI22D0BWP12T U133 ( .A1(n1227), .A2(n1226), .B1(n1227), .B2(n1226), .ZN(
        n36) );
  AO222D0BWP12T U134 ( .A1(pc_out[6]), .A2(n1361), .B1(n36), .B2(n1363), .C1(
        next_pc_in[6]), .C2(n1355), .Z(n2175) );
  MAOI22D0BWP12T U135 ( .A1(n1231), .A2(n1230), .B1(n1231), .B2(n1230), .ZN(
        n37) );
  AO222D0BWP12T U136 ( .A1(pc_out[8]), .A2(n1361), .B1(n37), .B2(n1363), .C1(
        next_pc_in[8]), .C2(n1355), .Z(n2177) );
  MAOI22D0BWP12T U137 ( .A1(n1237), .A2(n1236), .B1(n1237), .B2(n1236), .ZN(
        n38) );
  AO222D0BWP12T U138 ( .A1(pc_out[10]), .A2(n1361), .B1(n38), .B2(n1363), .C1(
        next_pc_in[10]), .C2(n1355), .Z(n2179) );
  MAOI22D0BWP12T U139 ( .A1(n1244), .A2(n1243), .B1(n1244), .B2(n1243), .ZN(
        n39) );
  AO222D0BWP12T U140 ( .A1(pc_out[12]), .A2(n1361), .B1(n39), .B2(n1363), .C1(
        next_pc_in[12]), .C2(n1355), .Z(n2181) );
  MAOI22D0BWP12T U141 ( .A1(n1324), .A2(n1323), .B1(n1324), .B2(n1323), .ZN(
        n40) );
  AO222D0BWP12T U142 ( .A1(pc_out[23]), .A2(n1361), .B1(n40), .B2(n1363), .C1(
        next_pc_in[23]), .C2(n1355), .Z(n2192) );
  AOI22D0BWP12T U143 ( .A1(r7[30]), .A2(n1200), .B1(r4[30]), .B2(n1199), .ZN(
        n41) );
  AOI22D0BWP12T U144 ( .A1(r6[30]), .A2(n1201), .B1(r2[30]), .B2(n1202), .ZN(
        n42) );
  AOI22D0BWP12T U145 ( .A1(r1[30]), .A2(n1203), .B1(r5[30]), .B2(n1204), .ZN(
        n43) );
  AOI22D0BWP12T U146 ( .A1(r0[30]), .A2(n1206), .B1(r3[30]), .B2(n1205), .ZN(
        n44) );
  ND4D0BWP12T U147 ( .A1(n41), .A2(n42), .A3(n43), .A4(n44), .ZN(n45) );
  AO22D0BWP12T U148 ( .A1(r9[30]), .A2(n1211), .B1(r10[30]), .B2(n1218), .Z(
        n46) );
  CKND0BWP12T U149 ( .I(r8[30]), .ZN(n47) );
  AOI22D0BWP12T U150 ( .A1(n[2011]), .A2(n1213), .B1(lr[30]), .B2(n1214), .ZN(
        n48) );
  CKND0BWP12T U151 ( .I(n1193), .ZN(n49) );
  CKND0BWP12T U152 ( .I(n1132), .ZN(n50) );
  AOI222D0BWP12T U153 ( .A1(n49), .A2(r12[30]), .B1(pc_out[30]), .B2(n1215), 
        .C1(n50), .C2(r11[30]), .ZN(n51) );
  OAI211D0BWP12T U154 ( .A1(n1136), .A2(n47), .B(n48), .C(n51), .ZN(n52) );
  AO211D0BWP12T U155 ( .A1(n1225), .A2(n45), .B(n46), .C(n52), .Z(regC_out[30]) );
  DCCKND8BWP12T U156 ( .I(readB_sel[4]), .ZN(n189) );
  NR2D3BWP12T U157 ( .A1(n175), .A2(n170), .ZN(n155) );
  RCAOI21D4BWP12T U158 ( .A1(n1331), .A2(n1330), .B(n1329), .ZN(n1336) );
  INVD1BWP12T U159 ( .I(n53), .ZN(n54) );
  INVD3BWP12T U160 ( .I(n1559), .ZN(n1948) );
  DCCKND4BWP12T U161 ( .I(n1989), .ZN(n1851) );
  NR4D1BWP12T U162 ( .A1(n1770), .A2(n1769), .A3(n1768), .A4(n1767), .ZN(n1778) );
  BUFFXD4BWP12T U163 ( .I(write1_in[28]), .Z(n1268) );
  TPNR2D2BWP12T U164 ( .A1(n1259), .A2(n1258), .ZN(n1262) );
  TPOAI22D1BWP12T U165 ( .A1(n1937), .A2(n1861), .B1(n1860), .B2(n1925), .ZN(
        n1868) );
  INR2XD2BWP12T U166 ( .A1(n144), .B1(n165), .ZN(n141) );
  ND3D4BWP12T U167 ( .A1(n147), .A2(readA_sel[0]), .A3(readA_sel[3]), .ZN(n165) );
  TPNR2D3BWP12T U168 ( .A1(n1247), .A2(n1246), .ZN(n1248) );
  TPND2D4BWP12T U169 ( .A1(n1244), .A2(n1243), .ZN(n1247) );
  BUFFXD4BWP12T U170 ( .I(write1_in[16]), .Z(n1232) );
  INR2D8BWP12T U171 ( .A1(n167), .B1(n164), .ZN(n150) );
  TPND2D3BWP12T U172 ( .A1(n1256), .A2(n1255), .ZN(n1259) );
  INR3D2BWP12T U173 ( .A1(n652), .B1(n651), .B2(n650), .ZN(n658) );
  INVD3BWP12T U174 ( .I(n155), .ZN(n1961) );
  INR2D8BWP12T U175 ( .A1(n204), .B1(n203), .ZN(n201) );
  TPAOI21D4BWP12T U176 ( .A1(write1_in[3]), .A2(n1330), .B(n95), .ZN(n107) );
  DCCKND4BWP12T U177 ( .I(n1995), .ZN(n1864) );
  TPAOI21D2BWP12T U178 ( .A1(write1_in[5]), .A2(n1330), .B(n94), .ZN(n373) );
  TPNR2D2BWP12T U179 ( .A1(n1338), .A2(n1334), .ZN(n1335) );
  TPAOI21D8BWP12T U180 ( .A1(n1327), .A2(n1330), .B(n1326), .ZN(n1338) );
  TPND2D2BWP12T U181 ( .A1(n108), .A2(n430), .ZN(n106) );
  TPND2D3BWP12T U182 ( .A1(n1249), .A2(n1248), .ZN(n1252) );
  TPNR2D4BWP12T U183 ( .A1(n1252), .A2(n1251), .ZN(n1255) );
  CKND2D2BWP12T U184 ( .A1(n1358), .A2(n1357), .ZN(n1360) );
  NR2XD3BWP12T U185 ( .A1(n1343), .A2(n1342), .ZN(n1358) );
  BUFFXD8BWP12T U186 ( .I(n536), .Z(n1780) );
  INR2XD2BWP12T U187 ( .A1(n381), .B1(n1354), .ZN(n1349) );
  XOR2XD2BWP12T U188 ( .A1(n1321), .A2(n1320), .Z(n1322) );
  INR2XD2BWP12T U189 ( .A1(n204), .B1(n213), .ZN(n183) );
  INR2XD2BWP12T U190 ( .A1(n214), .B1(n213), .ZN(n215) );
  INR2XD2BWP12T U191 ( .A1(n204), .B1(n211), .ZN(n187) );
  ND4D1BWP12T U192 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(
        regB_out[23]) );
  ND4D2BWP12T U193 ( .A1(n645), .A2(n644), .A3(n643), .A4(n642), .ZN(
        regA_out[22]) );
  ND4D1BWP12T U194 ( .A1(n268), .A2(n267), .A3(n266), .A4(n265), .ZN(
        regB_out[22]) );
  ND4D1BWP12T U195 ( .A1(n233), .A2(n232), .A3(n231), .A4(n230), .ZN(
        regB_out[24]) );
  ND4D1BWP12T U196 ( .A1(n777), .A2(n776), .A3(n775), .A4(n774), .ZN(
        regB_out[27]) );
  ND4D1BWP12T U197 ( .A1(n598), .A2(n597), .A3(n596), .A4(n595), .ZN(
        regB_out[25]) );
  INR2XD2BWP12T U198 ( .A1(n216), .B1(n213), .ZN(n185) );
  INR2XD2BWP12T U199 ( .A1(n209), .B1(n213), .ZN(n210) );
  INR2XD2BWP12T U200 ( .A1(n204), .B1(n218), .ZN(n205) );
  INR2XD2BWP12T U201 ( .A1(readB_sel[0]), .B1(n199), .ZN(n200) );
  INR2D2BWP12T U202 ( .A1(n214), .B1(n203), .ZN(n188) );
  IND2XD1BWP12T U203 ( .A1(write1_sel[4]), .B1(write1_en), .ZN(n85) );
  ND2D1BWP12T U204 ( .A1(n135), .A2(n109), .ZN(n453) );
  INVD1BWP12T U205 ( .I(n453), .ZN(n1299) );
  BUFFD2BWP12T U206 ( .I(write1_in[18]), .Z(n1238) );
  INR2D1BWP12T U207 ( .A1(write2_en), .B1(write2_sel[4]), .ZN(n58) );
  AN2XD1BWP12T U208 ( .A1(write2_sel[0]), .A2(n58), .Z(n87) );
  INVD1BWP12T U209 ( .I(write2_sel[3]), .ZN(n68) );
  AN2XD1BWP12T U210 ( .A1(n87), .A2(n68), .Z(n137) );
  INR2D1BWP12T U211 ( .A1(write2_sel[2]), .B1(write2_sel[1]), .ZN(n110) );
  CKND2D1BWP12T U212 ( .A1(n137), .A2(n110), .ZN(n57) );
  INVD1BWP12T U213 ( .I(reset), .ZN(n138) );
  ND2D1BWP12T U214 ( .A1(n453), .A2(n138), .ZN(n56) );
  NR2D1BWP12T U215 ( .A1(n57), .A2(n56), .ZN(n1298) );
  AO222D0BWP12T U216 ( .A1(n1299), .A2(n1238), .B1(n1297), .B2(r5[18]), .C1(
        write2_in[18]), .C2(n1298), .Z(n2475) );
  ND2D1BWP12T U217 ( .A1(n109), .A2(n130), .ZN(n444) );
  INVD1BWP12T U218 ( .I(n444), .ZN(n1281) );
  INR2D1BWP12T U219 ( .A1(n58), .B1(write2_sel[0]), .ZN(n69) );
  AN2XD1BWP12T U220 ( .A1(n69), .A2(write2_sel[3]), .Z(n131) );
  CKND2D1BWP12T U221 ( .A1(n131), .A2(n110), .ZN(n61) );
  INVD1BWP12T U222 ( .I(n61), .ZN(n59) );
  ND2D1BWP12T U223 ( .A1(n444), .A2(n138), .ZN(n60) );
  NR2D1BWP12T U224 ( .A1(n59), .A2(n60), .ZN(n1279) );
  NR2D1BWP12T U225 ( .A1(n61), .A2(n60), .ZN(n1280) );
  AO222D0BWP12T U226 ( .A1(n1281), .A2(n1238), .B1(n1279), .B2(r12[18]), .C1(
        write2_in[18]), .C2(n1280), .Z(n2251) );
  INR2D1BWP12T U227 ( .A1(n93), .B1(reset), .ZN(n79) );
  INVD1BWP12T U228 ( .I(n63), .ZN(n1317) );
  ND2D1BWP12T U229 ( .A1(n63), .A2(n138), .ZN(n66) );
  ND2D1BWP12T U230 ( .A1(write2_sel[2]), .A2(write2_sel[1]), .ZN(n99) );
  NR2D1BWP12T U231 ( .A1(n66), .A2(n64), .ZN(n820) );
  INVD1BWP12T U232 ( .I(n64), .ZN(n65) );
  NR2D1BWP12T U233 ( .A1(n66), .A2(n65), .ZN(n819) );
  AO222D0BWP12T U234 ( .A1(n1317), .A2(n1238), .B1(n820), .B2(write2_in[18]), 
        .C1(n819), .C2(tmp1[18]), .Z(n2155) );
  INR2D1BWP12T U235 ( .A1(n67), .B1(write1_sel[0]), .ZN(n119) );
  ND2D1BWP12T U236 ( .A1(n119), .A2(n109), .ZN(n471) );
  INVD1BWP12T U237 ( .I(n471), .ZN(n1296) );
  AN2XD1BWP12T U238 ( .A1(n69), .A2(n68), .Z(n120) );
  CKND2D1BWP12T U239 ( .A1(n120), .A2(n110), .ZN(n71) );
  ND2D1BWP12T U240 ( .A1(n471), .A2(n138), .ZN(n70) );
  NR2D1BWP12T U241 ( .A1(n71), .A2(n70), .ZN(n1295) );
  AO222D0BWP12T U242 ( .A1(n1296), .A2(n1238), .B1(n1294), .B2(r4[18]), .C1(
        write2_in[18]), .C2(n1295), .Z(n2507) );
  ND2D1BWP12T U243 ( .A1(n119), .A2(n79), .ZN(n468) );
  INVD1BWP12T U244 ( .I(n468), .ZN(n1284) );
  INVD1BWP12T U245 ( .I(n99), .ZN(n80) );
  ND2D1BWP12T U246 ( .A1(n120), .A2(n80), .ZN(n73) );
  ND2D1BWP12T U247 ( .A1(n468), .A2(n138), .ZN(n72) );
  NR2D1BWP12T U248 ( .A1(n73), .A2(n72), .ZN(n1283) );
  AO222D0BWP12T U249 ( .A1(n1284), .A2(n1238), .B1(n1282), .B2(r6[18]), .C1(
        write2_in[18]), .C2(n1283), .Z(n2443) );
  IND2D1BWP12T U250 ( .A1(write1_sel[2]), .B1(write1_sel[1]), .ZN(n126) );
  INVD1BWP12T U251 ( .I(n126), .ZN(n88) );
  ND2D1BWP12T U252 ( .A1(n88), .A2(n138), .ZN(n124) );
  CKND0BWP12T U253 ( .I(n130), .ZN(n74) );
  NR2D1BWP12T U254 ( .A1(n124), .A2(n74), .ZN(n1314) );
  INVD1BWP12T U255 ( .I(write2_sel[1]), .ZN(n89) );
  NR3D1BWP12T U256 ( .A1(n89), .A2(reset), .A3(write2_sel[2]), .ZN(n125) );
  CKND2D1BWP12T U257 ( .A1(n131), .A2(n125), .ZN(n76) );
  TPND2D0BWP12T U258 ( .A1(n88), .A2(n130), .ZN(n75) );
  INVD1BWP12T U259 ( .I(n448), .ZN(n1313) );
  AN3XD1BWP12T U260 ( .A1(n76), .A2(n138), .A3(n75), .Z(n1312) );
  AO222D0BWP12T U261 ( .A1(n1314), .A2(n1238), .B1(n1313), .B2(write2_in[18]), 
        .C1(n1312), .C2(r10[18]), .Z(n2315) );
  ND2D1BWP12T U262 ( .A1(n135), .A2(n79), .ZN(n441) );
  INVD1BWP12T U263 ( .I(n441), .ZN(n1305) );
  ND2D1BWP12T U264 ( .A1(n137), .A2(n80), .ZN(n78) );
  ND2D1BWP12T U265 ( .A1(n441), .A2(n138), .ZN(n77) );
  NR2D1BWP12T U266 ( .A1(n78), .A2(n77), .ZN(n1304) );
  AO222D0BWP12T U267 ( .A1(n1305), .A2(n1238), .B1(n1303), .B2(r7[18]), .C1(
        write2_in[18]), .C2(n1304), .Z(n2411) );
  ND2D1BWP12T U268 ( .A1(n79), .A2(n130), .ZN(n478) );
  INVD1BWP12T U269 ( .I(n478), .ZN(n1287) );
  ND2D1BWP12T U270 ( .A1(n131), .A2(n80), .ZN(n83) );
  INVD1BWP12T U271 ( .I(n83), .ZN(n81) );
  ND2D1BWP12T U272 ( .A1(n478), .A2(n138), .ZN(n82) );
  NR2D1BWP12T U273 ( .A1(n81), .A2(n82), .ZN(n1285) );
  NR2D1BWP12T U274 ( .A1(n83), .A2(n82), .ZN(n1286) );
  AO222D0BWP12T U275 ( .A1(n1287), .A2(n1238), .B1(n1285), .B2(lr[18]), .C1(
        write2_in[18]), .C2(n1286), .Z(n2219) );
  CKND2D1BWP12T U276 ( .A1(write1_sel[3]), .A2(write1_sel[0]), .ZN(n84) );
  NR2D1BWP12T U277 ( .A1(n85), .A2(n84), .ZN(n113) );
  CKND0BWP12T U278 ( .I(n113), .ZN(n86) );
  NR2D1BWP12T U279 ( .A1(n86), .A2(n124), .ZN(n1308) );
  ND2D1BWP12T U280 ( .A1(n87), .A2(write2_sel[3]), .ZN(n100) );
  INVD1BWP12T U281 ( .I(n100), .ZN(n114) );
  TPND2D0BWP12T U282 ( .A1(n113), .A2(n88), .ZN(n90) );
  AN3XD1BWP12T U283 ( .A1(n114), .A2(n125), .A3(n90), .Z(n1307) );
  NR2D0BWP12T U284 ( .A1(n89), .A2(write2_sel[2]), .ZN(n92) );
  INVD1BWP12T U285 ( .I(n90), .ZN(n91) );
  AOI211D1BWP12T U286 ( .A1(n114), .A2(n92), .B(reset), .C(n91), .ZN(n1306) );
  AO222D0BWP12T U287 ( .A1(n1308), .A2(n1238), .B1(n1307), .B2(write2_in[18]), 
        .C1(n1306), .C2(r11[18]), .Z(n2283) );
  AO222D0BWP12T U288 ( .A1(n1317), .A2(write1_in[21]), .B1(n820), .B2(
        write2_in[21]), .C1(n819), .C2(tmp1[21]), .Z(n2158) );
  AO222D0BWP12T U289 ( .A1(n1305), .A2(write1_in[21]), .B1(n1303), .B2(r7[21]), 
        .C1(write2_in[21]), .C2(n1304), .Z(n2414) );
  AO222D0BWP12T U290 ( .A1(n1299), .A2(write1_in[21]), .B1(n1297), .B2(r5[21]), 
        .C1(write2_in[21]), .C2(n1298), .Z(n2478) );
  AO222D0BWP12T U291 ( .A1(n1284), .A2(write1_in[21]), .B1(n1282), .B2(r6[21]), 
        .C1(write2_in[21]), .C2(n1283), .Z(n2446) );
  ND2D1BWP12T U292 ( .A1(n113), .A2(n93), .ZN(n1328) );
  INVD1BWP12T U293 ( .I(n1328), .ZN(n1330) );
  AN2XD0BWP12T U294 ( .A1(write2_in[5]), .A2(n1328), .Z(n94) );
  AN2XD0BWP12T U295 ( .A1(write2_in[3]), .A2(n1328), .Z(n95) );
  CKND2D0BWP12T U296 ( .A1(write2_in[2]), .A2(n1328), .ZN(n96) );
  IOA21D1BWP12T U297 ( .A1(write1_in[2]), .A2(n1330), .B(n96), .ZN(n108) );
  CKND2D0BWP12T U298 ( .A1(write2_in[1]), .A2(n1328), .ZN(n97) );
  IOA21D2BWP12T U299 ( .A1(write1_in[1]), .A2(n1330), .B(n97), .ZN(n430) );
  TPNR2D1BWP12T U300 ( .A1(n107), .A2(n106), .ZN(n105) );
  CKND2D0BWP12T U301 ( .A1(write2_in[4]), .A2(n1328), .ZN(n98) );
  IOA21D2BWP12T U302 ( .A1(write1_in[4]), .A2(n1330), .B(n98), .ZN(n104) );
  CKND2D2BWP12T U303 ( .A1(n105), .A2(n104), .ZN(n372) );
  OAI21D1BWP12T U304 ( .A1(n100), .A2(n99), .B(n1328), .ZN(n101) );
  INVD1BWP12T U305 ( .I(n101), .ZN(n431) );
  OR2XD1BWP12T U306 ( .A1(n431), .A2(reset), .Z(n1334) );
  INVD2BWP12T U307 ( .I(n1334), .ZN(n1363) );
  NR2D1BWP12T U308 ( .A1(n101), .A2(reset), .ZN(n103) );
  INVD1BWP12T U309 ( .I(n103), .ZN(n102) );
  NR2D1BWP12T U310 ( .A1(next_pc_en_BAR), .A2(n102), .ZN(n1362) );
  BUFFD1BWP12T U311 ( .I(n1362), .Z(n1355) );
  AN2D1BWP12T U312 ( .A1(next_pc_en_BAR), .A2(n103), .Z(n1361) );
  AO222D0BWP12T U313 ( .A1(n1308), .A2(write1_in[21]), .B1(n1307), .B2(
        write2_in[21]), .C1(n1306), .C2(r11[21]), .Z(n2286) );
  AO222D0BWP12T U314 ( .A1(n1314), .A2(write1_in[21]), .B1(n1313), .B2(
        write2_in[21]), .C1(n1312), .C2(r10[21]), .Z(n2318) );
  AO222D0BWP12T U315 ( .A1(n1281), .A2(write1_in[21]), .B1(n1279), .B2(r12[21]), .C1(write2_in[21]), .C2(n1280), .Z(n2254) );
  AO222D0BWP12T U316 ( .A1(n1287), .A2(write1_in[21]), .B1(n1285), .B2(lr[21]), 
        .C1(write2_in[21]), .C2(n1286), .Z(n2222) );
  AO222D0BWP12T U317 ( .A1(n1296), .A2(write1_in[21]), .B1(n1294), .B2(r4[21]), 
        .C1(write2_in[21]), .C2(n1295), .Z(n2510) );
  AO222D0BWP12T U318 ( .A1(n1317), .A2(write1_in[12]), .B1(n820), .B2(
        write2_in[12]), .C1(n819), .C2(tmp1[12]), .Z(n2149) );
  AO222D0BWP12T U319 ( .A1(n1317), .A2(write1_in[11]), .B1(n820), .B2(
        write2_in[11]), .C1(n819), .C2(tmp1[11]), .Z(n2148) );
  AO222D0BWP12T U320 ( .A1(n1296), .A2(write1_in[0]), .B1(n1294), .B2(r4[0]), 
        .C1(write2_in[0]), .C2(n1295), .Z(n2489) );
  AO222D0BWP12T U321 ( .A1(n1287), .A2(write1_in[0]), .B1(n1285), .B2(lr[0]), 
        .C1(write2_in[0]), .C2(n1286), .Z(n2201) );
  ND2D1BWP12T U322 ( .A1(n113), .A2(n109), .ZN(n451) );
  INVD1BWP12T U323 ( .I(n451), .ZN(n1316) );
  CKND2D1BWP12T U324 ( .A1(n114), .A2(n110), .ZN(n112) );
  ND2D1BWP12T U325 ( .A1(n451), .A2(n138), .ZN(n111) );
  AO222D0BWP12T U326 ( .A1(n1316), .A2(write1_in[0]), .B1(n421), .B2(n[2041]), 
        .C1(write2_in[0]), .C2(n1315), .Z(spin[0]) );
  INR3D0BWP12T U327 ( .A1(n138), .B1(write1_sel[2]), .B2(write1_sel[1]), .ZN(
        n134) );
  ND2D1BWP12T U328 ( .A1(n113), .A2(n134), .ZN(n465) );
  INVD1BWP12T U329 ( .I(n465), .ZN(n1293) );
  NR2D1BWP12T U330 ( .A1(write2_sel[2]), .A2(write2_sel[1]), .ZN(n136) );
  CKND2D1BWP12T U331 ( .A1(n114), .A2(n136), .ZN(n116) );
  ND2D1BWP12T U332 ( .A1(n465), .A2(n138), .ZN(n115) );
  NR2D1BWP12T U333 ( .A1(n116), .A2(n115), .ZN(n1292) );
  AO222D0BWP12T U334 ( .A1(n1293), .A2(write1_in[0]), .B1(n1291), .B2(r9[0]), 
        .C1(write2_in[0]), .C2(n1292), .Z(n2329) );
  ND2D1BWP12T U335 ( .A1(n119), .A2(n134), .ZN(n482) );
  INVD1BWP12T U336 ( .I(n482), .ZN(n1278) );
  CKND2D1BWP12T U337 ( .A1(n120), .A2(n136), .ZN(n118) );
  ND2D1BWP12T U338 ( .A1(n482), .A2(n138), .ZN(n117) );
  NR2D1BWP12T U339 ( .A1(n118), .A2(n117), .ZN(n1277) );
  AO222D0BWP12T U340 ( .A1(n1278), .A2(write1_in[0]), .B1(n1276), .B2(r0[0]), 
        .C1(write2_in[0]), .C2(n1277), .Z(n2617) );
  AO222D0BWP12T U341 ( .A1(n1308), .A2(write1_in[0]), .B1(n1307), .B2(
        write2_in[0]), .C1(n1306), .C2(r11[0]), .Z(n2265) );
  INVD1BWP12T U342 ( .I(n119), .ZN(n121) );
  NR2D1BWP12T U343 ( .A1(n121), .A2(n124), .ZN(n1275) );
  CKND2D1BWP12T U344 ( .A1(n120), .A2(n125), .ZN(n122) );
  NR2D1BWP12T U345 ( .A1(n121), .A2(n126), .ZN(n123) );
  NR2D1BWP12T U346 ( .A1(n122), .A2(n123), .ZN(n1274) );
  AO222D0BWP12T U347 ( .A1(n1275), .A2(write1_in[0]), .B1(n1274), .B2(
        write2_in[0]), .C1(n1273), .C2(r2[0]), .Z(n2553) );
  AO222D0BWP12T U348 ( .A1(n1305), .A2(write1_in[0]), .B1(n1303), .B2(r7[0]), 
        .C1(write2_in[0]), .C2(n1304), .Z(n2393) );
  AO222D0BWP12T U349 ( .A1(n1317), .A2(write1_in[0]), .B1(n820), .B2(
        write2_in[0]), .C1(n819), .C2(tmp1[0]), .Z(n2136) );
  INVD1BWP12T U350 ( .I(n135), .ZN(n127) );
  NR2D1BWP12T U351 ( .A1(n127), .A2(n124), .ZN(n1311) );
  CKND2D1BWP12T U352 ( .A1(n137), .A2(n125), .ZN(n128) );
  NR2D1BWP12T U353 ( .A1(n127), .A2(n126), .ZN(n129) );
  NR2D1BWP12T U354 ( .A1(n128), .A2(n129), .ZN(n1310) );
  AO222D0BWP12T U355 ( .A1(n1311), .A2(write1_in[0]), .B1(n1310), .B2(
        write2_in[0]), .C1(n1309), .C2(r3[0]), .Z(n2521) );
  ND2D1BWP12T U356 ( .A1(n134), .A2(n130), .ZN(n459) );
  INVD1BWP12T U357 ( .I(n459), .ZN(n1290) );
  CKND2D1BWP12T U358 ( .A1(n131), .A2(n136), .ZN(n133) );
  ND2D1BWP12T U359 ( .A1(n459), .A2(n138), .ZN(n132) );
  NR2D1BWP12T U360 ( .A1(n133), .A2(n132), .ZN(n1289) );
  AO222D0BWP12T U361 ( .A1(n1290), .A2(write1_in[0]), .B1(n1288), .B2(r8[0]), 
        .C1(write2_in[0]), .C2(n1289), .Z(n2361) );
  AO222D0BWP12T U362 ( .A1(n1281), .A2(write1_in[0]), .B1(n1279), .B2(r12[0]), 
        .C1(write2_in[0]), .C2(n1280), .Z(n2233) );
  AO222D0BWP12T U363 ( .A1(n1314), .A2(write1_in[0]), .B1(n1313), .B2(
        write2_in[0]), .C1(n1312), .C2(r10[0]), .Z(n2297) );
  ND2D1BWP12T U364 ( .A1(n135), .A2(n134), .ZN(n462) );
  INVD1BWP12T U365 ( .I(n462), .ZN(n1302) );
  CKND2D1BWP12T U366 ( .A1(n137), .A2(n136), .ZN(n140) );
  ND2D1BWP12T U367 ( .A1(n462), .A2(n138), .ZN(n139) );
  NR2D1BWP12T U368 ( .A1(n140), .A2(n139), .ZN(n1301) );
  AO222D0BWP12T U369 ( .A1(n1302), .A2(write1_in[0]), .B1(n1300), .B2(r1[0]), 
        .C1(write2_in[0]), .C2(n1301), .Z(n2585) );
  AO222D0BWP12T U370 ( .A1(n1299), .A2(write1_in[0]), .B1(n1297), .B2(r5[0]), 
        .C1(write2_in[0]), .C2(n1298), .Z(n2457) );
  AO222D0BWP12T U371 ( .A1(n1284), .A2(write1_in[0]), .B1(n1282), .B2(r6[0]), 
        .C1(write2_in[0]), .C2(n1283), .Z(n2425) );
  INVD0BWP12T U372 ( .I(pc_out[13]), .ZN(n143) );
  ND2D1BWP12T U373 ( .A1(readA_sel[2]), .A2(readA_sel[1]), .ZN(n172) );
  INVD2BWP12T U374 ( .I(readA_sel[4]), .ZN(n147) );
  IND2XD2BWP12T U375 ( .A1(readA_sel[2]), .B1(readA_sel[1]), .ZN(n170) );
  INVD1BWP12T U376 ( .I(n170), .ZN(n145) );
  INR2D4BWP12T U377 ( .A1(n145), .B1(n165), .ZN(n1559) );
  INVD1BWP12T U378 ( .I(r11[13]), .ZN(n142) );
  OAI22D1BWP12T U379 ( .A1(n143), .A2(n1949), .B1(n1948), .B2(n142), .ZN(n162)
         );
  INVD1BWP12T U380 ( .I(lr[13]), .ZN(n1180) );
  INR2D4BWP12T U381 ( .A1(readA_sel[3]), .B1(readA_sel[0]), .ZN(n153) );
  CKND2D4BWP12T U382 ( .A1(n153), .A2(n147), .ZN(n164) );
  INR2D2BWP12T U383 ( .A1(n144), .B1(n164), .ZN(n1561) );
  INVD3BWP12T U384 ( .I(n1561), .ZN(n1953) );
  INR2D4BWP12T U385 ( .A1(n145), .B1(n164), .ZN(n1560) );
  INVD3BWP12T U386 ( .I(n1560), .ZN(n1952) );
  INVD1BWP12T U387 ( .I(r10[13]), .ZN(n146) );
  OAI22D1BWP12T U388 ( .A1(n1180), .A2(n1953), .B1(n1952), .B2(n146), .ZN(n161) );
  NR2D1BWP12T U389 ( .A1(readA_sel[0]), .A2(readA_sel[3]), .ZN(n148) );
  CKND2D2BWP12T U390 ( .A1(n148), .A2(n147), .ZN(n175) );
  INVD1BWP12T U391 ( .I(n175), .ZN(n149) );
  INR2D2BWP12T U392 ( .A1(readA_sel[2]), .B1(readA_sel[1]), .ZN(n167) );
  CKND2D2BWP12T U393 ( .A1(n149), .A2(n167), .ZN(n1458) );
  DCCKND8BWP12T U394 ( .I(n1458), .ZN(n1957) );
  BUFFXD8BWP12T U395 ( .I(n521), .Z(n1809) );
  AOI22D1BWP12T U396 ( .A1(n150), .A2(r12[13]), .B1(n1809), .B2(tmp1[13]), 
        .ZN(n154) );
  IOA21D1BWP12T U397 ( .A1(n1957), .A2(r4[13]), .B(n154), .ZN(n160) );
  INVD1BWP12T U398 ( .I(r2[13]), .ZN(n158) );
  TPNR2D2BWP12T U399 ( .A1(readA_sel[2]), .A2(readA_sel[1]), .ZN(n176) );
  TPNR2D1BWP12T U400 ( .A1(readA_sel[4]), .A2(readA_sel[3]), .ZN(n156) );
  CKND2D2BWP12T U401 ( .A1(n156), .A2(readA_sel[0]), .ZN(n173) );
  INR2XD2BWP12T U402 ( .A1(n176), .B1(n173), .ZN(n1555) );
  INVD1BWP12T U403 ( .I(r1[13]), .ZN(n157) );
  OAI22D1BWP12T U404 ( .A1(n1961), .A2(n158), .B1(n1959), .B2(n157), .ZN(n159)
         );
  NR4D0BWP12T U405 ( .A1(n162), .A2(n161), .A3(n160), .A4(n159), .ZN(n182) );
  INR2D8BWP12T U406 ( .A1(n176), .B1(n165), .ZN(n1591) );
  NR2D1BWP12T U407 ( .A1(n175), .A2(n172), .ZN(n163) );
  BUFFD3BWP12T U408 ( .I(n163), .Z(n1590) );
  AOI22D1BWP12T U409 ( .A1(r9[13]), .A2(n1591), .B1(n1590), .B2(r6[13]), .ZN(
        n180) );
  INR2D2BWP12T U410 ( .A1(n176), .B1(n164), .ZN(n1593) );
  INR2D2BWP12T U411 ( .A1(n167), .B1(n165), .ZN(n166) );
  BUFFD2BWP12T U412 ( .I(n166), .Z(n1592) );
  AOI22D1BWP12T U413 ( .A1(r8[13]), .A2(n1593), .B1(n1592), .B2(n[2028]), .ZN(
        n179) );
  INVD1BWP12T U414 ( .I(n167), .ZN(n168) );
  NR2D1BWP12T U415 ( .A1(n173), .A2(n168), .ZN(n169) );
  BUFFD6BWP12T U416 ( .I(n169), .Z(n1594) );
  AOI22D1BWP12T U417 ( .A1(r5[13]), .A2(n1594), .B1(n171), .B2(r3[13]), .ZN(
        n178) );
  NR2D1BWP12T U418 ( .A1(n173), .A2(n172), .ZN(n174) );
  BUFFXD4BWP12T U419 ( .I(n174), .Z(n1596) );
  INR2XD2BWP12T U420 ( .A1(n176), .B1(n175), .ZN(n1595) );
  AOI22D1BWP12T U421 ( .A1(r7[13]), .A2(n1596), .B1(n1595), .B2(r0[13]), .ZN(
        n177) );
  AN4XD1BWP12T U422 ( .A1(n180), .A2(n179), .A3(n178), .A4(n177), .Z(n181) );
  NR2XD3BWP12T U423 ( .A1(readB_sel[1]), .A2(readB_sel[2]), .ZN(n204) );
  IND3D4BWP12T U424 ( .A1(readB_sel[3]), .B1(readB_sel[0]), .B2(n189), .ZN(
        n213) );
  INR2D1BWP12T U425 ( .A1(readB_sel[2]), .B1(readB_sel[1]), .ZN(n209) );
  IND3D2BWP12T U426 ( .A1(readB_sel[0]), .B1(readB_sel[3]), .B2(n189), .ZN(
        n211) );
  INR2D1BWP12T U427 ( .A1(n209), .B1(n211), .ZN(n184) );
  BUFFD6BWP12T U428 ( .I(n184), .Z(n1992) );
  AOI22D1BWP12T U429 ( .A1(r1[23]), .A2(n183), .B1(n1992), .B2(r12[23]), .ZN(
        n195) );
  INR2D2BWP12T U430 ( .A1(readB_sel[1]), .B1(readB_sel[2]), .ZN(n216) );
  INR2D1BWP12T U431 ( .A1(n214), .B1(n211), .ZN(n186) );
  BUFFD6BWP12T U432 ( .I(n186), .Z(n1993) );
  AOI22D1BWP12T U433 ( .A1(r3[23]), .A2(n185), .B1(n1993), .B2(lr[23]), .ZN(
        n194) );
  ND3XD4BWP12T U434 ( .A1(n189), .A2(readB_sel[3]), .A3(readB_sel[0]), .ZN(
        n203) );
  AOI22D1BWP12T U435 ( .A1(r8[23]), .A2(n187), .B1(n1994), .B2(n[2018]), .ZN(
        n193) );
  TPNR2D2BWP12T U436 ( .A1(readB_sel[3]), .A2(readB_sel[0]), .ZN(n190) );
  TPND2D3BWP12T U437 ( .A1(n190), .A2(n189), .ZN(n218) );
  INVD1BWP12T U438 ( .I(n214), .ZN(n191) );
  NR2D3BWP12T U439 ( .A1(n218), .A2(n191), .ZN(n1995) );
  AOI22D1BWP12T U440 ( .A1(pc_out[23]), .A2(n188), .B1(n1995), .B2(r6[23]), 
        .ZN(n192) );
  AN4XD1BWP12T U441 ( .A1(n195), .A2(n194), .A3(n193), .A4(n192), .Z(n222) );
  INVD1BWP12T U442 ( .I(readB_sel[0]), .ZN(n198) );
  INVD1BWP12T U443 ( .I(readB_sel[3]), .ZN(n196) );
  INR2D1BWP12T U444 ( .A1(readB_sel[4]), .B1(n196), .ZN(n197) );
  TPND2D2BWP12T U445 ( .A1(n214), .A2(n197), .ZN(n199) );
  INR2XD2BWP12T U446 ( .A1(n198), .B1(n199), .ZN(n2000) );
  AOI22D1BWP12T U447 ( .A1(tmp1[23]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[23]), .ZN(n208) );
  INVD1BWP12T U448 ( .I(n209), .ZN(n202) );
  BUFFD3BWP12T U449 ( .I(n536), .Z(n2001) );
  AOI22D1BWP12T U450 ( .A1(r9[23]), .A2(n201), .B1(n2001), .B2(r4[23]), .ZN(
        n207) );
  INR2D1BWP12T U451 ( .A1(n216), .B1(n203), .ZN(n537) );
  BUFFD2BWP12T U452 ( .I(n537), .Z(n1470) );
  AOI22D1BWP12T U453 ( .A1(r11[23]), .A2(n1470), .B1(n205), .B2(r0[23]), .ZN(
        n206) );
  AN3XD1BWP12T U454 ( .A1(n208), .A2(n207), .A3(n206), .Z(n221) );
  INR2D1BWP12T U455 ( .A1(n216), .B1(n211), .ZN(n212) );
  BUFFXD4BWP12T U456 ( .I(n212), .Z(n1988) );
  AOI22D1BWP12T U457 ( .A1(r5[23]), .A2(n210), .B1(n1988), .B2(r10[23]), .ZN(
        n220) );
  INVD1BWP12T U458 ( .I(n216), .ZN(n217) );
  TPNR2D2BWP12T U459 ( .A1(n218), .A2(n217), .ZN(n1989) );
  AOI22D1BWP12T U460 ( .A1(r7[23]), .A2(n215), .B1(n1989), .B2(r2[23]), .ZN(
        n219) );
  AOI22D1BWP12T U461 ( .A1(r1[24]), .A2(n183), .B1(n1992), .B2(r12[24]), .ZN(
        n226) );
  AOI22D1BWP12T U462 ( .A1(r3[24]), .A2(n185), .B1(n1993), .B2(lr[24]), .ZN(
        n225) );
  AOI22D1BWP12T U463 ( .A1(r8[24]), .A2(n187), .B1(n1994), .B2(n[2017]), .ZN(
        n224) );
  AOI22D1BWP12T U464 ( .A1(pc_out[24]), .A2(n188), .B1(n1995), .B2(r6[24]), 
        .ZN(n223) );
  AN4XD1BWP12T U465 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .Z(n233) );
  AOI22D1BWP12T U466 ( .A1(tmp1[24]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[24]), .ZN(n229) );
  AOI22D0BWP12T U467 ( .A1(r9[24]), .A2(n201), .B1(n2001), .B2(r4[24]), .ZN(
        n228) );
  AOI22D1BWP12T U468 ( .A1(r11[24]), .A2(n1470), .B1(n205), .B2(r0[24]), .ZN(
        n227) );
  AN3XD1BWP12T U469 ( .A1(n229), .A2(n228), .A3(n227), .Z(n232) );
  AOI22D1BWP12T U470 ( .A1(r5[24]), .A2(n210), .B1(n1988), .B2(r10[24]), .ZN(
        n231) );
  AOI22D1BWP12T U471 ( .A1(r7[24]), .A2(n215), .B1(n1989), .B2(r2[24]), .ZN(
        n230) );
  INVD1BWP12T U472 ( .I(r4[26]), .ZN(n236) );
  BUFFXD8BWP12T U473 ( .I(n521), .Z(n1486) );
  AOI22D1BWP12T U474 ( .A1(n150), .A2(r12[26]), .B1(n1486), .B2(tmp1[26]), 
        .ZN(n235) );
  AOI22D1BWP12T U475 ( .A1(r2[26]), .A2(n155), .B1(n1555), .B2(r1[26]), .ZN(
        n234) );
  AOI22D1BWP12T U476 ( .A1(r9[26]), .A2(n1591), .B1(n1590), .B2(r6[26]), .ZN(
        n240) );
  AOI22D1BWP12T U477 ( .A1(r8[26]), .A2(n1593), .B1(n1592), .B2(n[2015]), .ZN(
        n239) );
  AOI22D1BWP12T U478 ( .A1(r5[26]), .A2(n1594), .B1(n171), .B2(r3[26]), .ZN(
        n238) );
  AOI22D1BWP12T U479 ( .A1(r7[26]), .A2(n1596), .B1(n1595), .B2(r0[26]), .ZN(
        n237) );
  AN4XD1BWP12T U480 ( .A1(n240), .A2(n239), .A3(n238), .A4(n237), .Z(n243) );
  AOI22D1BWP12T U481 ( .A1(pc_out[26]), .A2(n141), .B1(n1559), .B2(r11[26]), 
        .ZN(n242) );
  AOI22D1BWP12T U482 ( .A1(lr[26]), .A2(n1561), .B1(n1560), .B2(r10[26]), .ZN(
        n241) );
  ND4D2BWP12T U483 ( .A1(n244), .A2(n243), .A3(n242), .A4(n241), .ZN(
        regA_out[26]) );
  INVD1BWP12T U484 ( .I(tmp1[8]), .ZN(n245) );
  CKND3BWP12T U485 ( .I(n2000), .ZN(n1847) );
  MOAI22D0BWP12T U486 ( .A1(n245), .A2(n1847), .B1(n200), .B2(immediate2_in[8]), .ZN(n251) );
  AOI22D1BWP12T U487 ( .A1(r9[8]), .A2(n201), .B1(n1780), .B2(r4[8]), .ZN(n247) );
  BUFFD2BWP12T U488 ( .I(n537), .Z(n2002) );
  AOI22D1BWP12T U489 ( .A1(r11[8]), .A2(n2002), .B1(n205), .B2(r0[8]), .ZN(
        n246) );
  ND2D1BWP12T U490 ( .A1(n247), .A2(n246), .ZN(n250) );
  INVD1BWP12T U491 ( .I(r5[8]), .ZN(n1756) );
  INVD4BWP12T U492 ( .I(n210), .ZN(n1846) );
  INVD4BWP12T U493 ( .I(n1988), .ZN(n1845) );
  INVD1BWP12T U494 ( .I(r10[8]), .ZN(n1742) );
  OAI22D1BWP12T U495 ( .A1(n1756), .A2(n1846), .B1(n1845), .B2(n1742), .ZN(
        n249) );
  DCCKND8BWP12T U496 ( .I(n215), .ZN(n1852) );
  INVD1BWP12T U497 ( .I(r7[8]), .ZN(n1758) );
  INVD1BWP12T U498 ( .I(r2[8]), .ZN(n1746) );
  OAI22D1BWP12T U499 ( .A1(n1852), .A2(n1758), .B1(n1851), .B2(n1746), .ZN(
        n248) );
  NR4D0BWP12T U500 ( .A1(n251), .A2(n250), .A3(n249), .A4(n248), .ZN(n257) );
  INVD1BWP12T U501 ( .I(r1[8]), .ZN(n1745) );
  INVD3BWP12T U502 ( .I(n183), .ZN(n1859) );
  INVD4BWP12T U503 ( .I(n1992), .ZN(n1858) );
  INVD1BWP12T U504 ( .I(r12[8]), .ZN(n960) );
  OAI22D1BWP12T U505 ( .A1(n1745), .A2(n1859), .B1(n1858), .B2(n960), .ZN(n255) );
  INVD1BWP12T U506 ( .I(r3[8]), .ZN(n1755) );
  INVD4BWP12T U507 ( .I(n1993), .ZN(n1860) );
  INVD1BWP12T U508 ( .I(lr[8]), .ZN(n1743) );
  OAI22D1BWP12T U509 ( .A1(n1755), .A2(n1861), .B1(n1860), .B2(n1743), .ZN(
        n254) );
  INVD3BWP12T U510 ( .I(n187), .ZN(n1863) );
  INVD1BWP12T U511 ( .I(r8[8]), .ZN(n1754) );
  DCCKND8BWP12T U512 ( .I(n1994), .ZN(n1862) );
  INVD1BWP12T U513 ( .I(n[2033]), .ZN(n1753) );
  OAI22D1BWP12T U514 ( .A1(n1863), .A2(n1754), .B1(n1862), .B2(n1753), .ZN(
        n253) );
  INVD6BWP12T U515 ( .I(n188), .ZN(n1865) );
  INVD1BWP12T U516 ( .I(pc_out[8]), .ZN(n1741) );
  INVD1BWP12T U517 ( .I(r6[8]), .ZN(n1751) );
  OAI22D1BWP12T U518 ( .A1(n1865), .A2(n1741), .B1(n1864), .B2(n1751), .ZN(
        n252) );
  NR4D0BWP12T U519 ( .A1(n255), .A2(n254), .A3(n253), .A4(n252), .ZN(n256) );
  CKND2D1BWP12T U520 ( .A1(n257), .A2(n256), .ZN(regB_out[8]) );
  AOI22D1BWP12T U521 ( .A1(r1[22]), .A2(n183), .B1(n1992), .B2(r12[22]), .ZN(
        n261) );
  AOI22D1BWP12T U522 ( .A1(r3[22]), .A2(n185), .B1(n1993), .B2(lr[22]), .ZN(
        n260) );
  AOI22D1BWP12T U523 ( .A1(r8[22]), .A2(n187), .B1(n1994), .B2(n[2019]), .ZN(
        n259) );
  AOI22D1BWP12T U524 ( .A1(pc_out[22]), .A2(n188), .B1(n1995), .B2(r6[22]), 
        .ZN(n258) );
  AN4XD1BWP12T U525 ( .A1(n261), .A2(n260), .A3(n259), .A4(n258), .Z(n268) );
  AOI22D1BWP12T U526 ( .A1(tmp1[22]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[22]), .ZN(n264) );
  AOI22D1BWP12T U527 ( .A1(r9[22]), .A2(n201), .B1(n2001), .B2(r4[22]), .ZN(
        n263) );
  AOI22D1BWP12T U528 ( .A1(r11[22]), .A2(n1470), .B1(n205), .B2(r0[22]), .ZN(
        n262) );
  AN3XD1BWP12T U529 ( .A1(n264), .A2(n263), .A3(n262), .Z(n267) );
  AOI22D1BWP12T U530 ( .A1(r5[22]), .A2(n210), .B1(n1988), .B2(r10[22]), .ZN(
        n266) );
  AOI22D1BWP12T U531 ( .A1(r7[22]), .A2(n215), .B1(n1989), .B2(r2[22]), .ZN(
        n265) );
  INVD1BWP12T U532 ( .I(tmp1[10]), .ZN(n269) );
  MOAI22D0BWP12T U533 ( .A1(n269), .A2(n1847), .B1(n200), .B2(
        immediate2_in[10]), .ZN(n275) );
  AOI22D1BWP12T U534 ( .A1(r9[10]), .A2(n201), .B1(n1780), .B2(r4[10]), .ZN(
        n271) );
  AOI22D1BWP12T U535 ( .A1(r11[10]), .A2(n2002), .B1(n205), .B2(r0[10]), .ZN(
        n270) );
  ND2D1BWP12T U536 ( .A1(n271), .A2(n270), .ZN(n274) );
  INVD1BWP12T U537 ( .I(r5[10]), .ZN(n1694) );
  INVD1BWP12T U538 ( .I(r10[10]), .ZN(n1680) );
  OAI22D1BWP12T U539 ( .A1(n1694), .A2(n1846), .B1(n1845), .B2(n1680), .ZN(
        n273) );
  INVD1BWP12T U540 ( .I(r7[10]), .ZN(n1696) );
  INVD1BWP12T U541 ( .I(r2[10]), .ZN(n1684) );
  OAI22D1BWP12T U542 ( .A1(n1852), .A2(n1696), .B1(n1851), .B2(n1684), .ZN(
        n272) );
  NR4D0BWP12T U543 ( .A1(n275), .A2(n274), .A3(n273), .A4(n272), .ZN(n281) );
  INVD1BWP12T U544 ( .I(r1[10]), .ZN(n1683) );
  INVD1BWP12T U545 ( .I(r12[10]), .ZN(n400) );
  OAI22D0BWP12T U546 ( .A1(n1683), .A2(n1859), .B1(n1858), .B2(n400), .ZN(n279) );
  INVD1BWP12T U547 ( .I(r3[10]), .ZN(n1693) );
  INVD1BWP12T U548 ( .I(lr[10]), .ZN(n1681) );
  OAI22D1BWP12T U549 ( .A1(n1693), .A2(n1861), .B1(n1860), .B2(n1681), .ZN(
        n278) );
  INVD1BWP12T U550 ( .I(r8[10]), .ZN(n1692) );
  INVD1BWP12T U551 ( .I(n[2031]), .ZN(n1691) );
  OAI22D1BWP12T U552 ( .A1(n1863), .A2(n1692), .B1(n1862), .B2(n1691), .ZN(
        n277) );
  INVD1BWP12T U553 ( .I(pc_out[10]), .ZN(n1679) );
  INVD1BWP12T U554 ( .I(r6[10]), .ZN(n1689) );
  OAI22D1BWP12T U555 ( .A1(n1865), .A2(n1679), .B1(n1864), .B2(n1689), .ZN(
        n276) );
  NR4D0BWP12T U556 ( .A1(n279), .A2(n278), .A3(n277), .A4(n276), .ZN(n280) );
  CKND2D1BWP12T U557 ( .A1(n281), .A2(n280), .ZN(regB_out[10]) );
  INVD1BWP12T U558 ( .I(tmp1[12]), .ZN(n282) );
  MOAI22D0BWP12T U559 ( .A1(n282), .A2(n1847), .B1(n200), .B2(
        immediate2_in[12]), .ZN(n288) );
  AOI22D1BWP12T U560 ( .A1(r9[12]), .A2(n201), .B1(n1780), .B2(r4[12]), .ZN(
        n284) );
  AOI22D1BWP12T U561 ( .A1(r11[12]), .A2(n2002), .B1(n205), .B2(r0[12]), .ZN(
        n283) );
  ND2D1BWP12T U562 ( .A1(n284), .A2(n283), .ZN(n287) );
  INVD1BWP12T U563 ( .I(r5[12]), .ZN(n1645) );
  INVD1BWP12T U564 ( .I(r10[12]), .ZN(n1631) );
  OAI22D1BWP12T U565 ( .A1(n1645), .A2(n1846), .B1(n1845), .B2(n1631), .ZN(
        n286) );
  INVD1BWP12T U566 ( .I(r7[12]), .ZN(n1647) );
  INVD1BWP12T U567 ( .I(r2[12]), .ZN(n1635) );
  OAI22D1BWP12T U568 ( .A1(n1852), .A2(n1647), .B1(n1851), .B2(n1635), .ZN(
        n285) );
  NR4D0BWP12T U569 ( .A1(n288), .A2(n287), .A3(n286), .A4(n285), .ZN(n294) );
  INVD1BWP12T U570 ( .I(r1[12]), .ZN(n1634) );
  INVD1BWP12T U571 ( .I(r12[12]), .ZN(n887) );
  OAI22D1BWP12T U572 ( .A1(n1634), .A2(n1859), .B1(n1858), .B2(n887), .ZN(n292) );
  INVD1BWP12T U573 ( .I(r3[12]), .ZN(n1644) );
  INVD1BWP12T U574 ( .I(lr[12]), .ZN(n1632) );
  OAI22D1BWP12T U575 ( .A1(n1644), .A2(n1861), .B1(n1860), .B2(n1632), .ZN(
        n291) );
  INVD1BWP12T U576 ( .I(r8[12]), .ZN(n1643) );
  INVD1BWP12T U577 ( .I(n[2029]), .ZN(n1642) );
  OAI22D1BWP12T U578 ( .A1(n1863), .A2(n1643), .B1(n1862), .B2(n1642), .ZN(
        n290) );
  INVD1BWP12T U579 ( .I(pc_out[12]), .ZN(n1630) );
  INVD1BWP12T U580 ( .I(r6[12]), .ZN(n1640) );
  OAI22D1BWP12T U581 ( .A1(n1865), .A2(n1630), .B1(n1864), .B2(n1640), .ZN(
        n289) );
  NR4D0BWP12T U582 ( .A1(n292), .A2(n291), .A3(n290), .A4(n289), .ZN(n293) );
  ND2D1BWP12T U583 ( .A1(n294), .A2(n293), .ZN(regB_out[12]) );
  AOI22D1BWP12T U584 ( .A1(r1[21]), .A2(n183), .B1(n1992), .B2(r12[21]), .ZN(
        n298) );
  AOI22D1BWP12T U585 ( .A1(r3[21]), .A2(n185), .B1(n1993), .B2(lr[21]), .ZN(
        n297) );
  AOI22D1BWP12T U586 ( .A1(r8[21]), .A2(n187), .B1(n1994), .B2(n[2020]), .ZN(
        n296) );
  AOI22D1BWP12T U587 ( .A1(pc_out[21]), .A2(n188), .B1(n1995), .B2(r6[21]), 
        .ZN(n295) );
  AN4XD1BWP12T U588 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .Z(n305) );
  AOI22D1BWP12T U589 ( .A1(tmp1[21]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[21]), .ZN(n301) );
  AOI22D1BWP12T U590 ( .A1(r9[21]), .A2(n201), .B1(n2001), .B2(r4[21]), .ZN(
        n300) );
  AOI22D1BWP12T U591 ( .A1(r11[21]), .A2(n1470), .B1(n205), .B2(r0[21]), .ZN(
        n299) );
  AN3XD1BWP12T U592 ( .A1(n301), .A2(n300), .A3(n299), .Z(n304) );
  AOI22D1BWP12T U593 ( .A1(r5[21]), .A2(n210), .B1(n1988), .B2(r10[21]), .ZN(
        n303) );
  AOI22D1BWP12T U594 ( .A1(r7[21]), .A2(n215), .B1(n1989), .B2(r2[21]), .ZN(
        n302) );
  ND4D2BWP12T U595 ( .A1(n305), .A2(n304), .A3(n303), .A4(n302), .ZN(
        regB_out[21]) );
  NR2D1BWP12T U596 ( .A1(readD_sel[1]), .A2(readD_sel[0]), .ZN(n319) );
  INVD1BWP12T U597 ( .I(n319), .ZN(n310) );
  IND2D1BWP12T U598 ( .A1(readD_sel[2]), .B1(readD_sel[3]), .ZN(n309) );
  NR2D1BWP12T U599 ( .A1(n310), .A2(n309), .ZN(n726) );
  IND2D1BWP12T U600 ( .A1(readD_sel[3]), .B1(readD_sel[2]), .ZN(n308) );
  NR2D1BWP12T U601 ( .A1(n310), .A2(n308), .ZN(n725) );
  AOI22D0BWP12T U602 ( .A1(r8[9]), .A2(n726), .B1(n725), .B2(r4[9]), .ZN(n307)
         );
  ND2D1BWP12T U603 ( .A1(readD_sel[3]), .A2(readD_sel[2]), .ZN(n321) );
  IND2D1BWP12T U604 ( .A1(readD_sel[1]), .B1(readD_sel[0]), .ZN(n315) );
  NR2D1BWP12T U605 ( .A1(n321), .A2(n315), .ZN(n728) );
  IND2D1BWP12T U606 ( .A1(readD_sel[0]), .B1(readD_sel[1]), .ZN(n317) );
  NR2D1BWP12T U607 ( .A1(n309), .A2(n317), .ZN(n727) );
  AOI22D0BWP12T U608 ( .A1(n[2032]), .A2(n728), .B1(n727), .B2(r10[9]), .ZN(
        n306) );
  CKND2D1BWP12T U609 ( .A1(n307), .A2(n306), .ZN(n326) );
  ND2D1BWP12T U610 ( .A1(readD_sel[1]), .A2(readD_sel[0]), .ZN(n320) );
  NR2D1BWP12T U611 ( .A1(n320), .A2(n308), .ZN(n732) );
  NR2D1BWP12T U612 ( .A1(n315), .A2(n308), .ZN(n731) );
  AOI22D0BWP12T U613 ( .A1(r7[9]), .A2(n732), .B1(n731), .B2(r5[9]), .ZN(n314)
         );
  NR2D1BWP12T U614 ( .A1(n321), .A2(n317), .ZN(n734) );
  NR2D1BWP12T U615 ( .A1(n309), .A2(n315), .ZN(n733) );
  AOI22D0BWP12T U616 ( .A1(lr[9]), .A2(n734), .B1(n733), .B2(r9[9]), .ZN(n313)
         );
  NR2D1BWP12T U617 ( .A1(n317), .A2(n308), .ZN(n736) );
  NR2D1BWP12T U618 ( .A1(n309), .A2(n320), .ZN(n735) );
  AOI22D0BWP12T U619 ( .A1(r6[9]), .A2(n736), .B1(n735), .B2(r11[9]), .ZN(n312) );
  NR2D1BWP12T U620 ( .A1(n321), .A2(n310), .ZN(n737) );
  CKND2D0BWP12T U621 ( .A1(n737), .A2(r12[9]), .ZN(n311) );
  ND4D1BWP12T U622 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .ZN(n325) );
  INVD1BWP12T U623 ( .I(r1[9]), .ZN(n1727) );
  NR2D1BWP12T U624 ( .A1(readD_sel[3]), .A2(readD_sel[2]), .ZN(n318) );
  INVD1BWP12T U625 ( .I(n318), .ZN(n316) );
  OR2XD1BWP12T U626 ( .A1(n315), .A2(n316), .Z(n748) );
  NR2D1BWP12T U627 ( .A1(n320), .A2(n316), .ZN(n743) );
  NR2D1BWP12T U628 ( .A1(n317), .A2(n316), .ZN(n742) );
  AOI22D0BWP12T U629 ( .A1(r3[9]), .A2(n743), .B1(n742), .B2(r2[9]), .ZN(n323)
         );
  AN2XD1BWP12T U630 ( .A1(n319), .A2(n318), .Z(n745) );
  NR2D1BWP12T U631 ( .A1(n321), .A2(n320), .ZN(n744) );
  AOI22D0BWP12T U632 ( .A1(n745), .A2(r0[9]), .B1(pc_out[9]), .B2(n744), .ZN(
        n322) );
  OAI211D0BWP12T U633 ( .A1(n1727), .A2(n748), .B(n323), .C(n322), .ZN(n324)
         );
  INVD1BWP12T U634 ( .I(readD_sel[4]), .ZN(n749) );
  OA31D0BWP12T U635 ( .A1(n326), .A2(n325), .A3(n324), .B(n749), .Z(
        regD_out[9]) );
  AOI22D0BWP12T U636 ( .A1(r8[10]), .A2(n726), .B1(n725), .B2(r4[10]), .ZN(
        n328) );
  AOI22D0BWP12T U637 ( .A1(n[2031]), .A2(n728), .B1(n727), .B2(r10[10]), .ZN(
        n327) );
  CKND2D1BWP12T U638 ( .A1(n328), .A2(n327), .ZN(n337) );
  AOI22D0BWP12T U639 ( .A1(r7[10]), .A2(n732), .B1(n731), .B2(r5[10]), .ZN(
        n332) );
  AOI22D0BWP12T U640 ( .A1(lr[10]), .A2(n734), .B1(n733), .B2(r9[10]), .ZN(
        n331) );
  AOI22D0BWP12T U641 ( .A1(r6[10]), .A2(n736), .B1(n735), .B2(r11[10]), .ZN(
        n330) );
  CKND2D0BWP12T U642 ( .A1(n737), .A2(r12[10]), .ZN(n329) );
  ND4D1BWP12T U643 ( .A1(n332), .A2(n331), .A3(n330), .A4(n329), .ZN(n336) );
  AOI22D0BWP12T U644 ( .A1(r3[10]), .A2(n743), .B1(n742), .B2(r2[10]), .ZN(
        n334) );
  AOI22D0BWP12T U645 ( .A1(n745), .A2(r0[10]), .B1(pc_out[10]), .B2(n744), 
        .ZN(n333) );
  OAI211D0BWP12T U646 ( .A1(n1683), .A2(n748), .B(n334), .C(n333), .ZN(n335)
         );
  OA31D0BWP12T U647 ( .A1(n337), .A2(n336), .A3(n335), .B(n749), .Z(
        regD_out[10]) );
  AOI22D0BWP12T U648 ( .A1(r8[11]), .A2(n726), .B1(n725), .B2(r4[11]), .ZN(
        n339) );
  AOI22D0BWP12T U649 ( .A1(n[2030]), .A2(n728), .B1(n727), .B2(r10[11]), .ZN(
        n338) );
  CKND2D1BWP12T U650 ( .A1(n339), .A2(n338), .ZN(n348) );
  AOI22D0BWP12T U651 ( .A1(r7[11]), .A2(n732), .B1(n731), .B2(r5[11]), .ZN(
        n343) );
  AOI22D0BWP12T U652 ( .A1(lr[11]), .A2(n734), .B1(n733), .B2(r9[11]), .ZN(
        n342) );
  AOI22D0BWP12T U653 ( .A1(r6[11]), .A2(n736), .B1(n735), .B2(r11[11]), .ZN(
        n341) );
  CKND2D0BWP12T U654 ( .A1(n737), .A2(r12[11]), .ZN(n340) );
  ND4D1BWP12T U655 ( .A1(n343), .A2(n342), .A3(n341), .A4(n340), .ZN(n347) );
  INVD1BWP12T U656 ( .I(r1[11]), .ZN(n1659) );
  AOI22D0BWP12T U657 ( .A1(r3[11]), .A2(n743), .B1(n742), .B2(r2[11]), .ZN(
        n345) );
  AOI22D0BWP12T U658 ( .A1(n745), .A2(r0[11]), .B1(pc_out[11]), .B2(n744), 
        .ZN(n344) );
  OAI211D0BWP12T U659 ( .A1(n1659), .A2(n748), .B(n345), .C(n344), .ZN(n346)
         );
  OA31D0BWP12T U660 ( .A1(n348), .A2(n347), .A3(n346), .B(n749), .Z(
        regD_out[11]) );
  AOI22D0BWP12T U661 ( .A1(r8[12]), .A2(n726), .B1(n725), .B2(r4[12]), .ZN(
        n350) );
  AOI22D0BWP12T U662 ( .A1(n[2029]), .A2(n728), .B1(n727), .B2(r10[12]), .ZN(
        n349) );
  CKND2D1BWP12T U663 ( .A1(n350), .A2(n349), .ZN(n359) );
  AOI22D0BWP12T U664 ( .A1(r7[12]), .A2(n732), .B1(n731), .B2(r5[12]), .ZN(
        n354) );
  AOI22D0BWP12T U665 ( .A1(lr[12]), .A2(n734), .B1(n733), .B2(r9[12]), .ZN(
        n353) );
  AOI22D0BWP12T U666 ( .A1(r6[12]), .A2(n736), .B1(n735), .B2(r11[12]), .ZN(
        n352) );
  CKND2D0BWP12T U667 ( .A1(n737), .A2(r12[12]), .ZN(n351) );
  ND4D1BWP12T U668 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .ZN(n358) );
  AOI22D0BWP12T U669 ( .A1(r3[12]), .A2(n743), .B1(n742), .B2(r2[12]), .ZN(
        n356) );
  AOI22D0BWP12T U670 ( .A1(n745), .A2(r0[12]), .B1(pc_out[12]), .B2(n744), 
        .ZN(n355) );
  OAI211D0BWP12T U671 ( .A1(n1634), .A2(n748), .B(n356), .C(n355), .ZN(n357)
         );
  OA31D0BWP12T U672 ( .A1(n359), .A2(n358), .A3(n357), .B(n749), .Z(
        regD_out[12]) );
  AN2XD0BWP12T U673 ( .A1(write2_in[28]), .A2(n1328), .Z(n360) );
  TPAOI21D1BWP12T U674 ( .A1(n1268), .A2(n1330), .B(n360), .ZN(n1353) );
  INVD1BWP12T U675 ( .I(n1353), .ZN(n381) );
  CKND2D0BWP12T U676 ( .A1(write2_in[25]), .A2(n1328), .ZN(n361) );
  IOA21D2BWP12T U677 ( .A1(write1_in[25]), .A2(n1330), .B(n361), .ZN(n1357) );
  BUFFD6BWP12T U678 ( .I(write1_in[24]), .Z(n1254) );
  CKAN2D1BWP12T U679 ( .A1(write2_in[24]), .A2(n1328), .Z(n362) );
  TPAOI21D8BWP12T U680 ( .A1(n1254), .A2(n1330), .B(n362), .ZN(n1342) );
  BUFFD2BWP12T U681 ( .I(write1_in[23]), .Z(n1253) );
  AN2XD0BWP12T U682 ( .A1(write2_in[23]), .A2(n1328), .Z(n363) );
  TPAOI21D4BWP12T U683 ( .A1(n1253), .A2(n1330), .B(n363), .ZN(n1323) );
  TPNR2D2BWP12T U684 ( .A1(n1342), .A2(n1323), .ZN(n364) );
  TPND2D2BWP12T U685 ( .A1(n1357), .A2(n364), .ZN(n379) );
  BUFFXD8BWP12T U686 ( .I(write1_in[26]), .Z(n1263) );
  AN2XD0BWP12T U687 ( .A1(write2_in[26]), .A2(n1328), .Z(n365) );
  AOI21D1BWP12T U688 ( .A1(n1263), .A2(n1330), .B(n365), .ZN(n1359) );
  BUFFD2BWP12T U689 ( .I(write1_in[20]), .Z(n1245) );
  CKND2D0BWP12T U690 ( .A1(write2_in[20]), .A2(n1328), .ZN(n366) );
  IOA21D1BWP12T U691 ( .A1(n1245), .A2(n1330), .B(n366), .ZN(n1270) );
  CKND2D0BWP12T U692 ( .A1(write2_in[16]), .A2(n1328), .ZN(n367) );
  IOA21D1BWP12T U693 ( .A1(n1232), .A2(n1330), .B(n367), .ZN(n1256) );
  CKND2D0BWP12T U694 ( .A1(write2_in[12]), .A2(n1328), .ZN(n368) );
  IOA21D1BWP12T U695 ( .A1(write1_in[12]), .A2(n1330), .B(n368), .ZN(n1244) );
  AN2XD0BWP12T U696 ( .A1(write2_in[9]), .A2(n1328), .Z(n369) );
  AOI21D1BWP12T U697 ( .A1(write1_in[9]), .A2(n1330), .B(n369), .ZN(n1235) );
  AN2XD0BWP12T U698 ( .A1(write2_in[7]), .A2(n1328), .Z(n370) );
  AOI21D1BWP12T U699 ( .A1(write1_in[7]), .A2(n1330), .B(n370), .ZN(n1229) );
  CKND2D0BWP12T U700 ( .A1(write2_in[6]), .A2(n1328), .ZN(n371) );
  IOA21D1BWP12T U701 ( .A1(write1_in[6]), .A2(n1330), .B(n371), .ZN(n1227) );
  TPNR2D1BWP12T U702 ( .A1(n373), .A2(n372), .ZN(n1226) );
  TPND2D1BWP12T U703 ( .A1(n1227), .A2(n1226), .ZN(n1228) );
  TPNR2D1BWP12T U704 ( .A1(n1229), .A2(n1228), .ZN(n1230) );
  TPND2D1BWP12T U705 ( .A1(n1231), .A2(n1230), .ZN(n1234) );
  NR2D2BWP12T U706 ( .A1(n1235), .A2(n1234), .ZN(n1237) );
  TPND2D2BWP12T U707 ( .A1(n1237), .A2(n1236), .ZN(n1240) );
  TPNR2D3BWP12T U708 ( .A1(n1241), .A2(n1240), .ZN(n1243) );
  AN2XD0BWP12T U709 ( .A1(write2_in[13]), .A2(n1328), .Z(n374) );
  AOI21D1BWP12T U710 ( .A1(write1_in[13]), .A2(n1330), .B(n374), .ZN(n1246) );
  BUFFD2BWP12T U711 ( .I(write1_in[15]), .Z(n1233) );
  AN2XD0BWP12T U712 ( .A1(write2_in[15]), .A2(n1328), .Z(n375) );
  TPAOI21D4BWP12T U713 ( .A1(n1233), .A2(n1330), .B(n375), .ZN(n1251) );
  AN2XD0BWP12T U714 ( .A1(write2_in[17]), .A2(n1328), .Z(n376) );
  AOI21D1BWP12T U715 ( .A1(n54), .A2(n1330), .B(n376), .ZN(n1258) );
  CKND2D0BWP12T U716 ( .A1(write2_in[18]), .A2(n1328), .ZN(n377) );
  IOA21D1BWP12T U717 ( .A1(n1238), .A2(n1330), .B(n377), .ZN(n1261) );
  TPND2D2BWP12T U718 ( .A1(n1262), .A2(n1261), .ZN(n1266) );
  BUFFD2BWP12T U719 ( .I(write1_in[19]), .Z(n1242) );
  AN2XD0BWP12T U720 ( .A1(write2_in[19]), .A2(n1328), .Z(n378) );
  AOI21D1BWP12T U721 ( .A1(n1242), .A2(n1330), .B(n378), .ZN(n1265) );
  TPNR2D2BWP12T U722 ( .A1(n1266), .A2(n1265), .ZN(n1269) );
  TPND2D2BWP12T U723 ( .A1(n1270), .A2(n1269), .ZN(n1272) );
  TPNR2D3BWP12T U724 ( .A1(n1272), .A2(n1271), .ZN(n1319) );
  BUFFD3BWP12T U725 ( .I(write1_in[22]), .Z(n1250) );
  TPND2D3BWP12T U726 ( .A1(n1319), .A2(n1318), .ZN(n1324) );
  TPNR3D2BWP12T U727 ( .A1(n379), .A2(n1359), .A3(n1324), .ZN(n1321) );
  BUFFXD8BWP12T U728 ( .I(write1_in[27]), .Z(n1264) );
  CKND2D0BWP12T U729 ( .A1(write2_in[27]), .A2(n1328), .ZN(n380) );
  IOA21D2BWP12T U730 ( .A1(n1264), .A2(n1330), .B(n380), .ZN(n1320) );
  TPND2D2BWP12T U731 ( .A1(n1321), .A2(n1320), .ZN(n1354) );
  BUFFD2BWP12T U732 ( .I(write1_in[29]), .Z(n1267) );
  MUX2D1BWP12T U733 ( .I0(n1267), .I1(write2_in[29]), .S(n1328), .Z(n1346) );
  AOI22D1BWP12T U734 ( .A1(next_pc_in[29]), .A2(n1355), .B1(n1361), .B2(
        pc_out[29]), .ZN(n382) );
  RCOAI21D1BWP12T U735 ( .A1(n383), .A2(n1334), .B(n382), .ZN(n2198) );
  AO222D0BWP12T U736 ( .A1(n1316), .A2(n1238), .B1(n421), .B2(n[2023]), .C1(
        write2_in[18]), .C2(n1315), .Z(spin[18]) );
  AO222D0BWP12T U737 ( .A1(n1316), .A2(write1_in[21]), .B1(n421), .B2(n[2020]), 
        .C1(write2_in[21]), .C2(n1315), .Z(spin[21]) );
  INVD1BWP12T U738 ( .I(r9[12]), .ZN(n1641) );
  INVD1BWP12T U739 ( .I(n1291), .ZN(n466) );
  INVD1BWP12T U740 ( .I(write1_in[12]), .ZN(n387) );
  INVD1BWP12T U741 ( .I(write2_in[12]), .ZN(n388) );
  INVD1BWP12T U742 ( .I(n1292), .ZN(n464) );
  OAI222D0BWP12T U743 ( .A1(n1641), .A2(n466), .B1(n387), .B2(n465), .C1(n388), 
        .C2(n464), .ZN(n2341) );
  INVD1BWP12T U744 ( .I(n1282), .ZN(n469) );
  INVD1BWP12T U745 ( .I(n1283), .ZN(n467) );
  OAI222D0BWP12T U746 ( .A1(n1640), .A2(n469), .B1(n387), .B2(n468), .C1(n388), 
        .C2(n467), .ZN(n2437) );
  INVD1BWP12T U747 ( .I(n1300), .ZN(n463) );
  INVD1BWP12T U748 ( .I(n1301), .ZN(n461) );
  OAI222D0BWP12T U749 ( .A1(n1634), .A2(n463), .B1(n387), .B2(n462), .C1(n388), 
        .C2(n461), .ZN(n2597) );
  INVD0BWP12T U750 ( .I(r4[12]), .ZN(n384) );
  INVD1BWP12T U751 ( .I(n1294), .ZN(n472) );
  INVD1BWP12T U752 ( .I(n1295), .ZN(n470) );
  OAI222D0BWP12T U753 ( .A1(n384), .A2(n472), .B1(n387), .B2(n471), .C1(n388), 
        .C2(n470), .ZN(n2501) );
  INVD1BWP12T U754 ( .I(n1307), .ZN(n476) );
  INVD1BWP12T U755 ( .I(n1308), .ZN(n475) );
  INVD1BWP12T U756 ( .I(n1306), .ZN(n474) );
  INVD1BWP12T U757 ( .I(r11[12]), .ZN(n1629) );
  OAI222D0BWP12T U758 ( .A1(n388), .A2(n476), .B1(n387), .B2(n475), .C1(n474), 
        .C2(n1629), .ZN(n2277) );
  AOI21D0BWP12T U759 ( .A1(n421), .A2(n[2029]), .B(reset), .ZN(n386) );
  CKND2D0BWP12T U760 ( .A1(write2_in[12]), .A2(n1315), .ZN(n385) );
  OAI211D0BWP12T U761 ( .A1(n451), .A2(n387), .B(n386), .C(n385), .ZN(spin[12]) );
  INVD1BWP12T U762 ( .I(n1285), .ZN(n479) );
  INVD1BWP12T U763 ( .I(n1286), .ZN(n477) );
  OAI222D0BWP12T U764 ( .A1(n1632), .A2(n479), .B1(n387), .B2(n478), .C1(n388), 
        .C2(n477), .ZN(n2213) );
  INVD1BWP12T U765 ( .I(n1279), .ZN(n445) );
  INVD1BWP12T U766 ( .I(n1280), .ZN(n443) );
  OAI222D0BWP12T U767 ( .A1(n887), .A2(n445), .B1(n387), .B2(n444), .C1(n388), 
        .C2(n443), .ZN(n2245) );
  INVD1BWP12T U768 ( .I(n1274), .ZN(n488) );
  INVD1BWP12T U769 ( .I(n1275), .ZN(n486) );
  INVD1BWP12T U770 ( .I(n1273), .ZN(n485) );
  OAI222D0BWP12T U771 ( .A1(n388), .A2(n488), .B1(n387), .B2(n486), .C1(n485), 
        .C2(n1635), .ZN(n2565) );
  INVD1BWP12T U772 ( .I(n1314), .ZN(n447) );
  INVD1BWP12T U773 ( .I(n1312), .ZN(n446) );
  OAI222D0BWP12T U774 ( .A1(n388), .A2(n448), .B1(n387), .B2(n447), .C1(n446), 
        .C2(n1631), .ZN(n2309) );
  INVD1BWP12T U775 ( .I(r0[12]), .ZN(n1646) );
  INVD1BWP12T U776 ( .I(n1276), .ZN(n484) );
  INVD1BWP12T U777 ( .I(n1277), .ZN(n480) );
  OAI222D0BWP12T U778 ( .A1(n1646), .A2(n484), .B1(n387), .B2(n482), .C1(n388), 
        .C2(n480), .ZN(n2629) );
  INVD1BWP12T U779 ( .I(n1288), .ZN(n460) );
  INVD1BWP12T U780 ( .I(n1289), .ZN(n458) );
  OAI222D0BWP12T U781 ( .A1(n1643), .A2(n460), .B1(n387), .B2(n459), .C1(n388), 
        .C2(n458), .ZN(n2373) );
  INVD1BWP12T U782 ( .I(n1303), .ZN(n442) );
  INVD1BWP12T U783 ( .I(n1304), .ZN(n440) );
  OAI222D0BWP12T U784 ( .A1(n1647), .A2(n442), .B1(n387), .B2(n441), .C1(n388), 
        .C2(n440), .ZN(n2405) );
  INVD1BWP12T U785 ( .I(n1297), .ZN(n454) );
  INVD1BWP12T U786 ( .I(n1298), .ZN(n452) );
  OAI222D0BWP12T U787 ( .A1(n1645), .A2(n454), .B1(n387), .B2(n453), .C1(n388), 
        .C2(n452), .ZN(n2469) );
  INVD1BWP12T U788 ( .I(n1310), .ZN(n457) );
  INVD1BWP12T U789 ( .I(n1311), .ZN(n456) );
  INVD1BWP12T U790 ( .I(n1309), .ZN(n455) );
  OAI222D0BWP12T U791 ( .A1(n388), .A2(n457), .B1(n387), .B2(n456), .C1(n455), 
        .C2(n1644), .ZN(n2533) );
  CKND0BWP12T U792 ( .I(r4[11]), .ZN(n389) );
  INVD1BWP12T U793 ( .I(write1_in[11]), .ZN(n408) );
  INVD1BWP12T U794 ( .I(write2_in[11]), .ZN(n407) );
  OAI222D0BWP12T U795 ( .A1(n389), .A2(n472), .B1(n408), .B2(n471), .C1(n407), 
        .C2(n470), .ZN(n2500) );
  AOI21D0BWP12T U796 ( .A1(n421), .A2(n[2030]), .B(reset), .ZN(n391) );
  CKND2D0BWP12T U797 ( .A1(write2_in[11]), .A2(n1315), .ZN(n390) );
  OAI211D0BWP12T U798 ( .A1(n451), .A2(n408), .B(n391), .C(n390), .ZN(spin[11]) );
  INVD1BWP12T U799 ( .I(r7[7]), .ZN(n1786) );
  INVD1BWP12T U800 ( .I(write1_in[7]), .ZN(n403) );
  INVD1BWP12T U801 ( .I(write2_in[7]), .ZN(n404) );
  OAI222D0BWP12T U802 ( .A1(n1786), .A2(n442), .B1(n403), .B2(n441), .C1(n404), 
        .C2(n440), .ZN(n2400) );
  INVD1BWP12T U803 ( .I(r10[7]), .ZN(n1783) );
  OAI222D0BWP12T U804 ( .A1(n404), .A2(n448), .B1(n403), .B2(n447), .C1(n446), 
        .C2(n1783), .ZN(n2304) );
  INVD0BWP12T U805 ( .I(r4[10]), .ZN(n1155) );
  INVD1BWP12T U806 ( .I(write1_in[10]), .ZN(n406) );
  INVD1BWP12T U807 ( .I(write2_in[10]), .ZN(n405) );
  OAI222D0BWP12T U808 ( .A1(n1155), .A2(n472), .B1(n406), .B2(n471), .C1(n405), 
        .C2(n470), .ZN(n2499) );
  INVD1BWP12T U809 ( .I(r12[11]), .ZN(n1121) );
  OAI222D0BWP12T U810 ( .A1(n1121), .A2(n445), .B1(n408), .B2(n444), .C1(n407), 
        .C2(n443), .ZN(n2244) );
  INVD1BWP12T U811 ( .I(r7[5]), .ZN(n1915) );
  INVD1BWP12T U812 ( .I(write1_in[5]), .ZN(n402) );
  INVD1BWP12T U813 ( .I(write2_in[5]), .ZN(n401) );
  OAI222D0BWP12T U814 ( .A1(n1915), .A2(n442), .B1(n402), .B2(n441), .C1(n401), 
        .C2(n440), .ZN(n2398) );
  OAI222D0BWP12T U815 ( .A1(n405), .A2(n488), .B1(n406), .B2(n486), .C1(n485), 
        .C2(n1684), .ZN(n2563) );
  INVD1BWP12T U816 ( .I(r2[11]), .ZN(n1660) );
  OAI222D0BWP12T U817 ( .A1(n407), .A2(n488), .B1(n408), .B2(n486), .C1(n485), 
        .C2(n1660), .ZN(n2564) );
  CKND0BWP12T U818 ( .I(r4[7]), .ZN(n392) );
  OAI222D0BWP12T U819 ( .A1(n392), .A2(n472), .B1(n403), .B2(n471), .C1(n404), 
        .C2(n470), .ZN(n2496) );
  AOI21D0BWP12T U820 ( .A1(n421), .A2(n[2031]), .B(reset), .ZN(n394) );
  CKND2D0BWP12T U821 ( .A1(write2_in[10]), .A2(n1315), .ZN(n393) );
  OAI211D0BWP12T U822 ( .A1(n451), .A2(n406), .B(n394), .C(n393), .ZN(spin[10]) );
  INVD1BWP12T U823 ( .I(r5[5]), .ZN(n1913) );
  OAI222D0BWP12T U824 ( .A1(n1913), .A2(n454), .B1(n402), .B2(n453), .C1(n401), 
        .C2(n452), .ZN(n2462) );
  CKND0BWP12T U825 ( .I(r4[5]), .ZN(n395) );
  OAI222D0BWP12T U826 ( .A1(n395), .A2(n472), .B1(n402), .B2(n471), .C1(n401), 
        .C2(n470), .ZN(n2494) );
  INVD1BWP12T U827 ( .I(r5[7]), .ZN(n1784) );
  OAI222D0BWP12T U828 ( .A1(n1784), .A2(n454), .B1(n403), .B2(n453), .C1(n404), 
        .C2(n452), .ZN(n2464) );
  INVD1BWP12T U829 ( .I(r12[7]), .ZN(n1791) );
  OAI222D0BWP12T U830 ( .A1(n1791), .A2(n445), .B1(n403), .B2(n444), .C1(n404), 
        .C2(n443), .ZN(n2240) );
  OAI222D0BWP12T U831 ( .A1(n1694), .A2(n454), .B1(n406), .B2(n453), .C1(n405), 
        .C2(n452), .ZN(n2467) );
  INVD1BWP12T U832 ( .I(r5[11]), .ZN(n1670) );
  OAI222D0BWP12T U833 ( .A1(n1670), .A2(n454), .B1(n408), .B2(n453), .C1(n407), 
        .C2(n452), .ZN(n2468) );
  AOI21D0BWP12T U834 ( .A1(n421), .A2(n[2034]), .B(reset), .ZN(n397) );
  CKND2D0BWP12T U835 ( .A1(write2_in[7]), .A2(n1315), .ZN(n396) );
  OAI211D0BWP12T U836 ( .A1(n451), .A2(n403), .B(n397), .C(n396), .ZN(spin[7])
         );
  INVD1BWP12T U837 ( .I(r3[11]), .ZN(n1669) );
  OAI222D0BWP12T U838 ( .A1(n407), .A2(n457), .B1(n408), .B2(n456), .C1(n455), 
        .C2(n1669), .ZN(n2532) );
  OAI222D0BWP12T U839 ( .A1(n405), .A2(n457), .B1(n406), .B2(n456), .C1(n455), 
        .C2(n1693), .ZN(n2531) );
  INVD1BWP12T U840 ( .I(r8[5]), .ZN(n1911) );
  OAI222D0BWP12T U841 ( .A1(n1911), .A2(n460), .B1(n402), .B2(n459), .C1(n401), 
        .C2(n458), .ZN(n2366) );
  INVD1BWP12T U842 ( .I(r10[11]), .ZN(n1656) );
  OAI222D0BWP12T U843 ( .A1(n407), .A2(n448), .B1(n408), .B2(n447), .C1(n446), 
        .C2(n1656), .ZN(n2308) );
  INVD1BWP12T U844 ( .I(r8[7]), .ZN(n1796) );
  OAI222D0BWP12T U845 ( .A1(n1796), .A2(n460), .B1(n403), .B2(n459), .C1(n404), 
        .C2(n458), .ZN(n2368) );
  OAI222D0BWP12T U846 ( .A1(n405), .A2(n448), .B1(n406), .B2(n447), .C1(n446), 
        .C2(n1680), .ZN(n2307) );
  INVD1BWP12T U847 ( .I(r3[5]), .ZN(n1912) );
  OAI222D0BWP12T U848 ( .A1(n401), .A2(n457), .B1(n402), .B2(n456), .C1(n455), 
        .C2(n1912), .ZN(n2526) );
  OAI222D0BWP12T U849 ( .A1(n1692), .A2(n460), .B1(n406), .B2(n459), .C1(n405), 
        .C2(n458), .ZN(n2371) );
  INVD1BWP12T U850 ( .I(r10[5]), .ZN(n1899) );
  OAI222D0BWP12T U851 ( .A1(n401), .A2(n448), .B1(n402), .B2(n447), .C1(n446), 
        .C2(n1899), .ZN(n2302) );
  AOI21D0BWP12T U852 ( .A1(n421), .A2(n[2036]), .B(reset), .ZN(n399) );
  CKND2D0BWP12T U853 ( .A1(write2_in[5]), .A2(n1315), .ZN(n398) );
  OAI211D0BWP12T U854 ( .A1(n451), .A2(n402), .B(n399), .C(n398), .ZN(spin[5])
         );
  INVD1BWP12T U855 ( .I(r12[5]), .ZN(n1838) );
  OAI222D0BWP12T U856 ( .A1(n1838), .A2(n445), .B1(n402), .B2(n444), .C1(n401), 
        .C2(n443), .ZN(n2238) );
  INVD1BWP12T U857 ( .I(r8[11]), .ZN(n1668) );
  OAI222D0BWP12T U858 ( .A1(n1668), .A2(n460), .B1(n408), .B2(n459), .C1(n407), 
        .C2(n458), .ZN(n2372) );
  INVD1BWP12T U859 ( .I(r3[7]), .ZN(n1794) );
  OAI222D0BWP12T U860 ( .A1(n404), .A2(n457), .B1(n403), .B2(n456), .C1(n455), 
        .C2(n1794), .ZN(n2528) );
  INVD1BWP12T U861 ( .I(r0[5]), .ZN(n1914) );
  OAI222D0BWP12T U862 ( .A1(n1914), .A2(n484), .B1(n402), .B2(n482), .C1(n401), 
        .C2(n480), .ZN(n2622) );
  INVD1BWP12T U863 ( .I(r1[7]), .ZN(n1792) );
  OAI222D0BWP12T U864 ( .A1(n1792), .A2(n463), .B1(n403), .B2(n462), .C1(n404), 
        .C2(n461), .ZN(n2592) );
  INVD1BWP12T U865 ( .I(r9[10]), .ZN(n1690) );
  OAI222D0BWP12T U866 ( .A1(n1690), .A2(n466), .B1(n406), .B2(n465), .C1(n405), 
        .C2(n464), .ZN(n2339) );
  INVD1BWP12T U867 ( .I(r11[10]), .ZN(n1678) );
  OAI222D0BWP12T U868 ( .A1(n405), .A2(n476), .B1(n406), .B2(n475), .C1(n474), 
        .C2(n1678), .ZN(n2275) );
  INVD1BWP12T U869 ( .I(lr[7]), .ZN(n1793) );
  OAI222D0BWP12T U870 ( .A1(n1793), .A2(n479), .B1(n403), .B2(n478), .C1(n404), 
        .C2(n477), .ZN(n2208) );
  INVD1BWP12T U871 ( .I(r11[11]), .ZN(n1654) );
  OAI222D0BWP12T U872 ( .A1(n407), .A2(n476), .B1(n408), .B2(n475), .C1(n474), 
        .C2(n1654), .ZN(n2276) );
  OAI222D0BWP12T U873 ( .A1(n1683), .A2(n463), .B1(n406), .B2(n462), .C1(n405), 
        .C2(n461), .ZN(n2595) );
  INVD1BWP12T U874 ( .I(r9[11]), .ZN(n1666) );
  OAI222D0BWP12T U875 ( .A1(n1666), .A2(n466), .B1(n408), .B2(n465), .C1(n407), 
        .C2(n464), .ZN(n2340) );
  INVD1BWP12T U876 ( .I(r0[10]), .ZN(n1695) );
  OAI222D0BWP12T U877 ( .A1(n1695), .A2(n484), .B1(n406), .B2(n482), .C1(n405), 
        .C2(n480), .ZN(n2627) );
  OAI222D0BWP12T U878 ( .A1(n1681), .A2(n479), .B1(n406), .B2(n478), .C1(n405), 
        .C2(n477), .ZN(n2211) );
  INVD1BWP12T U879 ( .I(r11[7]), .ZN(n1765) );
  OAI222D0BWP12T U880 ( .A1(n404), .A2(n476), .B1(n403), .B2(n475), .C1(n474), 
        .C2(n1765), .ZN(n2272) );
  INVD1BWP12T U881 ( .I(lr[11]), .ZN(n1657) );
  OAI222D0BWP12T U882 ( .A1(n1657), .A2(n479), .B1(n408), .B2(n478), .C1(n407), 
        .C2(n477), .ZN(n2212) );
  INVD1BWP12T U883 ( .I(r0[11]), .ZN(n1671) );
  OAI222D0BWP12T U884 ( .A1(n1671), .A2(n484), .B1(n408), .B2(n482), .C1(n407), 
        .C2(n480), .ZN(n2628) );
  INVD1BWP12T U885 ( .I(r9[7]), .ZN(n1771) );
  OAI222D0BWP12T U886 ( .A1(n1771), .A2(n466), .B1(n403), .B2(n465), .C1(n404), 
        .C2(n464), .ZN(n2336) );
  INVD1BWP12T U887 ( .I(r6[11]), .ZN(n1665) );
  OAI222D0BWP12T U888 ( .A1(n1665), .A2(n469), .B1(n408), .B2(n468), .C1(n407), 
        .C2(n467), .ZN(n2436) );
  INVD1BWP12T U889 ( .I(lr[5]), .ZN(n1900) );
  OAI222D0BWP12T U890 ( .A1(n1900), .A2(n479), .B1(n402), .B2(n478), .C1(n401), 
        .C2(n477), .ZN(n2206) );
  INVD1BWP12T U891 ( .I(r0[7]), .ZN(n1772) );
  OAI222D0BWP12T U892 ( .A1(n1772), .A2(n484), .B1(n403), .B2(n482), .C1(n404), 
        .C2(n480), .ZN(n2624) );
  INVD1BWP12T U893 ( .I(r2[5]), .ZN(n1903) );
  OAI222D0BWP12T U894 ( .A1(n401), .A2(n488), .B1(n402), .B2(n486), .C1(n485), 
        .C2(n1903), .ZN(n2558) );
  INVD1BWP12T U895 ( .I(r6[5]), .ZN(n1908) );
  OAI222D0BWP12T U896 ( .A1(n1908), .A2(n469), .B1(n402), .B2(n468), .C1(n401), 
        .C2(n467), .ZN(n2430) );
  INVD1BWP12T U897 ( .I(r9[5]), .ZN(n1909) );
  OAI222D0BWP12T U898 ( .A1(n1909), .A2(n466), .B1(n402), .B2(n465), .C1(n401), 
        .C2(n464), .ZN(n2334) );
  INVD1BWP12T U899 ( .I(r6[7]), .ZN(n1797) );
  OAI222D0BWP12T U900 ( .A1(n1797), .A2(n469), .B1(n403), .B2(n468), .C1(n404), 
        .C2(n467), .ZN(n2432) );
  INVD1BWP12T U901 ( .I(r11[5]), .ZN(n1897) );
  OAI222D0BWP12T U902 ( .A1(n401), .A2(n476), .B1(n402), .B2(n475), .C1(n474), 
        .C2(n1897), .ZN(n2270) );
  OAI222D0BWP12T U903 ( .A1(n400), .A2(n445), .B1(n406), .B2(n444), .C1(n405), 
        .C2(n443), .ZN(n2243) );
  OAI222D0BWP12T U904 ( .A1(n1696), .A2(n442), .B1(n406), .B2(n441), .C1(n405), 
        .C2(n440), .ZN(n2403) );
  OAI222D0BWP12T U905 ( .A1(n1659), .A2(n463), .B1(n408), .B2(n462), .C1(n407), 
        .C2(n461), .ZN(n2596) );
  INVD1BWP12T U906 ( .I(r1[5]), .ZN(n1902) );
  OAI222D0BWP12T U907 ( .A1(n1902), .A2(n463), .B1(n402), .B2(n462), .C1(n401), 
        .C2(n461), .ZN(n2590) );
  INVD1BWP12T U908 ( .I(r2[7]), .ZN(n1785) );
  OAI222D0BWP12T U909 ( .A1(n404), .A2(n488), .B1(n403), .B2(n486), .C1(n485), 
        .C2(n1785), .ZN(n2560) );
  OAI222D0BWP12T U910 ( .A1(n1689), .A2(n469), .B1(n406), .B2(n468), .C1(n405), 
        .C2(n467), .ZN(n2435) );
  INVD1BWP12T U911 ( .I(r7[11]), .ZN(n1672) );
  OAI222D0BWP12T U912 ( .A1(n1672), .A2(n442), .B1(n408), .B2(n441), .C1(n407), 
        .C2(n440), .ZN(n2404) );
  INVD1BWP12T U913 ( .I(lr[1]), .ZN(n1925) );
  INVD1BWP12T U914 ( .I(write1_in[1]), .ZN(n434) );
  INVD1BWP12T U915 ( .I(write2_in[1]), .ZN(n435) );
  OAI222D0BWP12T U916 ( .A1(n1925), .A2(n479), .B1(n434), .B2(n478), .C1(n435), 
        .C2(n477), .ZN(n2202) );
  INVD1BWP12T U917 ( .I(write1_in[8]), .ZN(n436) );
  INVD1BWP12T U918 ( .I(write2_in[8]), .ZN(n437) );
  OAI222D0BWP12T U919 ( .A1(n1751), .A2(n469), .B1(n436), .B2(n468), .C1(n437), 
        .C2(n467), .ZN(n2433) );
  INVD1BWP12T U920 ( .I(r7[1]), .ZN(n1940) );
  OAI222D0BWP12T U921 ( .A1(n1940), .A2(n442), .B1(n434), .B2(n441), .C1(n435), 
        .C2(n440), .ZN(n2394) );
  INVD1BWP12T U922 ( .I(r9[4]), .ZN(n1884) );
  INVD1BWP12T U923 ( .I(write1_in[4]), .ZN(n433) );
  INVD1BWP12T U924 ( .I(write2_in[4]), .ZN(n432) );
  OAI222D0BWP12T U925 ( .A1(n1884), .A2(n466), .B1(n433), .B2(n465), .C1(n432), 
        .C2(n464), .ZN(n2333) );
  AOI21D0BWP12T U926 ( .A1(n421), .A2(n[2040]), .B(reset), .ZN(n410) );
  CKND2D0BWP12T U927 ( .A1(write2_in[1]), .A2(n1315), .ZN(n409) );
  OAI211D0BWP12T U928 ( .A1(n451), .A2(n434), .B(n410), .C(n409), .ZN(spin[1])
         );
  INVD1BWP12T U929 ( .I(write1_in[3]), .ZN(n427) );
  AOI21D0BWP12T U930 ( .A1(n421), .A2(n[2038]), .B(reset), .ZN(n412) );
  CKND2D0BWP12T U931 ( .A1(write2_in[3]), .A2(n1315), .ZN(n411) );
  OAI211D0BWP12T U932 ( .A1(n451), .A2(n427), .B(n412), .C(n411), .ZN(spin[3])
         );
  AOI21D0BWP12T U933 ( .A1(n421), .A2(n[2037]), .B(reset), .ZN(n414) );
  CKND2D0BWP12T U934 ( .A1(write2_in[4]), .A2(n1315), .ZN(n413) );
  OAI211D0BWP12T U935 ( .A1(n451), .A2(n433), .B(n414), .C(n413), .ZN(spin[4])
         );
  INVD1BWP12T U936 ( .I(r9[3]), .ZN(n810) );
  INVD1BWP12T U937 ( .I(write2_in[3]), .ZN(n426) );
  OAI222D0BWP12T U938 ( .A1(n810), .A2(n466), .B1(n427), .B2(n465), .C1(n426), 
        .C2(n464), .ZN(n2332) );
  INVD1BWP12T U939 ( .I(write1_in[9]), .ZN(n424) );
  INVD1BWP12T U940 ( .I(write2_in[9]), .ZN(n425) );
  OAI222D0BWP12T U941 ( .A1(n1727), .A2(n463), .B1(n424), .B2(n462), .C1(n425), 
        .C2(n461), .ZN(n2594) );
  INVD1BWP12T U942 ( .I(r6[9]), .ZN(n1732) );
  OAI222D0BWP12T U943 ( .A1(n1732), .A2(n469), .B1(n424), .B2(n468), .C1(n425), 
        .C2(n467), .ZN(n2434) );
  INVD1BWP12T U944 ( .I(r7[3]), .ZN(n822) );
  OAI222D0BWP12T U945 ( .A1(n822), .A2(n442), .B1(n427), .B2(n441), .C1(n426), 
        .C2(n440), .ZN(n2396) );
  AO222D0BWP12T U946 ( .A1(n1317), .A2(write1_in[10]), .B1(n820), .B2(
        write2_in[10]), .C1(n819), .C2(tmp1[10]), .Z(n2147) );
  INVD1BWP12T U947 ( .I(r6[1]), .ZN(n1933) );
  OAI222D0BWP12T U948 ( .A1(n1933), .A2(n469), .B1(n434), .B2(n468), .C1(n435), 
        .C2(n467), .ZN(n2426) );
  INVD1BWP12T U949 ( .I(r9[8]), .ZN(n1752) );
  OAI222D0BWP12T U950 ( .A1(n1752), .A2(n466), .B1(n436), .B2(n465), .C1(n437), 
        .C2(n464), .ZN(n2337) );
  OAI222D0BWP12T U951 ( .A1(n1754), .A2(n460), .B1(n436), .B2(n459), .C1(n437), 
        .C2(n458), .ZN(n2369) );
  INVD1BWP12T U952 ( .I(r5[4]), .ZN(n1888) );
  OAI222D0BWP12T U953 ( .A1(n1888), .A2(n454), .B1(n433), .B2(n453), .C1(n432), 
        .C2(n452), .ZN(n2461) );
  INVD1BWP12T U954 ( .I(r9[9]), .ZN(n1707) );
  OAI222D0BWP12T U955 ( .A1(n1707), .A2(n466), .B1(n424), .B2(n465), .C1(n425), 
        .C2(n464), .ZN(n2338) );
  CKND0BWP12T U956 ( .I(r4[8]), .ZN(n415) );
  OAI222D0BWP12T U957 ( .A1(n415), .A2(n472), .B1(n436), .B2(n471), .C1(n437), 
        .C2(n470), .ZN(n2497) );
  INVD1BWP12T U958 ( .I(r0[1]), .ZN(n1939) );
  OAI222D0BWP12T U959 ( .A1(n1939), .A2(n484), .B1(n434), .B2(n482), .C1(n435), 
        .C2(n480), .ZN(n2618) );
  CKND0BWP12T U960 ( .I(r4[9]), .ZN(n416) );
  OAI222D0BWP12T U961 ( .A1(n416), .A2(n472), .B1(n424), .B2(n471), .C1(n425), 
        .C2(n470), .ZN(n2498) );
  INVD1BWP12T U962 ( .I(r0[9]), .ZN(n1708) );
  OAI222D0BWP12T U963 ( .A1(n1708), .A2(n484), .B1(n424), .B2(n482), .C1(n425), 
        .C2(n480), .ZN(n2626) );
  INVD1BWP12T U964 ( .I(r6[4]), .ZN(n1883) );
  OAI222D0BWP12T U965 ( .A1(n1883), .A2(n469), .B1(n433), .B2(n468), .C1(n432), 
        .C2(n467), .ZN(n2429) );
  INVD1BWP12T U966 ( .I(r8[9]), .ZN(n1731) );
  OAI222D0BWP12T U967 ( .A1(n1731), .A2(n460), .B1(n424), .B2(n459), .C1(n425), 
        .C2(n458), .ZN(n2370) );
  INVD1BWP12T U968 ( .I(r6[3]), .ZN(n827) );
  OAI222D0BWP12T U969 ( .A1(n827), .A2(n469), .B1(n427), .B2(n468), .C1(n426), 
        .C2(n467), .ZN(n2428) );
  INVD1BWP12T U970 ( .I(r5[3]), .ZN(n825) );
  OAI222D0BWP12T U971 ( .A1(n825), .A2(n454), .B1(n427), .B2(n453), .C1(n426), 
        .C2(n452), .ZN(n2460) );
  INVD1BWP12T U972 ( .I(r7[4]), .ZN(n1890) );
  OAI222D0BWP12T U973 ( .A1(n1890), .A2(n442), .B1(n433), .B2(n441), .C1(n432), 
        .C2(n440), .ZN(n2397) );
  AO222D0BWP12T U974 ( .A1(n1317), .A2(write1_in[5]), .B1(n820), .B2(
        write2_in[5]), .C1(n819), .C2(tmp1[5]), .Z(n2142) );
  INVD1BWP12T U975 ( .I(r0[8]), .ZN(n1757) );
  OAI222D0BWP12T U976 ( .A1(n1757), .A2(n484), .B1(n436), .B2(n482), .C1(n437), 
        .C2(n480), .ZN(n2625) );
  INVD1BWP12T U977 ( .I(r0[4]), .ZN(n1889) );
  OAI222D0BWP12T U978 ( .A1(n1889), .A2(n484), .B1(n433), .B2(n482), .C1(n432), 
        .C2(n480), .ZN(n2621) );
  INVD1BWP12T U979 ( .I(r5[1]), .ZN(n1938) );
  OAI222D0BWP12T U980 ( .A1(n1938), .A2(n454), .B1(n434), .B2(n453), .C1(n435), 
        .C2(n452), .ZN(n2458) );
  INVD1BWP12T U981 ( .I(r8[4]), .ZN(n1886) );
  OAI222D0BWP12T U982 ( .A1(n1886), .A2(n460), .B1(n433), .B2(n459), .C1(n432), 
        .C2(n458), .ZN(n2365) );
  CKND0BWP12T U983 ( .I(r4[4]), .ZN(n417) );
  OAI222D0BWP12T U984 ( .A1(n417), .A2(n472), .B1(n433), .B2(n471), .C1(n432), 
        .C2(n470), .ZN(n2493) );
  INVD1BWP12T U985 ( .I(r0[3]), .ZN(n831) );
  OAI222D0BWP12T U986 ( .A1(n831), .A2(n484), .B1(n427), .B2(n482), .C1(n426), 
        .C2(n480), .ZN(n2620) );
  INVD1BWP12T U987 ( .I(r8[3]), .ZN(n812) );
  OAI222D0BWP12T U988 ( .A1(n812), .A2(n460), .B1(n427), .B2(n459), .C1(n426), 
        .C2(n458), .ZN(n2364) );
  CKND0BWP12T U989 ( .I(r4[3]), .ZN(n821) );
  OAI222D0BWP12T U990 ( .A1(n821), .A2(n472), .B1(n427), .B2(n471), .C1(n426), 
        .C2(n470), .ZN(n2492) );
  OAI222D0BWP12T U991 ( .A1(n1758), .A2(n442), .B1(n436), .B2(n441), .C1(n437), 
        .C2(n440), .ZN(n2401) );
  AO222D0BWP12T U992 ( .A1(n1317), .A2(write1_in[7]), .B1(n820), .B2(
        write2_in[7]), .C1(n819), .C2(tmp1[7]), .Z(n2144) );
  AOI21D0BWP12T U993 ( .A1(n421), .A2(n[2033]), .B(reset), .ZN(n419) );
  CKND2D0BWP12T U994 ( .A1(write2_in[8]), .A2(n1315), .ZN(n418) );
  OAI211D0BWP12T U995 ( .A1(n451), .A2(n436), .B(n419), .C(n418), .ZN(spin[8])
         );
  INVD1BWP12T U996 ( .I(r8[1]), .ZN(n1936) );
  OAI222D0BWP12T U997 ( .A1(n1936), .A2(n460), .B1(n434), .B2(n459), .C1(n435), 
        .C2(n458), .ZN(n2362) );
  INVD1BWP12T U998 ( .I(r5[9]), .ZN(n1719) );
  OAI222D0BWP12T U999 ( .A1(n1719), .A2(n454), .B1(n424), .B2(n453), .C1(n425), 
        .C2(n452), .ZN(n2466) );
  CKND0BWP12T U1000 ( .I(r4[1]), .ZN(n420) );
  OAI222D0BWP12T U1001 ( .A1(n420), .A2(n472), .B1(n434), .B2(n471), .C1(n435), 
        .C2(n470), .ZN(n2490) );
  AOI21D0BWP12T U1002 ( .A1(n421), .A2(n[2032]), .B(reset), .ZN(n423) );
  CKND2D0BWP12T U1003 ( .A1(write2_in[9]), .A2(n1315), .ZN(n422) );
  OAI211D0BWP12T U1004 ( .A1(n451), .A2(n424), .B(n423), .C(n422), .ZN(spin[9]) );
  OAI222D0BWP12T U1005 ( .A1(n1756), .A2(n454), .B1(n436), .B2(n453), .C1(n437), .C2(n452), .ZN(n2465) );
  INVD1BWP12T U1006 ( .I(r7[9]), .ZN(n1721) );
  OAI222D0BWP12T U1007 ( .A1(n1721), .A2(n442), .B1(n424), .B2(n441), .C1(n425), .C2(n440), .ZN(n2402) );
  INVD1BWP12T U1008 ( .I(r11[3]), .ZN(n802) );
  OAI222D0BWP12T U1009 ( .A1(n426), .A2(n476), .B1(n427), .B2(n475), .C1(n474), 
        .C2(n802), .ZN(n2268) );
  INVD1BWP12T U1010 ( .I(r2[4]), .ZN(n1878) );
  OAI222D0BWP12T U1011 ( .A1(n432), .A2(n488), .B1(n433), .B2(n486), .C1(n485), 
        .C2(n1878), .ZN(n2557) );
  INVD1BWP12T U1012 ( .I(r10[3]), .ZN(n803) );
  OAI222D0BWP12T U1013 ( .A1(n426), .A2(n448), .B1(n427), .B2(n447), .C1(n446), 
        .C2(n803), .ZN(n2300) );
  INVD1BWP12T U1014 ( .I(r3[3]), .ZN(n830) );
  OAI222D0BWP12T U1015 ( .A1(n426), .A2(n457), .B1(n427), .B2(n456), .C1(n455), 
        .C2(n830), .ZN(n2524) );
  INVD1BWP12T U1016 ( .I(r11[9]), .ZN(n1703) );
  OAI222D0BWP12T U1017 ( .A1(n425), .A2(n476), .B1(n424), .B2(n475), .C1(n474), 
        .C2(n1703), .ZN(n2274) );
  INVD1BWP12T U1018 ( .I(r2[3]), .ZN(n828) );
  OAI222D0BWP12T U1019 ( .A1(n426), .A2(n488), .B1(n427), .B2(n486), .C1(n485), 
        .C2(n828), .ZN(n2556) );
  INVD1BWP12T U1020 ( .I(lr[3]), .ZN(n804) );
  OAI222D0BWP12T U1021 ( .A1(n804), .A2(n479), .B1(n427), .B2(n478), .C1(n426), 
        .C2(n477), .ZN(n2204) );
  INVD1BWP12T U1022 ( .I(r12[1]), .ZN(n1857) );
  OAI222D0BWP12T U1023 ( .A1(n1857), .A2(n445), .B1(n434), .B2(n444), .C1(n435), .C2(n443), .ZN(n2234) );
  INVD1BWP12T U1024 ( .I(r1[3]), .ZN(n824) );
  OAI222D0BWP12T U1025 ( .A1(n824), .A2(n463), .B1(n427), .B2(n462), .C1(n426), 
        .C2(n461), .ZN(n2588) );
  OAI222D0BWP12T U1026 ( .A1(n960), .A2(n445), .B1(n436), .B2(n444), .C1(n437), 
        .C2(n443), .ZN(n2241) );
  INVD1BWP12T U1027 ( .I(r9[1]), .ZN(n1934) );
  OAI222D0BWP12T U1028 ( .A1(n1934), .A2(n466), .B1(n434), .B2(n465), .C1(n435), .C2(n464), .ZN(n2330) );
  OAI222D0BWP12T U1029 ( .A1(n437), .A2(n488), .B1(n436), .B2(n486), .C1(n485), 
        .C2(n1746), .ZN(n2561) );
  INVD1BWP12T U1030 ( .I(r3[1]), .ZN(n1937) );
  OAI222D0BWP12T U1031 ( .A1(n435), .A2(n457), .B1(n434), .B2(n456), .C1(n455), 
        .C2(n1937), .ZN(n2522) );
  INVD1BWP12T U1032 ( .I(r12[9]), .ZN(n1726) );
  OAI222D0BWP12T U1033 ( .A1(n1726), .A2(n445), .B1(n424), .B2(n444), .C1(n425), .C2(n443), .ZN(n2242) );
  INVD1BWP12T U1034 ( .I(r11[4]), .ZN(n1872) );
  OAI222D0BWP12T U1035 ( .A1(n432), .A2(n476), .B1(n433), .B2(n475), .C1(n474), 
        .C2(n1872), .ZN(n2269) );
  INVD1BWP12T U1036 ( .I(r1[1]), .ZN(n1927) );
  OAI222D0BWP12T U1037 ( .A1(n1927), .A2(n463), .B1(n434), .B2(n462), .C1(n435), .C2(n461), .ZN(n2586) );
  INVD1BWP12T U1038 ( .I(lr[4]), .ZN(n1875) );
  OAI222D0BWP12T U1039 ( .A1(n1875), .A2(n479), .B1(n433), .B2(n478), .C1(n432), .C2(n477), .ZN(n2205) );
  INVD1BWP12T U1040 ( .I(lr[9]), .ZN(n1728) );
  OAI222D0BWP12T U1041 ( .A1(n1728), .A2(n479), .B1(n424), .B2(n478), .C1(n425), .C2(n477), .ZN(n2210) );
  INVD1BWP12T U1042 ( .I(r10[1]), .ZN(n1924) );
  OAI222D0BWP12T U1043 ( .A1(n435), .A2(n448), .B1(n434), .B2(n447), .C1(n446), 
        .C2(n1924), .ZN(n2298) );
  INVD1BWP12T U1044 ( .I(r3[9]), .ZN(n1729) );
  OAI222D0BWP12T U1045 ( .A1(n425), .A2(n457), .B1(n424), .B2(n456), .C1(n455), 
        .C2(n1729), .ZN(n2530) );
  OAI222D0BWP12T U1046 ( .A1(n1743), .A2(n479), .B1(n436), .B2(n478), .C1(n437), .C2(n477), .ZN(n2209) );
  INVD1BWP12T U1047 ( .I(r11[8]), .ZN(n1740) );
  OAI222D0BWP12T U1048 ( .A1(n437), .A2(n476), .B1(n436), .B2(n475), .C1(n474), 
        .C2(n1740), .ZN(n2273) );
  INVD1BWP12T U1049 ( .I(r3[4]), .ZN(n1887) );
  OAI222D0BWP12T U1050 ( .A1(n432), .A2(n457), .B1(n433), .B2(n456), .C1(n455), 
        .C2(n1887), .ZN(n2525) );
  INVD1BWP12T U1051 ( .I(r10[4]), .ZN(n1874) );
  OAI222D0BWP12T U1052 ( .A1(n432), .A2(n448), .B1(n433), .B2(n447), .C1(n446), 
        .C2(n1874), .ZN(n2301) );
  INVD1BWP12T U1053 ( .I(r1[4]), .ZN(n1877) );
  OAI222D0BWP12T U1054 ( .A1(n1877), .A2(n463), .B1(n433), .B2(n462), .C1(n432), .C2(n461), .ZN(n2589) );
  OAI222D0BWP12T U1055 ( .A1(n437), .A2(n457), .B1(n436), .B2(n456), .C1(n455), 
        .C2(n1755), .ZN(n2529) );
  INVD1BWP12T U1056 ( .I(r2[9]), .ZN(n1720) );
  OAI222D0BWP12T U1057 ( .A1(n425), .A2(n488), .B1(n424), .B2(n486), .C1(n485), 
        .C2(n1720), .ZN(n2562) );
  INVD1BWP12T U1058 ( .I(r10[9]), .ZN(n1718) );
  OAI222D0BWP12T U1059 ( .A1(n425), .A2(n448), .B1(n424), .B2(n447), .C1(n446), 
        .C2(n1718), .ZN(n2306) );
  INVD1BWP12T U1060 ( .I(r12[3]), .ZN(n606) );
  OAI222D0BWP12T U1061 ( .A1(n606), .A2(n445), .B1(n427), .B2(n444), .C1(n426), 
        .C2(n443), .ZN(n2236) );
  AOI21D0BWP12T U1062 ( .A1(n1355), .A2(next_pc_in[1]), .B(reset), .ZN(n429)
         );
  TPND2D0BWP12T U1063 ( .A1(n1361), .A2(pc_out[1]), .ZN(n428) );
  OAI211D0BWP12T U1064 ( .A1(n431), .A2(n430), .B(n429), .C(n428), .ZN(n2170)
         );
  INVD1BWP12T U1065 ( .I(r11[1]), .ZN(n1922) );
  OAI222D0BWP12T U1066 ( .A1(n435), .A2(n476), .B1(n434), .B2(n475), .C1(n474), 
        .C2(n1922), .ZN(n2266) );
  OAI222D0BWP12T U1067 ( .A1(n1745), .A2(n463), .B1(n436), .B2(n462), .C1(n437), .C2(n461), .ZN(n2593) );
  INVD1BWP12T U1068 ( .I(r12[4]), .ZN(n544) );
  OAI222D0BWP12T U1069 ( .A1(n544), .A2(n445), .B1(n433), .B2(n444), .C1(n432), 
        .C2(n443), .ZN(n2237) );
  INVD1BWP12T U1070 ( .I(r2[1]), .ZN(n1928) );
  OAI222D0BWP12T U1071 ( .A1(n435), .A2(n488), .B1(n434), .B2(n486), .C1(n485), 
        .C2(n1928), .ZN(n2554) );
  OAI222D0BWP12T U1072 ( .A1(n437), .A2(n448), .B1(n436), .B2(n447), .C1(n446), 
        .C2(n1742), .ZN(n2305) );
  INVD1BWP12T U1073 ( .I(write1_in[2]), .ZN(n487) );
  AOI21D0BWP12T U1074 ( .A1(n421), .A2(n[2039]), .B(reset), .ZN(n439) );
  CKND2D0BWP12T U1075 ( .A1(write2_in[2]), .A2(n1315), .ZN(n438) );
  OAI211D0BWP12T U1076 ( .A1(n451), .A2(n487), .B(n439), .C(n438), .ZN(spin[2]) );
  INVD1BWP12T U1077 ( .I(r12[2]), .ZN(n760) );
  INVD1BWP12T U1078 ( .I(write2_in[2]), .ZN(n489) );
  OAI222D0BWP12T U1079 ( .A1(n760), .A2(n445), .B1(n487), .B2(n444), .C1(n489), 
        .C2(n443), .ZN(n2235) );
  AO222D0BWP12T U1080 ( .A1(n1317), .A2(write1_in[8]), .B1(n820), .B2(
        write2_in[8]), .C1(n819), .C2(tmp1[8]), .Z(n2145) );
  INVD1BWP12T U1081 ( .I(write2_in[6]), .ZN(n481) );
  INVD1BWP12T U1082 ( .I(write1_in[6]), .ZN(n483) );
  INVD1BWP12T U1083 ( .I(r3[6]), .ZN(n1821) );
  OAI222D0BWP12T U1084 ( .A1(n481), .A2(n457), .B1(n483), .B2(n456), .C1(n455), 
        .C2(n1821), .ZN(n2527) );
  INVD1BWP12T U1085 ( .I(r7[2]), .ZN(n1980) );
  OAI222D0BWP12T U1086 ( .A1(n1980), .A2(n442), .B1(n487), .B2(n441), .C1(n489), .C2(n440), .ZN(n2395) );
  INVD1BWP12T U1087 ( .I(r7[6]), .ZN(n1824) );
  OAI222D0BWP12T U1088 ( .A1(n1824), .A2(n442), .B1(n483), .B2(n441), .C1(n481), .C2(n440), .ZN(n2399) );
  INVD1BWP12T U1089 ( .I(r8[6]), .ZN(n1820) );
  OAI222D0BWP12T U1090 ( .A1(n1820), .A2(n460), .B1(n483), .B2(n459), .C1(n481), .C2(n458), .ZN(n2367) );
  INVD1BWP12T U1091 ( .I(r12[6]), .ZN(n1110) );
  OAI222D0BWP12T U1092 ( .A1(n1110), .A2(n445), .B1(n483), .B2(n444), .C1(n481), .C2(n443), .ZN(n2239) );
  INVD1BWP12T U1093 ( .I(r10[2]), .ZN(n1951) );
  OAI222D0BWP12T U1094 ( .A1(n489), .A2(n448), .B1(n487), .B2(n447), .C1(n446), 
        .C2(n1951), .ZN(n2299) );
  INVD1BWP12T U1095 ( .I(r10[6]), .ZN(n1807) );
  OAI222D0BWP12T U1096 ( .A1(n481), .A2(n448), .B1(n483), .B2(n447), .C1(n446), 
        .C2(n1807), .ZN(n2303) );
  AOI21D0BWP12T U1097 ( .A1(n421), .A2(n[2035]), .B(reset), .ZN(n450) );
  CKND2D0BWP12T U1098 ( .A1(write2_in[6]), .A2(n1315), .ZN(n449) );
  OAI211D0BWP12T U1099 ( .A1(n451), .A2(n483), .B(n450), .C(n449), .ZN(spin[6]) );
  INVD1BWP12T U1100 ( .I(r5[6]), .ZN(n1822) );
  OAI222D0BWP12T U1101 ( .A1(n1822), .A2(n454), .B1(n483), .B2(n453), .C1(n481), .C2(n452), .ZN(n2463) );
  INVD1BWP12T U1102 ( .I(r5[2]), .ZN(n1977) );
  OAI222D0BWP12T U1103 ( .A1(n1977), .A2(n454), .B1(n487), .B2(n453), .C1(n489), .C2(n452), .ZN(n2459) );
  INVD1BWP12T U1104 ( .I(r9[2]), .ZN(n1968) );
  OAI222D0BWP12T U1105 ( .A1(n1968), .A2(n466), .B1(n487), .B2(n465), .C1(n489), .C2(n464), .ZN(n2331) );
  INVD1BWP12T U1106 ( .I(r0[2]), .ZN(n1978) );
  OAI222D0BWP12T U1107 ( .A1(n1978), .A2(n484), .B1(n487), .B2(n482), .C1(n489), .C2(n480), .ZN(n2619) );
  INVD1BWP12T U1108 ( .I(r3[2]), .ZN(n1974) );
  OAI222D0BWP12T U1109 ( .A1(n489), .A2(n457), .B1(n487), .B2(n456), .C1(n455), 
        .C2(n1974), .ZN(n2523) );
  CKND0BWP12T U1110 ( .I(r4[2]), .ZN(n850) );
  OAI222D0BWP12T U1111 ( .A1(n850), .A2(n472), .B1(n487), .B2(n471), .C1(n489), 
        .C2(n470), .ZN(n2491) );
  INVD1BWP12T U1112 ( .I(lr[2]), .ZN(n1954) );
  OAI222D0BWP12T U1113 ( .A1(n1954), .A2(n479), .B1(n487), .B2(n478), .C1(n489), .C2(n477), .ZN(n2203) );
  INVD1BWP12T U1114 ( .I(r1[6]), .ZN(n1811) );
  OAI222D0BWP12T U1115 ( .A1(n1811), .A2(n463), .B1(n483), .B2(n462), .C1(n481), .C2(n461), .ZN(n2591) );
  INVD1BWP12T U1116 ( .I(r8[2]), .ZN(n1972) );
  OAI222D0BWP12T U1117 ( .A1(n1972), .A2(n460), .B1(n487), .B2(n459), .C1(n489), .C2(n458), .ZN(n2363) );
  INVD1BWP12T U1118 ( .I(r6[2]), .ZN(n1966) );
  OAI222D0BWP12T U1119 ( .A1(n1966), .A2(n469), .B1(n487), .B2(n468), .C1(n489), .C2(n467), .ZN(n2427) );
  INVD1BWP12T U1120 ( .I(r1[2]), .ZN(n1958) );
  OAI222D0BWP12T U1121 ( .A1(n1958), .A2(n463), .B1(n487), .B2(n462), .C1(n489), .C2(n461), .ZN(n2587) );
  AO222D0BWP12T U1122 ( .A1(n1317), .A2(write1_in[1]), .B1(n820), .B2(
        write2_in[1]), .C1(n819), .C2(tmp1[1]), .Z(n2138) );
  INVD1BWP12T U1123 ( .I(r9[6]), .ZN(n1818) );
  OAI222D0BWP12T U1124 ( .A1(n1818), .A2(n466), .B1(n483), .B2(n465), .C1(n481), .C2(n464), .ZN(n2335) );
  INVD1BWP12T U1125 ( .I(r11[6]), .ZN(n1805) );
  OAI222D0BWP12T U1126 ( .A1(n481), .A2(n476), .B1(n483), .B2(n475), .C1(n474), 
        .C2(n1805), .ZN(n2271) );
  AO222D0BWP12T U1127 ( .A1(n1317), .A2(write1_in[3]), .B1(n820), .B2(
        write2_in[3]), .C1(n819), .C2(tmp1[3]), .Z(n2140) );
  INVD1BWP12T U1128 ( .I(r6[6]), .ZN(n1817) );
  OAI222D0BWP12T U1129 ( .A1(n1817), .A2(n469), .B1(n483), .B2(n468), .C1(n481), .C2(n467), .ZN(n2431) );
  CKND0BWP12T U1130 ( .I(r4[6]), .ZN(n473) );
  OAI222D0BWP12T U1131 ( .A1(n473), .A2(n472), .B1(n483), .B2(n471), .C1(n481), 
        .C2(n470), .ZN(n2495) );
  INVD1BWP12T U1132 ( .I(r11[2]), .ZN(n1947) );
  OAI222D0BWP12T U1133 ( .A1(n489), .A2(n476), .B1(n487), .B2(n475), .C1(n474), 
        .C2(n1947), .ZN(n2267) );
  INVD1BWP12T U1134 ( .I(lr[6]), .ZN(n1808) );
  OAI222D0BWP12T U1135 ( .A1(n1808), .A2(n479), .B1(n483), .B2(n478), .C1(n481), .C2(n477), .ZN(n2207) );
  INVD1BWP12T U1136 ( .I(r2[6]), .ZN(n1812) );
  OAI222D0BWP12T U1137 ( .A1(n481), .A2(n488), .B1(n483), .B2(n486), .C1(n485), 
        .C2(n1812), .ZN(n2559) );
  INVD1BWP12T U1138 ( .I(r0[6]), .ZN(n1823) );
  OAI222D0BWP12T U1139 ( .A1(n1823), .A2(n484), .B1(n483), .B2(n482), .C1(n481), .C2(n480), .ZN(n2623) );
  AO222D0BWP12T U1140 ( .A1(n1317), .A2(write1_in[9]), .B1(n820), .B2(
        write2_in[9]), .C1(n819), .C2(tmp1[9]), .Z(n2146) );
  INVD1BWP12T U1141 ( .I(r2[2]), .ZN(n1960) );
  OAI222D0BWP12T U1142 ( .A1(n489), .A2(n488), .B1(n487), .B2(n486), .C1(n485), 
        .C2(n1960), .ZN(n2555) );
  AO222D0BWP12T U1143 ( .A1(n1317), .A2(write1_in[6]), .B1(n820), .B2(
        write2_in[6]), .C1(n819), .C2(tmp1[6]), .Z(n2143) );
  INVD1BWP12T U1144 ( .I(pc_out[20]), .ZN(n490) );
  INVD1BWP12T U1145 ( .I(r11[20]), .ZN(n1027) );
  OAI22D1BWP12T U1146 ( .A1(n490), .A2(n1949), .B1(n1948), .B2(n1027), .ZN(
        n498) );
  INVD1BWP12T U1147 ( .I(lr[20]), .ZN(n492) );
  INVD1BWP12T U1148 ( .I(r10[20]), .ZN(n491) );
  OAI22D1BWP12T U1149 ( .A1(n492), .A2(n1953), .B1(n1952), .B2(n491), .ZN(n497) );
  INVD1BWP12T U1150 ( .I(r2[20]), .ZN(n494) );
  INVD1BWP12T U1151 ( .I(r1[20]), .ZN(n493) );
  OAI22D1BWP12T U1152 ( .A1(n1961), .A2(n494), .B1(n1959), .B2(n493), .ZN(n495) );
  NR4D0BWP12T U1153 ( .A1(n498), .A2(n497), .A3(n496), .A4(n495), .ZN(n504) );
  AOI22D1BWP12T U1154 ( .A1(r9[20]), .A2(n1591), .B1(n1590), .B2(r6[20]), .ZN(
        n502) );
  AOI22D1BWP12T U1155 ( .A1(r8[20]), .A2(n1593), .B1(n1592), .B2(n[2021]), 
        .ZN(n501) );
  AOI22D1BWP12T U1156 ( .A1(r5[20]), .A2(n1594), .B1(n171), .B2(r3[20]), .ZN(
        n500) );
  AOI22D1BWP12T U1157 ( .A1(r7[20]), .A2(n1596), .B1(n1595), .B2(r0[20]), .ZN(
        n499) );
  AN4XD1BWP12T U1158 ( .A1(n502), .A2(n501), .A3(n500), .A4(n499), .Z(n503) );
  CKND2D1BWP12T U1159 ( .A1(n504), .A2(n503), .ZN(regA_out[20]) );
  INVD0BWP12T U1160 ( .I(pc_out[14]), .ZN(n506) );
  INVD1BWP12T U1161 ( .I(r11[14]), .ZN(n505) );
  OAI22D1BWP12T U1162 ( .A1(n506), .A2(n1949), .B1(n1948), .B2(n505), .ZN(n512) );
  INVD1BWP12T U1163 ( .I(lr[14]), .ZN(n1087) );
  INVD1BWP12T U1164 ( .I(r10[14]), .ZN(n1085) );
  OAI22D1BWP12T U1165 ( .A1(n1087), .A2(n1953), .B1(n1952), .B2(n1085), .ZN(
        n511) );
  AOI22D1BWP12T U1166 ( .A1(n150), .A2(r12[14]), .B1(n1809), .B2(tmp1[14]), 
        .ZN(n507) );
  IOA21D1BWP12T U1167 ( .A1(n1957), .A2(r4[14]), .B(n507), .ZN(n510) );
  INVD1BWP12T U1168 ( .I(r2[14]), .ZN(n624) );
  INVD1BWP12T U1169 ( .I(r1[14]), .ZN(n508) );
  OAI22D1BWP12T U1170 ( .A1(n1961), .A2(n624), .B1(n1959), .B2(n508), .ZN(n509) );
  NR4D0BWP12T U1171 ( .A1(n512), .A2(n511), .A3(n510), .A4(n509), .ZN(n518) );
  AOI22D1BWP12T U1172 ( .A1(r9[14]), .A2(n1591), .B1(n1590), .B2(r6[14]), .ZN(
        n516) );
  AOI22D1BWP12T U1173 ( .A1(r8[14]), .A2(n1593), .B1(n1592), .B2(n[2027]), 
        .ZN(n515) );
  AOI22D1BWP12T U1174 ( .A1(r5[14]), .A2(n1594), .B1(n171), .B2(r3[14]), .ZN(
        n514) );
  AOI22D1BWP12T U1175 ( .A1(r7[14]), .A2(n1596), .B1(n1595), .B2(r0[14]), .ZN(
        n513) );
  AN4XD1BWP12T U1176 ( .A1(n516), .A2(n515), .A3(n514), .A4(n513), .Z(n517) );
  CKND2D1BWP12T U1177 ( .A1(n518), .A2(n517), .ZN(regA_out[14]) );
  INVD1BWP12T U1178 ( .I(pc_out[0]), .ZN(n520) );
  INVD1BWP12T U1179 ( .I(r11[0]), .ZN(n519) );
  OAI22D1BWP12T U1180 ( .A1(n520), .A2(n1949), .B1(n1948), .B2(n519), .ZN(n528) );
  INVD1BWP12T U1181 ( .I(lr[0]), .ZN(n995) );
  INVD1BWP12T U1182 ( .I(r10[0]), .ZN(n994) );
  OAI22D1BWP12T U1183 ( .A1(n995), .A2(n1953), .B1(n1952), .B2(n994), .ZN(n527) );
  BUFFXD3BWP12T U1184 ( .I(n521), .Z(n1955) );
  AOI22D1BWP12T U1185 ( .A1(n150), .A2(r12[0]), .B1(n1955), .B2(tmp1[0]), .ZN(
        n522) );
  IOA21D1BWP12T U1186 ( .A1(n1957), .A2(r4[0]), .B(n522), .ZN(n526) );
  INVD1BWP12T U1187 ( .I(r2[0]), .ZN(n524) );
  INVD1BWP12T U1188 ( .I(r1[0]), .ZN(n523) );
  OAI22D1BWP12T U1189 ( .A1(n1961), .A2(n524), .B1(n1959), .B2(n523), .ZN(n525) );
  NR4D0BWP12T U1190 ( .A1(n528), .A2(n527), .A3(n526), .A4(n525), .ZN(n534) );
  AOI22D1BWP12T U1191 ( .A1(r9[0]), .A2(n1591), .B1(n1590), .B2(r6[0]), .ZN(
        n532) );
  AOI22D1BWP12T U1192 ( .A1(r8[0]), .A2(n1593), .B1(n1592), .B2(n[2041]), .ZN(
        n531) );
  AOI22D1BWP12T U1193 ( .A1(r5[0]), .A2(n1594), .B1(n171), .B2(r3[0]), .ZN(
        n530) );
  AOI22D1BWP12T U1194 ( .A1(r7[0]), .A2(n1596), .B1(n1595), .B2(r0[0]), .ZN(
        n529) );
  AN4XD1BWP12T U1195 ( .A1(n532), .A2(n531), .A3(n530), .A4(n529), .Z(n533) );
  CKND2D1BWP12T U1196 ( .A1(n534), .A2(n533), .ZN(regA_out[0]) );
  OAI22D1BWP12T U1197 ( .A1(n1888), .A2(n1846), .B1(n1845), .B2(n1874), .ZN(
        n543) );
  INVD1BWP12T U1198 ( .I(tmp1[4]), .ZN(n535) );
  MOAI22D0BWP12T U1199 ( .A1(n535), .A2(n1847), .B1(n200), .B2(
        immediate2_in[4]), .ZN(n542) );
  AOI22D1BWP12T U1200 ( .A1(r9[4]), .A2(n201), .B1(n1780), .B2(r4[4]), .ZN(
        n539) );
  AOI22D1BWP12T U1201 ( .A1(r11[4]), .A2(n537), .B1(n205), .B2(r0[4]), .ZN(
        n538) );
  ND2D1BWP12T U1202 ( .A1(n539), .A2(n538), .ZN(n541) );
  NR4D0BWP12T U1203 ( .A1(n543), .A2(n542), .A3(n541), .A4(n540), .ZN(n550) );
  OAI22D1BWP12T U1204 ( .A1(n1877), .A2(n1859), .B1(n1858), .B2(n544), .ZN(
        n548) );
  OAI22D1BWP12T U1205 ( .A1(n1887), .A2(n1861), .B1(n1860), .B2(n1875), .ZN(
        n547) );
  INVD1BWP12T U1206 ( .I(n[2037]), .ZN(n1885) );
  OAI22D1BWP12T U1207 ( .A1(n1863), .A2(n1886), .B1(n1862), .B2(n1885), .ZN(
        n546) );
  INVD1BWP12T U1208 ( .I(pc_out[4]), .ZN(n1873) );
  OAI22D1BWP12T U1209 ( .A1(n1865), .A2(n1873), .B1(n1864), .B2(n1883), .ZN(
        n545) );
  NR4D0BWP12T U1210 ( .A1(n548), .A2(n547), .A3(n546), .A4(n545), .ZN(n549) );
  CKND2D1BWP12T U1211 ( .A1(n550), .A2(n549), .ZN(regB_out[4]) );
  INVD0BWP12T U1212 ( .I(tmp1[11]), .ZN(n551) );
  MOAI22D0BWP12T U1213 ( .A1(n551), .A2(n1847), .B1(n200), .B2(
        immediate2_in[11]), .ZN(n557) );
  AOI22D1BWP12T U1214 ( .A1(r9[11]), .A2(n201), .B1(n1780), .B2(r4[11]), .ZN(
        n553) );
  AOI22D1BWP12T U1215 ( .A1(r11[11]), .A2(n2002), .B1(n205), .B2(r0[11]), .ZN(
        n552) );
  ND2D1BWP12T U1216 ( .A1(n553), .A2(n552), .ZN(n556) );
  OAI22D1BWP12T U1217 ( .A1(n1670), .A2(n1846), .B1(n1845), .B2(n1656), .ZN(
        n555) );
  OAI22D1BWP12T U1218 ( .A1(n1852), .A2(n1672), .B1(n1851), .B2(n1660), .ZN(
        n554) );
  NR4D0BWP12T U1219 ( .A1(n557), .A2(n556), .A3(n555), .A4(n554), .ZN(n563) );
  OAI22D1BWP12T U1220 ( .A1(n1659), .A2(n1859), .B1(n1858), .B2(n1121), .ZN(
        n561) );
  OAI22D1BWP12T U1221 ( .A1(n1669), .A2(n1861), .B1(n1860), .B2(n1657), .ZN(
        n560) );
  INVD1BWP12T U1222 ( .I(n[2030]), .ZN(n1667) );
  OAI22D1BWP12T U1223 ( .A1(n1863), .A2(n1668), .B1(n1862), .B2(n1667), .ZN(
        n559) );
  INVD1BWP12T U1224 ( .I(pc_out[11]), .ZN(n1655) );
  OAI22D1BWP12T U1225 ( .A1(n1865), .A2(n1655), .B1(n1864), .B2(n1665), .ZN(
        n558) );
  NR4D0BWP12T U1226 ( .A1(n561), .A2(n560), .A3(n559), .A4(n558), .ZN(n562) );
  CKND2D1BWP12T U1227 ( .A1(n563), .A2(n562), .ZN(regB_out[11]) );
  INVD1BWP12T U1228 ( .I(tmp1[6]), .ZN(n564) );
  MOAI22D0BWP12T U1229 ( .A1(n564), .A2(n1847), .B1(n200), .B2(
        immediate2_in[6]), .ZN(n570) );
  AOI22D1BWP12T U1230 ( .A1(r9[6]), .A2(n201), .B1(n1780), .B2(r4[6]), .ZN(
        n566) );
  AOI22D1BWP12T U1231 ( .A1(r11[6]), .A2(n537), .B1(n205), .B2(r0[6]), .ZN(
        n565) );
  ND2D1BWP12T U1232 ( .A1(n566), .A2(n565), .ZN(n569) );
  OAI22D1BWP12T U1233 ( .A1(n1822), .A2(n1846), .B1(n1845), .B2(n1807), .ZN(
        n568) );
  OAI22D1BWP12T U1234 ( .A1(n1852), .A2(n1824), .B1(n1851), .B2(n1812), .ZN(
        n567) );
  NR4D0BWP12T U1235 ( .A1(n570), .A2(n569), .A3(n568), .A4(n567), .ZN(n576) );
  OAI22D1BWP12T U1236 ( .A1(n1811), .A2(n1859), .B1(n1858), .B2(n1110), .ZN(
        n574) );
  OAI22D1BWP12T U1237 ( .A1(n1821), .A2(n1861), .B1(n1860), .B2(n1808), .ZN(
        n573) );
  INVD1BWP12T U1238 ( .I(n[2035]), .ZN(n1819) );
  OAI22D1BWP12T U1239 ( .A1(n1863), .A2(n1820), .B1(n1862), .B2(n1819), .ZN(
        n572) );
  INVD1BWP12T U1240 ( .I(pc_out[6]), .ZN(n1806) );
  OAI22D1BWP12T U1241 ( .A1(n1865), .A2(n1806), .B1(n1864), .B2(n1817), .ZN(
        n571) );
  NR4D0BWP12T U1242 ( .A1(n574), .A2(n573), .A3(n572), .A4(n571), .ZN(n575) );
  CKND2D1BWP12T U1243 ( .A1(n576), .A2(n575), .ZN(regB_out[6]) );
  INVD1BWP12T U1244 ( .I(r4[28]), .ZN(n579) );
  AOI22D1BWP12T U1245 ( .A1(n150), .A2(r12[28]), .B1(n1486), .B2(tmp1[28]), 
        .ZN(n578) );
  AOI22D1BWP12T U1246 ( .A1(r2[28]), .A2(n155), .B1(n1555), .B2(r1[28]), .ZN(
        n577) );
  OA211D1BWP12T U1247 ( .A1(n579), .A2(n1458), .B(n578), .C(n577), .Z(n587) );
  AOI22D1BWP12T U1248 ( .A1(r9[28]), .A2(n1591), .B1(n1590), .B2(r6[28]), .ZN(
        n583) );
  AOI22D1BWP12T U1249 ( .A1(r8[28]), .A2(n1593), .B1(n1592), .B2(n[2013]), 
        .ZN(n582) );
  AOI22D1BWP12T U1250 ( .A1(r5[28]), .A2(n1594), .B1(n171), .B2(r3[28]), .ZN(
        n581) );
  AOI22D1BWP12T U1251 ( .A1(r7[28]), .A2(n1596), .B1(n1595), .B2(r0[28]), .ZN(
        n580) );
  AN4XD1BWP12T U1252 ( .A1(n583), .A2(n582), .A3(n581), .A4(n580), .Z(n586) );
  AOI22D1BWP12T U1253 ( .A1(pc_out[28]), .A2(n141), .B1(n1559), .B2(r11[28]), 
        .ZN(n585) );
  AOI22D1BWP12T U1254 ( .A1(lr[28]), .A2(n1561), .B1(n1560), .B2(r10[28]), 
        .ZN(n584) );
  AOI22D1BWP12T U1255 ( .A1(r1[25]), .A2(n183), .B1(n1992), .B2(r12[25]), .ZN(
        n591) );
  AOI22D1BWP12T U1256 ( .A1(r3[25]), .A2(n185), .B1(n1993), .B2(lr[25]), .ZN(
        n590) );
  AOI22D1BWP12T U1257 ( .A1(r8[25]), .A2(n187), .B1(n1994), .B2(n[2016]), .ZN(
        n589) );
  AOI22D1BWP12T U1258 ( .A1(pc_out[25]), .A2(n188), .B1(n1995), .B2(r6[25]), 
        .ZN(n588) );
  AN4XD1BWP12T U1259 ( .A1(n591), .A2(n590), .A3(n589), .A4(n588), .Z(n598) );
  AOI22D1BWP12T U1260 ( .A1(tmp1[25]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[25]), .ZN(n594) );
  AOI22D0BWP12T U1261 ( .A1(r9[25]), .A2(n201), .B1(n2001), .B2(r4[25]), .ZN(
        n593) );
  AOI22D1BWP12T U1262 ( .A1(r11[25]), .A2(n1470), .B1(n205), .B2(r0[25]), .ZN(
        n592) );
  AN3XD1BWP12T U1263 ( .A1(n594), .A2(n593), .A3(n592), .Z(n597) );
  AOI22D1BWP12T U1264 ( .A1(r5[25]), .A2(n210), .B1(n1988), .B2(r10[25]), .ZN(
        n596) );
  AOI22D1BWP12T U1265 ( .A1(r7[25]), .A2(n215), .B1(n1989), .B2(r2[25]), .ZN(
        n595) );
  OAI22D1BWP12T U1266 ( .A1(n825), .A2(n1846), .B1(n1845), .B2(n803), .ZN(n605) );
  INVD1BWP12T U1267 ( .I(tmp1[3]), .ZN(n599) );
  MOAI22D0BWP12T U1268 ( .A1(n599), .A2(n1847), .B1(n200), .B2(
        immediate2_in[3]), .ZN(n604) );
  AOI22D1BWP12T U1269 ( .A1(r9[3]), .A2(n201), .B1(n1780), .B2(r4[3]), .ZN(
        n601) );
  AOI22D1BWP12T U1270 ( .A1(r11[3]), .A2(n537), .B1(n205), .B2(r0[3]), .ZN(
        n600) );
  ND2D1BWP12T U1271 ( .A1(n601), .A2(n600), .ZN(n603) );
  NR4D0BWP12T U1272 ( .A1(n605), .A2(n604), .A3(n603), .A4(n602), .ZN(n612) );
  OAI22D1BWP12T U1273 ( .A1(n824), .A2(n1859), .B1(n1858), .B2(n606), .ZN(n610) );
  OAI22D1BWP12T U1274 ( .A1(n830), .A2(n1861), .B1(n1860), .B2(n804), .ZN(n609) );
  INVD1BWP12T U1275 ( .I(n[2038]), .ZN(n811) );
  OAI22D1BWP12T U1276 ( .A1(n1863), .A2(n812), .B1(n1862), .B2(n811), .ZN(n608) );
  INVD1BWP12T U1277 ( .I(pc_out[3]), .ZN(n836) );
  NR4D0BWP12T U1278 ( .A1(n610), .A2(n609), .A3(n608), .A4(n607), .ZN(n611) );
  ND2D1BWP12T U1279 ( .A1(n612), .A2(n611), .ZN(regB_out[3]) );
  INVD1BWP12T U1280 ( .I(r4[30]), .ZN(n615) );
  AOI22D1BWP12T U1281 ( .A1(n150), .A2(r12[30]), .B1(n1486), .B2(tmp1[30]), 
        .ZN(n614) );
  AOI22D1BWP12T U1282 ( .A1(r2[30]), .A2(n155), .B1(n1555), .B2(r1[30]), .ZN(
        n613) );
  AOI22D1BWP12T U1283 ( .A1(r8[30]), .A2(n1593), .B1(n1592), .B2(n[2011]), 
        .ZN(n619) );
  AOI22D1BWP12T U1284 ( .A1(r9[30]), .A2(n1591), .B1(n1590), .B2(r6[30]), .ZN(
        n618) );
  AOI22D1BWP12T U1285 ( .A1(r5[30]), .A2(n1594), .B1(n171), .B2(r3[30]), .ZN(
        n617) );
  AOI22D1BWP12T U1286 ( .A1(r7[30]), .A2(n1596), .B1(n1595), .B2(r0[30]), .ZN(
        n616) );
  INVD1BWP12T U1287 ( .I(tmp1[14]), .ZN(n620) );
  MOAI22D0BWP12T U1288 ( .A1(n620), .A2(n1847), .B1(n200), .B2(
        immediate2_in[14]), .ZN(n628) );
  AOI22D1BWP12T U1289 ( .A1(r9[14]), .A2(n201), .B1(n1780), .B2(r4[14]), .ZN(
        n622) );
  AOI22D1BWP12T U1290 ( .A1(r11[14]), .A2(n2002), .B1(n205), .B2(r0[14]), .ZN(
        n621) );
  ND2D1BWP12T U1291 ( .A1(n622), .A2(n621), .ZN(n627) );
  INVD1BWP12T U1292 ( .I(r5[14]), .ZN(n623) );
  OAI22D1BWP12T U1293 ( .A1(n623), .A2(n1846), .B1(n1845), .B2(n1085), .ZN(
        n626) );
  NR4D0BWP12T U1294 ( .A1(n628), .A2(n627), .A3(n626), .A4(n625), .ZN(n634) );
  AOI22D1BWP12T U1295 ( .A1(r1[14]), .A2(n183), .B1(n1992), .B2(r12[14]), .ZN(
        n632) );
  AOI22D1BWP12T U1296 ( .A1(r3[14]), .A2(n185), .B1(n1993), .B2(lr[14]), .ZN(
        n631) );
  AOI22D1BWP12T U1297 ( .A1(r8[14]), .A2(n187), .B1(n1994), .B2(n[2027]), .ZN(
        n630) );
  AOI22D1BWP12T U1298 ( .A1(pc_out[14]), .A2(n188), .B1(n1995), .B2(r6[14]), 
        .ZN(n629) );
  AN4XD1BWP12T U1299 ( .A1(n632), .A2(n631), .A3(n630), .A4(n629), .Z(n633) );
  CKND2D1BWP12T U1300 ( .A1(n634), .A2(n633), .ZN(regB_out[14]) );
  INVD1BWP12T U1301 ( .I(r4[22]), .ZN(n637) );
  AOI22D1BWP12T U1302 ( .A1(n150), .A2(r12[22]), .B1(n1486), .B2(tmp1[22]), 
        .ZN(n636) );
  AOI22D1BWP12T U1303 ( .A1(r2[22]), .A2(n155), .B1(n1555), .B2(r1[22]), .ZN(
        n635) );
  OA211D1BWP12T U1304 ( .A1(n637), .A2(n1458), .B(n636), .C(n635), .Z(n645) );
  AOI22D1BWP12T U1305 ( .A1(r9[22]), .A2(n1591), .B1(n1590), .B2(r6[22]), .ZN(
        n641) );
  AOI22D1BWP12T U1306 ( .A1(r8[22]), .A2(n1593), .B1(n1592), .B2(n[2019]), 
        .ZN(n640) );
  AOI22D1BWP12T U1307 ( .A1(r5[22]), .A2(n1594), .B1(n171), .B2(r3[22]), .ZN(
        n639) );
  AOI22D1BWP12T U1308 ( .A1(r7[22]), .A2(n1596), .B1(n1595), .B2(r0[22]), .ZN(
        n638) );
  AN4XD1BWP12T U1309 ( .A1(n641), .A2(n640), .A3(n639), .A4(n638), .Z(n644) );
  AOI22D1BWP12T U1310 ( .A1(pc_out[22]), .A2(n141), .B1(n1559), .B2(r11[22]), 
        .ZN(n643) );
  AOI22D1BWP12T U1311 ( .A1(lr[22]), .A2(n1561), .B1(n1560), .B2(r10[22]), 
        .ZN(n642) );
  AOI22D1BWP12T U1312 ( .A1(r5[0]), .A2(n210), .B1(n1988), .B2(r10[0]), .ZN(
        n647) );
  AOI22D1BWP12T U1313 ( .A1(r7[0]), .A2(n215), .B1(n1989), .B2(r2[0]), .ZN(
        n646) );
  ND2D1BWP12T U1314 ( .A1(n647), .A2(n646), .ZN(n651) );
  AOI22D1BWP12T U1315 ( .A1(r9[0]), .A2(n201), .B1(n1780), .B2(r4[0]), .ZN(
        n649) );
  AOI22D1BWP12T U1316 ( .A1(r11[0]), .A2(n537), .B1(n205), .B2(r0[0]), .ZN(
        n648) );
  ND2D1BWP12T U1317 ( .A1(n649), .A2(n648), .ZN(n650) );
  AOI22D1BWP12T U1318 ( .A1(r1[0]), .A2(n183), .B1(n1992), .B2(r12[0]), .ZN(
        n656) );
  AOI22D1BWP12T U1319 ( .A1(r3[0]), .A2(n185), .B1(n1993), .B2(lr[0]), .ZN(
        n655) );
  AOI22D1BWP12T U1320 ( .A1(r8[0]), .A2(n187), .B1(n1994), .B2(n[2041]), .ZN(
        n654) );
  AOI22D1BWP12T U1321 ( .A1(pc_out[0]), .A2(n188), .B1(n1995), .B2(r6[0]), 
        .ZN(n653) );
  AN4XD1BWP12T U1322 ( .A1(n656), .A2(n655), .A3(n654), .A4(n653), .Z(n657) );
  TPND2D1BWP12T U1323 ( .A1(n658), .A2(n657), .ZN(regB_out[0]) );
  AOI22D0BWP12T U1324 ( .A1(r8[7]), .A2(n726), .B1(n725), .B2(r4[7]), .ZN(n660) );
  AOI22D0BWP12T U1325 ( .A1(n[2034]), .A2(n728), .B1(n727), .B2(r10[7]), .ZN(
        n659) );
  CKND2D1BWP12T U1326 ( .A1(n660), .A2(n659), .ZN(n669) );
  AOI22D0BWP12T U1327 ( .A1(r7[7]), .A2(n732), .B1(n731), .B2(r5[7]), .ZN(n664) );
  AOI22D0BWP12T U1328 ( .A1(lr[7]), .A2(n734), .B1(n733), .B2(r9[7]), .ZN(n663) );
  AOI22D0BWP12T U1329 ( .A1(r6[7]), .A2(n736), .B1(n735), .B2(r11[7]), .ZN(
        n662) );
  CKND2D0BWP12T U1330 ( .A1(n737), .A2(r12[7]), .ZN(n661) );
  ND4D1BWP12T U1331 ( .A1(n664), .A2(n663), .A3(n662), .A4(n661), .ZN(n668) );
  AOI22D0BWP12T U1332 ( .A1(r3[7]), .A2(n743), .B1(n742), .B2(r2[7]), .ZN(n666) );
  AOI22D0BWP12T U1333 ( .A1(n745), .A2(r0[7]), .B1(pc_out[7]), .B2(n744), .ZN(
        n665) );
  OAI211D0BWP12T U1334 ( .A1(n1792), .A2(n748), .B(n666), .C(n665), .ZN(n667)
         );
  OA31D0BWP12T U1335 ( .A1(n669), .A2(n668), .A3(n667), .B(n749), .Z(
        regD_out[7]) );
  AOI22D0BWP12T U1336 ( .A1(r8[5]), .A2(n726), .B1(n725), .B2(r4[5]), .ZN(n671) );
  AOI22D0BWP12T U1337 ( .A1(n[2036]), .A2(n728), .B1(n727), .B2(r10[5]), .ZN(
        n670) );
  CKND2D1BWP12T U1338 ( .A1(n671), .A2(n670), .ZN(n680) );
  AOI22D0BWP12T U1339 ( .A1(r7[5]), .A2(n732), .B1(n731), .B2(r5[5]), .ZN(n675) );
  AOI22D0BWP12T U1340 ( .A1(lr[5]), .A2(n734), .B1(n733), .B2(r9[5]), .ZN(n674) );
  AOI22D0BWP12T U1341 ( .A1(r6[5]), .A2(n736), .B1(n735), .B2(r11[5]), .ZN(
        n673) );
  CKND2D0BWP12T U1342 ( .A1(n737), .A2(r12[5]), .ZN(n672) );
  ND4D1BWP12T U1343 ( .A1(n675), .A2(n674), .A3(n673), .A4(n672), .ZN(n679) );
  AOI22D0BWP12T U1344 ( .A1(r3[5]), .A2(n743), .B1(n742), .B2(r2[5]), .ZN(n677) );
  AOI22D0BWP12T U1345 ( .A1(n745), .A2(r0[5]), .B1(pc_out[5]), .B2(n744), .ZN(
        n676) );
  OAI211D0BWP12T U1346 ( .A1(n1902), .A2(n748), .B(n677), .C(n676), .ZN(n678)
         );
  OA31D0BWP12T U1347 ( .A1(n680), .A2(n679), .A3(n678), .B(n749), .Z(
        regD_out[5]) );
  AOI22D0BWP12T U1348 ( .A1(r8[2]), .A2(n726), .B1(n725), .B2(r4[2]), .ZN(n682) );
  AOI22D0BWP12T U1349 ( .A1(n[2039]), .A2(n728), .B1(n727), .B2(r10[2]), .ZN(
        n681) );
  CKND2D1BWP12T U1350 ( .A1(n682), .A2(n681), .ZN(n691) );
  AOI22D0BWP12T U1351 ( .A1(r7[2]), .A2(n732), .B1(n731), .B2(r5[2]), .ZN(n686) );
  AOI22D0BWP12T U1352 ( .A1(lr[2]), .A2(n734), .B1(n733), .B2(r9[2]), .ZN(n685) );
  AOI22D0BWP12T U1353 ( .A1(r6[2]), .A2(n736), .B1(n735), .B2(r11[2]), .ZN(
        n684) );
  CKND2D0BWP12T U1354 ( .A1(n737), .A2(r12[2]), .ZN(n683) );
  ND4D1BWP12T U1355 ( .A1(n686), .A2(n685), .A3(n684), .A4(n683), .ZN(n690) );
  AOI22D0BWP12T U1356 ( .A1(r3[2]), .A2(n743), .B1(n742), .B2(r2[2]), .ZN(n688) );
  AOI22D0BWP12T U1357 ( .A1(n745), .A2(r0[2]), .B1(pc_out[2]), .B2(n744), .ZN(
        n687) );
  OAI211D0BWP12T U1358 ( .A1(n1958), .A2(n748), .B(n688), .C(n687), .ZN(n689)
         );
  OA31D0BWP12T U1359 ( .A1(n691), .A2(n690), .A3(n689), .B(n749), .Z(
        regD_out[2]) );
  AOI22D0BWP12T U1360 ( .A1(r8[6]), .A2(n726), .B1(n725), .B2(r4[6]), .ZN(n693) );
  AOI22D0BWP12T U1361 ( .A1(n[2035]), .A2(n728), .B1(n727), .B2(r10[6]), .ZN(
        n692) );
  CKND2D1BWP12T U1362 ( .A1(n693), .A2(n692), .ZN(n702) );
  AOI22D0BWP12T U1363 ( .A1(r7[6]), .A2(n732), .B1(n731), .B2(r5[6]), .ZN(n697) );
  AOI22D0BWP12T U1364 ( .A1(lr[6]), .A2(n734), .B1(n733), .B2(r9[6]), .ZN(n696) );
  AOI22D0BWP12T U1365 ( .A1(r6[6]), .A2(n736), .B1(n735), .B2(r11[6]), .ZN(
        n695) );
  CKND2D0BWP12T U1366 ( .A1(n737), .A2(r12[6]), .ZN(n694) );
  ND4D1BWP12T U1367 ( .A1(n697), .A2(n696), .A3(n695), .A4(n694), .ZN(n701) );
  AOI22D0BWP12T U1368 ( .A1(r3[6]), .A2(n743), .B1(n742), .B2(r2[6]), .ZN(n699) );
  AOI22D0BWP12T U1369 ( .A1(n745), .A2(r0[6]), .B1(pc_out[6]), .B2(n744), .ZN(
        n698) );
  OAI211D0BWP12T U1370 ( .A1(n1811), .A2(n748), .B(n699), .C(n698), .ZN(n700)
         );
  OA31D0BWP12T U1371 ( .A1(n702), .A2(n701), .A3(n700), .B(n749), .Z(
        regD_out[6]) );
  AOI22D0BWP12T U1372 ( .A1(r8[4]), .A2(n726), .B1(n725), .B2(r4[4]), .ZN(n704) );
  AOI22D0BWP12T U1373 ( .A1(n[2037]), .A2(n728), .B1(n727), .B2(r10[4]), .ZN(
        n703) );
  CKND2D1BWP12T U1374 ( .A1(n704), .A2(n703), .ZN(n713) );
  AOI22D0BWP12T U1375 ( .A1(r7[4]), .A2(n732), .B1(n731), .B2(r5[4]), .ZN(n708) );
  AOI22D0BWP12T U1376 ( .A1(lr[4]), .A2(n734), .B1(n733), .B2(r9[4]), .ZN(n707) );
  AOI22D0BWP12T U1377 ( .A1(r6[4]), .A2(n736), .B1(n735), .B2(r11[4]), .ZN(
        n706) );
  CKND2D0BWP12T U1378 ( .A1(n737), .A2(r12[4]), .ZN(n705) );
  ND4D1BWP12T U1379 ( .A1(n708), .A2(n707), .A3(n706), .A4(n705), .ZN(n712) );
  AOI22D0BWP12T U1380 ( .A1(r3[4]), .A2(n743), .B1(n742), .B2(r2[4]), .ZN(n710) );
  AOI22D0BWP12T U1381 ( .A1(n745), .A2(r0[4]), .B1(pc_out[4]), .B2(n744), .ZN(
        n709) );
  OAI211D0BWP12T U1382 ( .A1(n1877), .A2(n748), .B(n710), .C(n709), .ZN(n711)
         );
  OA31D0BWP12T U1383 ( .A1(n713), .A2(n712), .A3(n711), .B(n749), .Z(
        regD_out[4]) );
  AOI22D0BWP12T U1384 ( .A1(r8[3]), .A2(n726), .B1(n725), .B2(r4[3]), .ZN(n715) );
  AOI22D0BWP12T U1385 ( .A1(n[2038]), .A2(n728), .B1(n727), .B2(r10[3]), .ZN(
        n714) );
  CKND2D1BWP12T U1386 ( .A1(n715), .A2(n714), .ZN(n724) );
  AOI22D0BWP12T U1387 ( .A1(r7[3]), .A2(n732), .B1(n731), .B2(r5[3]), .ZN(n719) );
  AOI22D0BWP12T U1388 ( .A1(lr[3]), .A2(n734), .B1(n733), .B2(r9[3]), .ZN(n718) );
  AOI22D0BWP12T U1389 ( .A1(r6[3]), .A2(n736), .B1(n735), .B2(r11[3]), .ZN(
        n717) );
  CKND2D0BWP12T U1390 ( .A1(n737), .A2(r12[3]), .ZN(n716) );
  ND4D1BWP12T U1391 ( .A1(n719), .A2(n718), .A3(n717), .A4(n716), .ZN(n723) );
  AOI22D0BWP12T U1392 ( .A1(r3[3]), .A2(n743), .B1(n742), .B2(r2[3]), .ZN(n721) );
  AOI22D0BWP12T U1393 ( .A1(n745), .A2(r0[3]), .B1(pc_out[3]), .B2(n744), .ZN(
        n720) );
  OAI211D0BWP12T U1394 ( .A1(n824), .A2(n748), .B(n721), .C(n720), .ZN(n722)
         );
  OA31D0BWP12T U1395 ( .A1(n724), .A2(n723), .A3(n722), .B(n749), .Z(
        regD_out[3]) );
  AOI22D0BWP12T U1396 ( .A1(r8[8]), .A2(n726), .B1(n725), .B2(r4[8]), .ZN(n730) );
  AOI22D0BWP12T U1397 ( .A1(n[2033]), .A2(n728), .B1(n727), .B2(r10[8]), .ZN(
        n729) );
  CKND2D1BWP12T U1398 ( .A1(n730), .A2(n729), .ZN(n752) );
  AOI22D0BWP12T U1399 ( .A1(r7[8]), .A2(n732), .B1(n731), .B2(r5[8]), .ZN(n741) );
  AOI22D0BWP12T U1400 ( .A1(lr[8]), .A2(n734), .B1(n733), .B2(r9[8]), .ZN(n740) );
  AOI22D0BWP12T U1401 ( .A1(r6[8]), .A2(n736), .B1(n735), .B2(r11[8]), .ZN(
        n739) );
  CKND2D0BWP12T U1402 ( .A1(n737), .A2(r12[8]), .ZN(n738) );
  ND4D1BWP12T U1403 ( .A1(n741), .A2(n740), .A3(n739), .A4(n738), .ZN(n751) );
  AOI22D0BWP12T U1404 ( .A1(r3[8]), .A2(n743), .B1(n742), .B2(r2[8]), .ZN(n747) );
  AOI22D0BWP12T U1405 ( .A1(n745), .A2(r0[8]), .B1(pc_out[8]), .B2(n744), .ZN(
        n746) );
  OAI211D0BWP12T U1406 ( .A1(n1745), .A2(n748), .B(n747), .C(n746), .ZN(n750)
         );
  OA31D0BWP12T U1407 ( .A1(n752), .A2(n751), .A3(n750), .B(n749), .Z(
        regD_out[8]) );
  OAI22D1BWP12T U1408 ( .A1(n1977), .A2(n1846), .B1(n1845), .B2(n1951), .ZN(
        n759) );
  INVD1BWP12T U1409 ( .I(tmp1[2]), .ZN(n753) );
  MOAI22D0BWP12T U1410 ( .A1(n753), .A2(n1847), .B1(n200), .B2(
        immediate2_in[2]), .ZN(n758) );
  AOI22D1BWP12T U1411 ( .A1(r9[2]), .A2(n201), .B1(n536), .B2(r4[2]), .ZN(n755) );
  AOI22D1BWP12T U1412 ( .A1(r11[2]), .A2(n537), .B1(n205), .B2(r0[2]), .ZN(
        n754) );
  ND2D1BWP12T U1413 ( .A1(n755), .A2(n754), .ZN(n757) );
  TPOAI22D1BWP12T U1414 ( .A1(n1852), .A2(n1980), .B1(n1851), .B2(n1960), .ZN(
        n756) );
  NR4D0BWP12T U1415 ( .A1(n759), .A2(n758), .A3(n757), .A4(n756), .ZN(n766) );
  OAI22D1BWP12T U1416 ( .A1(n1958), .A2(n1859), .B1(n1858), .B2(n760), .ZN(
        n764) );
  OAI22D1BWP12T U1417 ( .A1(n1974), .A2(n1861), .B1(n1860), .B2(n1954), .ZN(
        n763) );
  INVD1BWP12T U1418 ( .I(n[2039]), .ZN(n1970) );
  OAI22D1BWP12T U1419 ( .A1(n1863), .A2(n1972), .B1(n1862), .B2(n1970), .ZN(
        n762) );
  INVD1BWP12T U1420 ( .I(pc_out[2]), .ZN(n1950) );
  TPOAI22D1BWP12T U1421 ( .A1(n1865), .A2(n1950), .B1(n1864), .B2(n1966), .ZN(
        n761) );
  NR4D0BWP12T U1422 ( .A1(n764), .A2(n763), .A3(n762), .A4(n761), .ZN(n765) );
  ND2D1BWP12T U1423 ( .A1(n766), .A2(n765), .ZN(regB_out[2]) );
  AOI22D1BWP12T U1424 ( .A1(r1[27]), .A2(n183), .B1(n1992), .B2(r12[27]), .ZN(
        n770) );
  AOI22D1BWP12T U1425 ( .A1(r3[27]), .A2(n185), .B1(n1993), .B2(lr[27]), .ZN(
        n769) );
  AOI22D1BWP12T U1426 ( .A1(r8[27]), .A2(n187), .B1(n1994), .B2(n[2014]), .ZN(
        n768) );
  AOI22D1BWP12T U1427 ( .A1(pc_out[27]), .A2(n188), .B1(n1995), .B2(r6[27]), 
        .ZN(n767) );
  AN4XD1BWP12T U1428 ( .A1(n770), .A2(n769), .A3(n768), .A4(n767), .Z(n777) );
  AOI22D1BWP12T U1429 ( .A1(tmp1[27]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[27]), .ZN(n773) );
  AOI22D0BWP12T U1430 ( .A1(r9[27]), .A2(n201), .B1(n2001), .B2(r4[27]), .ZN(
        n772) );
  AOI22D1BWP12T U1431 ( .A1(r11[27]), .A2(n1470), .B1(n205), .B2(r0[27]), .ZN(
        n771) );
  AN3XD1BWP12T U1432 ( .A1(n773), .A2(n772), .A3(n771), .Z(n776) );
  AOI22D1BWP12T U1433 ( .A1(r5[27]), .A2(n210), .B1(n1988), .B2(r10[27]), .ZN(
        n775) );
  AOI22D1BWP12T U1434 ( .A1(r7[27]), .A2(n215), .B1(n1989), .B2(r2[27]), .ZN(
        n774) );
  INVD1BWP12T U1435 ( .I(r4[23]), .ZN(n780) );
  AOI22D1BWP12T U1436 ( .A1(n150), .A2(r12[23]), .B1(n1486), .B2(tmp1[23]), 
        .ZN(n779) );
  AOI22D1BWP12T U1437 ( .A1(r2[23]), .A2(n155), .B1(n1555), .B2(r1[23]), .ZN(
        n778) );
  OA211D1BWP12T U1438 ( .A1(n780), .A2(n1458), .B(n779), .C(n778), .Z(n788) );
  AOI22D1BWP12T U1439 ( .A1(r9[23]), .A2(n1591), .B1(n1590), .B2(r6[23]), .ZN(
        n784) );
  AOI22D1BWP12T U1440 ( .A1(r8[23]), .A2(n1593), .B1(n1592), .B2(n[2018]), 
        .ZN(n783) );
  AOI22D1BWP12T U1441 ( .A1(r5[23]), .A2(n1594), .B1(n171), .B2(r3[23]), .ZN(
        n782) );
  AOI22D1BWP12T U1442 ( .A1(r7[23]), .A2(n1596), .B1(n1595), .B2(r0[23]), .ZN(
        n781) );
  AN4XD1BWP12T U1443 ( .A1(n784), .A2(n783), .A3(n782), .A4(n781), .Z(n787) );
  AOI22D1BWP12T U1444 ( .A1(pc_out[23]), .A2(n141), .B1(n1559), .B2(r11[23]), 
        .ZN(n786) );
  AOI22D1BWP12T U1445 ( .A1(lr[23]), .A2(n1561), .B1(n1560), .B2(r10[23]), 
        .ZN(n785) );
  ND4D2BWP12T U1446 ( .A1(n788), .A2(n787), .A3(n786), .A4(n785), .ZN(
        regA_out[23]) );
  INR2D2BWP12T U1447 ( .A1(next_cpsr_in[0]), .B1(reset), .ZN(cpsrin[0]) );
  INVD1BWP12T U1448 ( .I(lr[21]), .ZN(n791) );
  AOI22D1BWP12T U1449 ( .A1(pc_out[21]), .A2(n141), .B1(n1559), .B2(r11[21]), 
        .ZN(n790) );
  CKND2D1BWP12T U1450 ( .A1(n1560), .A2(r10[21]), .ZN(n789) );
  OA211D1BWP12T U1451 ( .A1(n1953), .A2(n791), .B(n790), .C(n789), .Z(n801) );
  INVD1BWP12T U1452 ( .I(r4[21]), .ZN(n794) );
  AOI22D1BWP12T U1453 ( .A1(n150), .A2(r12[21]), .B1(n1486), .B2(tmp1[21]), 
        .ZN(n793) );
  AOI22D1BWP12T U1454 ( .A1(r2[21]), .A2(n155), .B1(n1555), .B2(r1[21]), .ZN(
        n792) );
  OA211D1BWP12T U1455 ( .A1(n794), .A2(n1458), .B(n793), .C(n792), .Z(n800) );
  AOI22D1BWP12T U1456 ( .A1(r9[21]), .A2(n1591), .B1(n1590), .B2(r6[21]), .ZN(
        n798) );
  AOI22D1BWP12T U1457 ( .A1(r8[21]), .A2(n1593), .B1(n1592), .B2(n[2020]), 
        .ZN(n797) );
  AOI22D1BWP12T U1458 ( .A1(r5[21]), .A2(n1594), .B1(n171), .B2(r3[21]), .ZN(
        n796) );
  AOI22D1BWP12T U1459 ( .A1(r7[21]), .A2(n1596), .B1(n1595), .B2(r0[21]), .ZN(
        n795) );
  AN4XD1BWP12T U1460 ( .A1(n798), .A2(n797), .A3(n796), .A4(n795), .Z(n799) );
  ND3D2BWP12T U1461 ( .A1(n801), .A2(n800), .A3(n799), .ZN(regA_out[21]) );
  AO222D0BWP12T U1462 ( .A1(n1284), .A2(n1268), .B1(n1282), .B2(r6[28]), .C1(
        write2_in[28]), .C2(n1283), .Z(n2453) );
  AO222D0BWP12T U1463 ( .A1(n1302), .A2(n1268), .B1(n1300), .B2(r1[28]), .C1(
        write2_in[28]), .C2(n1301), .Z(n2613) );
  AO222D0BWP12T U1464 ( .A1(n1278), .A2(n1268), .B1(n1276), .B2(r0[28]), .C1(
        write2_in[28]), .C2(n1277), .Z(n2645) );
  AO222D0BWP12T U1465 ( .A1(n1296), .A2(n1268), .B1(n1294), .B2(r4[28]), .C1(
        write2_in[28]), .C2(n1295), .Z(n2517) );
  AO222D0BWP12T U1466 ( .A1(n1281), .A2(n1268), .B1(n1279), .B2(r12[28]), .C1(
        write2_in[28]), .C2(n1280), .Z(n2261) );
  AO222D0BWP12T U1467 ( .A1(n1299), .A2(n1268), .B1(n1297), .B2(r5[28]), .C1(
        write2_in[28]), .C2(n1298), .Z(n2485) );
  OAI22D1BWP12T U1468 ( .A1(n836), .A2(n1949), .B1(n1948), .B2(n802), .ZN(n809) );
  OAI22D1BWP12T U1469 ( .A1(n804), .A2(n1953), .B1(n1952), .B2(n803), .ZN(n808) );
  AOI22D1BWP12T U1470 ( .A1(n150), .A2(r12[3]), .B1(n1955), .B2(tmp1[3]), .ZN(
        n805) );
  IOA21D1BWP12T U1471 ( .A1(n1957), .A2(r4[3]), .B(n805), .ZN(n807) );
  OAI22D1BWP12T U1472 ( .A1(n1961), .A2(n828), .B1(n1959), .B2(n824), .ZN(n806) );
  NR4D1BWP12T U1473 ( .A1(n809), .A2(n808), .A3(n807), .A4(n806), .ZN(n818) );
  INVD3BWP12T U1474 ( .I(n1590), .ZN(n1967) );
  TPOAI22D1BWP12T U1475 ( .A1(n1969), .A2(n810), .B1(n1967), .B2(n827), .ZN(
        n816) );
  INVD3BWP12T U1476 ( .I(n1593), .ZN(n1973) );
  DCCKND4BWP12T U1477 ( .I(n1592), .ZN(n1971) );
  OAI22D1BWP12T U1478 ( .A1(n1973), .A2(n812), .B1(n1971), .B2(n811), .ZN(n815) );
  INVD2BWP12T U1479 ( .I(n1594), .ZN(n1976) );
  INVD2BWP12T U1480 ( .I(n171), .ZN(n1975) );
  OAI22D1BWP12T U1481 ( .A1(n825), .A2(n1976), .B1(n1975), .B2(n830), .ZN(n814) );
  INVD2BWP12T U1482 ( .I(n1596), .ZN(n1981) );
  INVD2BWP12T U1483 ( .I(n1595), .ZN(n1979) );
  OAI22D1BWP12T U1484 ( .A1(n1981), .A2(n822), .B1(n1979), .B2(n831), .ZN(n813) );
  NR4D1BWP12T U1485 ( .A1(n816), .A2(n815), .A3(n814), .A4(n813), .ZN(n817) );
  ND2D4BWP12T U1486 ( .A1(n818), .A2(n817), .ZN(regA_out[3]) );
  AO222D1BWP12T U1487 ( .A1(n1317), .A2(write1_in[2]), .B1(n820), .B2(
        write2_in[2]), .C1(n819), .C2(tmp1[2]), .Z(n2139) );
  IND2D1BWP12T U1488 ( .A1(readC_sel[0]), .B1(readC_sel[1]), .ZN(n842) );
  INVD1BWP12T U1489 ( .I(readC_sel[4]), .ZN(n1225) );
  ND3D1BWP12T U1490 ( .A1(readC_sel[2]), .A2(readC_sel[3]), .A3(n1225), .ZN(
        n844) );
  NR2D1BWP12T U1491 ( .A1(n842), .A2(n844), .ZN(n1214) );
  CKND0BWP12T U1492 ( .I(readC_sel[3]), .ZN(n823) );
  TPND2D0BWP12T U1493 ( .A1(readC_sel[2]), .A2(n823), .ZN(n826) );
  ND2D1BWP12T U1494 ( .A1(readC_sel[1]), .A2(readC_sel[0]), .ZN(n840) );
  OR2XD1BWP12T U1495 ( .A1(n826), .A2(n840), .Z(n1157) );
  OR2XD1BWP12T U1496 ( .A1(readC_sel[0]), .A2(readC_sel[1]), .Z(n843) );
  OR2XD1BWP12T U1497 ( .A1(n826), .A2(n843), .Z(n1156) );
  OAI22D0BWP12T U1498 ( .A1(n822), .A2(n1157), .B1(n1156), .B2(n821), .ZN(n835) );
  IND2D1BWP12T U1499 ( .A1(readC_sel[1]), .B1(readC_sel[0]), .ZN(n845) );
  OR2XD1BWP12T U1500 ( .A1(n845), .A2(n826), .Z(n1159) );
  INVD1BWP12T U1501 ( .I(readC_sel[2]), .ZN(n839) );
  TPND2D0BWP12T U1502 ( .A1(n839), .A2(n823), .ZN(n829) );
  OR2XD1BWP12T U1503 ( .A1(n845), .A2(n829), .Z(n1158) );
  OAI22D0BWP12T U1504 ( .A1(n825), .A2(n1159), .B1(n1158), .B2(n824), .ZN(n834) );
  OR2XD1BWP12T U1505 ( .A1(n842), .A2(n829), .Z(n1161) );
  OR2XD1BWP12T U1506 ( .A1(n826), .A2(n842), .Z(n1160) );
  OAI22D0BWP12T U1507 ( .A1(n1161), .A2(n828), .B1(n1160), .B2(n827), .ZN(n833) );
  OR2XD1BWP12T U1508 ( .A1(n829), .A2(n843), .Z(n1163) );
  OR2XD1BWP12T U1509 ( .A1(n829), .A2(n840), .Z(n1162) );
  OAI22D0BWP12T U1510 ( .A1(n831), .A2(n1163), .B1(n1162), .B2(n830), .ZN(n832) );
  NR4D0BWP12T U1511 ( .A1(n835), .A2(n834), .A3(n833), .A4(n832), .ZN(n837) );
  OR2XD1BWP12T U1512 ( .A1(n840), .A2(n844), .Z(n906) );
  OAI22D0BWP12T U1513 ( .A1(n837), .A2(readC_sel[4]), .B1(n906), .B2(n836), 
        .ZN(n838) );
  AOI21D0BWP12T U1514 ( .A1(lr[3]), .A2(n1214), .B(n838), .ZN(n849) );
  ND3D1BWP12T U1515 ( .A1(readC_sel[3]), .A2(n1225), .A3(n839), .ZN(n841) );
  OR2XD1BWP12T U1516 ( .A1(n845), .A2(n841), .Z(n1074) );
  INVD1BWP12T U1517 ( .I(n1074), .ZN(n1211) );
  OR2XD1BWP12T U1518 ( .A1(n840), .A2(n841), .Z(n1132) );
  INVD1BWP12T U1519 ( .I(n1132), .ZN(n1217) );
  AOI22D0BWP12T U1520 ( .A1(r9[3]), .A2(n1211), .B1(n1217), .B2(r11[3]), .ZN(
        n848) );
  NR2D1BWP12T U1521 ( .A1(n843), .A2(n841), .ZN(n1212) );
  OR2XD1BWP12T U1522 ( .A1(n842), .A2(n841), .Z(n1099) );
  INVD1BWP12T U1523 ( .I(n1099), .ZN(n1218) );
  AOI22D0BWP12T U1524 ( .A1(r8[3]), .A2(n1212), .B1(n1218), .B2(r10[3]), .ZN(
        n847) );
  NR2D1BWP12T U1525 ( .A1(n843), .A2(n844), .ZN(n1216) );
  NR2D1BWP12T U1526 ( .A1(n845), .A2(n844), .ZN(n1213) );
  AOI22D0BWP12T U1527 ( .A1(r12[3]), .A2(n1216), .B1(n1213), .B2(n[2038]), 
        .ZN(n846) );
  ND4D1BWP12T U1528 ( .A1(n849), .A2(n848), .A3(n847), .A4(n846), .ZN(
        regC_out[3]) );
  OAI22D0BWP12T U1529 ( .A1(n1980), .A2(n1157), .B1(n1156), .B2(n850), .ZN(
        n854) );
  OAI22D0BWP12T U1530 ( .A1(n1977), .A2(n1159), .B1(n1158), .B2(n1958), .ZN(
        n853) );
  OAI22D0BWP12T U1531 ( .A1(n1161), .A2(n1960), .B1(n1160), .B2(n1966), .ZN(
        n852) );
  OAI22D0BWP12T U1532 ( .A1(n1978), .A2(n1163), .B1(n1162), .B2(n1974), .ZN(
        n851) );
  NR4D0BWP12T U1533 ( .A1(n854), .A2(n853), .A3(n852), .A4(n851), .ZN(n855) );
  OAI22D0BWP12T U1534 ( .A1(n855), .A2(readC_sel[4]), .B1(n906), .B2(n1950), 
        .ZN(n856) );
  AOI21D0BWP12T U1535 ( .A1(lr[2]), .A2(n1214), .B(n856), .ZN(n860) );
  AOI22D0BWP12T U1536 ( .A1(r9[2]), .A2(n1211), .B1(n1217), .B2(r11[2]), .ZN(
        n859) );
  AOI22D0BWP12T U1537 ( .A1(r8[2]), .A2(n1212), .B1(n1218), .B2(r10[2]), .ZN(
        n858) );
  AOI22D0BWP12T U1538 ( .A1(r12[2]), .A2(n1216), .B1(n1213), .B2(n[2039]), 
        .ZN(n857) );
  ND4D1BWP12T U1539 ( .A1(n860), .A2(n859), .A3(n858), .A4(n857), .ZN(
        regC_out[2]) );
  AOI22D0BWP12T U1540 ( .A1(r12[25]), .A2(n1216), .B1(n1211), .B2(r9[25]), 
        .ZN(n872) );
  AOI22D0BWP12T U1541 ( .A1(lr[25]), .A2(n1214), .B1(n1213), .B2(n[2016]), 
        .ZN(n871) );
  AOI22D0BWP12T U1542 ( .A1(r10[25]), .A2(n1218), .B1(n1217), .B2(r11[25]), 
        .ZN(n870) );
  AOI22D0BWP12T U1543 ( .A1(r7[25]), .A2(n1200), .B1(n1199), .B2(r4[25]), .ZN(
        n864) );
  AOI22D0BWP12T U1544 ( .A1(r2[25]), .A2(n1202), .B1(n1201), .B2(r6[25]), .ZN(
        n863) );
  AOI22D0BWP12T U1545 ( .A1(r5[25]), .A2(n1204), .B1(n1203), .B2(r1[25]), .ZN(
        n862) );
  AOI22D0BWP12T U1546 ( .A1(r0[25]), .A2(n1206), .B1(n1205), .B2(r3[25]), .ZN(
        n861) );
  ND4D1BWP12T U1547 ( .A1(n864), .A2(n863), .A3(n862), .A4(n861), .ZN(n868) );
  CKND0BWP12T U1548 ( .I(pc_out[25]), .ZN(n866) );
  INVD1BWP12T U1549 ( .I(n1212), .ZN(n1136) );
  CKND0BWP12T U1550 ( .I(r8[25]), .ZN(n865) );
  OAI22D0BWP12T U1551 ( .A1(n866), .A2(n906), .B1(n1136), .B2(n865), .ZN(n867)
         );
  AOI21D0BWP12T U1552 ( .A1(n868), .A2(n1225), .B(n867), .ZN(n869) );
  ND4D1BWP12T U1553 ( .A1(n872), .A2(n871), .A3(n870), .A4(n869), .ZN(
        regC_out[25]) );
  AOI22D0BWP12T U1554 ( .A1(r8[4]), .A2(n1212), .B1(n1218), .B2(r10[4]), .ZN(
        n882) );
  AOI22D0BWP12T U1555 ( .A1(r12[4]), .A2(n1216), .B1(n1213), .B2(n[2037]), 
        .ZN(n881) );
  AOI22D0BWP12T U1556 ( .A1(r9[4]), .A2(n1211), .B1(n1217), .B2(r11[4]), .ZN(
        n880) );
  AOI22D0BWP12T U1557 ( .A1(r7[4]), .A2(n1200), .B1(n1199), .B2(r4[4]), .ZN(
        n876) );
  AOI22D0BWP12T U1558 ( .A1(r2[4]), .A2(n1202), .B1(n1201), .B2(r6[4]), .ZN(
        n875) );
  AOI22D0BWP12T U1559 ( .A1(r5[4]), .A2(n1204), .B1(n1203), .B2(r1[4]), .ZN(
        n874) );
  AOI22D0BWP12T U1560 ( .A1(r0[4]), .A2(n1206), .B1(n1205), .B2(r3[4]), .ZN(
        n873) );
  ND4D1BWP12T U1561 ( .A1(n876), .A2(n875), .A3(n874), .A4(n873), .ZN(n878) );
  INVD1BWP12T U1562 ( .I(n1214), .ZN(n1181) );
  OAI22D0BWP12T U1563 ( .A1(n1873), .A2(n906), .B1(n1181), .B2(n1875), .ZN(
        n877) );
  AOI21D0BWP12T U1564 ( .A1(n878), .A2(n1225), .B(n877), .ZN(n879) );
  ND4D1BWP12T U1565 ( .A1(n882), .A2(n881), .A3(n880), .A4(n879), .ZN(
        regC_out[4]) );
  AOI22D0BWP12T U1566 ( .A1(r8[12]), .A2(n1212), .B1(n1211), .B2(r9[12]), .ZN(
        n893) );
  AOI22D0BWP12T U1567 ( .A1(lr[12]), .A2(n1214), .B1(n1213), .B2(n[2029]), 
        .ZN(n892) );
  AOI22D0BWP12T U1568 ( .A1(r10[12]), .A2(n1218), .B1(n1217), .B2(r11[12]), 
        .ZN(n891) );
  AOI22D0BWP12T U1569 ( .A1(r7[12]), .A2(n1200), .B1(n1199), .B2(r4[12]), .ZN(
        n886) );
  AOI22D0BWP12T U1570 ( .A1(r2[12]), .A2(n1202), .B1(n1201), .B2(r6[12]), .ZN(
        n885) );
  AOI22D0BWP12T U1571 ( .A1(r5[12]), .A2(n1204), .B1(n1203), .B2(r1[12]), .ZN(
        n884) );
  AOI22D0BWP12T U1572 ( .A1(r0[12]), .A2(n1206), .B1(n1205), .B2(r3[12]), .ZN(
        n883) );
  ND4D1BWP12T U1573 ( .A1(n886), .A2(n885), .A3(n884), .A4(n883), .ZN(n889) );
  INVD1BWP12T U1574 ( .I(n1216), .ZN(n1193) );
  OAI22D0BWP12T U1575 ( .A1(n1630), .A2(n906), .B1(n1193), .B2(n887), .ZN(n888) );
  AOI21D0BWP12T U1576 ( .A1(n889), .A2(n1225), .B(n888), .ZN(n890) );
  ND4D1BWP12T U1577 ( .A1(n893), .A2(n892), .A3(n891), .A4(n890), .ZN(
        regC_out[12]) );
  AOI22D0BWP12T U1578 ( .A1(r8[26]), .A2(n1212), .B1(n1211), .B2(r9[26]), .ZN(
        n905) );
  AOI22D0BWP12T U1579 ( .A1(lr[26]), .A2(n1214), .B1(n1216), .B2(r12[26]), 
        .ZN(n904) );
  AOI22D0BWP12T U1580 ( .A1(r10[26]), .A2(n1218), .B1(n1217), .B2(r11[26]), 
        .ZN(n903) );
  AOI22D0BWP12T U1581 ( .A1(r7[26]), .A2(n1200), .B1(n1199), .B2(r4[26]), .ZN(
        n897) );
  AOI22D0BWP12T U1582 ( .A1(r2[26]), .A2(n1202), .B1(n1201), .B2(r6[26]), .ZN(
        n896) );
  AOI22D0BWP12T U1583 ( .A1(r5[26]), .A2(n1204), .B1(n1203), .B2(r1[26]), .ZN(
        n895) );
  AOI22D0BWP12T U1584 ( .A1(r0[26]), .A2(n1206), .B1(n1205), .B2(r3[26]), .ZN(
        n894) );
  ND4D1BWP12T U1585 ( .A1(n897), .A2(n896), .A3(n895), .A4(n894), .ZN(n901) );
  CKND0BWP12T U1586 ( .I(pc_out[26]), .ZN(n899) );
  CKND0BWP12T U1587 ( .I(n[2015]), .ZN(n898) );
  INVD1BWP12T U1588 ( .I(n1213), .ZN(n1168) );
  OAI22D0BWP12T U1589 ( .A1(n899), .A2(n906), .B1(n898), .B2(n1168), .ZN(n900)
         );
  AOI21D0BWP12T U1590 ( .A1(n901), .A2(n1225), .B(n900), .ZN(n902) );
  ND4D1BWP12T U1591 ( .A1(n905), .A2(n904), .A3(n903), .A4(n902), .ZN(
        regC_out[26]) );
  INVD1BWP12T U1592 ( .I(n906), .ZN(n1215) );
  AOI22D0BWP12T U1593 ( .A1(pc_out[24]), .A2(n1215), .B1(n1212), .B2(r8[24]), 
        .ZN(n920) );
  AOI22D0BWP12T U1594 ( .A1(r9[24]), .A2(n1211), .B1(n1217), .B2(r11[24]), 
        .ZN(n919) );
  AOI22D0BWP12T U1595 ( .A1(r7[24]), .A2(n1200), .B1(n1199), .B2(r4[24]), .ZN(
        n910) );
  AOI22D0BWP12T U1596 ( .A1(r2[24]), .A2(n1202), .B1(n1201), .B2(r6[24]), .ZN(
        n909) );
  AOI22D0BWP12T U1597 ( .A1(r5[24]), .A2(n1204), .B1(n1203), .B2(r1[24]), .ZN(
        n908) );
  AOI22D0BWP12T U1598 ( .A1(r0[24]), .A2(n1206), .B1(n1205), .B2(r3[24]), .ZN(
        n907) );
  ND4D1BWP12T U1599 ( .A1(n910), .A2(n909), .A3(n908), .A4(n907), .ZN(n917) );
  CKND0BWP12T U1600 ( .I(r12[24]), .ZN(n912) );
  CKND0BWP12T U1601 ( .I(r10[24]), .ZN(n911) );
  OAI22D0BWP12T U1602 ( .A1(n1193), .A2(n912), .B1(n911), .B2(n1099), .ZN(n916) );
  CKND0BWP12T U1603 ( .I(n[2017]), .ZN(n914) );
  CKND0BWP12T U1604 ( .I(lr[24]), .ZN(n913) );
  OAI22D0BWP12T U1605 ( .A1(n914), .A2(n1168), .B1(n1181), .B2(n913), .ZN(n915) );
  AOI211D0BWP12T U1606 ( .A1(n917), .A2(n1225), .B(n916), .C(n915), .ZN(n918)
         );
  ND3D1BWP12T U1607 ( .A1(n920), .A2(n919), .A3(n918), .ZN(regC_out[24]) );
  AOI22D0BWP12T U1608 ( .A1(pc_out[27]), .A2(n1215), .B1(n1212), .B2(r8[27]), 
        .ZN(n932) );
  AOI22D0BWP12T U1609 ( .A1(lr[27]), .A2(n1214), .B1(n1216), .B2(r12[27]), 
        .ZN(n931) );
  AOI22D0BWP12T U1610 ( .A1(r9[27]), .A2(n1211), .B1(n1218), .B2(r10[27]), 
        .ZN(n930) );
  AOI22D0BWP12T U1611 ( .A1(r7[27]), .A2(n1200), .B1(n1199), .B2(r4[27]), .ZN(
        n924) );
  AOI22D0BWP12T U1612 ( .A1(r2[27]), .A2(n1202), .B1(n1201), .B2(r6[27]), .ZN(
        n923) );
  AOI22D0BWP12T U1613 ( .A1(r5[27]), .A2(n1204), .B1(n1203), .B2(r1[27]), .ZN(
        n922) );
  AOI22D0BWP12T U1614 ( .A1(r0[27]), .A2(n1206), .B1(n1205), .B2(r3[27]), .ZN(
        n921) );
  ND4D1BWP12T U1615 ( .A1(n924), .A2(n923), .A3(n922), .A4(n921), .ZN(n928) );
  CKND0BWP12T U1616 ( .I(n[2014]), .ZN(n926) );
  CKND0BWP12T U1617 ( .I(r11[27]), .ZN(n925) );
  OAI22D0BWP12T U1618 ( .A1(n926), .A2(n1168), .B1(n1132), .B2(n925), .ZN(n927) );
  AOI21D0BWP12T U1619 ( .A1(n928), .A2(n1225), .B(n927), .ZN(n929) );
  ND4D1BWP12T U1620 ( .A1(n932), .A2(n931), .A3(n930), .A4(n929), .ZN(
        regC_out[27]) );
  AOI22D0BWP12T U1621 ( .A1(pc_out[29]), .A2(n1215), .B1(n1212), .B2(r8[29]), 
        .ZN(n944) );
  AOI22D0BWP12T U1622 ( .A1(lr[29]), .A2(n1214), .B1(n1216), .B2(r12[29]), 
        .ZN(n943) );
  AOI22D0BWP12T U1623 ( .A1(r10[29]), .A2(n1218), .B1(n1217), .B2(r11[29]), 
        .ZN(n942) );
  AOI22D0BWP12T U1624 ( .A1(r7[29]), .A2(n1200), .B1(n1199), .B2(r4[29]), .ZN(
        n936) );
  AOI22D0BWP12T U1625 ( .A1(r2[29]), .A2(n1202), .B1(n1201), .B2(r6[29]), .ZN(
        n935) );
  AOI22D0BWP12T U1626 ( .A1(r5[29]), .A2(n1204), .B1(n1203), .B2(r1[29]), .ZN(
        n934) );
  AOI22D0BWP12T U1627 ( .A1(r0[29]), .A2(n1206), .B1(n1205), .B2(r3[29]), .ZN(
        n933) );
  ND4D1BWP12T U1628 ( .A1(n936), .A2(n935), .A3(n934), .A4(n933), .ZN(n940) );
  CKND0BWP12T U1629 ( .I(n[2012]), .ZN(n938) );
  CKND0BWP12T U1630 ( .I(r9[29]), .ZN(n937) );
  OAI22D0BWP12T U1631 ( .A1(n938), .A2(n1168), .B1(n1074), .B2(n937), .ZN(n939) );
  AOI21D0BWP12T U1632 ( .A1(n940), .A2(n1225), .B(n939), .ZN(n941) );
  ND4D1BWP12T U1633 ( .A1(n944), .A2(n943), .A3(n942), .A4(n941), .ZN(
        regC_out[29]) );
  AOI22D0BWP12T U1634 ( .A1(pc_out[15]), .A2(n1215), .B1(n1218), .B2(r10[15]), 
        .ZN(n955) );
  AOI22D0BWP12T U1635 ( .A1(n[2026]), .A2(n1213), .B1(n1216), .B2(r12[15]), 
        .ZN(n954) );
  AOI22D0BWP12T U1636 ( .A1(r9[15]), .A2(n1211), .B1(n1217), .B2(r11[15]), 
        .ZN(n953) );
  AOI22D0BWP12T U1637 ( .A1(r7[15]), .A2(n1200), .B1(n1199), .B2(r4[15]), .ZN(
        n948) );
  AOI22D0BWP12T U1638 ( .A1(r2[15]), .A2(n1202), .B1(n1201), .B2(r6[15]), .ZN(
        n947) );
  AOI22D0BWP12T U1639 ( .A1(r5[15]), .A2(n1204), .B1(n1203), .B2(r1[15]), .ZN(
        n946) );
  AOI22D0BWP12T U1640 ( .A1(r0[15]), .A2(n1206), .B1(n1205), .B2(r3[15]), .ZN(
        n945) );
  ND4D1BWP12T U1641 ( .A1(n948), .A2(n947), .A3(n946), .A4(n945), .ZN(n951) );
  INVD1BWP12T U1642 ( .I(lr[15]), .ZN(n1582) );
  CKND0BWP12T U1643 ( .I(r8[15]), .ZN(n949) );
  OAI22D0BWP12T U1644 ( .A1(n1181), .A2(n1582), .B1(n949), .B2(n1136), .ZN(
        n950) );
  AOI21D0BWP12T U1645 ( .A1(n951), .A2(n1225), .B(n950), .ZN(n952) );
  ND4D1BWP12T U1646 ( .A1(n955), .A2(n954), .A3(n953), .A4(n952), .ZN(
        regC_out[15]) );
  AOI22D0BWP12T U1647 ( .A1(pc_out[8]), .A2(n1215), .B1(n1211), .B2(r9[8]), 
        .ZN(n966) );
  AOI22D0BWP12T U1648 ( .A1(lr[8]), .A2(n1214), .B1(n1213), .B2(n[2033]), .ZN(
        n965) );
  AOI22D0BWP12T U1649 ( .A1(r10[8]), .A2(n1218), .B1(n1217), .B2(r11[8]), .ZN(
        n964) );
  AOI22D0BWP12T U1650 ( .A1(r7[8]), .A2(n1200), .B1(n1199), .B2(r4[8]), .ZN(
        n959) );
  AOI22D0BWP12T U1651 ( .A1(r2[8]), .A2(n1202), .B1(n1201), .B2(r6[8]), .ZN(
        n958) );
  AOI22D0BWP12T U1652 ( .A1(r5[8]), .A2(n1204), .B1(n1203), .B2(r1[8]), .ZN(
        n957) );
  AOI22D0BWP12T U1653 ( .A1(r0[8]), .A2(n1206), .B1(n1205), .B2(r3[8]), .ZN(
        n956) );
  ND4D1BWP12T U1654 ( .A1(n959), .A2(n958), .A3(n957), .A4(n956), .ZN(n962) );
  OAI22D0BWP12T U1655 ( .A1(n1193), .A2(n960), .B1(n1754), .B2(n1136), .ZN(
        n961) );
  AOI21D0BWP12T U1656 ( .A1(n962), .A2(n1225), .B(n961), .ZN(n963) );
  ND4D1BWP12T U1657 ( .A1(n966), .A2(n965), .A3(n964), .A4(n963), .ZN(
        regC_out[8]) );
  AOI22D0BWP12T U1658 ( .A1(n[2040]), .A2(n1213), .B1(n1218), .B2(r10[1]), 
        .ZN(n977) );
  AOI22D0BWP12T U1659 ( .A1(r9[1]), .A2(n1211), .B1(n1217), .B2(r11[1]), .ZN(
        n976) );
  OAI22D0BWP12T U1660 ( .A1(n1181), .A2(n1925), .B1(n1936), .B2(n1136), .ZN(
        n968) );
  NR2D0BWP12T U1661 ( .A1(n1857), .A2(n1193), .ZN(n967) );
  AOI211D0BWP12T U1662 ( .A1(pc_out[1]), .A2(n1215), .B(n968), .C(n967), .ZN(
        n975) );
  AOI22D0BWP12T U1663 ( .A1(r7[1]), .A2(n1200), .B1(n1199), .B2(r4[1]), .ZN(
        n972) );
  AOI22D0BWP12T U1664 ( .A1(r2[1]), .A2(n1202), .B1(n1201), .B2(r6[1]), .ZN(
        n971) );
  AOI22D0BWP12T U1665 ( .A1(r5[1]), .A2(n1204), .B1(n1203), .B2(r1[1]), .ZN(
        n970) );
  AOI22D0BWP12T U1666 ( .A1(r0[1]), .A2(n1206), .B1(n1205), .B2(r3[1]), .ZN(
        n969) );
  ND4D1BWP12T U1667 ( .A1(n972), .A2(n971), .A3(n970), .A4(n969), .ZN(n973) );
  CKND2D0BWP12T U1668 ( .A1(n973), .A2(n1225), .ZN(n974) );
  ND4D1BWP12T U1669 ( .A1(n977), .A2(n976), .A3(n975), .A4(n974), .ZN(
        regC_out[1]) );
  AOI22D0BWP12T U1670 ( .A1(pc_out[18]), .A2(n1215), .B1(n1211), .B2(r9[18]), 
        .ZN(n989) );
  AOI22D0BWP12T U1671 ( .A1(lr[18]), .A2(n1214), .B1(n1213), .B2(n[2023]), 
        .ZN(n988) );
  AOI22D0BWP12T U1672 ( .A1(r10[18]), .A2(n1218), .B1(n1217), .B2(r11[18]), 
        .ZN(n987) );
  AOI22D0BWP12T U1673 ( .A1(r7[18]), .A2(n1200), .B1(n1199), .B2(r4[18]), .ZN(
        n981) );
  AOI22D0BWP12T U1674 ( .A1(r2[18]), .A2(n1202), .B1(n1201), .B2(r6[18]), .ZN(
        n980) );
  AOI22D0BWP12T U1675 ( .A1(r5[18]), .A2(n1204), .B1(n1203), .B2(r1[18]), .ZN(
        n979) );
  AOI22D0BWP12T U1676 ( .A1(r0[18]), .A2(n1206), .B1(n1205), .B2(r3[18]), .ZN(
        n978) );
  ND4D1BWP12T U1677 ( .A1(n981), .A2(n980), .A3(n979), .A4(n978), .ZN(n985) );
  CKND0BWP12T U1678 ( .I(r12[18]), .ZN(n983) );
  CKND0BWP12T U1679 ( .I(r8[18]), .ZN(n982) );
  TPOAI22D0BWP12T U1680 ( .A1(n1193), .A2(n983), .B1(n982), .B2(n1136), .ZN(
        n984) );
  AOI21D0BWP12T U1681 ( .A1(n985), .A2(n1225), .B(n984), .ZN(n986) );
  ND4D1BWP12T U1682 ( .A1(n989), .A2(n988), .A3(n987), .A4(n986), .ZN(
        regC_out[18]) );
  AOI22D0BWP12T U1683 ( .A1(pc_out[0]), .A2(n1215), .B1(n1212), .B2(r8[0]), 
        .ZN(n1001) );
  AOI22D0BWP12T U1684 ( .A1(n[2041]), .A2(n1213), .B1(n1216), .B2(r12[0]), 
        .ZN(n1000) );
  AOI22D0BWP12T U1685 ( .A1(r9[0]), .A2(n1211), .B1(n1217), .B2(r11[0]), .ZN(
        n999) );
  AOI22D0BWP12T U1686 ( .A1(r7[0]), .A2(n1200), .B1(n1199), .B2(r4[0]), .ZN(
        n993) );
  AOI22D0BWP12T U1687 ( .A1(r2[0]), .A2(n1202), .B1(n1201), .B2(r6[0]), .ZN(
        n992) );
  AOI22D0BWP12T U1688 ( .A1(r5[0]), .A2(n1204), .B1(n1203), .B2(r1[0]), .ZN(
        n991) );
  AOI22D0BWP12T U1689 ( .A1(r0[0]), .A2(n1206), .B1(n1205), .B2(r3[0]), .ZN(
        n990) );
  ND4D1BWP12T U1690 ( .A1(n993), .A2(n992), .A3(n991), .A4(n990), .ZN(n997) );
  OAI22D0BWP12T U1691 ( .A1(n1181), .A2(n995), .B1(n994), .B2(n1099), .ZN(n996) );
  AOI21D0BWP12T U1692 ( .A1(n997), .A2(n1225), .B(n996), .ZN(n998) );
  ND4D1BWP12T U1693 ( .A1(n1001), .A2(n1000), .A3(n999), .A4(n998), .ZN(
        regC_out[0]) );
  AOI22D0BWP12T U1694 ( .A1(pc_out[5]), .A2(n1215), .B1(n1212), .B2(r8[5]), 
        .ZN(n1011) );
  AOI22D0BWP12T U1695 ( .A1(r12[5]), .A2(n1216), .B1(n1213), .B2(n[2036]), 
        .ZN(n1010) );
  AOI22D0BWP12T U1696 ( .A1(r10[5]), .A2(n1218), .B1(n1217), .B2(r11[5]), .ZN(
        n1009) );
  AOI22D0BWP12T U1697 ( .A1(r7[5]), .A2(n1200), .B1(n1199), .B2(r4[5]), .ZN(
        n1005) );
  AOI22D0BWP12T U1698 ( .A1(r2[5]), .A2(n1202), .B1(n1201), .B2(r6[5]), .ZN(
        n1004) );
  AOI22D0BWP12T U1699 ( .A1(r5[5]), .A2(n1204), .B1(n1203), .B2(r1[5]), .ZN(
        n1003) );
  AOI22D0BWP12T U1700 ( .A1(r0[5]), .A2(n1206), .B1(n1205), .B2(r3[5]), .ZN(
        n1002) );
  ND4D1BWP12T U1701 ( .A1(n1005), .A2(n1004), .A3(n1003), .A4(n1002), .ZN(
        n1007) );
  OAI22D0BWP12T U1702 ( .A1(n1181), .A2(n1900), .B1(n1909), .B2(n1074), .ZN(
        n1006) );
  AOI21D0BWP12T U1703 ( .A1(n1007), .A2(n1225), .B(n1006), .ZN(n1008) );
  ND4D1BWP12T U1704 ( .A1(n1011), .A2(n1010), .A3(n1009), .A4(n1008), .ZN(
        regC_out[5]) );
  AOI22D0BWP12T U1705 ( .A1(pc_out[19]), .A2(n1215), .B1(n1212), .B2(r8[19]), 
        .ZN(n1022) );
  AOI22D0BWP12T U1706 ( .A1(n[2022]), .A2(n1213), .B1(n1216), .B2(r12[19]), 
        .ZN(n1021) );
  AOI22D0BWP12T U1707 ( .A1(r10[19]), .A2(n1218), .B1(n1217), .B2(r11[19]), 
        .ZN(n1020) );
  AOI22D0BWP12T U1708 ( .A1(r7[19]), .A2(n1200), .B1(n1199), .B2(r4[19]), .ZN(
        n1015) );
  AOI22D0BWP12T U1709 ( .A1(r2[19]), .A2(n1202), .B1(n1201), .B2(r6[19]), .ZN(
        n1014) );
  AOI22D0BWP12T U1710 ( .A1(r5[19]), .A2(n1204), .B1(n1203), .B2(r1[19]), .ZN(
        n1013) );
  AOI22D0BWP12T U1711 ( .A1(r0[19]), .A2(n1206), .B1(n1205), .B2(r3[19]), .ZN(
        n1012) );
  ND4D1BWP12T U1712 ( .A1(n1015), .A2(n1014), .A3(n1013), .A4(n1012), .ZN(
        n1018) );
  INVD1BWP12T U1713 ( .I(lr[19]), .ZN(n1485) );
  CKND0BWP12T U1714 ( .I(r9[19]), .ZN(n1016) );
  OAI22D0BWP12T U1715 ( .A1(n1181), .A2(n1485), .B1(n1016), .B2(n1074), .ZN(
        n1017) );
  AOI21D0BWP12T U1716 ( .A1(n1018), .A2(n1225), .B(n1017), .ZN(n1019) );
  ND4D1BWP12T U1717 ( .A1(n1022), .A2(n1021), .A3(n1020), .A4(n1019), .ZN(
        regC_out[19]) );
  AOI22D0BWP12T U1718 ( .A1(pc_out[20]), .A2(n1215), .B1(n1212), .B2(r8[20]), 
        .ZN(n1034) );
  AOI22D0BWP12T U1719 ( .A1(lr[20]), .A2(n1214), .B1(n1216), .B2(r12[20]), 
        .ZN(n1033) );
  AOI22D0BWP12T U1720 ( .A1(r9[20]), .A2(n1211), .B1(n1218), .B2(r10[20]), 
        .ZN(n1032) );
  AOI22D0BWP12T U1721 ( .A1(r7[20]), .A2(n1200), .B1(n1199), .B2(r4[20]), .ZN(
        n1026) );
  AOI22D0BWP12T U1722 ( .A1(r2[20]), .A2(n1202), .B1(n1201), .B2(r6[20]), .ZN(
        n1025) );
  AOI22D0BWP12T U1723 ( .A1(r5[20]), .A2(n1204), .B1(n1203), .B2(r1[20]), .ZN(
        n1024) );
  AOI22D0BWP12T U1724 ( .A1(r0[20]), .A2(n1206), .B1(n1205), .B2(r3[20]), .ZN(
        n1023) );
  ND4D1BWP12T U1725 ( .A1(n1026), .A2(n1025), .A3(n1024), .A4(n1023), .ZN(
        n1030) );
  CKND0BWP12T U1726 ( .I(n[2021]), .ZN(n1028) );
  OAI22D0BWP12T U1727 ( .A1(n1028), .A2(n1168), .B1(n1132), .B2(n1027), .ZN(
        n1029) );
  AOI21D0BWP12T U1728 ( .A1(n1030), .A2(n1225), .B(n1029), .ZN(n1031) );
  ND4D1BWP12T U1729 ( .A1(n1034), .A2(n1033), .A3(n1032), .A4(n1031), .ZN(
        regC_out[20]) );
  CKND0BWP12T U1730 ( .I(r8[23]), .ZN(n1040) );
  AOI22D0BWP12T U1731 ( .A1(r7[23]), .A2(n1200), .B1(n1199), .B2(r4[23]), .ZN(
        n1038) );
  AOI22D0BWP12T U1732 ( .A1(r2[23]), .A2(n1202), .B1(n1201), .B2(r6[23]), .ZN(
        n1037) );
  AOI22D0BWP12T U1733 ( .A1(r5[23]), .A2(n1204), .B1(n1203), .B2(r1[23]), .ZN(
        n1036) );
  AOI22D0BWP12T U1734 ( .A1(r0[23]), .A2(n1206), .B1(n1205), .B2(r3[23]), .ZN(
        n1035) );
  ND4D1BWP12T U1735 ( .A1(n1038), .A2(n1037), .A3(n1036), .A4(n1035), .ZN(
        n1039) );
  MOAI22D0BWP12T U1736 ( .A1(n1136), .A2(n1040), .B1(n1039), .B2(n1225), .ZN(
        n1041) );
  AOI21D0BWP12T U1737 ( .A1(lr[23]), .A2(n1214), .B(n1041), .ZN(n1045) );
  AOI22D0BWP12T U1738 ( .A1(r9[23]), .A2(n1211), .B1(n1217), .B2(r11[23]), 
        .ZN(n1044) );
  AOI22D0BWP12T U1739 ( .A1(pc_out[23]), .A2(n1215), .B1(n1218), .B2(r10[23]), 
        .ZN(n1043) );
  AOI22D0BWP12T U1740 ( .A1(n[2018]), .A2(n1213), .B1(n1216), .B2(r12[23]), 
        .ZN(n1042) );
  ND4D1BWP12T U1741 ( .A1(n1045), .A2(n1044), .A3(n1043), .A4(n1042), .ZN(
        regC_out[23]) );
  AOI22D0BWP12T U1742 ( .A1(r12[31]), .A2(n1216), .B1(n1215), .B2(pc_out[31]), 
        .ZN(n1057) );
  AOI22D0BWP12T U1743 ( .A1(lr[31]), .A2(n1214), .B1(n1213), .B2(n[2010]), 
        .ZN(n1056) );
  AOI22D0BWP12T U1744 ( .A1(r8[31]), .A2(n1212), .B1(n1217), .B2(r11[31]), 
        .ZN(n1055) );
  AOI22D0BWP12T U1745 ( .A1(r7[31]), .A2(n1200), .B1(n1199), .B2(r4[31]), .ZN(
        n1049) );
  AOI22D0BWP12T U1746 ( .A1(r2[31]), .A2(n1202), .B1(n1201), .B2(r6[31]), .ZN(
        n1048) );
  AOI22D0BWP12T U1747 ( .A1(r5[31]), .A2(n1204), .B1(n1203), .B2(r1[31]), .ZN(
        n1047) );
  AOI22D0BWP12T U1748 ( .A1(r0[31]), .A2(n1206), .B1(n1205), .B2(r3[31]), .ZN(
        n1046) );
  ND4D1BWP12T U1749 ( .A1(n1049), .A2(n1048), .A3(n1047), .A4(n1046), .ZN(
        n1053) );
  CKND0BWP12T U1750 ( .I(r9[31]), .ZN(n1051) );
  CKND0BWP12T U1751 ( .I(r10[31]), .ZN(n1050) );
  OAI22D0BWP12T U1752 ( .A1(n1074), .A2(n1051), .B1(n1050), .B2(n1099), .ZN(
        n1052) );
  AOI21D0BWP12T U1753 ( .A1(n1053), .A2(n1225), .B(n1052), .ZN(n1054) );
  ND4D1BWP12T U1754 ( .A1(n1057), .A2(n1056), .A3(n1055), .A4(n1054), .ZN(
        regC_out[31]) );
  AOI22D0BWP12T U1755 ( .A1(r8[28]), .A2(n1212), .B1(n1218), .B2(r10[28]), 
        .ZN(n1069) );
  AOI22D0BWP12T U1756 ( .A1(n[2013]), .A2(n1213), .B1(n1215), .B2(pc_out[28]), 
        .ZN(n1068) );
  AOI22D0BWP12T U1757 ( .A1(r9[28]), .A2(n1211), .B1(n1217), .B2(r11[28]), 
        .ZN(n1067) );
  AOI22D0BWP12T U1758 ( .A1(r7[28]), .A2(n1200), .B1(n1199), .B2(r4[28]), .ZN(
        n1061) );
  AOI22D0BWP12T U1759 ( .A1(r2[28]), .A2(n1202), .B1(n1201), .B2(r6[28]), .ZN(
        n1060) );
  AOI22D0BWP12T U1760 ( .A1(r5[28]), .A2(n1204), .B1(n1203), .B2(r1[28]), .ZN(
        n1059) );
  AOI22D0BWP12T U1761 ( .A1(r0[28]), .A2(n1206), .B1(n1205), .B2(r3[28]), .ZN(
        n1058) );
  ND4D1BWP12T U1762 ( .A1(n1061), .A2(n1060), .A3(n1059), .A4(n1058), .ZN(
        n1065) );
  CKND0BWP12T U1763 ( .I(lr[28]), .ZN(n1063) );
  CKND0BWP12T U1764 ( .I(r12[28]), .ZN(n1062) );
  TPOAI22D0BWP12T U1765 ( .A1(n1181), .A2(n1063), .B1(n1062), .B2(n1193), .ZN(
        n1064) );
  AOI21D0BWP12T U1766 ( .A1(n1065), .A2(n1225), .B(n1064), .ZN(n1066) );
  ND4D1BWP12T U1767 ( .A1(n1069), .A2(n1068), .A3(n1067), .A4(n1066), .ZN(
        regC_out[28]) );
  AOI22D0BWP12T U1768 ( .A1(r12[9]), .A2(n1216), .B1(n1215), .B2(pc_out[9]), 
        .ZN(n1080) );
  AOI22D0BWP12T U1769 ( .A1(lr[9]), .A2(n1214), .B1(n1213), .B2(n[2032]), .ZN(
        n1079) );
  AOI22D0BWP12T U1770 ( .A1(r10[9]), .A2(n1218), .B1(n1217), .B2(r11[9]), .ZN(
        n1078) );
  AOI22D0BWP12T U1771 ( .A1(r7[9]), .A2(n1200), .B1(n1199), .B2(r4[9]), .ZN(
        n1073) );
  AOI22D0BWP12T U1772 ( .A1(r2[9]), .A2(n1202), .B1(n1201), .B2(r6[9]), .ZN(
        n1072) );
  AOI22D0BWP12T U1773 ( .A1(r5[9]), .A2(n1204), .B1(n1203), .B2(r1[9]), .ZN(
        n1071) );
  AOI22D0BWP12T U1774 ( .A1(r0[9]), .A2(n1206), .B1(n1205), .B2(r3[9]), .ZN(
        n1070) );
  ND4D1BWP12T U1775 ( .A1(n1073), .A2(n1072), .A3(n1071), .A4(n1070), .ZN(
        n1076) );
  OAI22D0BWP12T U1776 ( .A1(n1136), .A2(n1731), .B1(n1707), .B2(n1074), .ZN(
        n1075) );
  AOI21D0BWP12T U1777 ( .A1(n1076), .A2(n1225), .B(n1075), .ZN(n1077) );
  ND4D1BWP12T U1778 ( .A1(n1080), .A2(n1079), .A3(n1078), .A4(n1077), .ZN(
        regC_out[9]) );
  AOI22D0BWP12T U1779 ( .A1(r12[14]), .A2(n1216), .B1(n1215), .B2(pc_out[14]), 
        .ZN(n1094) );
  AOI22D0BWP12T U1780 ( .A1(r9[14]), .A2(n1211), .B1(n1217), .B2(r11[14]), 
        .ZN(n1093) );
  AOI22D0BWP12T U1781 ( .A1(r7[14]), .A2(n1200), .B1(n1199), .B2(r4[14]), .ZN(
        n1084) );
  AOI22D0BWP12T U1782 ( .A1(r2[14]), .A2(n1202), .B1(n1201), .B2(r6[14]), .ZN(
        n1083) );
  AOI22D0BWP12T U1783 ( .A1(r5[14]), .A2(n1204), .B1(n1203), .B2(r1[14]), .ZN(
        n1082) );
  AOI22D0BWP12T U1784 ( .A1(r0[14]), .A2(n1206), .B1(n1205), .B2(r3[14]), .ZN(
        n1081) );
  ND4D1BWP12T U1785 ( .A1(n1084), .A2(n1083), .A3(n1082), .A4(n1081), .ZN(
        n1091) );
  CKND0BWP12T U1786 ( .I(r8[14]), .ZN(n1086) );
  OAI22D0BWP12T U1787 ( .A1(n1136), .A2(n1086), .B1(n1085), .B2(n1099), .ZN(
        n1090) );
  CKND0BWP12T U1788 ( .I(n[2027]), .ZN(n1088) );
  OAI22D0BWP12T U1789 ( .A1(n1088), .A2(n1168), .B1(n1181), .B2(n1087), .ZN(
        n1089) );
  AOI211D0BWP12T U1790 ( .A1(n1091), .A2(n1225), .B(n1090), .C(n1089), .ZN(
        n1092) );
  ND3D1BWP12T U1791 ( .A1(n1094), .A2(n1093), .A3(n1092), .ZN(regC_out[14]) );
  AOI22D0BWP12T U1792 ( .A1(n[2034]), .A2(n1213), .B1(n1215), .B2(pc_out[7]), 
        .ZN(n1105) );
  AOI22D0BWP12T U1793 ( .A1(r9[7]), .A2(n1211), .B1(n1217), .B2(r11[7]), .ZN(
        n1104) );
  AOI22D0BWP12T U1794 ( .A1(r7[7]), .A2(n1200), .B1(n1199), .B2(r4[7]), .ZN(
        n1098) );
  AOI22D0BWP12T U1795 ( .A1(r2[7]), .A2(n1202), .B1(n1201), .B2(r6[7]), .ZN(
        n1097) );
  AOI22D0BWP12T U1796 ( .A1(r5[7]), .A2(n1204), .B1(n1203), .B2(r1[7]), .ZN(
        n1096) );
  AOI22D0BWP12T U1797 ( .A1(r0[7]), .A2(n1206), .B1(n1205), .B2(r3[7]), .ZN(
        n1095) );
  ND4D1BWP12T U1798 ( .A1(n1098), .A2(n1097), .A3(n1096), .A4(n1095), .ZN(
        n1102) );
  OAI22D0BWP12T U1799 ( .A1(n1193), .A2(n1791), .B1(n1796), .B2(n1136), .ZN(
        n1101) );
  OAI22D0BWP12T U1800 ( .A1(n1181), .A2(n1793), .B1(n1783), .B2(n1099), .ZN(
        n1100) );
  AOI211D0BWP12T U1801 ( .A1(n1102), .A2(n1225), .B(n1101), .C(n1100), .ZN(
        n1103) );
  ND3D1BWP12T U1802 ( .A1(n1105), .A2(n1104), .A3(n1103), .ZN(regC_out[7]) );
  AOI22D0BWP12T U1803 ( .A1(r8[6]), .A2(n1212), .B1(n1211), .B2(r9[6]), .ZN(
        n1116) );
  AOI22D0BWP12T U1804 ( .A1(lr[6]), .A2(n1214), .B1(n1215), .B2(pc_out[6]), 
        .ZN(n1115) );
  AOI22D0BWP12T U1805 ( .A1(r10[6]), .A2(n1218), .B1(n1217), .B2(r11[6]), .ZN(
        n1114) );
  AOI22D0BWP12T U1806 ( .A1(r7[6]), .A2(n1200), .B1(n1199), .B2(r4[6]), .ZN(
        n1109) );
  AOI22D0BWP12T U1807 ( .A1(r2[6]), .A2(n1202), .B1(n1201), .B2(r6[6]), .ZN(
        n1108) );
  AOI22D0BWP12T U1808 ( .A1(r5[6]), .A2(n1204), .B1(n1203), .B2(r1[6]), .ZN(
        n1107) );
  AOI22D0BWP12T U1809 ( .A1(r0[6]), .A2(n1206), .B1(n1205), .B2(r3[6]), .ZN(
        n1106) );
  ND4D1BWP12T U1810 ( .A1(n1109), .A2(n1108), .A3(n1107), .A4(n1106), .ZN(
        n1112) );
  OAI22D0BWP12T U1811 ( .A1(n1819), .A2(n1168), .B1(n1193), .B2(n1110), .ZN(
        n1111) );
  AOI21D0BWP12T U1812 ( .A1(n1112), .A2(n1225), .B(n1111), .ZN(n1113) );
  ND4D1BWP12T U1813 ( .A1(n1116), .A2(n1115), .A3(n1114), .A4(n1113), .ZN(
        regC_out[6]) );
  AOI22D0BWP12T U1814 ( .A1(r8[11]), .A2(n1212), .B1(n1211), .B2(r9[11]), .ZN(
        n1127) );
  AOI22D0BWP12T U1815 ( .A1(lr[11]), .A2(n1214), .B1(n1215), .B2(pc_out[11]), 
        .ZN(n1126) );
  AOI22D0BWP12T U1816 ( .A1(r10[11]), .A2(n1218), .B1(n1217), .B2(r11[11]), 
        .ZN(n1125) );
  AOI22D0BWP12T U1817 ( .A1(r7[11]), .A2(n1200), .B1(n1199), .B2(r4[11]), .ZN(
        n1120) );
  AOI22D0BWP12T U1818 ( .A1(r2[11]), .A2(n1202), .B1(n1201), .B2(r6[11]), .ZN(
        n1119) );
  AOI22D0BWP12T U1819 ( .A1(r5[11]), .A2(n1204), .B1(n1203), .B2(r1[11]), .ZN(
        n1118) );
  AOI22D0BWP12T U1820 ( .A1(r0[11]), .A2(n1206), .B1(n1205), .B2(r3[11]), .ZN(
        n1117) );
  ND4D1BWP12T U1821 ( .A1(n1120), .A2(n1119), .A3(n1118), .A4(n1117), .ZN(
        n1123) );
  OAI22D0BWP12T U1822 ( .A1(n1667), .A2(n1168), .B1(n1193), .B2(n1121), .ZN(
        n1122) );
  AOI21D0BWP12T U1823 ( .A1(n1123), .A2(n1225), .B(n1122), .ZN(n1124) );
  ND4D1BWP12T U1824 ( .A1(n1127), .A2(n1126), .A3(n1125), .A4(n1124), .ZN(
        regC_out[11]) );
  AOI22D0BWP12T U1825 ( .A1(r12[22]), .A2(n1216), .B1(n1215), .B2(pc_out[22]), 
        .ZN(n1143) );
  AOI22D0BWP12T U1826 ( .A1(r9[22]), .A2(n1211), .B1(n1218), .B2(r10[22]), 
        .ZN(n1142) );
  AOI22D0BWP12T U1827 ( .A1(r7[22]), .A2(n1200), .B1(n1199), .B2(r4[22]), .ZN(
        n1131) );
  AOI22D0BWP12T U1828 ( .A1(r2[22]), .A2(n1202), .B1(n1201), .B2(r6[22]), .ZN(
        n1130) );
  AOI22D0BWP12T U1829 ( .A1(r5[22]), .A2(n1204), .B1(n1203), .B2(r1[22]), .ZN(
        n1129) );
  AOI22D0BWP12T U1830 ( .A1(r0[22]), .A2(n1206), .B1(n1205), .B2(r3[22]), .ZN(
        n1128) );
  ND4D1BWP12T U1831 ( .A1(n1131), .A2(n1130), .A3(n1129), .A4(n1128), .ZN(
        n1140) );
  CKND0BWP12T U1832 ( .I(lr[22]), .ZN(n1134) );
  CKND0BWP12T U1833 ( .I(r11[22]), .ZN(n1133) );
  OAI22D0BWP12T U1834 ( .A1(n1181), .A2(n1134), .B1(n1133), .B2(n1132), .ZN(
        n1139) );
  CKND0BWP12T U1835 ( .I(n[2019]), .ZN(n1137) );
  CKND0BWP12T U1836 ( .I(r8[22]), .ZN(n1135) );
  OAI22D0BWP12T U1837 ( .A1(n1137), .A2(n1168), .B1(n1136), .B2(n1135), .ZN(
        n1138) );
  AOI211D0BWP12T U1838 ( .A1(n1140), .A2(n1225), .B(n1139), .C(n1138), .ZN(
        n1141) );
  ND3D1BWP12T U1839 ( .A1(n1143), .A2(n1142), .A3(n1141), .ZN(regC_out[22]) );
  AOI22D0BWP12T U1840 ( .A1(r8[17]), .A2(n1212), .B1(n1218), .B2(r10[17]), 
        .ZN(n1154) );
  AOI22D0BWP12T U1841 ( .A1(r12[17]), .A2(n1216), .B1(n1215), .B2(pc_out[17]), 
        .ZN(n1153) );
  AOI22D0BWP12T U1842 ( .A1(r9[17]), .A2(n1211), .B1(n1217), .B2(r11[17]), 
        .ZN(n1152) );
  AOI22D0BWP12T U1843 ( .A1(r7[17]), .A2(n1200), .B1(n1199), .B2(r4[17]), .ZN(
        n1147) );
  AOI22D0BWP12T U1844 ( .A1(r2[17]), .A2(n1202), .B1(n1201), .B2(r6[17]), .ZN(
        n1146) );
  AOI22D0BWP12T U1845 ( .A1(r5[17]), .A2(n1204), .B1(n1203), .B2(r1[17]), .ZN(
        n1145) );
  AOI22D0BWP12T U1846 ( .A1(r0[17]), .A2(n1206), .B1(n1205), .B2(r3[17]), .ZN(
        n1144) );
  ND4D1BWP12T U1847 ( .A1(n1147), .A2(n1146), .A3(n1145), .A4(n1144), .ZN(
        n1150) );
  CKND0BWP12T U1848 ( .I(n[2024]), .ZN(n1148) );
  INVD1BWP12T U1849 ( .I(lr[17]), .ZN(n1525) );
  OAI22D0BWP12T U1850 ( .A1(n1148), .A2(n1168), .B1(n1181), .B2(n1525), .ZN(
        n1149) );
  AOI21D0BWP12T U1851 ( .A1(n1150), .A2(n1225), .B(n1149), .ZN(n1151) );
  ND4D1BWP12T U1852 ( .A1(n1154), .A2(n1153), .A3(n1152), .A4(n1151), .ZN(
        regC_out[17]) );
  OAI22D0BWP12T U1853 ( .A1(n1696), .A2(n1157), .B1(n1156), .B2(n1155), .ZN(
        n1167) );
  OAI22D0BWP12T U1854 ( .A1(n1694), .A2(n1159), .B1(n1158), .B2(n1683), .ZN(
        n1166) );
  OAI22D0BWP12T U1855 ( .A1(n1161), .A2(n1684), .B1(n1160), .B2(n1689), .ZN(
        n1165) );
  OAI22D0BWP12T U1856 ( .A1(n1695), .A2(n1163), .B1(n1162), .B2(n1693), .ZN(
        n1164) );
  NR4D0BWP12T U1857 ( .A1(n1167), .A2(n1166), .A3(n1165), .A4(n1164), .ZN(
        n1169) );
  OAI22D0BWP12T U1858 ( .A1(n1169), .A2(readC_sel[4]), .B1(n1168), .B2(n1691), 
        .ZN(n1170) );
  AOI21D0BWP12T U1859 ( .A1(lr[10]), .A2(n1214), .B(n1170), .ZN(n1174) );
  AOI22D0BWP12T U1860 ( .A1(r9[10]), .A2(n1211), .B1(n1217), .B2(r11[10]), 
        .ZN(n1173) );
  AOI22D0BWP12T U1861 ( .A1(r8[10]), .A2(n1212), .B1(n1218), .B2(r10[10]), 
        .ZN(n1172) );
  AOI22D0BWP12T U1862 ( .A1(r12[10]), .A2(n1216), .B1(n1215), .B2(pc_out[10]), 
        .ZN(n1171) );
  ND4D1BWP12T U1863 ( .A1(n1174), .A2(n1173), .A3(n1172), .A4(n1171), .ZN(
        regC_out[10]) );
  AOI22D0BWP12T U1864 ( .A1(r7[13]), .A2(n1200), .B1(n1199), .B2(r4[13]), .ZN(
        n1178) );
  AOI22D0BWP12T U1865 ( .A1(r2[13]), .A2(n1202), .B1(n1201), .B2(r6[13]), .ZN(
        n1177) );
  AOI22D0BWP12T U1866 ( .A1(r5[13]), .A2(n1204), .B1(n1203), .B2(r1[13]), .ZN(
        n1176) );
  AOI22D0BWP12T U1867 ( .A1(r0[13]), .A2(n1206), .B1(n1205), .B2(r3[13]), .ZN(
        n1175) );
  ND4D1BWP12T U1868 ( .A1(n1178), .A2(n1177), .A3(n1176), .A4(n1175), .ZN(
        n1179) );
  MOAI22D0BWP12T U1869 ( .A1(n1181), .A2(n1180), .B1(n1179), .B2(n1225), .ZN(
        n1182) );
  AOI21D0BWP12T U1870 ( .A1(n[2028]), .A2(n1213), .B(n1182), .ZN(n1186) );
  AOI22D0BWP12T U1871 ( .A1(r10[13]), .A2(n1218), .B1(n1217), .B2(r11[13]), 
        .ZN(n1185) );
  AOI22D0BWP12T U1872 ( .A1(r8[13]), .A2(n1212), .B1(n1211), .B2(r9[13]), .ZN(
        n1184) );
  AOI22D0BWP12T U1873 ( .A1(r12[13]), .A2(n1216), .B1(n1215), .B2(pc_out[13]), 
        .ZN(n1183) );
  ND4D1BWP12T U1874 ( .A1(n1186), .A2(n1185), .A3(n1184), .A4(n1183), .ZN(
        regC_out[13]) );
  CKND0BWP12T U1875 ( .I(r12[16]), .ZN(n1192) );
  AOI22D0BWP12T U1876 ( .A1(r7[16]), .A2(n1200), .B1(n1199), .B2(r4[16]), .ZN(
        n1190) );
  AOI22D0BWP12T U1877 ( .A1(r2[16]), .A2(n1202), .B1(n1201), .B2(r6[16]), .ZN(
        n1189) );
  AOI22D0BWP12T U1878 ( .A1(r5[16]), .A2(n1204), .B1(n1203), .B2(r1[16]), .ZN(
        n1188) );
  AOI22D0BWP12T U1879 ( .A1(r0[16]), .A2(n1206), .B1(n1205), .B2(r3[16]), .ZN(
        n1187) );
  ND4D1BWP12T U1880 ( .A1(n1190), .A2(n1189), .A3(n1188), .A4(n1187), .ZN(
        n1191) );
  MOAI22D0BWP12T U1881 ( .A1(n1193), .A2(n1192), .B1(n1191), .B2(n1225), .ZN(
        n1194) );
  AOI21D0BWP12T U1882 ( .A1(lr[16]), .A2(n1214), .B(n1194), .ZN(n1198) );
  AOI22D0BWP12T U1883 ( .A1(r9[16]), .A2(n1211), .B1(n1217), .B2(r11[16]), 
        .ZN(n1197) );
  AOI22D0BWP12T U1884 ( .A1(r8[16]), .A2(n1212), .B1(n1218), .B2(r10[16]), 
        .ZN(n1196) );
  AOI22D0BWP12T U1885 ( .A1(n[2025]), .A2(n1213), .B1(n1215), .B2(pc_out[16]), 
        .ZN(n1195) );
  ND4D1BWP12T U1886 ( .A1(n1198), .A2(n1197), .A3(n1196), .A4(n1195), .ZN(
        regC_out[16]) );
  AO222D1BWP12T U1887 ( .A1(n1317), .A2(write1_in[4]), .B1(n820), .B2(
        write2_in[4]), .C1(n819), .C2(tmp1[4]), .Z(n2141) );
  AOI22D0BWP12T U1888 ( .A1(r7[21]), .A2(n1200), .B1(n1199), .B2(r4[21]), .ZN(
        n1210) );
  AOI22D0BWP12T U1889 ( .A1(r2[21]), .A2(n1202), .B1(n1201), .B2(r6[21]), .ZN(
        n1209) );
  AOI22D0BWP12T U1890 ( .A1(r5[21]), .A2(n1204), .B1(n1203), .B2(r1[21]), .ZN(
        n1208) );
  AOI22D0BWP12T U1891 ( .A1(r0[21]), .A2(n1206), .B1(n1205), .B2(r3[21]), .ZN(
        n1207) );
  ND4D1BWP12T U1892 ( .A1(n1210), .A2(n1209), .A3(n1208), .A4(n1207), .ZN(
        n1224) );
  AOI22D0BWP12T U1893 ( .A1(r8[21]), .A2(n1212), .B1(n1211), .B2(r9[21]), .ZN(
        n1222) );
  AOI22D0BWP12T U1894 ( .A1(lr[21]), .A2(n1214), .B1(n1213), .B2(n[2020]), 
        .ZN(n1221) );
  AOI22D0BWP12T U1895 ( .A1(r12[21]), .A2(n1216), .B1(n1215), .B2(pc_out[21]), 
        .ZN(n1220) );
  AOI22D0BWP12T U1896 ( .A1(r10[21]), .A2(n1218), .B1(n1217), .B2(r11[21]), 
        .ZN(n1219) );
  ND4D1BWP12T U1897 ( .A1(n1222), .A2(n1221), .A3(n1220), .A4(n1219), .ZN(
        n1223) );
  AO21D1BWP12T U1898 ( .A1(n1225), .A2(n1224), .B(n1223), .Z(regC_out[21]) );
  AO222D1BWP12T U1899 ( .A1(n1314), .A2(write1_in[13]), .B1(n1313), .B2(
        write2_in[13]), .C1(n1312), .C2(r10[13]), .Z(n2310) );
  AO222D1BWP12T U1900 ( .A1(n1308), .A2(write1_in[13]), .B1(n1307), .B2(
        write2_in[13]), .C1(n1306), .C2(r11[13]), .Z(n2278) );
  AO222D1BWP12T U1901 ( .A1(n1275), .A2(write1_in[13]), .B1(n1274), .B2(
        write2_in[13]), .C1(n1273), .C2(r2[13]), .Z(n2566) );
  AO222D1BWP12T U1902 ( .A1(n1311), .A2(write1_in[13]), .B1(n1310), .B2(
        write2_in[13]), .C1(n1309), .C2(r3[13]), .Z(n2534) );
  AO222D1BWP12T U1903 ( .A1(n1296), .A2(write1_in[13]), .B1(n1294), .B2(r4[13]), .C1(write2_in[13]), .C2(n1295), .Z(n2502) );
  AO222D1BWP12T U1904 ( .A1(n1302), .A2(write1_in[13]), .B1(n1300), .B2(r1[13]), .C1(write2_in[13]), .C2(n1301), .Z(n2598) );
  AO222D1BWP12T U1905 ( .A1(n1290), .A2(write1_in[13]), .B1(n1288), .B2(r8[13]), .C1(write2_in[13]), .C2(n1289), .Z(n2374) );
  AO222D1BWP12T U1906 ( .A1(n1293), .A2(write1_in[13]), .B1(n1291), .B2(r9[13]), .C1(write2_in[13]), .C2(n1292), .Z(n2342) );
  AO222D1BWP12T U1907 ( .A1(n1287), .A2(write1_in[13]), .B1(n1285), .B2(lr[13]), .C1(write2_in[13]), .C2(n1286), .Z(n2214) );
  AO222D1BWP12T U1908 ( .A1(n1305), .A2(write1_in[13]), .B1(n1303), .B2(r7[13]), .C1(write2_in[13]), .C2(n1304), .Z(n2406) );
  AO222D1BWP12T U1909 ( .A1(n1278), .A2(write1_in[13]), .B1(n1276), .B2(r0[13]), .C1(write2_in[13]), .C2(n1277), .Z(n2630) );
  AO222D1BWP12T U1910 ( .A1(n1299), .A2(write1_in[13]), .B1(n1297), .B2(r5[13]), .C1(write2_in[13]), .C2(n1298), .Z(n2470) );
  AO222D1BWP12T U1911 ( .A1(n1281), .A2(write1_in[13]), .B1(n1279), .B2(
        r12[13]), .C1(write2_in[13]), .C2(n1280), .Z(n2246) );
  AO222D1BWP12T U1912 ( .A1(n1284), .A2(write1_in[13]), .B1(n1282), .B2(r6[13]), .C1(write2_in[13]), .C2(n1283), .Z(n2438) );
  AO222D1BWP12T U1913 ( .A1(n1316), .A2(write1_in[13]), .B1(n421), .B2(n[2028]), .C1(write2_in[13]), .C2(n1315), .Z(spin[13]) );
  AO222D1BWP12T U1914 ( .A1(n1317), .A2(write1_in[13]), .B1(n820), .B2(
        write2_in[13]), .C1(n819), .C2(tmp1[13]), .Z(n2150) );
  AO222D1BWP12T U1915 ( .A1(n1290), .A2(write1_in[14]), .B1(n1288), .B2(r8[14]), .C1(write2_in[14]), .C2(n1289), .Z(n2375) );
  AO222D1BWP12T U1916 ( .A1(n1281), .A2(write1_in[14]), .B1(n1279), .B2(
        r12[14]), .C1(write2_in[14]), .C2(n1280), .Z(n2247) );
  AO222D1BWP12T U1917 ( .A1(n1293), .A2(write1_in[14]), .B1(n1291), .B2(r9[14]), .C1(write2_in[14]), .C2(n1292), .Z(n2343) );
  AO222D1BWP12T U1918 ( .A1(n1284), .A2(write1_in[14]), .B1(n1282), .B2(r6[14]), .C1(write2_in[14]), .C2(n1283), .Z(n2439) );
  AO222D1BWP12T U1919 ( .A1(n1287), .A2(write1_in[14]), .B1(n1285), .B2(lr[14]), .C1(write2_in[14]), .C2(n1286), .Z(n2215) );
  AO222D1BWP12T U1920 ( .A1(n1278), .A2(write1_in[14]), .B1(n1276), .B2(r0[14]), .C1(write2_in[14]), .C2(n1277), .Z(n2631) );
  AO222D1BWP12T U1921 ( .A1(n1275), .A2(write1_in[14]), .B1(n1274), .B2(
        write2_in[14]), .C1(n1273), .C2(r2[14]), .Z(n2567) );
  AO222D1BWP12T U1922 ( .A1(n1302), .A2(write1_in[14]), .B1(n1300), .B2(r1[14]), .C1(write2_in[14]), .C2(n1301), .Z(n2599) );
  AO222D1BWP12T U1923 ( .A1(n1296), .A2(write1_in[14]), .B1(n1294), .B2(r4[14]), .C1(write2_in[14]), .C2(n1295), .Z(n2503) );
  AO222D1BWP12T U1924 ( .A1(n1308), .A2(write1_in[14]), .B1(n1307), .B2(
        write2_in[14]), .C1(n1306), .C2(r11[14]), .Z(n2279) );
  AO222D1BWP12T U1925 ( .A1(n1311), .A2(write1_in[14]), .B1(n1310), .B2(
        write2_in[14]), .C1(n1309), .C2(r3[14]), .Z(n2535) );
  AO222D1BWP12T U1926 ( .A1(n1299), .A2(write1_in[14]), .B1(n1297), .B2(r5[14]), .C1(write2_in[14]), .C2(n1298), .Z(n2471) );
  AO222D1BWP12T U1927 ( .A1(n1305), .A2(write1_in[14]), .B1(n1303), .B2(r7[14]), .C1(write2_in[14]), .C2(n1304), .Z(n2407) );
  AO222D1BWP12T U1928 ( .A1(n1314), .A2(write1_in[14]), .B1(n1313), .B2(
        write2_in[14]), .C1(n1312), .C2(r10[14]), .Z(n2311) );
  AO222D1BWP12T U1929 ( .A1(n1316), .A2(write1_in[14]), .B1(n421), .B2(n[2027]), .C1(write2_in[14]), .C2(n1315), .Z(spin[14]) );
  AO222D1BWP12T U1930 ( .A1(n1317), .A2(write1_in[14]), .B1(n820), .B2(
        write2_in[14]), .C1(n819), .C2(tmp1[14]), .Z(n2151) );
  AO222D1BWP12T U1931 ( .A1(n1290), .A2(n1232), .B1(n1288), .B2(r8[16]), .C1(
        write2_in[16]), .C2(n1289), .Z(n2377) );
  AO222D1BWP12T U1932 ( .A1(n1293), .A2(n1232), .B1(n1291), .B2(r9[16]), .C1(
        write2_in[16]), .C2(n1292), .Z(n2345) );
  AO222D1BWP12T U1933 ( .A1(n1281), .A2(n1232), .B1(n1279), .B2(r12[16]), .C1(
        write2_in[16]), .C2(n1280), .Z(n2249) );
  AO222D1BWP12T U1934 ( .A1(n1302), .A2(n1232), .B1(n1300), .B2(r1[16]), .C1(
        write2_in[16]), .C2(n1301), .Z(n2601) );
  AO222D1BWP12T U1935 ( .A1(n1284), .A2(n1232), .B1(n1282), .B2(r6[16]), .C1(
        write2_in[16]), .C2(n1283), .Z(n2441) );
  AO222D1BWP12T U1936 ( .A1(n1299), .A2(n1232), .B1(n1297), .B2(r5[16]), .C1(
        write2_in[16]), .C2(n1298), .Z(n2473) );
  AO222D1BWP12T U1937 ( .A1(n1305), .A2(n1232), .B1(n1303), .B2(r7[16]), .C1(
        write2_in[16]), .C2(n1304), .Z(n2409) );
  AO222D1BWP12T U1938 ( .A1(n1278), .A2(n1232), .B1(n1276), .B2(r0[16]), .C1(
        write2_in[16]), .C2(n1277), .Z(n2633) );
  AO222D1BWP12T U1939 ( .A1(n1296), .A2(n1232), .B1(n1294), .B2(r4[16]), .C1(
        write2_in[16]), .C2(n1295), .Z(n2505) );
  AO222D1BWP12T U1940 ( .A1(n1287), .A2(n1232), .B1(n1285), .B2(lr[16]), .C1(
        write2_in[16]), .C2(n1286), .Z(n2217) );
  AO222D1BWP12T U1941 ( .A1(n1275), .A2(n1232), .B1(n1274), .B2(write2_in[16]), 
        .C1(n1273), .C2(r2[16]), .Z(n2569) );
  AO222D1BWP12T U1942 ( .A1(n1308), .A2(n1232), .B1(n1307), .B2(write2_in[16]), 
        .C1(n1306), .C2(r11[16]), .Z(n2281) );
  AO222D1BWP12T U1943 ( .A1(n1314), .A2(n1232), .B1(n1313), .B2(write2_in[16]), 
        .C1(n1312), .C2(r10[16]), .Z(n2313) );
  AO222D1BWP12T U1944 ( .A1(n1311), .A2(n1232), .B1(n1310), .B2(write2_in[16]), 
        .C1(n1309), .C2(r3[16]), .Z(n2537) );
  AO222D1BWP12T U1945 ( .A1(n1316), .A2(n1232), .B1(n421), .B2(n[2025]), .C1(
        write2_in[16]), .C2(n1315), .Z(spin[16]) );
  AO222D1BWP12T U1946 ( .A1(n1317), .A2(n1232), .B1(n820), .B2(write2_in[16]), 
        .C1(n819), .C2(tmp1[16]), .Z(n2153) );
  AO222D1BWP12T U1947 ( .A1(n1287), .A2(n1233), .B1(n1285), .B2(lr[15]), .C1(
        write2_in[15]), .C2(n1286), .Z(n2216) );
  AO222D1BWP12T U1948 ( .A1(n1296), .A2(n1233), .B1(n1294), .B2(r4[15]), .C1(
        write2_in[15]), .C2(n1295), .Z(n2504) );
  AO222D1BWP12T U1949 ( .A1(n1299), .A2(n1233), .B1(n1297), .B2(r5[15]), .C1(
        write2_in[15]), .C2(n1298), .Z(n2472) );
  AO222D1BWP12T U1950 ( .A1(n1290), .A2(n1233), .B1(n1288), .B2(r8[15]), .C1(
        write2_in[15]), .C2(n1289), .Z(n2376) );
  AO222D1BWP12T U1951 ( .A1(n1302), .A2(n1233), .B1(n1300), .B2(r1[15]), .C1(
        write2_in[15]), .C2(n1301), .Z(n2600) );
  AO222D1BWP12T U1952 ( .A1(n1305), .A2(n1233), .B1(n1303), .B2(r7[15]), .C1(
        write2_in[15]), .C2(n1304), .Z(n2408) );
  AO222D1BWP12T U1953 ( .A1(n1293), .A2(n1233), .B1(n1291), .B2(r9[15]), .C1(
        write2_in[15]), .C2(n1292), .Z(n2344) );
  AO222D1BWP12T U1954 ( .A1(n1284), .A2(n1233), .B1(n1282), .B2(r6[15]), .C1(
        write2_in[15]), .C2(n1283), .Z(n2440) );
  AO222D1BWP12T U1955 ( .A1(n1281), .A2(n1233), .B1(n1279), .B2(r12[15]), .C1(
        write2_in[15]), .C2(n1280), .Z(n2248) );
  AO222D1BWP12T U1956 ( .A1(n1278), .A2(n1233), .B1(n1276), .B2(r0[15]), .C1(
        write2_in[15]), .C2(n1277), .Z(n2632) );
  AO222D1BWP12T U1957 ( .A1(n1275), .A2(n1233), .B1(n1274), .B2(write2_in[15]), 
        .C1(n1273), .C2(r2[15]), .Z(n2568) );
  AO222D1BWP12T U1958 ( .A1(n1308), .A2(n1233), .B1(n1307), .B2(write2_in[15]), 
        .C1(n1306), .C2(r11[15]), .Z(n2280) );
  AO222D1BWP12T U1959 ( .A1(n1314), .A2(n1233), .B1(n1313), .B2(write2_in[15]), 
        .C1(n1312), .C2(r10[15]), .Z(n2312) );
  AO222D1BWP12T U1960 ( .A1(n1311), .A2(n1233), .B1(n1310), .B2(write2_in[15]), 
        .C1(n1309), .C2(r3[15]), .Z(n2536) );
  AO222D1BWP12T U1961 ( .A1(n1316), .A2(n1233), .B1(n421), .B2(n[2026]), .C1(
        write2_in[15]), .C2(n1315), .Z(spin[15]) );
  AO222D1BWP12T U1962 ( .A1(n1317), .A2(n1233), .B1(n820), .B2(write2_in[15]), 
        .C1(n819), .C2(tmp1[15]), .Z(n2152) );
  AO222D1BWP12T U1963 ( .A1(n1290), .A2(n1238), .B1(n1288), .B2(r8[18]), .C1(
        write2_in[18]), .C2(n1289), .Z(n2379) );
  AO222D1BWP12T U1964 ( .A1(n1302), .A2(n1238), .B1(n1300), .B2(r1[18]), .C1(
        write2_in[18]), .C2(n1301), .Z(n2603) );
  AO222D1BWP12T U1965 ( .A1(n1278), .A2(n1238), .B1(n1276), .B2(r0[18]), .C1(
        write2_in[18]), .C2(n1277), .Z(n2635) );
  AO222D1BWP12T U1966 ( .A1(n1293), .A2(n1238), .B1(n1291), .B2(r9[18]), .C1(
        write2_in[18]), .C2(n1292), .Z(n2347) );
  AO222D1BWP12T U1967 ( .A1(n1311), .A2(n1238), .B1(n1310), .B2(write2_in[18]), 
        .C1(n1309), .C2(r3[18]), .Z(n2539) );
  AO222D1BWP12T U1968 ( .A1(n1275), .A2(n1238), .B1(n1274), .B2(write2_in[18]), 
        .C1(n1273), .C2(r2[18]), .Z(n2571) );
  AO222D1BWP12T U1969 ( .A1(n1290), .A2(n55), .B1(n1288), .B2(r8[17]), .C1(
        write2_in[17]), .C2(n1289), .Z(n2378) );
  AO222D1BWP12T U1970 ( .A1(n1287), .A2(n55), .B1(n1285), .B2(lr[17]), .C1(
        write2_in[17]), .C2(n1286), .Z(n2218) );
  AO222D1BWP12T U1971 ( .A1(n1293), .A2(n55), .B1(n1291), .B2(r9[17]), .C1(
        write2_in[17]), .C2(n1292), .Z(n2346) );
  AO222D1BWP12T U1972 ( .A1(n1296), .A2(n55), .B1(n1294), .B2(r4[17]), .C1(
        write2_in[17]), .C2(n1295), .Z(n2506) );
  AO222D1BWP12T U1973 ( .A1(n1302), .A2(n55), .B1(n1300), .B2(r1[17]), .C1(
        write2_in[17]), .C2(n1301), .Z(n2602) );
  AO222D1BWP12T U1974 ( .A1(n1299), .A2(n55), .B1(n1297), .B2(r5[17]), .C1(
        write2_in[17]), .C2(n1298), .Z(n2474) );
  AO222D1BWP12T U1975 ( .A1(n1284), .A2(n55), .B1(n1282), .B2(r6[17]), .C1(
        write2_in[17]), .C2(n1283), .Z(n2442) );
  AO222D1BWP12T U1976 ( .A1(n1305), .A2(n55), .B1(n1303), .B2(r7[17]), .C1(
        write2_in[17]), .C2(n1304), .Z(n2410) );
  AO222D1BWP12T U1977 ( .A1(n1278), .A2(n55), .B1(n1276), .B2(r0[17]), .C1(
        write2_in[17]), .C2(n1277), .Z(n2634) );
  AO222D1BWP12T U1978 ( .A1(n1281), .A2(n55), .B1(n1279), .B2(r12[17]), .C1(
        write2_in[17]), .C2(n1280), .Z(n2250) );
  AO222D1BWP12T U1979 ( .A1(n1308), .A2(n55), .B1(n1307), .B2(write2_in[17]), 
        .C1(n1306), .C2(r11[17]), .Z(n2282) );
  AO222D1BWP12T U1980 ( .A1(n1275), .A2(n55), .B1(n1274), .B2(write2_in[17]), 
        .C1(n1273), .C2(r2[17]), .Z(n2570) );
  AO222D1BWP12T U1981 ( .A1(n1314), .A2(n55), .B1(n1313), .B2(write2_in[17]), 
        .C1(n1312), .C2(r10[17]), .Z(n2314) );
  AO222D1BWP12T U1982 ( .A1(n1311), .A2(n55), .B1(n1310), .B2(write2_in[17]), 
        .C1(n1309), .C2(r3[17]), .Z(n2538) );
  AO222D1BWP12T U1983 ( .A1(n1316), .A2(n55), .B1(n421), .B2(n[2024]), .C1(
        write2_in[17]), .C2(n1315), .Z(spin[17]) );
  AO222D1BWP12T U1984 ( .A1(n1317), .A2(n55), .B1(n820), .B2(write2_in[17]), 
        .C1(n819), .C2(tmp1[17]), .Z(n2154) );
  AO222D1BWP12T U1985 ( .A1(n1287), .A2(n1242), .B1(n1285), .B2(lr[19]), .C1(
        write2_in[19]), .C2(n1286), .Z(n2220) );
  AO222D1BWP12T U1986 ( .A1(n1299), .A2(n1242), .B1(n1297), .B2(r5[19]), .C1(
        write2_in[19]), .C2(n1298), .Z(n2476) );
  AO222D1BWP12T U1987 ( .A1(n1290), .A2(n1242), .B1(n1288), .B2(r8[19]), .C1(
        write2_in[19]), .C2(n1289), .Z(n2380) );
  AO222D1BWP12T U1988 ( .A1(n1293), .A2(n1242), .B1(n1291), .B2(r9[19]), .C1(
        write2_in[19]), .C2(n1292), .Z(n2348) );
  AO222D1BWP12T U1989 ( .A1(n1281), .A2(n1242), .B1(n1279), .B2(r12[19]), .C1(
        write2_in[19]), .C2(n1280), .Z(n2252) );
  AO222D1BWP12T U1990 ( .A1(n1302), .A2(n1242), .B1(n1300), .B2(r1[19]), .C1(
        write2_in[19]), .C2(n1301), .Z(n2604) );
  AO222D1BWP12T U1991 ( .A1(n1305), .A2(n1242), .B1(n1303), .B2(r7[19]), .C1(
        write2_in[19]), .C2(n1304), .Z(n2412) );
  AO222D1BWP12T U1992 ( .A1(n1278), .A2(n1242), .B1(n1276), .B2(r0[19]), .C1(
        write2_in[19]), .C2(n1277), .Z(n2636) );
  AO222D1BWP12T U1993 ( .A1(n1296), .A2(n1242), .B1(n1294), .B2(r4[19]), .C1(
        write2_in[19]), .C2(n1295), .Z(n2508) );
  AO222D1BWP12T U1994 ( .A1(n1284), .A2(n1242), .B1(n1282), .B2(r6[19]), .C1(
        write2_in[19]), .C2(n1283), .Z(n2444) );
  AO222D1BWP12T U1995 ( .A1(n1308), .A2(n1242), .B1(n1307), .B2(write2_in[19]), 
        .C1(n1306), .C2(r11[19]), .Z(n2284) );
  AO222D1BWP12T U1996 ( .A1(n1314), .A2(n1242), .B1(n1313), .B2(write2_in[19]), 
        .C1(n1312), .C2(r10[19]), .Z(n2316) );
  AO222D1BWP12T U1997 ( .A1(n1275), .A2(n1242), .B1(n1274), .B2(write2_in[19]), 
        .C1(n1273), .C2(r2[19]), .Z(n2572) );
  AO222D1BWP12T U1998 ( .A1(n1311), .A2(n1242), .B1(n1310), .B2(write2_in[19]), 
        .C1(n1309), .C2(r3[19]), .Z(n2540) );
  AO222D1BWP12T U1999 ( .A1(n1316), .A2(n1242), .B1(n421), .B2(n[2022]), .C1(
        write2_in[19]), .C2(n1315), .Z(spin[19]) );
  AO222D1BWP12T U2000 ( .A1(n1317), .A2(n1242), .B1(n820), .B2(write2_in[19]), 
        .C1(n819), .C2(tmp1[19]), .Z(n2156) );
  AO222D1BWP12T U2001 ( .A1(n1293), .A2(n1245), .B1(n1291), .B2(r9[20]), .C1(
        write2_in[20]), .C2(n1292), .Z(n2349) );
  AO222D1BWP12T U2002 ( .A1(n1287), .A2(n1245), .B1(n1285), .B2(lr[20]), .C1(
        write2_in[20]), .C2(n1286), .Z(n2221) );
  AO222D1BWP12T U2003 ( .A1(n1302), .A2(n1245), .B1(n1300), .B2(r1[20]), .C1(
        write2_in[20]), .C2(n1301), .Z(n2605) );
  AO222D1BWP12T U2004 ( .A1(n1299), .A2(n1245), .B1(n1297), .B2(r5[20]), .C1(
        write2_in[20]), .C2(n1298), .Z(n2477) );
  AO222D1BWP12T U2005 ( .A1(n1290), .A2(n1245), .B1(n1288), .B2(r8[20]), .C1(
        write2_in[20]), .C2(n1289), .Z(n2381) );
  AO222D1BWP12T U2006 ( .A1(n1281), .A2(n1245), .B1(n1279), .B2(r12[20]), .C1(
        write2_in[20]), .C2(n1280), .Z(n2253) );
  AO222D1BWP12T U2007 ( .A1(n1284), .A2(n1245), .B1(n1282), .B2(r6[20]), .C1(
        write2_in[20]), .C2(n1283), .Z(n2445) );
  AO222D1BWP12T U2008 ( .A1(n1296), .A2(n1245), .B1(n1294), .B2(r4[20]), .C1(
        write2_in[20]), .C2(n1295), .Z(n2509) );
  AO222D1BWP12T U2009 ( .A1(n1278), .A2(n1245), .B1(n1276), .B2(r0[20]), .C1(
        write2_in[20]), .C2(n1277), .Z(n2637) );
  AO222D1BWP12T U2010 ( .A1(n1305), .A2(n1245), .B1(n1303), .B2(r7[20]), .C1(
        write2_in[20]), .C2(n1304), .Z(n2413) );
  AO222D1BWP12T U2011 ( .A1(n1314), .A2(n1245), .B1(n1313), .B2(write2_in[20]), 
        .C1(n1312), .C2(r10[20]), .Z(n2317) );
  AO222D1BWP12T U2012 ( .A1(n1275), .A2(n1245), .B1(n1274), .B2(write2_in[20]), 
        .C1(n1273), .C2(r2[20]), .Z(n2573) );
  AO222D1BWP12T U2013 ( .A1(n1308), .A2(n1245), .B1(n1307), .B2(write2_in[20]), 
        .C1(n1306), .C2(r11[20]), .Z(n2285) );
  AO222D1BWP12T U2014 ( .A1(n1311), .A2(n1245), .B1(n1310), .B2(write2_in[20]), 
        .C1(n1309), .C2(r3[20]), .Z(n2541) );
  AO222D1BWP12T U2015 ( .A1(n1316), .A2(n1245), .B1(n421), .B2(n[2021]), .C1(
        write2_in[20]), .C2(n1315), .Z(spin[20]) );
  AO222D1BWP12T U2016 ( .A1(n1317), .A2(n1245), .B1(n820), .B2(write2_in[20]), 
        .C1(n819), .C2(tmp1[20]), .Z(n2157) );
  AO222D1BWP12T U2017 ( .A1(n1302), .A2(write1_in[21]), .B1(n1300), .B2(r1[21]), .C1(write2_in[21]), .C2(n1301), .Z(n2606) );
  AO222D1BWP12T U2018 ( .A1(n1311), .A2(write1_in[21]), .B1(n1310), .B2(
        write2_in[21]), .C1(n1309), .C2(r3[21]), .Z(n2542) );
  AO222D1BWP12T U2019 ( .A1(n1290), .A2(write1_in[21]), .B1(n1288), .B2(r8[21]), .C1(write2_in[21]), .C2(n1289), .Z(n2382) );
  AO222D1BWP12T U2020 ( .A1(n1275), .A2(write1_in[21]), .B1(n1274), .B2(
        write2_in[21]), .C1(n1273), .C2(r2[21]), .Z(n2574) );
  AO222D1BWP12T U2021 ( .A1(n1293), .A2(write1_in[21]), .B1(n1291), .B2(r9[21]), .C1(write2_in[21]), .C2(n1292), .Z(n2350) );
  AO222D1BWP12T U2022 ( .A1(n1278), .A2(write1_in[21]), .B1(n1276), .B2(r0[21]), .C1(write2_in[21]), .C2(n1277), .Z(n2638) );
  AO222D1BWP12T U2023 ( .A1(n1290), .A2(n1250), .B1(n1288), .B2(r8[22]), .C1(
        write2_in[22]), .C2(n1289), .Z(n2383) );
  AO222D1BWP12T U2024 ( .A1(n1293), .A2(n1250), .B1(n1291), .B2(r9[22]), .C1(
        write2_in[22]), .C2(n1292), .Z(n2351) );
  AO222D1BWP12T U2025 ( .A1(n1287), .A2(n1250), .B1(n1285), .B2(lr[22]), .C1(
        write2_in[22]), .C2(n1286), .Z(n2223) );
  AO222D1BWP12T U2026 ( .A1(n1305), .A2(n1250), .B1(n1303), .B2(r7[22]), .C1(
        write2_in[22]), .C2(n1304), .Z(n2415) );
  AO222D1BWP12T U2027 ( .A1(n1299), .A2(n1250), .B1(n1297), .B2(r5[22]), .C1(
        write2_in[22]), .C2(n1298), .Z(n2479) );
  AO222D1BWP12T U2028 ( .A1(n1296), .A2(n1250), .B1(n1294), .B2(r4[22]), .C1(
        write2_in[22]), .C2(n1295), .Z(n2511) );
  AO222D1BWP12T U2029 ( .A1(n1302), .A2(n1250), .B1(n1300), .B2(r1[22]), .C1(
        write2_in[22]), .C2(n1301), .Z(n2607) );
  AO222D1BWP12T U2030 ( .A1(n1278), .A2(n1250), .B1(n1276), .B2(r0[22]), .C1(
        write2_in[22]), .C2(n1277), .Z(n2639) );
  AO222D1BWP12T U2031 ( .A1(n1281), .A2(n1250), .B1(n1279), .B2(r12[22]), .C1(
        write2_in[22]), .C2(n1280), .Z(n2255) );
  AO222D1BWP12T U2032 ( .A1(n1284), .A2(n1250), .B1(n1282), .B2(r6[22]), .C1(
        write2_in[22]), .C2(n1283), .Z(n2447) );
  AO222D1BWP12T U2033 ( .A1(n1311), .A2(n1250), .B1(n1310), .B2(write2_in[22]), 
        .C1(n1309), .C2(r3[22]), .Z(n2543) );
  AO222D1BWP12T U2034 ( .A1(n1308), .A2(n1250), .B1(n1307), .B2(write2_in[22]), 
        .C1(n1306), .C2(r11[22]), .Z(n2287) );
  AO222D1BWP12T U2035 ( .A1(n1314), .A2(n1250), .B1(n1313), .B2(write2_in[22]), 
        .C1(n1312), .C2(r10[22]), .Z(n2319) );
  AO222D1BWP12T U2036 ( .A1(n1275), .A2(n1250), .B1(n1274), .B2(write2_in[22]), 
        .C1(n1273), .C2(r2[22]), .Z(n2575) );
  AO222D1BWP12T U2037 ( .A1(n1316), .A2(n1250), .B1(n421), .B2(n[2019]), .C1(
        write2_in[22]), .C2(n1315), .Z(spin[22]) );
  AO222D1BWP12T U2038 ( .A1(n1317), .A2(n1250), .B1(n820), .B2(write2_in[22]), 
        .C1(n819), .C2(tmp1[22]), .Z(n2159) );
  AO222D1BWP12T U2039 ( .A1(n1290), .A2(n1253), .B1(n1288), .B2(r8[23]), .C1(
        write2_in[23]), .C2(n1289), .Z(n2384) );
  AO222D1BWP12T U2040 ( .A1(n1293), .A2(n1253), .B1(n1291), .B2(r9[23]), .C1(
        write2_in[23]), .C2(n1292), .Z(n2352) );
  AO222D1BWP12T U2041 ( .A1(n1305), .A2(n1253), .B1(n1303), .B2(r7[23]), .C1(
        write2_in[23]), .C2(n1304), .Z(n2416) );
  AO222D1BWP12T U2042 ( .A1(n1287), .A2(n1253), .B1(n1285), .B2(lr[23]), .C1(
        write2_in[23]), .C2(n1286), .Z(n2224) );
  AO222D1BWP12T U2043 ( .A1(n1281), .A2(n1253), .B1(n1279), .B2(r12[23]), .C1(
        write2_in[23]), .C2(n1280), .Z(n2256) );
  AO222D1BWP12T U2044 ( .A1(n1302), .A2(n1253), .B1(n1300), .B2(r1[23]), .C1(
        write2_in[23]), .C2(n1301), .Z(n2608) );
  AO222D1BWP12T U2045 ( .A1(n1299), .A2(n1253), .B1(n1297), .B2(r5[23]), .C1(
        write2_in[23]), .C2(n1298), .Z(n2480) );
  AO222D1BWP12T U2046 ( .A1(n1296), .A2(n1253), .B1(n1294), .B2(r4[23]), .C1(
        write2_in[23]), .C2(n1295), .Z(n2512) );
  AO222D1BWP12T U2047 ( .A1(n1278), .A2(n1253), .B1(n1276), .B2(r0[23]), .C1(
        write2_in[23]), .C2(n1277), .Z(n2640) );
  AO222D1BWP12T U2048 ( .A1(n1284), .A2(n1253), .B1(n1282), .B2(r6[23]), .C1(
        write2_in[23]), .C2(n1283), .Z(n2448) );
  AO222D1BWP12T U2049 ( .A1(n1311), .A2(n1253), .B1(n1310), .B2(write2_in[23]), 
        .C1(n1309), .C2(r3[23]), .Z(n2544) );
  AO222D1BWP12T U2050 ( .A1(n1314), .A2(n1253), .B1(n1313), .B2(write2_in[23]), 
        .C1(n1312), .C2(r10[23]), .Z(n2320) );
  AO222D1BWP12T U2051 ( .A1(n1275), .A2(n1253), .B1(n1274), .B2(write2_in[23]), 
        .C1(n1273), .C2(r2[23]), .Z(n2576) );
  AO222D1BWP12T U2052 ( .A1(n1308), .A2(n1253), .B1(n1307), .B2(write2_in[23]), 
        .C1(n1306), .C2(r11[23]), .Z(n2288) );
  AO222D1BWP12T U2053 ( .A1(n1316), .A2(n1253), .B1(n421), .B2(n[2018]), .C1(
        write2_in[23]), .C2(n1315), .Z(spin[23]) );
  AO222D1BWP12T U2054 ( .A1(n1317), .A2(n1253), .B1(n820), .B2(write2_in[23]), 
        .C1(n819), .C2(tmp1[23]), .Z(n2160) );
  AO222D1BWP12T U2055 ( .A1(n1281), .A2(n1254), .B1(n1279), .B2(r12[24]), .C1(
        write2_in[24]), .C2(n1280), .Z(n2257) );
  AO222D1BWP12T U2056 ( .A1(n1293), .A2(n1254), .B1(n1291), .B2(r9[24]), .C1(
        write2_in[24]), .C2(n1292), .Z(n2353) );
  AO222D1BWP12T U2057 ( .A1(n1287), .A2(n1254), .B1(n1285), .B2(lr[24]), .C1(
        write2_in[24]), .C2(n1286), .Z(n2225) );
  AO222D1BWP12T U2058 ( .A1(n1290), .A2(n1254), .B1(n1288), .B2(r8[24]), .C1(
        write2_in[24]), .C2(n1289), .Z(n2385) );
  AO222D1BWP12T U2059 ( .A1(n1296), .A2(n1254), .B1(n1294), .B2(r4[24]), .C1(
        write2_in[24]), .C2(n1295), .Z(n2513) );
  AO222D1BWP12T U2060 ( .A1(n1302), .A2(n1254), .B1(n1300), .B2(r1[24]), .C1(
        write2_in[24]), .C2(n1301), .Z(n2609) );
  AO222D1BWP12T U2061 ( .A1(n1278), .A2(n1254), .B1(n1276), .B2(r0[24]), .C1(
        write2_in[24]), .C2(n1277), .Z(n2641) );
  AO222D1BWP12T U2062 ( .A1(n1299), .A2(n1254), .B1(n1297), .B2(r5[24]), .C1(
        write2_in[24]), .C2(n1298), .Z(n2481) );
  AO222D1BWP12T U2063 ( .A1(n1305), .A2(n1254), .B1(n1303), .B2(r7[24]), .C1(
        write2_in[24]), .C2(n1304), .Z(n2417) );
  AO222D1BWP12T U2064 ( .A1(n1284), .A2(n1254), .B1(n1282), .B2(r6[24]), .C1(
        write2_in[24]), .C2(n1283), .Z(n2449) );
  AO222D1BWP12T U2065 ( .A1(n1314), .A2(n1254), .B1(n1313), .B2(write2_in[24]), 
        .C1(n1312), .C2(r10[24]), .Z(n2321) );
  AO222D1BWP12T U2066 ( .A1(n1275), .A2(n1254), .B1(n1274), .B2(write2_in[24]), 
        .C1(n1273), .C2(r2[24]), .Z(n2577) );
  AO222D1BWP12T U2067 ( .A1(n1308), .A2(n1254), .B1(n1307), .B2(write2_in[24]), 
        .C1(n1306), .C2(r11[24]), .Z(n2289) );
  AO222D1BWP12T U2068 ( .A1(n1311), .A2(n1254), .B1(n1310), .B2(write2_in[24]), 
        .C1(n1309), .C2(r3[24]), .Z(n2545) );
  AO222D1BWP12T U2069 ( .A1(n1316), .A2(n1254), .B1(n421), .B2(n[2017]), .C1(
        write2_in[24]), .C2(n1315), .Z(spin[24]) );
  AO222D1BWP12T U2070 ( .A1(n1317), .A2(n1254), .B1(n820), .B2(write2_in[24]), 
        .C1(n819), .C2(tmp1[24]), .Z(n2161) );
  AO222D1BWP12T U2071 ( .A1(n1290), .A2(write1_in[25]), .B1(n1288), .B2(r8[25]), .C1(write2_in[25]), .C2(n1289), .Z(n2386) );
  AO222D1BWP12T U2072 ( .A1(n1305), .A2(write1_in[25]), .B1(n1303), .B2(r7[25]), .C1(write2_in[25]), .C2(n1304), .Z(n2418) );
  AO222D1BWP12T U2073 ( .A1(n1299), .A2(write1_in[25]), .B1(n1297), .B2(r5[25]), .C1(write2_in[25]), .C2(n1298), .Z(n2482) );
  AO222D1BWP12T U2074 ( .A1(n1293), .A2(write1_in[25]), .B1(n1291), .B2(r9[25]), .C1(write2_in[25]), .C2(n1292), .Z(n2354) );
  AO222D1BWP12T U2075 ( .A1(n1296), .A2(write1_in[25]), .B1(n1294), .B2(r4[25]), .C1(write2_in[25]), .C2(n1295), .Z(n2514) );
  AO222D1BWP12T U2076 ( .A1(n1281), .A2(write1_in[25]), .B1(n1279), .B2(
        r12[25]), .C1(write2_in[25]), .C2(n1280), .Z(n2258) );
  AO222D1BWP12T U2077 ( .A1(n1287), .A2(write1_in[25]), .B1(n1285), .B2(lr[25]), .C1(write2_in[25]), .C2(n1286), .Z(n2226) );
  AO222D1BWP12T U2078 ( .A1(n1278), .A2(write1_in[25]), .B1(n1276), .B2(r0[25]), .C1(write2_in[25]), .C2(n1277), .Z(n2642) );
  AO222D1BWP12T U2079 ( .A1(n1302), .A2(write1_in[25]), .B1(n1300), .B2(r1[25]), .C1(write2_in[25]), .C2(n1301), .Z(n2610) );
  AO222D1BWP12T U2080 ( .A1(n1284), .A2(write1_in[25]), .B1(n1282), .B2(r6[25]), .C1(write2_in[25]), .C2(n1283), .Z(n2450) );
  AO222D1BWP12T U2081 ( .A1(n1308), .A2(write1_in[25]), .B1(n1307), .B2(
        write2_in[25]), .C1(n1306), .C2(r11[25]), .Z(n2290) );
  AO222D1BWP12T U2082 ( .A1(n1275), .A2(write1_in[25]), .B1(n1274), .B2(
        write2_in[25]), .C1(n1273), .C2(r2[25]), .Z(n2578) );
  AO222D1BWP12T U2083 ( .A1(n1311), .A2(write1_in[25]), .B1(n1310), .B2(
        write2_in[25]), .C1(n1309), .C2(r3[25]), .Z(n2546) );
  AO222D1BWP12T U2084 ( .A1(n1314), .A2(write1_in[25]), .B1(n1313), .B2(
        write2_in[25]), .C1(n1312), .C2(r10[25]), .Z(n2322) );
  AO222D1BWP12T U2085 ( .A1(n1316), .A2(write1_in[25]), .B1(n421), .B2(n[2016]), .C1(write2_in[25]), .C2(n1315), .Z(spin[25]) );
  AO222D1BWP12T U2086 ( .A1(n1317), .A2(write1_in[25]), .B1(n820), .B2(
        write2_in[25]), .C1(n819), .C2(tmp1[25]), .Z(n2162) );
  XOR2D1BWP12T U2087 ( .A1(n1256), .A2(n1255), .Z(n1257) );
  AO222D1BWP12T U2088 ( .A1(n1257), .A2(n1363), .B1(n1355), .B2(next_pc_in[16]), .C1(n1361), .C2(pc_out[16]), .Z(n2185) );
  CKXOR2D0BWP12T U2089 ( .A1(n1259), .A2(n1258), .Z(n1260) );
  AO222D1BWP12T U2090 ( .A1(n1260), .A2(n1363), .B1(n1355), .B2(next_pc_in[17]), .C1(n1361), .C2(pc_out[17]), .Z(n2186) );
  AO222D1BWP12T U2091 ( .A1(n1290), .A2(n1263), .B1(n1288), .B2(r8[26]), .C1(
        write2_in[26]), .C2(n1289), .Z(n2387) );
  AO222D1BWP12T U2092 ( .A1(n1284), .A2(n1263), .B1(n1282), .B2(r6[26]), .C1(
        write2_in[26]), .C2(n1283), .Z(n2451) );
  AO222D1BWP12T U2093 ( .A1(n1287), .A2(n1263), .B1(n1285), .B2(lr[26]), .C1(
        write2_in[26]), .C2(n1286), .Z(n2227) );
  AO222D1BWP12T U2094 ( .A1(n1293), .A2(n1263), .B1(n1291), .B2(r9[26]), .C1(
        write2_in[26]), .C2(n1292), .Z(n2355) );
  AO222D1BWP12T U2095 ( .A1(n1281), .A2(n1263), .B1(n1279), .B2(r12[26]), .C1(
        write2_in[26]), .C2(n1280), .Z(n2259) );
  AO222D1BWP12T U2096 ( .A1(n1302), .A2(n1263), .B1(n1300), .B2(r1[26]), .C1(
        write2_in[26]), .C2(n1301), .Z(n2611) );
  AO222D1BWP12T U2097 ( .A1(n1278), .A2(n1263), .B1(n1276), .B2(r0[26]), .C1(
        write2_in[26]), .C2(n1277), .Z(n2643) );
  AO222D1BWP12T U2098 ( .A1(n1305), .A2(n1263), .B1(n1303), .B2(r7[26]), .C1(
        write2_in[26]), .C2(n1304), .Z(n2419) );
  AO222D1BWP12T U2099 ( .A1(n1299), .A2(n1263), .B1(n1297), .B2(r5[26]), .C1(
        write2_in[26]), .C2(n1298), .Z(n2483) );
  AO222D1BWP12T U2100 ( .A1(n1296), .A2(n1263), .B1(n1294), .B2(r4[26]), .C1(
        write2_in[26]), .C2(n1295), .Z(n2515) );
  AO222D1BWP12T U2101 ( .A1(n1311), .A2(n1263), .B1(n1310), .B2(write2_in[26]), 
        .C1(n1309), .C2(r3[26]), .Z(n2547) );
  AO222D1BWP12T U2102 ( .A1(n1275), .A2(n1263), .B1(n1274), .B2(write2_in[26]), 
        .C1(n1273), .C2(r2[26]), .Z(n2579) );
  AO222D1BWP12T U2103 ( .A1(n1308), .A2(n1263), .B1(n1307), .B2(write2_in[26]), 
        .C1(n1306), .C2(r11[26]), .Z(n2291) );
  AO222D1BWP12T U2104 ( .A1(n1314), .A2(n1263), .B1(n1313), .B2(write2_in[26]), 
        .C1(n1312), .C2(r10[26]), .Z(n2323) );
  AO222D1BWP12T U2105 ( .A1(n1316), .A2(n1263), .B1(n421), .B2(n[2015]), .C1(
        write2_in[26]), .C2(n1315), .Z(spin[26]) );
  AO222D1BWP12T U2106 ( .A1(n1317), .A2(n1263), .B1(n820), .B2(write2_in[26]), 
        .C1(n819), .C2(tmp1[26]), .Z(n2163) );
  AO222D1BWP12T U2107 ( .A1(n1293), .A2(n1264), .B1(n1291), .B2(r9[27]), .C1(
        write2_in[27]), .C2(n1292), .Z(n2356) );
  AO222D1BWP12T U2108 ( .A1(n1287), .A2(n1264), .B1(n1285), .B2(lr[27]), .C1(
        write2_in[27]), .C2(n1286), .Z(n2228) );
  AO222D1BWP12T U2109 ( .A1(n1290), .A2(n1264), .B1(n1288), .B2(r8[27]), .C1(
        write2_in[27]), .C2(n1289), .Z(n2388) );
  AO222D1BWP12T U2110 ( .A1(n1302), .A2(n1264), .B1(n1300), .B2(r1[27]), .C1(
        write2_in[27]), .C2(n1301), .Z(n2612) );
  AO222D1BWP12T U2111 ( .A1(n1278), .A2(n1264), .B1(n1276), .B2(r0[27]), .C1(
        write2_in[27]), .C2(n1277), .Z(n2644) );
  AO222D1BWP12T U2112 ( .A1(n1296), .A2(n1264), .B1(n1294), .B2(r4[27]), .C1(
        write2_in[27]), .C2(n1295), .Z(n2516) );
  AO222D1BWP12T U2113 ( .A1(n1305), .A2(n1264), .B1(n1303), .B2(r7[27]), .C1(
        write2_in[27]), .C2(n1304), .Z(n2420) );
  AO222D1BWP12T U2114 ( .A1(n1299), .A2(n1264), .B1(n1297), .B2(r5[27]), .C1(
        write2_in[27]), .C2(n1298), .Z(n2484) );
  AO222D1BWP12T U2115 ( .A1(n1281), .A2(n1264), .B1(n1279), .B2(r12[27]), .C1(
        write2_in[27]), .C2(n1280), .Z(n2260) );
  AO222D1BWP12T U2116 ( .A1(n1284), .A2(n1264), .B1(n1282), .B2(r6[27]), .C1(
        write2_in[27]), .C2(n1283), .Z(n2452) );
  AO222D1BWP12T U2117 ( .A1(n1308), .A2(n1264), .B1(n1307), .B2(write2_in[27]), 
        .C1(n1306), .C2(r11[27]), .Z(n2292) );
  AO222D1BWP12T U2118 ( .A1(n1311), .A2(n1264), .B1(n1310), .B2(write2_in[27]), 
        .C1(n1309), .C2(r3[27]), .Z(n2548) );
  AO222D1BWP12T U2119 ( .A1(n1314), .A2(n1264), .B1(n1313), .B2(write2_in[27]), 
        .C1(n1312), .C2(r10[27]), .Z(n2324) );
  AO222D1BWP12T U2120 ( .A1(n1275), .A2(n1264), .B1(n1274), .B2(write2_in[27]), 
        .C1(n1273), .C2(r2[27]), .Z(n2580) );
  AO222D1BWP12T U2121 ( .A1(n1316), .A2(n1264), .B1(n421), .B2(n[2014]), .C1(
        write2_in[27]), .C2(n1315), .Z(spin[27]) );
  AO222D1BWP12T U2122 ( .A1(n1317), .A2(n1264), .B1(n820), .B2(write2_in[27]), 
        .C1(n819), .C2(tmp1[27]), .Z(n2164) );
  AO222D1BWP12T U2123 ( .A1(n1293), .A2(n1267), .B1(n1291), .B2(r9[29]), .C1(
        write2_in[29]), .C2(n1292), .Z(n2358) );
  AO222D1BWP12T U2124 ( .A1(n1290), .A2(n1267), .B1(n1288), .B2(r8[29]), .C1(
        write2_in[29]), .C2(n1289), .Z(n2390) );
  AO222D1BWP12T U2125 ( .A1(n1287), .A2(n1267), .B1(n1285), .B2(lr[29]), .C1(
        write2_in[29]), .C2(n1286), .Z(n2230) );
  AO222D1BWP12T U2126 ( .A1(n1302), .A2(n1267), .B1(n1300), .B2(r1[29]), .C1(
        write2_in[29]), .C2(n1301), .Z(n2614) );
  AO222D1BWP12T U2127 ( .A1(n1296), .A2(n1267), .B1(n1294), .B2(r4[29]), .C1(
        write2_in[29]), .C2(n1295), .Z(n2518) );
  AO222D1BWP12T U2128 ( .A1(n1299), .A2(n1267), .B1(n1297), .B2(r5[29]), .C1(
        write2_in[29]), .C2(n1298), .Z(n2486) );
  AO222D1BWP12T U2129 ( .A1(n1278), .A2(n1267), .B1(n1276), .B2(r0[29]), .C1(
        write2_in[29]), .C2(n1277), .Z(n2646) );
  AO222D1BWP12T U2130 ( .A1(n1305), .A2(n1267), .B1(n1303), .B2(r7[29]), .C1(
        write2_in[29]), .C2(n1304), .Z(n2422) );
  AO222D1BWP12T U2131 ( .A1(n1281), .A2(n1267), .B1(n1279), .B2(r12[29]), .C1(
        write2_in[29]), .C2(n1280), .Z(n2262) );
  AO222D1BWP12T U2132 ( .A1(n1284), .A2(n1267), .B1(n1282), .B2(r6[29]), .C1(
        write2_in[29]), .C2(n1283), .Z(n2454) );
  AO222D1BWP12T U2133 ( .A1(n1311), .A2(n1267), .B1(n1310), .B2(write2_in[29]), 
        .C1(n1309), .C2(r3[29]), .Z(n2550) );
  AO222D1BWP12T U2134 ( .A1(n1275), .A2(n1267), .B1(n1274), .B2(write2_in[29]), 
        .C1(n1273), .C2(r2[29]), .Z(n2582) );
  AO222D1BWP12T U2135 ( .A1(n1308), .A2(n1267), .B1(n1307), .B2(write2_in[29]), 
        .C1(n1306), .C2(r11[29]), .Z(n2294) );
  AO222D1BWP12T U2136 ( .A1(n1314), .A2(n1267), .B1(n1313), .B2(write2_in[29]), 
        .C1(n1312), .C2(r10[29]), .Z(n2326) );
  AO222D1BWP12T U2137 ( .A1(n1316), .A2(n1267), .B1(n421), .B2(n[2012]), .C1(
        write2_in[29]), .C2(n1315), .Z(spin[29]) );
  AO222D1BWP12T U2138 ( .A1(n1317), .A2(n1267), .B1(n820), .B2(write2_in[29]), 
        .C1(n819), .C2(tmp1[29]), .Z(n2166) );
  AO222D1BWP12T U2139 ( .A1(n1287), .A2(n1268), .B1(n1285), .B2(lr[28]), .C1(
        write2_in[28]), .C2(n1286), .Z(n2229) );
  AO222D1BWP12T U2140 ( .A1(n1305), .A2(n1268), .B1(n1303), .B2(r7[28]), .C1(
        write2_in[28]), .C2(n1304), .Z(n2421) );
  AO222D1BWP12T U2141 ( .A1(n1293), .A2(n1268), .B1(n1291), .B2(r9[28]), .C1(
        write2_in[28]), .C2(n1292), .Z(n2357) );
  AO222D1BWP12T U2142 ( .A1(n1290), .A2(n1268), .B1(n1288), .B2(r8[28]), .C1(
        write2_in[28]), .C2(n1289), .Z(n2389) );
  AO222D1BWP12T U2143 ( .A1(n1275), .A2(n1268), .B1(n1274), .B2(write2_in[28]), 
        .C1(n1273), .C2(r2[28]), .Z(n2581) );
  AO222D1BWP12T U2144 ( .A1(n1311), .A2(n1268), .B1(n1310), .B2(write2_in[28]), 
        .C1(n1309), .C2(r3[28]), .Z(n2549) );
  AO222D1BWP12T U2145 ( .A1(n1308), .A2(n1268), .B1(n1307), .B2(write2_in[28]), 
        .C1(n1306), .C2(r11[28]), .Z(n2293) );
  AO222D1BWP12T U2146 ( .A1(n1314), .A2(n1268), .B1(n1313), .B2(write2_in[28]), 
        .C1(n1312), .C2(r10[28]), .Z(n2325) );
  AO222D1BWP12T U2147 ( .A1(n1316), .A2(n1268), .B1(n421), .B2(n[2013]), .C1(
        write2_in[28]), .C2(n1315), .Z(spin[28]) );
  AO222D1BWP12T U2148 ( .A1(n1317), .A2(n1268), .B1(n820), .B2(write2_in[28]), 
        .C1(n819), .C2(tmp1[28]), .Z(n2165) );
  BUFFD6BWP12T U2149 ( .I(write1_in[30]), .Z(n1331) );
  AO222D1BWP12T U2150 ( .A1(n1290), .A2(n1331), .B1(n1288), .B2(r8[30]), .C1(
        write2_in[30]), .C2(n1289), .Z(n2391) );
  AO222D1BWP12T U2151 ( .A1(n1281), .A2(n1331), .B1(n1279), .B2(r12[30]), .C1(
        write2_in[30]), .C2(n1280), .Z(n2263) );
  AO222D1BWP12T U2152 ( .A1(n1293), .A2(n1331), .B1(n1291), .B2(r9[30]), .C1(
        write2_in[30]), .C2(n1292), .Z(n2359) );
  AO222D1BWP12T U2153 ( .A1(n1287), .A2(n1331), .B1(n1285), .B2(lr[30]), .C1(
        write2_in[30]), .C2(n1286), .Z(n2231) );
  AO222D1BWP12T U2154 ( .A1(n1296), .A2(n1331), .B1(n1294), .B2(r4[30]), .C1(
        write2_in[30]), .C2(n1295), .Z(n2519) );
  AO222D1BWP12T U2155 ( .A1(n1302), .A2(n1331), .B1(n1300), .B2(r1[30]), .C1(
        write2_in[30]), .C2(n1301), .Z(n2615) );
  AO222D1BWP12T U2156 ( .A1(n1278), .A2(n1331), .B1(n1276), .B2(r0[30]), .C1(
        write2_in[30]), .C2(n1277), .Z(n2647) );
  AO222D1BWP12T U2157 ( .A1(n1299), .A2(n1331), .B1(n1297), .B2(r5[30]), .C1(
        write2_in[30]), .C2(n1298), .Z(n2487) );
  AO222D1BWP12T U2158 ( .A1(n1305), .A2(n1331), .B1(n1303), .B2(r7[30]), .C1(
        write2_in[30]), .C2(n1304), .Z(n2423) );
  AO222D1BWP12T U2159 ( .A1(n1284), .A2(n1331), .B1(n1282), .B2(r6[30]), .C1(
        write2_in[30]), .C2(n1283), .Z(n2455) );
  AO222D1BWP12T U2160 ( .A1(n1308), .A2(n1331), .B1(n1307), .B2(write2_in[30]), 
        .C1(n1306), .C2(r11[30]), .Z(n2295) );
  AO222D1BWP12T U2161 ( .A1(n1275), .A2(n1331), .B1(n1274), .B2(write2_in[30]), 
        .C1(n1273), .C2(r2[30]), .Z(n2583) );
  AO222D1BWP12T U2162 ( .A1(n1314), .A2(n1331), .B1(n1313), .B2(write2_in[30]), 
        .C1(n1312), .C2(r10[30]), .Z(n2327) );
  AO222D1BWP12T U2163 ( .A1(n1311), .A2(n1331), .B1(n1310), .B2(write2_in[30]), 
        .C1(n1309), .C2(r3[30]), .Z(n2551) );
  AO222D1BWP12T U2164 ( .A1(n1316), .A2(n1331), .B1(n421), .B2(n[2011]), .C1(
        write2_in[30]), .C2(n1315), .Z(spin[30]) );
  AO222D1BWP12T U2165 ( .A1(n1317), .A2(n1331), .B1(n820), .B2(write2_in[30]), 
        .C1(n819), .C2(tmp1[30]), .Z(n2167) );
  BUFFD6BWP12T U2166 ( .I(write1_in[31]), .Z(n1327) );
  AO222D1BWP12T U2167 ( .A1(n1327), .A2(n1275), .B1(write2_in[31]), .B2(n1274), 
        .C1(n1273), .C2(r2[31]), .Z(n2584) );
  AO222D1BWP12T U2168 ( .A1(n1327), .A2(n1278), .B1(write2_in[31]), .B2(n1277), 
        .C1(r0[31]), .C2(n1276), .Z(n2648) );
  AO222D1BWP12T U2169 ( .A1(n1327), .A2(n1281), .B1(write2_in[31]), .B2(n1280), 
        .C1(r12[31]), .C2(n1279), .Z(n2264) );
  AO222D1BWP12T U2170 ( .A1(n1327), .A2(n1284), .B1(write2_in[31]), .B2(n1283), 
        .C1(r6[31]), .C2(n1282), .Z(n2456) );
  AO222D1BWP12T U2171 ( .A1(n1327), .A2(n1287), .B1(write2_in[31]), .B2(n1286), 
        .C1(lr[31]), .C2(n1285), .Z(n2232) );
  AO222D1BWP12T U2172 ( .A1(n1327), .A2(n1290), .B1(write2_in[31]), .B2(n1289), 
        .C1(r8[31]), .C2(n1288), .Z(n2392) );
  AO222D1BWP12T U2173 ( .A1(n1327), .A2(n1293), .B1(write2_in[31]), .B2(n1292), 
        .C1(r9[31]), .C2(n1291), .Z(n2360) );
  AO222D1BWP12T U2174 ( .A1(n1327), .A2(n1296), .B1(write2_in[31]), .B2(n1295), 
        .C1(r4[31]), .C2(n1294), .Z(n2520) );
  AO222D1BWP12T U2175 ( .A1(n1327), .A2(n1299), .B1(write2_in[31]), .B2(n1298), 
        .C1(r5[31]), .C2(n1297), .Z(n2488) );
  AO222D1BWP12T U2176 ( .A1(n1327), .A2(n1302), .B1(write2_in[31]), .B2(n1301), 
        .C1(r1[31]), .C2(n1300), .Z(n2616) );
  AO222D1BWP12T U2177 ( .A1(n1327), .A2(n1305), .B1(write2_in[31]), .B2(n1304), 
        .C1(r7[31]), .C2(n1303), .Z(n2424) );
  AO222D1BWP12T U2178 ( .A1(n1327), .A2(n1308), .B1(write2_in[31]), .B2(n1307), 
        .C1(n1306), .C2(r11[31]), .Z(n2296) );
  AO222D1BWP12T U2179 ( .A1(n1327), .A2(n1311), .B1(write2_in[31]), .B2(n1310), 
        .C1(n1309), .C2(r3[31]), .Z(n2552) );
  AO222D1BWP12T U2180 ( .A1(n1327), .A2(n1314), .B1(write2_in[31]), .B2(n1313), 
        .C1(n1312), .C2(r10[31]), .Z(n2328) );
  AO222D1BWP12T U2181 ( .A1(n1327), .A2(n1316), .B1(write2_in[31]), .B2(n1315), 
        .C1(n[2010]), .C2(n421), .Z(spin[31]) );
  AO222D1BWP12T U2182 ( .A1(n1327), .A2(n1317), .B1(write2_in[31]), .B2(n820), 
        .C1(n819), .C2(tmp1[31]), .Z(n2168) );
  AO222D1BWP12T U2183 ( .A1(n1322), .A2(n1363), .B1(n1355), .B2(next_pc_in[27]), .C1(n1361), .C2(pc_out[27]), .Z(n2196) );
  OR2D4BWP12T U2184 ( .A1(n1324), .A2(n1323), .Z(n1343) );
  XOR2D1BWP12T U2185 ( .A1(n1343), .A2(n1342), .Z(n1325) );
  AO222D1BWP12T U2186 ( .A1(n1325), .A2(n1363), .B1(n1355), .B2(next_pc_in[24]), .C1(n1361), .C2(pc_out[24]), .Z(n2193) );
  CKND2D2BWP12T U2187 ( .A1(n1349), .A2(n1346), .ZN(n1352) );
  AN2XD0BWP12T U2188 ( .A1(write2_in[31]), .A2(n1328), .Z(n1326) );
  AN2XD0BWP12T U2189 ( .A1(write2_in[30]), .A2(n1328), .Z(n1329) );
  INVD2BWP12T U2190 ( .I(n1336), .ZN(n1332) );
  TPND2D2BWP12T U2191 ( .A1(n1332), .A2(n1363), .ZN(n1348) );
  INVD1BWP12T U2192 ( .I(n1348), .ZN(n1333) );
  ND2D1BWP12T U2193 ( .A1(n1338), .A2(n1333), .ZN(n1341) );
  ND2D1BWP12T U2194 ( .A1(n1335), .A2(n1352), .ZN(n1340) );
  ND2D1BWP12T U2195 ( .A1(n1336), .A2(n1363), .ZN(n1351) );
  OA21D1BWP12T U2196 ( .A1(n1338), .A2(n1351), .B(n1337), .Z(n1339) );
  OAI211D1BWP12T U2197 ( .A1(n1352), .A2(n1341), .B(n1340), .C(n1339), .ZN(
        n2200) );
  XOR2D1BWP12T U2198 ( .A1(n1358), .A2(n1357), .Z(n1344) );
  AO222D1BWP12T U2199 ( .A1(n1344), .A2(n1363), .B1(n1362), .B2(next_pc_in[25]), .C1(n1361), .C2(pc_out[25]), .Z(n2194) );
  AOI22D1BWP12T U2200 ( .A1(next_pc_in[30]), .A2(n1355), .B1(n1361), .B2(
        pc_out[30]), .ZN(n1345) );
  RCIAO21D0BWP12T U2201 ( .A1(n1349), .A2(n1348), .B(n1347), .ZN(n1350) );
  OAI21D1BWP12T U2202 ( .A1(n1352), .A2(n1351), .B(n1350), .ZN(n2199) );
  XOR2D2BWP12T U2203 ( .A1(n1354), .A2(n1353), .Z(n1356) );
  AO222D1BWP12T U2204 ( .A1(n1356), .A2(n1363), .B1(n1355), .B2(next_pc_in[28]), .C1(n1361), .C2(pc_out[28]), .Z(n2197) );
  XOR2D2BWP12T U2205 ( .A1(n1360), .A2(n1359), .Z(n1364) );
  AO222D1BWP12T U2206 ( .A1(n1364), .A2(n1363), .B1(n1362), .B2(next_pc_in[26]), .C1(n1361), .C2(pc_out[26]), .Z(n2195) );
  AOI22D1BWP12T U2207 ( .A1(r1[26]), .A2(n183), .B1(n1992), .B2(r12[26]), .ZN(
        n1368) );
  AOI22D1BWP12T U2208 ( .A1(r3[26]), .A2(n185), .B1(n1993), .B2(lr[26]), .ZN(
        n1367) );
  AOI22D1BWP12T U2209 ( .A1(r8[26]), .A2(n187), .B1(n1994), .B2(n[2015]), .ZN(
        n1366) );
  AOI22D1BWP12T U2210 ( .A1(pc_out[26]), .A2(n188), .B1(n1995), .B2(r6[26]), 
        .ZN(n1365) );
  AN4XD1BWP12T U2211 ( .A1(n1368), .A2(n1367), .A3(n1366), .A4(n1365), .Z(
        n1375) );
  AOI22D1BWP12T U2212 ( .A1(tmp1[26]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[26]), .ZN(n1371) );
  AOI22D1BWP12T U2213 ( .A1(r9[26]), .A2(n201), .B1(n2001), .B2(r4[26]), .ZN(
        n1370) );
  AOI22D1BWP12T U2214 ( .A1(r11[26]), .A2(n1470), .B1(n205), .B2(r0[26]), .ZN(
        n1369) );
  AN3XD1BWP12T U2215 ( .A1(n1371), .A2(n1370), .A3(n1369), .Z(n1374) );
  AOI22D1BWP12T U2216 ( .A1(r5[26]), .A2(n210), .B1(n1988), .B2(r10[26]), .ZN(
        n1373) );
  AOI22D1BWP12T U2217 ( .A1(r7[26]), .A2(n215), .B1(n1989), .B2(r2[26]), .ZN(
        n1372) );
  ND4D1BWP12T U2218 ( .A1(n1375), .A2(n1374), .A3(n1373), .A4(n1372), .ZN(
        regB_out[26]) );
  AOI22D1BWP12T U2219 ( .A1(r1[28]), .A2(n183), .B1(n1992), .B2(r12[28]), .ZN(
        n1379) );
  AOI22D1BWP12T U2220 ( .A1(r3[28]), .A2(n185), .B1(n1993), .B2(lr[28]), .ZN(
        n1378) );
  AOI22D1BWP12T U2221 ( .A1(r8[28]), .A2(n187), .B1(n1994), .B2(n[2013]), .ZN(
        n1377) );
  AOI22D1BWP12T U2222 ( .A1(pc_out[28]), .A2(n188), .B1(n1995), .B2(r6[28]), 
        .ZN(n1376) );
  AN4XD1BWP12T U2223 ( .A1(n1379), .A2(n1378), .A3(n1377), .A4(n1376), .Z(
        n1386) );
  AOI22D1BWP12T U2224 ( .A1(tmp1[28]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[28]), .ZN(n1382) );
  AOI22D1BWP12T U2225 ( .A1(r9[28]), .A2(n201), .B1(n2001), .B2(r4[28]), .ZN(
        n1381) );
  AOI22D1BWP12T U2226 ( .A1(r11[28]), .A2(n1470), .B1(n205), .B2(r0[28]), .ZN(
        n1380) );
  AN3XD1BWP12T U2227 ( .A1(n1382), .A2(n1381), .A3(n1380), .Z(n1385) );
  AOI22D1BWP12T U2228 ( .A1(r5[28]), .A2(n210), .B1(n1988), .B2(r10[28]), .ZN(
        n1384) );
  AOI22D1BWP12T U2229 ( .A1(r7[28]), .A2(n215), .B1(n1989), .B2(r2[28]), .ZN(
        n1383) );
  ND4D1BWP12T U2230 ( .A1(n1386), .A2(n1385), .A3(n1384), .A4(n1383), .ZN(
        regB_out[28]) );
  AOI22D1BWP12T U2231 ( .A1(r1[29]), .A2(n183), .B1(n1992), .B2(r12[29]), .ZN(
        n1390) );
  AOI22D1BWP12T U2232 ( .A1(r3[29]), .A2(n185), .B1(n1993), .B2(lr[29]), .ZN(
        n1389) );
  AOI22D1BWP12T U2233 ( .A1(r8[29]), .A2(n187), .B1(n1994), .B2(n[2012]), .ZN(
        n1388) );
  AOI22D1BWP12T U2234 ( .A1(pc_out[29]), .A2(n188), .B1(n1995), .B2(r6[29]), 
        .ZN(n1387) );
  AN4XD1BWP12T U2235 ( .A1(n1390), .A2(n1389), .A3(n1388), .A4(n1387), .Z(
        n1397) );
  AOI22D1BWP12T U2236 ( .A1(tmp1[29]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[29]), .ZN(n1393) );
  AOI22D1BWP12T U2237 ( .A1(r9[29]), .A2(n201), .B1(n2001), .B2(r4[29]), .ZN(
        n1392) );
  AOI22D1BWP12T U2238 ( .A1(r11[29]), .A2(n1470), .B1(n205), .B2(r0[29]), .ZN(
        n1391) );
  AN3XD1BWP12T U2239 ( .A1(n1393), .A2(n1392), .A3(n1391), .Z(n1396) );
  AOI22D1BWP12T U2240 ( .A1(r5[29]), .A2(n210), .B1(n1988), .B2(r10[29]), .ZN(
        n1395) );
  AOI22D1BWP12T U2241 ( .A1(r7[29]), .A2(n215), .B1(n1989), .B2(r2[29]), .ZN(
        n1394) );
  ND4D1BWP12T U2242 ( .A1(n1397), .A2(n1396), .A3(n1395), .A4(n1394), .ZN(
        regB_out[29]) );
  AOI22D1BWP12T U2243 ( .A1(tmp1[30]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[30]), .ZN(n1400) );
  AOI22D1BWP12T U2244 ( .A1(r9[30]), .A2(n201), .B1(n2001), .B2(r4[30]), .ZN(
        n1399) );
  AOI22D1BWP12T U2245 ( .A1(r11[30]), .A2(n1470), .B1(n205), .B2(r0[30]), .ZN(
        n1398) );
  AOI22D1BWP12T U2246 ( .A1(r1[31]), .A2(n183), .B1(n1992), .B2(r12[31]), .ZN(
        n1404) );
  AOI22D1BWP12T U2247 ( .A1(r3[31]), .A2(n185), .B1(n1993), .B2(lr[31]), .ZN(
        n1403) );
  AOI22D1BWP12T U2248 ( .A1(r8[31]), .A2(n187), .B1(n1994), .B2(n[2010]), .ZN(
        n1402) );
  AOI22D1BWP12T U2249 ( .A1(pc_out[31]), .A2(n188), .B1(n1995), .B2(r6[31]), 
        .ZN(n1401) );
  AN4XD1BWP12T U2250 ( .A1(n1404), .A2(n1403), .A3(n1402), .A4(n1401), .Z(
        n1411) );
  AOI22D1BWP12T U2251 ( .A1(tmp1[31]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[31]), .ZN(n1407) );
  AOI22D0BWP12T U2252 ( .A1(r9[31]), .A2(n201), .B1(n2001), .B2(r4[31]), .ZN(
        n1406) );
  AOI22D1BWP12T U2253 ( .A1(r11[31]), .A2(n1470), .B1(n205), .B2(r0[31]), .ZN(
        n1405) );
  AN3XD1BWP12T U2254 ( .A1(n1407), .A2(n1406), .A3(n1405), .Z(n1410) );
  AOI22D1BWP12T U2255 ( .A1(r5[31]), .A2(n210), .B1(n1988), .B2(r10[31]), .ZN(
        n1409) );
  AOI22D1BWP12T U2256 ( .A1(r7[31]), .A2(n215), .B1(n1989), .B2(r2[31]), .ZN(
        n1408) );
  ND4D1BWP12T U2257 ( .A1(n1411), .A2(n1410), .A3(n1409), .A4(n1408), .ZN(
        regB_out[31]) );
  INVD1BWP12T U2258 ( .I(r4[29]), .ZN(n1414) );
  AOI22D1BWP12T U2259 ( .A1(n150), .A2(r12[29]), .B1(n1486), .B2(tmp1[29]), 
        .ZN(n1413) );
  AOI22D1BWP12T U2260 ( .A1(r2[29]), .A2(n155), .B1(n1555), .B2(r1[29]), .ZN(
        n1412) );
  OA211D1BWP12T U2261 ( .A1(n1414), .A2(n1458), .B(n1413), .C(n1412), .Z(n1422) );
  AOI22D1BWP12T U2262 ( .A1(r9[29]), .A2(n1591), .B1(n1590), .B2(r6[29]), .ZN(
        n1418) );
  AOI22D1BWP12T U2263 ( .A1(r8[29]), .A2(n1593), .B1(n1592), .B2(n[2012]), 
        .ZN(n1417) );
  AOI22D1BWP12T U2264 ( .A1(r5[29]), .A2(n1594), .B1(n171), .B2(r3[29]), .ZN(
        n1416) );
  AOI22D1BWP12T U2265 ( .A1(r7[29]), .A2(n1596), .B1(n1595), .B2(r0[29]), .ZN(
        n1415) );
  AN4XD1BWP12T U2266 ( .A1(n1418), .A2(n1417), .A3(n1416), .A4(n1415), .Z(
        n1421) );
  AOI22D1BWP12T U2267 ( .A1(pc_out[29]), .A2(n141), .B1(n1559), .B2(r11[29]), 
        .ZN(n1420) );
  AOI22D1BWP12T U2268 ( .A1(lr[29]), .A2(n1561), .B1(n1560), .B2(r10[29]), 
        .ZN(n1419) );
  ND4D1BWP12T U2269 ( .A1(n1422), .A2(n1421), .A3(n1420), .A4(n1419), .ZN(
        regA_out[29]) );
  INVD1BWP12T U2270 ( .I(r4[31]), .ZN(n1425) );
  AOI22D1BWP12T U2271 ( .A1(n150), .A2(r12[31]), .B1(n1486), .B2(tmp1[31]), 
        .ZN(n1424) );
  AOI22D1BWP12T U2272 ( .A1(r2[31]), .A2(n155), .B1(n1555), .B2(r1[31]), .ZN(
        n1423) );
  OA211D1BWP12T U2273 ( .A1(n1425), .A2(n1458), .B(n1424), .C(n1423), .Z(n1433) );
  AOI22D1BWP12T U2274 ( .A1(r9[31]), .A2(n1591), .B1(n1590), .B2(r6[31]), .ZN(
        n1429) );
  AOI22D1BWP12T U2275 ( .A1(r8[31]), .A2(n1593), .B1(n1592), .B2(n[2010]), 
        .ZN(n1428) );
  AOI22D1BWP12T U2276 ( .A1(r5[31]), .A2(n1594), .B1(n171), .B2(r3[31]), .ZN(
        n1427) );
  AOI22D1BWP12T U2277 ( .A1(r7[31]), .A2(n1596), .B1(n1595), .B2(r0[31]), .ZN(
        n1426) );
  AN4XD1BWP12T U2278 ( .A1(n1429), .A2(n1428), .A3(n1427), .A4(n1426), .Z(
        n1432) );
  AOI22D1BWP12T U2279 ( .A1(pc_out[31]), .A2(n141), .B1(n1559), .B2(r11[31]), 
        .ZN(n1431) );
  AOI22D1BWP12T U2280 ( .A1(lr[31]), .A2(n1561), .B1(n1560), .B2(r10[31]), 
        .ZN(n1430) );
  ND4D1BWP12T U2281 ( .A1(n1433), .A2(n1432), .A3(n1431), .A4(n1430), .ZN(
        regA_out[31]) );
  INVD1BWP12T U2282 ( .I(r4[25]), .ZN(n1436) );
  AOI22D1BWP12T U2283 ( .A1(n150), .A2(r12[25]), .B1(n1486), .B2(tmp1[25]), 
        .ZN(n1435) );
  AOI22D1BWP12T U2284 ( .A1(r2[25]), .A2(n155), .B1(n1555), .B2(r1[25]), .ZN(
        n1434) );
  OA211D1BWP12T U2285 ( .A1(n1436), .A2(n1458), .B(n1435), .C(n1434), .Z(n1444) );
  AOI22D1BWP12T U2286 ( .A1(r9[25]), .A2(n1591), .B1(n1590), .B2(r6[25]), .ZN(
        n1440) );
  AOI22D1BWP12T U2287 ( .A1(r8[25]), .A2(n1593), .B1(n1592), .B2(n[2016]), 
        .ZN(n1439) );
  AOI22D1BWP12T U2288 ( .A1(r5[25]), .A2(n1594), .B1(n171), .B2(r3[25]), .ZN(
        n1438) );
  AOI22D1BWP12T U2289 ( .A1(r7[25]), .A2(n1596), .B1(n1595), .B2(r0[25]), .ZN(
        n1437) );
  AN4XD1BWP12T U2290 ( .A1(n1440), .A2(n1439), .A3(n1438), .A4(n1437), .Z(
        n1443) );
  AOI22D1BWP12T U2291 ( .A1(pc_out[25]), .A2(n141), .B1(n1559), .B2(r11[25]), 
        .ZN(n1442) );
  AOI22D1BWP12T U2292 ( .A1(lr[25]), .A2(n1561), .B1(n1560), .B2(r10[25]), 
        .ZN(n1441) );
  ND4D1BWP12T U2293 ( .A1(n1444), .A2(n1443), .A3(n1442), .A4(n1441), .ZN(
        regA_out[25]) );
  INVD1BWP12T U2294 ( .I(r4[24]), .ZN(n1447) );
  AOI22D1BWP12T U2295 ( .A1(n150), .A2(r12[24]), .B1(n1486), .B2(tmp1[24]), 
        .ZN(n1446) );
  AOI22D1BWP12T U2296 ( .A1(r2[24]), .A2(n155), .B1(n1555), .B2(r1[24]), .ZN(
        n1445) );
  OA211D1BWP12T U2297 ( .A1(n1447), .A2(n1458), .B(n1446), .C(n1445), .Z(n1455) );
  AOI22D1BWP12T U2298 ( .A1(r9[24]), .A2(n1591), .B1(n1590), .B2(r6[24]), .ZN(
        n1451) );
  AOI22D1BWP12T U2299 ( .A1(r8[24]), .A2(n1593), .B1(n1592), .B2(n[2017]), 
        .ZN(n1450) );
  AOI22D1BWP12T U2300 ( .A1(r5[24]), .A2(n1594), .B1(n171), .B2(r3[24]), .ZN(
        n1449) );
  AOI22D1BWP12T U2301 ( .A1(r7[24]), .A2(n1596), .B1(n1595), .B2(r0[24]), .ZN(
        n1448) );
  AN4XD1BWP12T U2302 ( .A1(n1451), .A2(n1450), .A3(n1449), .A4(n1448), .Z(
        n1454) );
  AOI22D1BWP12T U2303 ( .A1(pc_out[24]), .A2(n141), .B1(n1559), .B2(r11[24]), 
        .ZN(n1453) );
  AOI22D1BWP12T U2304 ( .A1(lr[24]), .A2(n1561), .B1(n1560), .B2(r10[24]), 
        .ZN(n1452) );
  ND4D1BWP12T U2305 ( .A1(n1455), .A2(n1454), .A3(n1453), .A4(n1452), .ZN(
        regA_out[24]) );
  INVD1BWP12T U2306 ( .I(r4[27]), .ZN(n1459) );
  AOI22D1BWP12T U2307 ( .A1(n150), .A2(r12[27]), .B1(n1486), .B2(tmp1[27]), 
        .ZN(n1457) );
  AOI22D1BWP12T U2308 ( .A1(r2[27]), .A2(n155), .B1(n1555), .B2(r1[27]), .ZN(
        n1456) );
  OA211D1BWP12T U2309 ( .A1(n1459), .A2(n1458), .B(n1457), .C(n1456), .Z(n1467) );
  AOI22D1BWP12T U2310 ( .A1(r9[27]), .A2(n1591), .B1(n1590), .B2(r6[27]), .ZN(
        n1463) );
  AOI22D1BWP12T U2311 ( .A1(r8[27]), .A2(n1593), .B1(n1592), .B2(n[2014]), 
        .ZN(n1462) );
  AOI22D1BWP12T U2312 ( .A1(r5[27]), .A2(n1594), .B1(n171), .B2(r3[27]), .ZN(
        n1461) );
  AOI22D1BWP12T U2313 ( .A1(r7[27]), .A2(n1596), .B1(n1595), .B2(r0[27]), .ZN(
        n1460) );
  AN4XD1BWP12T U2314 ( .A1(n1463), .A2(n1462), .A3(n1461), .A4(n1460), .Z(
        n1466) );
  AOI22D1BWP12T U2315 ( .A1(pc_out[27]), .A2(n141), .B1(n1559), .B2(r11[27]), 
        .ZN(n1465) );
  AOI22D1BWP12T U2316 ( .A1(lr[27]), .A2(n1561), .B1(n1560), .B2(r10[27]), 
        .ZN(n1464) );
  ND4D1BWP12T U2317 ( .A1(n1467), .A2(n1466), .A3(n1465), .A4(n1464), .ZN(
        regA_out[27]) );
  AOI22D1BWP12T U2318 ( .A1(tmp1[20]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[20]), .ZN(n1475) );
  AOI22D1BWP12T U2319 ( .A1(r5[20]), .A2(n210), .B1(n1988), .B2(r10[20]), .ZN(
        n1469) );
  AOI22D1BWP12T U2320 ( .A1(r7[20]), .A2(n215), .B1(n1989), .B2(r2[20]), .ZN(
        n1468) );
  ND2D1BWP12T U2321 ( .A1(n1469), .A2(n1468), .ZN(n1474) );
  AOI22D1BWP12T U2322 ( .A1(r9[20]), .A2(n201), .B1(n2001), .B2(r4[20]), .ZN(
        n1472) );
  AOI22D1BWP12T U2323 ( .A1(r11[20]), .A2(n1470), .B1(n205), .B2(r0[20]), .ZN(
        n1471) );
  ND2D1BWP12T U2324 ( .A1(n1472), .A2(n1471), .ZN(n1473) );
  INR3D0BWP12T U2325 ( .A1(n1475), .B1(n1474), .B2(n1473), .ZN(n1481) );
  AOI22D1BWP12T U2326 ( .A1(r1[20]), .A2(n183), .B1(n1992), .B2(r12[20]), .ZN(
        n1479) );
  AOI22D1BWP12T U2327 ( .A1(r3[20]), .A2(n185), .B1(n1993), .B2(lr[20]), .ZN(
        n1478) );
  AOI22D1BWP12T U2328 ( .A1(r8[20]), .A2(n187), .B1(n1994), .B2(n[2021]), .ZN(
        n1477) );
  AOI22D1BWP12T U2329 ( .A1(pc_out[20]), .A2(n188), .B1(n1995), .B2(r6[20]), 
        .ZN(n1476) );
  AN4XD1BWP12T U2330 ( .A1(n1479), .A2(n1478), .A3(n1477), .A4(n1476), .Z(
        n1480) );
  ND2D1BWP12T U2331 ( .A1(n1481), .A2(n1480), .ZN(regB_out[20]) );
  INVD1BWP12T U2332 ( .I(pc_out[19]), .ZN(n1483) );
  INVD1BWP12T U2333 ( .I(r11[19]), .ZN(n1482) );
  INVD1BWP12T U2334 ( .I(r10[19]), .ZN(n1484) );
  OAI22D1BWP12T U2335 ( .A1(n1485), .A2(n1953), .B1(n1952), .B2(n1484), .ZN(
        n1491) );
  AOI22D1BWP12T U2336 ( .A1(n150), .A2(r12[19]), .B1(n1486), .B2(tmp1[19]), 
        .ZN(n1487) );
  IOA21D1BWP12T U2337 ( .A1(n1957), .A2(r4[19]), .B(n1487), .ZN(n1490) );
  INVD1BWP12T U2338 ( .I(r2[19]), .ZN(n1489) );
  INVD1BWP12T U2339 ( .I(r1[19]), .ZN(n1488) );
  AOI22D1BWP12T U2340 ( .A1(r9[19]), .A2(n1591), .B1(n1590), .B2(r6[19]), .ZN(
        n1495) );
  AOI22D1BWP12T U2341 ( .A1(r8[19]), .A2(n1593), .B1(n1592), .B2(n[2022]), 
        .ZN(n1494) );
  AOI22D1BWP12T U2342 ( .A1(r5[19]), .A2(n1594), .B1(n171), .B2(r3[19]), .ZN(
        n1493) );
  AOI22D1BWP12T U2343 ( .A1(r7[19]), .A2(n1596), .B1(n1595), .B2(r0[19]), .ZN(
        n1492) );
  AN4XD1BWP12T U2344 ( .A1(n1495), .A2(n1494), .A3(n1493), .A4(n1492), .Z(
        n1496) );
  ND2D1BWP12T U2345 ( .A1(n1497), .A2(n1496), .ZN(regA_out[19]) );
  AOI22D1BWP12T U2346 ( .A1(r9[18]), .A2(n1591), .B1(n1590), .B2(r6[18]), .ZN(
        n1501) );
  AOI22D1BWP12T U2347 ( .A1(r8[18]), .A2(n1593), .B1(n1592), .B2(n[2023]), 
        .ZN(n1500) );
  AOI22D1BWP12T U2348 ( .A1(r5[18]), .A2(n1594), .B1(n171), .B2(r3[18]), .ZN(
        n1499) );
  AOI22D1BWP12T U2349 ( .A1(r7[18]), .A2(n1596), .B1(n1595), .B2(r0[18]), .ZN(
        n1498) );
  AN4XD1BWP12T U2350 ( .A1(n1501), .A2(n1500), .A3(n1499), .A4(n1498), .Z(
        n1508) );
  AOI22D1BWP12T U2351 ( .A1(n150), .A2(r12[18]), .B1(n1809), .B2(tmp1[18]), 
        .ZN(n1504) );
  AOI22D1BWP12T U2352 ( .A1(r2[18]), .A2(n155), .B1(n1555), .B2(r1[18]), .ZN(
        n1503) );
  ND2D1BWP12T U2353 ( .A1(n1957), .A2(r4[18]), .ZN(n1502) );
  AN3XD1BWP12T U2354 ( .A1(n1504), .A2(n1503), .A3(n1502), .Z(n1507) );
  AOI22D1BWP12T U2355 ( .A1(pc_out[18]), .A2(n141), .B1(n1559), .B2(r11[18]), 
        .ZN(n1506) );
  AOI22D1BWP12T U2356 ( .A1(lr[18]), .A2(n1561), .B1(n1560), .B2(r10[18]), 
        .ZN(n1505) );
  ND4D1BWP12T U2357 ( .A1(n1508), .A2(n1507), .A3(n1506), .A4(n1505), .ZN(
        regA_out[18]) );
  AOI22D1BWP12T U2358 ( .A1(tmp1[18]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[18]), .ZN(n1511) );
  AOI22D1BWP12T U2359 ( .A1(r9[18]), .A2(n201), .B1(n1780), .B2(r4[18]), .ZN(
        n1510) );
  AOI22D1BWP12T U2360 ( .A1(r11[18]), .A2(n2002), .B1(n205), .B2(r0[18]), .ZN(
        n1509) );
  ND3D1BWP12T U2361 ( .A1(n1511), .A2(n1510), .A3(n1509), .ZN(n1515) );
  AOI22D1BWP12T U2362 ( .A1(r5[18]), .A2(n210), .B1(n1988), .B2(r10[18]), .ZN(
        n1513) );
  AOI22D1BWP12T U2363 ( .A1(r7[18]), .A2(n215), .B1(n1989), .B2(r2[18]), .ZN(
        n1512) );
  ND2D1BWP12T U2364 ( .A1(n1513), .A2(n1512), .ZN(n1514) );
  NR2D1BWP12T U2365 ( .A1(n1515), .A2(n1514), .ZN(n1521) );
  AOI22D1BWP12T U2366 ( .A1(r1[18]), .A2(n183), .B1(n1992), .B2(r12[18]), .ZN(
        n1519) );
  AOI22D1BWP12T U2367 ( .A1(r3[18]), .A2(n185), .B1(n1993), .B2(lr[18]), .ZN(
        n1518) );
  AOI22D1BWP12T U2368 ( .A1(r8[18]), .A2(n187), .B1(n1994), .B2(n[2023]), .ZN(
        n1517) );
  AOI22D1BWP12T U2369 ( .A1(pc_out[18]), .A2(n188), .B1(n1995), .B2(r6[18]), 
        .ZN(n1516) );
  AN4XD1BWP12T U2370 ( .A1(n1519), .A2(n1518), .A3(n1517), .A4(n1516), .Z(
        n1520) );
  ND2D1BWP12T U2371 ( .A1(n1521), .A2(n1520), .ZN(regB_out[18]) );
  INVD0BWP12T U2372 ( .I(pc_out[17]), .ZN(n1523) );
  INVD1BWP12T U2373 ( .I(r11[17]), .ZN(n1522) );
  OAI22D1BWP12T U2374 ( .A1(n1523), .A2(n1949), .B1(n1948), .B2(n1522), .ZN(
        n1531) );
  INVD1BWP12T U2375 ( .I(r10[17]), .ZN(n1524) );
  OAI22D1BWP12T U2376 ( .A1(n1525), .A2(n1953), .B1(n1952), .B2(n1524), .ZN(
        n1530) );
  INVD1BWP12T U2377 ( .I(r2[17]), .ZN(n1527) );
  INVD1BWP12T U2378 ( .I(r1[17]), .ZN(n1526) );
  OAI22D1BWP12T U2379 ( .A1(n1961), .A2(n1527), .B1(n1959), .B2(n1526), .ZN(
        n1528) );
  NR4D0BWP12T U2380 ( .A1(n1531), .A2(n1530), .A3(n1529), .A4(n1528), .ZN(
        n1537) );
  AOI22D1BWP12T U2381 ( .A1(r9[17]), .A2(n1591), .B1(n1590), .B2(r6[17]), .ZN(
        n1535) );
  AOI22D1BWP12T U2382 ( .A1(r8[17]), .A2(n1593), .B1(n1592), .B2(n[2024]), 
        .ZN(n1534) );
  AOI22D1BWP12T U2383 ( .A1(r5[17]), .A2(n1594), .B1(n171), .B2(r3[17]), .ZN(
        n1533) );
  AOI22D1BWP12T U2384 ( .A1(r7[17]), .A2(n1596), .B1(n1595), .B2(r0[17]), .ZN(
        n1532) );
  AN4XD1BWP12T U2385 ( .A1(n1535), .A2(n1534), .A3(n1533), .A4(n1532), .Z(
        n1536) );
  ND2D1BWP12T U2386 ( .A1(n1537), .A2(n1536), .ZN(regA_out[17]) );
  AOI22D1BWP12T U2387 ( .A1(tmp1[17]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[17]), .ZN(n1540) );
  AOI22D1BWP12T U2388 ( .A1(r9[17]), .A2(n201), .B1(n1780), .B2(r4[17]), .ZN(
        n1539) );
  AOI22D1BWP12T U2389 ( .A1(r11[17]), .A2(n2002), .B1(n205), .B2(r0[17]), .ZN(
        n1538) );
  ND3D1BWP12T U2390 ( .A1(n1540), .A2(n1539), .A3(n1538), .ZN(n1544) );
  AOI22D1BWP12T U2391 ( .A1(r5[17]), .A2(n210), .B1(n1988), .B2(r10[17]), .ZN(
        n1542) );
  AOI22D1BWP12T U2392 ( .A1(r7[17]), .A2(n215), .B1(n1989), .B2(r2[17]), .ZN(
        n1541) );
  ND2D1BWP12T U2393 ( .A1(n1542), .A2(n1541), .ZN(n1543) );
  NR2D1BWP12T U2394 ( .A1(n1544), .A2(n1543), .ZN(n1550) );
  AOI22D1BWP12T U2395 ( .A1(r1[17]), .A2(n183), .B1(n1992), .B2(r12[17]), .ZN(
        n1548) );
  AOI22D1BWP12T U2396 ( .A1(r3[17]), .A2(n185), .B1(n1993), .B2(lr[17]), .ZN(
        n1547) );
  AOI22D1BWP12T U2397 ( .A1(r8[17]), .A2(n187), .B1(n1994), .B2(n[2024]), .ZN(
        n1546) );
  AOI22D1BWP12T U2398 ( .A1(pc_out[17]), .A2(n188), .B1(n1995), .B2(r6[17]), 
        .ZN(n1545) );
  AN4XD1BWP12T U2399 ( .A1(n1548), .A2(n1547), .A3(n1546), .A4(n1545), .Z(
        n1549) );
  ND2D1BWP12T U2400 ( .A1(n1550), .A2(n1549), .ZN(regB_out[17]) );
  AOI22D1BWP12T U2401 ( .A1(r9[16]), .A2(n1591), .B1(n1590), .B2(r6[16]), .ZN(
        n1554) );
  AOI22D1BWP12T U2402 ( .A1(r8[16]), .A2(n1593), .B1(n1592), .B2(n[2025]), 
        .ZN(n1553) );
  AOI22D1BWP12T U2403 ( .A1(r5[16]), .A2(n1594), .B1(n171), .B2(r3[16]), .ZN(
        n1552) );
  AOI22D1BWP12T U2404 ( .A1(r7[16]), .A2(n1596), .B1(n1595), .B2(r0[16]), .ZN(
        n1551) );
  AN4XD1BWP12T U2405 ( .A1(n1554), .A2(n1553), .A3(n1552), .A4(n1551), .Z(
        n1565) );
  AOI22D1BWP12T U2406 ( .A1(n150), .A2(r12[16]), .B1(n1809), .B2(tmp1[16]), 
        .ZN(n1558) );
  AOI22D1BWP12T U2407 ( .A1(r2[16]), .A2(n155), .B1(n1555), .B2(r1[16]), .ZN(
        n1557) );
  ND2D1BWP12T U2408 ( .A1(n1957), .A2(r4[16]), .ZN(n1556) );
  AN3XD1BWP12T U2409 ( .A1(n1558), .A2(n1557), .A3(n1556), .Z(n1564) );
  AOI22D1BWP12T U2410 ( .A1(pc_out[16]), .A2(n141), .B1(n1559), .B2(r11[16]), 
        .ZN(n1563) );
  AOI22D1BWP12T U2411 ( .A1(lr[16]), .A2(n1561), .B1(n1560), .B2(r10[16]), 
        .ZN(n1562) );
  ND4D1BWP12T U2412 ( .A1(n1565), .A2(n1564), .A3(n1563), .A4(n1562), .ZN(
        regA_out[16]) );
  AOI22D1BWP12T U2413 ( .A1(tmp1[16]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[16]), .ZN(n1568) );
  AOI22D1BWP12T U2414 ( .A1(r9[16]), .A2(n201), .B1(n1780), .B2(r4[16]), .ZN(
        n1567) );
  AOI22D1BWP12T U2415 ( .A1(r11[16]), .A2(n2002), .B1(n205), .B2(r0[16]), .ZN(
        n1566) );
  ND3D1BWP12T U2416 ( .A1(n1568), .A2(n1567), .A3(n1566), .ZN(n1572) );
  AOI22D1BWP12T U2417 ( .A1(r5[16]), .A2(n210), .B1(n1988), .B2(r10[16]), .ZN(
        n1570) );
  AOI22D1BWP12T U2418 ( .A1(r7[16]), .A2(n215), .B1(n1989), .B2(r2[16]), .ZN(
        n1569) );
  ND2D1BWP12T U2419 ( .A1(n1570), .A2(n1569), .ZN(n1571) );
  NR2D1BWP12T U2420 ( .A1(n1572), .A2(n1571), .ZN(n1578) );
  AOI22D1BWP12T U2421 ( .A1(r1[16]), .A2(n183), .B1(n1992), .B2(r12[16]), .ZN(
        n1576) );
  AOI22D1BWP12T U2422 ( .A1(r3[16]), .A2(n185), .B1(n1993), .B2(lr[16]), .ZN(
        n1575) );
  AOI22D1BWP12T U2423 ( .A1(r8[16]), .A2(n187), .B1(n1994), .B2(n[2025]), .ZN(
        n1574) );
  AOI22D1BWP12T U2424 ( .A1(pc_out[16]), .A2(n188), .B1(n1995), .B2(r6[16]), 
        .ZN(n1573) );
  AN4XD1BWP12T U2425 ( .A1(n1576), .A2(n1575), .A3(n1574), .A4(n1573), .Z(
        n1577) );
  ND2D1BWP12T U2426 ( .A1(n1578), .A2(n1577), .ZN(regB_out[16]) );
  INVD0BWP12T U2427 ( .I(pc_out[15]), .ZN(n1580) );
  INVD1BWP12T U2428 ( .I(r11[15]), .ZN(n1579) );
  OAI22D1BWP12T U2429 ( .A1(n1580), .A2(n1949), .B1(n1948), .B2(n1579), .ZN(
        n1589) );
  INVD1BWP12T U2430 ( .I(r10[15]), .ZN(n1581) );
  OAI22D1BWP12T U2431 ( .A1(n1582), .A2(n1953), .B1(n1952), .B2(n1581), .ZN(
        n1588) );
  AOI22D1BWP12T U2432 ( .A1(n150), .A2(r12[15]), .B1(n1809), .B2(tmp1[15]), 
        .ZN(n1583) );
  IOA21D1BWP12T U2433 ( .A1(n1957), .A2(r4[15]), .B(n1583), .ZN(n1587) );
  INVD1BWP12T U2434 ( .I(r2[15]), .ZN(n1585) );
  INVD1BWP12T U2435 ( .I(r1[15]), .ZN(n1584) );
  OAI22D1BWP12T U2436 ( .A1(n1961), .A2(n1585), .B1(n1959), .B2(n1584), .ZN(
        n1586) );
  NR4D0BWP12T U2437 ( .A1(n1589), .A2(n1588), .A3(n1587), .A4(n1586), .ZN(
        n1602) );
  AOI22D1BWP12T U2438 ( .A1(r9[15]), .A2(n1591), .B1(n1590), .B2(r6[15]), .ZN(
        n1600) );
  AOI22D1BWP12T U2439 ( .A1(r8[15]), .A2(n1593), .B1(n1592), .B2(n[2026]), 
        .ZN(n1599) );
  AOI22D1BWP12T U2440 ( .A1(r5[15]), .A2(n1594), .B1(n171), .B2(r3[15]), .ZN(
        n1598) );
  AOI22D1BWP12T U2441 ( .A1(r7[15]), .A2(n1596), .B1(n1595), .B2(r0[15]), .ZN(
        n1597) );
  AN4XD1BWP12T U2442 ( .A1(n1600), .A2(n1599), .A3(n1598), .A4(n1597), .Z(
        n1601) );
  ND2D1BWP12T U2443 ( .A1(n1602), .A2(n1601), .ZN(regA_out[15]) );
  AOI22D1BWP12T U2444 ( .A1(tmp1[15]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[15]), .ZN(n1605) );
  AOI22D1BWP12T U2445 ( .A1(r9[15]), .A2(n201), .B1(n1780), .B2(r4[15]), .ZN(
        n1604) );
  AOI22D1BWP12T U2446 ( .A1(r11[15]), .A2(n2002), .B1(n205), .B2(r0[15]), .ZN(
        n1603) );
  ND3D1BWP12T U2447 ( .A1(n1605), .A2(n1604), .A3(n1603), .ZN(n1609) );
  AOI22D1BWP12T U2448 ( .A1(r5[15]), .A2(n210), .B1(n1988), .B2(r10[15]), .ZN(
        n1607) );
  AOI22D1BWP12T U2449 ( .A1(r7[15]), .A2(n215), .B1(n1989), .B2(r2[15]), .ZN(
        n1606) );
  ND2D1BWP12T U2450 ( .A1(n1607), .A2(n1606), .ZN(n1608) );
  NR2D1BWP12T U2451 ( .A1(n1609), .A2(n1608), .ZN(n1615) );
  AOI22D1BWP12T U2452 ( .A1(r1[15]), .A2(n183), .B1(n1992), .B2(r12[15]), .ZN(
        n1613) );
  AOI22D1BWP12T U2453 ( .A1(r3[15]), .A2(n185), .B1(n1993), .B2(lr[15]), .ZN(
        n1612) );
  AOI22D1BWP12T U2454 ( .A1(r8[15]), .A2(n187), .B1(n1994), .B2(n[2026]), .ZN(
        n1611) );
  AOI22D1BWP12T U2455 ( .A1(pc_out[15]), .A2(n188), .B1(n1995), .B2(r6[15]), 
        .ZN(n1610) );
  AN4XD1BWP12T U2456 ( .A1(n1613), .A2(n1612), .A3(n1611), .A4(n1610), .Z(
        n1614) );
  ND2D1BWP12T U2457 ( .A1(n1615), .A2(n1614), .ZN(regB_out[15]) );
  AOI22D1BWP12T U2458 ( .A1(tmp1[13]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[13]), .ZN(n1618) );
  AOI22D1BWP12T U2459 ( .A1(r9[13]), .A2(n201), .B1(n1780), .B2(r4[13]), .ZN(
        n1617) );
  AOI22D1BWP12T U2460 ( .A1(r11[13]), .A2(n2002), .B1(n205), .B2(r0[13]), .ZN(
        n1616) );
  ND3D1BWP12T U2461 ( .A1(n1618), .A2(n1617), .A3(n1616), .ZN(n1628) );
  AOI22D1BWP12T U2462 ( .A1(r1[13]), .A2(n183), .B1(n1992), .B2(r12[13]), .ZN(
        n1620) );
  AOI22D1BWP12T U2463 ( .A1(r8[13]), .A2(n187), .B1(n1994), .B2(n[2028]), .ZN(
        n1619) );
  ND2D1BWP12T U2464 ( .A1(n1620), .A2(n1619), .ZN(n1627) );
  AOI22D1BWP12T U2465 ( .A1(r3[13]), .A2(n185), .B1(n1993), .B2(lr[13]), .ZN(
        n1622) );
  AOI22D1BWP12T U2466 ( .A1(pc_out[13]), .A2(n188), .B1(n1995), .B2(r6[13]), 
        .ZN(n1621) );
  ND2D1BWP12T U2467 ( .A1(n1622), .A2(n1621), .ZN(n1626) );
  AOI22D1BWP12T U2468 ( .A1(r5[13]), .A2(n210), .B1(n1988), .B2(r10[13]), .ZN(
        n1624) );
  AOI22D1BWP12T U2469 ( .A1(r7[13]), .A2(n215), .B1(n1989), .B2(r2[13]), .ZN(
        n1623) );
  ND2D1BWP12T U2470 ( .A1(n1624), .A2(n1623), .ZN(n1625) );
  OR4XD1BWP12T U2471 ( .A1(n1628), .A2(n1627), .A3(n1626), .A4(n1625), .Z(
        regB_out[13]) );
  OAI22D1BWP12T U2472 ( .A1(n1630), .A2(n1949), .B1(n1948), .B2(n1629), .ZN(
        n1639) );
  OAI22D1BWP12T U2473 ( .A1(n1632), .A2(n1953), .B1(n1952), .B2(n1631), .ZN(
        n1638) );
  AOI22D1BWP12T U2474 ( .A1(n150), .A2(r12[12]), .B1(n1809), .B2(tmp1[12]), 
        .ZN(n1633) );
  IOA21D1BWP12T U2475 ( .A1(n1957), .A2(r4[12]), .B(n1633), .ZN(n1637) );
  OAI22D1BWP12T U2476 ( .A1(n1961), .A2(n1635), .B1(n1959), .B2(n1634), .ZN(
        n1636) );
  NR4D0BWP12T U2477 ( .A1(n1639), .A2(n1638), .A3(n1637), .A4(n1636), .ZN(
        n1653) );
  OAI22D1BWP12T U2478 ( .A1(n1969), .A2(n1641), .B1(n1967), .B2(n1640), .ZN(
        n1651) );
  OAI22D1BWP12T U2479 ( .A1(n1973), .A2(n1643), .B1(n1971), .B2(n1642), .ZN(
        n1650) );
  OAI22D1BWP12T U2480 ( .A1(n1645), .A2(n1976), .B1(n1975), .B2(n1644), .ZN(
        n1649) );
  OAI22D1BWP12T U2481 ( .A1(n1981), .A2(n1647), .B1(n1979), .B2(n1646), .ZN(
        n1648) );
  NR4D0BWP12T U2482 ( .A1(n1651), .A2(n1650), .A3(n1649), .A4(n1648), .ZN(
        n1652) );
  ND2D1BWP12T U2483 ( .A1(n1653), .A2(n1652), .ZN(regA_out[12]) );
  OAI22D1BWP12T U2484 ( .A1(n1655), .A2(n1949), .B1(n1948), .B2(n1654), .ZN(
        n1664) );
  OAI22D1BWP12T U2485 ( .A1(n1657), .A2(n1953), .B1(n1952), .B2(n1656), .ZN(
        n1663) );
  AOI22D1BWP12T U2486 ( .A1(n150), .A2(r12[11]), .B1(n1809), .B2(tmp1[11]), 
        .ZN(n1658) );
  IOA21D1BWP12T U2487 ( .A1(n1957), .A2(r4[11]), .B(n1658), .ZN(n1662) );
  OAI22D1BWP12T U2488 ( .A1(n1961), .A2(n1660), .B1(n1959), .B2(n1659), .ZN(
        n1661) );
  OAI22D1BWP12T U2489 ( .A1(n1969), .A2(n1666), .B1(n1967), .B2(n1665), .ZN(
        n1676) );
  OAI22D1BWP12T U2490 ( .A1(n1973), .A2(n1668), .B1(n1971), .B2(n1667), .ZN(
        n1675) );
  OAI22D1BWP12T U2491 ( .A1(n1670), .A2(n1976), .B1(n1975), .B2(n1669), .ZN(
        n1674) );
  OAI22D1BWP12T U2492 ( .A1(n1981), .A2(n1672), .B1(n1979), .B2(n1671), .ZN(
        n1673) );
  NR4D0BWP12T U2493 ( .A1(n1676), .A2(n1675), .A3(n1674), .A4(n1673), .ZN(
        n1677) );
  OAI22D1BWP12T U2494 ( .A1(n1679), .A2(n1949), .B1(n1948), .B2(n1678), .ZN(
        n1688) );
  OAI22D1BWP12T U2495 ( .A1(n1681), .A2(n1953), .B1(n1952), .B2(n1680), .ZN(
        n1687) );
  AOI22D1BWP12T U2496 ( .A1(n150), .A2(r12[10]), .B1(n1809), .B2(tmp1[10]), 
        .ZN(n1682) );
  IOA21D1BWP12T U2497 ( .A1(n1957), .A2(r4[10]), .B(n1682), .ZN(n1686) );
  OAI22D1BWP12T U2498 ( .A1(n1961), .A2(n1684), .B1(n1959), .B2(n1683), .ZN(
        n1685) );
  NR4D0BWP12T U2499 ( .A1(n1688), .A2(n1687), .A3(n1686), .A4(n1685), .ZN(
        n1702) );
  OAI22D1BWP12T U2500 ( .A1(n1973), .A2(n1692), .B1(n1971), .B2(n1691), .ZN(
        n1699) );
  OAI22D1BWP12T U2501 ( .A1(n1694), .A2(n1976), .B1(n1975), .B2(n1693), .ZN(
        n1698) );
  OAI22D1BWP12T U2502 ( .A1(n1981), .A2(n1696), .B1(n1979), .B2(n1695), .ZN(
        n1697) );
  NR4D0BWP12T U2503 ( .A1(n1700), .A2(n1699), .A3(n1698), .A4(n1697), .ZN(
        n1701) );
  ND2D1BWP12T U2504 ( .A1(n1702), .A2(n1701), .ZN(regA_out[10]) );
  INVD1BWP12T U2505 ( .I(pc_out[9]), .ZN(n1733) );
  AOI22D1BWP12T U2506 ( .A1(n150), .A2(r12[9]), .B1(n1809), .B2(tmp1[9]), .ZN(
        n1704) );
  IOA21D1BWP12T U2507 ( .A1(n1957), .A2(r4[9]), .B(n1704), .ZN(n1706) );
  OAI22D1BWP12T U2508 ( .A1(n1961), .A2(n1720), .B1(n1959), .B2(n1727), .ZN(
        n1705) );
  OAI22D1BWP12T U2509 ( .A1(n1969), .A2(n1707), .B1(n1967), .B2(n1732), .ZN(
        n1712) );
  INVD1BWP12T U2510 ( .I(n[2032]), .ZN(n1730) );
  OAI22D1BWP12T U2511 ( .A1(n1981), .A2(n1721), .B1(n1979), .B2(n1708), .ZN(
        n1709) );
  NR4D0BWP12T U2512 ( .A1(n1712), .A2(n1711), .A3(n1710), .A4(n1709), .ZN(
        n1713) );
  ND2D1BWP12T U2513 ( .A1(n1714), .A2(n1713), .ZN(regA_out[9]) );
  INVD0BWP12T U2514 ( .I(tmp1[9]), .ZN(n1715) );
  MOAI22D0BWP12T U2515 ( .A1(n1715), .A2(n1847), .B1(n200), .B2(
        immediate2_in[9]), .ZN(n1725) );
  AOI22D1BWP12T U2516 ( .A1(r9[9]), .A2(n201), .B1(n1780), .B2(r4[9]), .ZN(
        n1717) );
  AOI22D1BWP12T U2517 ( .A1(r11[9]), .A2(n2002), .B1(n205), .B2(r0[9]), .ZN(
        n1716) );
  ND2D1BWP12T U2518 ( .A1(n1717), .A2(n1716), .ZN(n1724) );
  OAI22D1BWP12T U2519 ( .A1(n1719), .A2(n1846), .B1(n1845), .B2(n1718), .ZN(
        n1723) );
  OAI22D1BWP12T U2520 ( .A1(n1852), .A2(n1721), .B1(n1851), .B2(n1720), .ZN(
        n1722) );
  NR4D0BWP12T U2521 ( .A1(n1725), .A2(n1724), .A3(n1723), .A4(n1722), .ZN(
        n1739) );
  OAI22D1BWP12T U2522 ( .A1(n1727), .A2(n1859), .B1(n1858), .B2(n1726), .ZN(
        n1737) );
  OAI22D1BWP12T U2523 ( .A1(n1729), .A2(n1861), .B1(n1860), .B2(n1728), .ZN(
        n1736) );
  OAI22D1BWP12T U2524 ( .A1(n1863), .A2(n1731), .B1(n1862), .B2(n1730), .ZN(
        n1735) );
  OAI22D1BWP12T U2525 ( .A1(n1865), .A2(n1733), .B1(n1864), .B2(n1732), .ZN(
        n1734) );
  NR4D0BWP12T U2526 ( .A1(n1737), .A2(n1736), .A3(n1735), .A4(n1734), .ZN(
        n1738) );
  ND2D1BWP12T U2527 ( .A1(n1739), .A2(n1738), .ZN(regB_out[9]) );
  OAI22D1BWP12T U2528 ( .A1(n1741), .A2(n1949), .B1(n1948), .B2(n1740), .ZN(
        n1750) );
  OAI22D1BWP12T U2529 ( .A1(n1743), .A2(n1953), .B1(n1952), .B2(n1742), .ZN(
        n1749) );
  AOI22D1BWP12T U2530 ( .A1(n150), .A2(r12[8]), .B1(n1809), .B2(tmp1[8]), .ZN(
        n1744) );
  IOA21D1BWP12T U2531 ( .A1(n1957), .A2(r4[8]), .B(n1744), .ZN(n1748) );
  OAI22D1BWP12T U2532 ( .A1(n1961), .A2(n1746), .B1(n1959), .B2(n1745), .ZN(
        n1747) );
  NR4D0BWP12T U2533 ( .A1(n1750), .A2(n1749), .A3(n1748), .A4(n1747), .ZN(
        n1764) );
  OAI22D1BWP12T U2534 ( .A1(n1969), .A2(n1752), .B1(n1967), .B2(n1751), .ZN(
        n1762) );
  OAI22D1BWP12T U2535 ( .A1(n1973), .A2(n1754), .B1(n1971), .B2(n1753), .ZN(
        n1761) );
  OAI22D1BWP12T U2536 ( .A1(n1756), .A2(n1976), .B1(n1975), .B2(n1755), .ZN(
        n1760) );
  OAI22D1BWP12T U2537 ( .A1(n1981), .A2(n1758), .B1(n1979), .B2(n1757), .ZN(
        n1759) );
  NR4D0BWP12T U2538 ( .A1(n1762), .A2(n1761), .A3(n1760), .A4(n1759), .ZN(
        n1763) );
  ND2D1BWP12T U2539 ( .A1(n1764), .A2(n1763), .ZN(regA_out[8]) );
  INVD1BWP12T U2540 ( .I(pc_out[7]), .ZN(n1798) );
  OAI22D1BWP12T U2541 ( .A1(n1798), .A2(n1949), .B1(n1948), .B2(n1765), .ZN(
        n1770) );
  OAI22D1BWP12T U2542 ( .A1(n1793), .A2(n1953), .B1(n1952), .B2(n1783), .ZN(
        n1769) );
  AOI22D1BWP12T U2543 ( .A1(n150), .A2(r12[7]), .B1(n1809), .B2(tmp1[7]), .ZN(
        n1766) );
  IOA21D1BWP12T U2544 ( .A1(n1957), .A2(r4[7]), .B(n1766), .ZN(n1768) );
  OAI22D1BWP12T U2545 ( .A1(n1961), .A2(n1785), .B1(n1959), .B2(n1792), .ZN(
        n1767) );
  OAI22D1BWP12T U2546 ( .A1(n1969), .A2(n1771), .B1(n1967), .B2(n1797), .ZN(
        n1776) );
  INVD1BWP12T U2547 ( .I(n[2034]), .ZN(n1795) );
  OAI22D1BWP12T U2548 ( .A1(n1973), .A2(n1796), .B1(n1971), .B2(n1795), .ZN(
        n1775) );
  OAI22D1BWP12T U2549 ( .A1(n1784), .A2(n1976), .B1(n1975), .B2(n1794), .ZN(
        n1774) );
  OAI22D1BWP12T U2550 ( .A1(n1981), .A2(n1786), .B1(n1979), .B2(n1772), .ZN(
        n1773) );
  NR4D0BWP12T U2551 ( .A1(n1776), .A2(n1775), .A3(n1774), .A4(n1773), .ZN(
        n1777) );
  ND2D1BWP12T U2552 ( .A1(n1778), .A2(n1777), .ZN(regA_out[7]) );
  INVD0BWP12T U2553 ( .I(tmp1[7]), .ZN(n1779) );
  MOAI22D0BWP12T U2554 ( .A1(n1779), .A2(n1847), .B1(n200), .B2(
        immediate2_in[7]), .ZN(n1790) );
  AOI22D1BWP12T U2555 ( .A1(r9[7]), .A2(n201), .B1(n1780), .B2(r4[7]), .ZN(
        n1782) );
  AOI22D1BWP12T U2556 ( .A1(r11[7]), .A2(n537), .B1(n205), .B2(r0[7]), .ZN(
        n1781) );
  ND2D1BWP12T U2557 ( .A1(n1782), .A2(n1781), .ZN(n1789) );
  OAI22D1BWP12T U2558 ( .A1(n1784), .A2(n1846), .B1(n1845), .B2(n1783), .ZN(
        n1788) );
  OAI22D1BWP12T U2559 ( .A1(n1852), .A2(n1786), .B1(n1851), .B2(n1785), .ZN(
        n1787) );
  NR4D0BWP12T U2560 ( .A1(n1790), .A2(n1789), .A3(n1788), .A4(n1787), .ZN(
        n1804) );
  OAI22D1BWP12T U2561 ( .A1(n1792), .A2(n1859), .B1(n1858), .B2(n1791), .ZN(
        n1802) );
  OAI22D1BWP12T U2562 ( .A1(n1794), .A2(n1861), .B1(n1860), .B2(n1793), .ZN(
        n1801) );
  OAI22D1BWP12T U2563 ( .A1(n1863), .A2(n1796), .B1(n1862), .B2(n1795), .ZN(
        n1800) );
  OAI22D1BWP12T U2564 ( .A1(n1865), .A2(n1798), .B1(n1864), .B2(n1797), .ZN(
        n1799) );
  NR4D0BWP12T U2565 ( .A1(n1802), .A2(n1801), .A3(n1800), .A4(n1799), .ZN(
        n1803) );
  ND2D1BWP12T U2566 ( .A1(n1804), .A2(n1803), .ZN(regB_out[7]) );
  OAI22D1BWP12T U2567 ( .A1(n1806), .A2(n1949), .B1(n1948), .B2(n1805), .ZN(
        n1816) );
  OAI22D1BWP12T U2568 ( .A1(n1808), .A2(n1953), .B1(n1952), .B2(n1807), .ZN(
        n1815) );
  AOI22D1BWP12T U2569 ( .A1(n150), .A2(r12[6]), .B1(n1809), .B2(tmp1[6]), .ZN(
        n1810) );
  IOA21D1BWP12T U2570 ( .A1(n1957), .A2(r4[6]), .B(n1810), .ZN(n1814) );
  OAI22D1BWP12T U2571 ( .A1(n1961), .A2(n1812), .B1(n1959), .B2(n1811), .ZN(
        n1813) );
  NR4D0BWP12T U2572 ( .A1(n1816), .A2(n1815), .A3(n1814), .A4(n1813), .ZN(
        n1830) );
  OAI22D1BWP12T U2573 ( .A1(n1969), .A2(n1818), .B1(n1967), .B2(n1817), .ZN(
        n1828) );
  OAI22D1BWP12T U2574 ( .A1(n1973), .A2(n1820), .B1(n1971), .B2(n1819), .ZN(
        n1827) );
  OAI22D1BWP12T U2575 ( .A1(n1822), .A2(n1976), .B1(n1975), .B2(n1821), .ZN(
        n1826) );
  OAI22D1BWP12T U2576 ( .A1(n1981), .A2(n1824), .B1(n1979), .B2(n1823), .ZN(
        n1825) );
  NR4D0BWP12T U2577 ( .A1(n1828), .A2(n1827), .A3(n1826), .A4(n1825), .ZN(
        n1829) );
  ND2D1BWP12T U2578 ( .A1(n1830), .A2(n1829), .ZN(regA_out[6]) );
  INVD0BWP12T U2579 ( .I(tmp1[5]), .ZN(n1831) );
  MOAI22D0BWP12T U2580 ( .A1(n1831), .A2(n1847), .B1(n200), .B2(
        immediate2_in[5]), .ZN(n1837) );
  AOI22D1BWP12T U2581 ( .A1(r9[5]), .A2(n201), .B1(n1780), .B2(r4[5]), .ZN(
        n1833) );
  AOI22D1BWP12T U2582 ( .A1(r11[5]), .A2(n537), .B1(n205), .B2(r0[5]), .ZN(
        n1832) );
  ND2D1BWP12T U2583 ( .A1(n1833), .A2(n1832), .ZN(n1836) );
  OAI22D1BWP12T U2584 ( .A1(n1913), .A2(n1846), .B1(n1845), .B2(n1899), .ZN(
        n1835) );
  NR4D0BWP12T U2585 ( .A1(n1837), .A2(n1836), .A3(n1835), .A4(n1834), .ZN(
        n1844) );
  OAI22D1BWP12T U2586 ( .A1(n1902), .A2(n1859), .B1(n1858), .B2(n1838), .ZN(
        n1842) );
  OAI22D1BWP12T U2587 ( .A1(n1912), .A2(n1861), .B1(n1860), .B2(n1900), .ZN(
        n1841) );
  INVD1BWP12T U2588 ( .I(n[2036]), .ZN(n1910) );
  OAI22D1BWP12T U2589 ( .A1(n1863), .A2(n1911), .B1(n1862), .B2(n1910), .ZN(
        n1840) );
  INVD1BWP12T U2590 ( .I(pc_out[5]), .ZN(n1898) );
  OAI22D1BWP12T U2591 ( .A1(n1865), .A2(n1898), .B1(n1864), .B2(n1908), .ZN(
        n1839) );
  NR4D0BWP12T U2592 ( .A1(n1842), .A2(n1841), .A3(n1840), .A4(n1839), .ZN(
        n1843) );
  ND2D1BWP12T U2593 ( .A1(n1844), .A2(n1843), .ZN(regB_out[5]) );
  OAI22D1BWP12T U2594 ( .A1(n1938), .A2(n1846), .B1(n1845), .B2(n1924), .ZN(
        n1856) );
  INVD1BWP12T U2595 ( .I(tmp1[1]), .ZN(n1848) );
  AOI22D1BWP12T U2596 ( .A1(r9[1]), .A2(n201), .B1(n536), .B2(r4[1]), .ZN(
        n1850) );
  NR4D0BWP12T U2597 ( .A1(n1856), .A2(n1855), .A3(n1854), .A4(n1853), .ZN(
        n1871) );
  TPOAI22D1BWP12T U2598 ( .A1(n1927), .A2(n1859), .B1(n1858), .B2(n1857), .ZN(
        n1869) );
  INVD1BWP12T U2599 ( .I(n[2040]), .ZN(n1935) );
  TPOAI22D1BWP12T U2600 ( .A1(n1863), .A2(n1936), .B1(n1862), .B2(n1935), .ZN(
        n1867) );
  INVD1BWP12T U2601 ( .I(pc_out[1]), .ZN(n1923) );
  TPOAI22D1BWP12T U2602 ( .A1(n1865), .A2(n1923), .B1(n1864), .B2(n1933), .ZN(
        n1866) );
  OAI22D1BWP12T U2603 ( .A1(n1873), .A2(n1949), .B1(n1948), .B2(n1872), .ZN(
        n1882) );
  OAI22D1BWP12T U2604 ( .A1(n1875), .A2(n1953), .B1(n1952), .B2(n1874), .ZN(
        n1881) );
  AOI22D1BWP12T U2605 ( .A1(n150), .A2(r12[4]), .B1(n1955), .B2(tmp1[4]), .ZN(
        n1876) );
  IOA21D1BWP12T U2606 ( .A1(n1957), .A2(r4[4]), .B(n1876), .ZN(n1880) );
  OAI22D1BWP12T U2607 ( .A1(n1961), .A2(n1878), .B1(n1959), .B2(n1877), .ZN(
        n1879) );
  NR4D0BWP12T U2608 ( .A1(n1882), .A2(n1881), .A3(n1880), .A4(n1879), .ZN(
        n1896) );
  OAI22D1BWP12T U2609 ( .A1(n1969), .A2(n1884), .B1(n1967), .B2(n1883), .ZN(
        n1894) );
  OAI22D1BWP12T U2610 ( .A1(n1973), .A2(n1886), .B1(n1971), .B2(n1885), .ZN(
        n1893) );
  OAI22D1BWP12T U2611 ( .A1(n1888), .A2(n1976), .B1(n1975), .B2(n1887), .ZN(
        n1892) );
  OAI22D1BWP12T U2612 ( .A1(n1981), .A2(n1890), .B1(n1979), .B2(n1889), .ZN(
        n1891) );
  NR4D0BWP12T U2613 ( .A1(n1894), .A2(n1893), .A3(n1892), .A4(n1891), .ZN(
        n1895) );
  ND2D1BWP12T U2614 ( .A1(n1896), .A2(n1895), .ZN(regA_out[4]) );
  OAI22D1BWP12T U2615 ( .A1(n1898), .A2(n1949), .B1(n1948), .B2(n1897), .ZN(
        n1907) );
  OAI22D1BWP12T U2616 ( .A1(n1900), .A2(n1953), .B1(n1952), .B2(n1899), .ZN(
        n1906) );
  AOI22D1BWP12T U2617 ( .A1(n150), .A2(r12[5]), .B1(n1955), .B2(tmp1[5]), .ZN(
        n1901) );
  IOA21D1BWP12T U2618 ( .A1(n1957), .A2(r4[5]), .B(n1901), .ZN(n1905) );
  OAI22D1BWP12T U2619 ( .A1(n1961), .A2(n1903), .B1(n1959), .B2(n1902), .ZN(
        n1904) );
  NR4D1BWP12T U2620 ( .A1(n1907), .A2(n1906), .A3(n1905), .A4(n1904), .ZN(
        n1921) );
  OAI22D1BWP12T U2621 ( .A1(n1969), .A2(n1909), .B1(n1967), .B2(n1908), .ZN(
        n1919) );
  OAI22D1BWP12T U2622 ( .A1(n1973), .A2(n1911), .B1(n1971), .B2(n1910), .ZN(
        n1918) );
  OAI22D1BWP12T U2623 ( .A1(n1913), .A2(n1976), .B1(n1975), .B2(n1912), .ZN(
        n1917) );
  OAI22D1BWP12T U2624 ( .A1(n1981), .A2(n1915), .B1(n1979), .B2(n1914), .ZN(
        n1916) );
  NR4D0BWP12T U2625 ( .A1(n1919), .A2(n1918), .A3(n1917), .A4(n1916), .ZN(
        n1920) );
  ND2D1BWP12T U2626 ( .A1(n1921), .A2(n1920), .ZN(regA_out[5]) );
  OAI22D1BWP12T U2627 ( .A1(n1923), .A2(n1949), .B1(n1948), .B2(n1922), .ZN(
        n1932) );
  OAI22D1BWP12T U2628 ( .A1(n1925), .A2(n1953), .B1(n1952), .B2(n1924), .ZN(
        n1931) );
  AOI22D1BWP12T U2629 ( .A1(n150), .A2(r12[1]), .B1(n1955), .B2(tmp1[1]), .ZN(
        n1926) );
  IOA21D1BWP12T U2630 ( .A1(n1957), .A2(r4[1]), .B(n1926), .ZN(n1930) );
  OAI22D1BWP12T U2631 ( .A1(n1961), .A2(n1928), .B1(n1959), .B2(n1927), .ZN(
        n1929) );
  NR4D1BWP12T U2632 ( .A1(n1932), .A2(n1931), .A3(n1930), .A4(n1929), .ZN(
        n1946) );
  OAI22D1BWP12T U2633 ( .A1(n1969), .A2(n1934), .B1(n1967), .B2(n1933), .ZN(
        n1944) );
  OAI22D1BWP12T U2634 ( .A1(n1973), .A2(n1936), .B1(n1971), .B2(n1935), .ZN(
        n1943) );
  OAI22D1BWP12T U2635 ( .A1(n1938), .A2(n1976), .B1(n1975), .B2(n1937), .ZN(
        n1942) );
  OAI22D1BWP12T U2636 ( .A1(n1981), .A2(n1940), .B1(n1979), .B2(n1939), .ZN(
        n1941) );
  NR4D0BWP12T U2637 ( .A1(n1944), .A2(n1943), .A3(n1942), .A4(n1941), .ZN(
        n1945) );
  ND2D1BWP12T U2638 ( .A1(n1946), .A2(n1945), .ZN(regA_out[1]) );
  OAI22D1BWP12T U2639 ( .A1(n1950), .A2(n1949), .B1(n1948), .B2(n1947), .ZN(
        n1965) );
  OAI22D1BWP12T U2640 ( .A1(n1954), .A2(n1953), .B1(n1952), .B2(n1951), .ZN(
        n1964) );
  AOI22D1BWP12T U2641 ( .A1(n150), .A2(r12[2]), .B1(n1955), .B2(tmp1[2]), .ZN(
        n1956) );
  IOA21D1BWP12T U2642 ( .A1(n1957), .A2(r4[2]), .B(n1956), .ZN(n1963) );
  OAI22D1BWP12T U2643 ( .A1(n1961), .A2(n1960), .B1(n1959), .B2(n1958), .ZN(
        n1962) );
  NR4D0BWP12T U2644 ( .A1(n1965), .A2(n1964), .A3(n1963), .A4(n1962), .ZN(
        n1987) );
  OAI22D1BWP12T U2645 ( .A1(n1969), .A2(n1968), .B1(n1967), .B2(n1966), .ZN(
        n1985) );
  OAI22D1BWP12T U2646 ( .A1(n1973), .A2(n1972), .B1(n1971), .B2(n1970), .ZN(
        n1984) );
  OAI22D1BWP12T U2647 ( .A1(n1977), .A2(n1976), .B1(n1975), .B2(n1974), .ZN(
        n1983) );
  OAI22D1BWP12T U2648 ( .A1(n1981), .A2(n1980), .B1(n1979), .B2(n1978), .ZN(
        n1982) );
  NR4D0BWP12T U2649 ( .A1(n1985), .A2(n1984), .A3(n1983), .A4(n1982), .ZN(
        n1986) );
  ND2D1BWP12T U2650 ( .A1(n1987), .A2(n1986), .ZN(regA_out[2]) );
  INR2D1BWP12T U2651 ( .A1(next_cpsr_in[3]), .B1(reset), .ZN(cpsrin[3]) );
  INR2D1BWP12T U2652 ( .A1(next_cpsr_in[1]), .B1(reset), .ZN(cpsrin[1]) );
  AOI22D1BWP12T U2653 ( .A1(r5[19]), .A2(n210), .B1(n1988), .B2(r10[19]), .ZN(
        n1991) );
  AOI22D1BWP12T U2654 ( .A1(r7[19]), .A2(n215), .B1(n1989), .B2(r2[19]), .ZN(
        n1990) );
  ND2D1BWP12T U2655 ( .A1(n1991), .A2(n1990), .ZN(n2008) );
  AOI22D1BWP12T U2656 ( .A1(r1[19]), .A2(n183), .B1(n1992), .B2(r12[19]), .ZN(
        n1999) );
  AOI22D1BWP12T U2657 ( .A1(r3[19]), .A2(n185), .B1(n1993), .B2(lr[19]), .ZN(
        n1998) );
  AOI22D1BWP12T U2658 ( .A1(r8[19]), .A2(n187), .B1(n1994), .B2(n[2022]), .ZN(
        n1997) );
  AOI22D1BWP12T U2659 ( .A1(pc_out[19]), .A2(n188), .B1(n1995), .B2(r6[19]), 
        .ZN(n1996) );
  AN4XD1BWP12T U2660 ( .A1(n1999), .A2(n1998), .A3(n1997), .A4(n1996), .Z(
        n2007) );
  AOI22D1BWP12T U2661 ( .A1(tmp1[19]), .A2(n2000), .B1(n200), .B2(
        immediate2_in[19]), .ZN(n2005) );
  AOI22D1BWP12T U2662 ( .A1(r9[19]), .A2(n201), .B1(n2001), .B2(r4[19]), .ZN(
        n2004) );
  AOI22D1BWP12T U2663 ( .A1(r11[19]), .A2(n2002), .B1(n205), .B2(r0[19]), .ZN(
        n2003) );
  AN3XD1BWP12T U2664 ( .A1(n2005), .A2(n2004), .A3(n2003), .Z(n2006) );
  IND3D1BWP12T U2665 ( .A1(n2008), .B1(n2007), .B2(n2006), .ZN(regB_out[19])
         );
endmodule


module ALU_VARIABLE ( a, b, op, c_in, result, c_out, z, n, v );
  input [31:0] a;
  input [31:0] b;
  input [3:0] op;
  output [31:0] result;
  input c_in;
  output c_out, z, n, v;
  wire   mult_x_18_n1029, mult_x_18_n1025, mult_x_18_n1021, mult_x_18_n1017,
         mult_x_18_n1013, mult_x_18_n1009, mult_x_18_n1005, mult_x_18_n998,
         mult_x_18_n997, mult_x_18_n994, mult_x_18_n993, mult_x_18_n990,
         mult_x_18_n989, mult_x_18_n986, mult_x_18_n985, mult_x_18_n982,
         mult_x_18_n981, mult_x_18_n978, mult_x_18_n977, mult_x_18_n974,
         mult_x_18_n973, mult_x_18_n969, mult_x_18_n967, mult_x_18_n965,
         mult_x_18_n964, mult_x_18_n963, mult_x_18_n961, mult_x_18_n960,
         mult_x_18_n959, mult_x_18_n958, mult_x_18_n957, mult_x_18_n956,
         mult_x_18_n955, mult_x_18_n954, mult_x_18_n953, mult_x_18_n952,
         mult_x_18_n951, mult_x_18_n950, mult_x_18_n949, mult_x_18_n948,
         mult_x_18_n947, mult_x_18_n946, mult_x_18_n945, mult_x_18_n944,
         mult_x_18_n942, mult_x_18_n941, mult_x_18_n940, mult_x_18_n939,
         mult_x_18_n938, mult_x_18_n937, mult_x_18_n936, mult_x_18_n935,
         mult_x_18_n934, mult_x_18_n933, mult_x_18_n932, mult_x_18_n931,
         mult_x_18_n930, mult_x_18_n929, mult_x_18_n928, mult_x_18_n927,
         mult_x_18_n926, mult_x_18_n925, mult_x_18_n924, mult_x_18_n923,
         mult_x_18_n922, mult_x_18_n921, mult_x_18_n920, mult_x_18_n919,
         mult_x_18_n918, mult_x_18_n917, mult_x_18_n913, mult_x_18_n912,
         mult_x_18_n911, mult_x_18_n910, mult_x_18_n909, mult_x_18_n908,
         mult_x_18_n907, mult_x_18_n906, mult_x_18_n905, mult_x_18_n904,
         mult_x_18_n903, mult_x_18_n902, mult_x_18_n901, mult_x_18_n900,
         mult_x_18_n899, mult_x_18_n898, mult_x_18_n897, mult_x_18_n896,
         mult_x_18_n895, mult_x_18_n894, mult_x_18_n893, mult_x_18_n892,
         mult_x_18_n890, mult_x_18_n889, mult_x_18_n888, mult_x_18_n886,
         mult_x_18_n884, mult_x_18_n882, mult_x_18_n881, mult_x_18_n880,
         mult_x_18_n878, mult_x_18_n877, mult_x_18_n876, mult_x_18_n874,
         mult_x_18_n873, mult_x_18_n872, mult_x_18_n871, mult_x_18_n870,
         mult_x_18_n869, mult_x_18_n866, mult_x_18_n865, mult_x_18_n864,
         mult_x_18_n863, mult_x_18_n862, mult_x_18_n861, mult_x_18_n860,
         mult_x_18_n859, mult_x_18_n858, mult_x_18_n857, mult_x_18_n856,
         mult_x_18_n855, mult_x_18_n854, mult_x_18_n853, mult_x_18_n852,
         mult_x_18_n851, mult_x_18_n850, mult_x_18_n849, mult_x_18_n848,
         mult_x_18_n846, mult_x_18_n845, mult_x_18_n844, mult_x_18_n843,
         mult_x_18_n842, mult_x_18_n841, mult_x_18_n840, mult_x_18_n839,
         mult_x_18_n838, mult_x_18_n837, mult_x_18_n836, mult_x_18_n835,
         mult_x_18_n834, mult_x_18_n833, mult_x_18_n832, mult_x_18_n831,
         mult_x_18_n830, mult_x_18_n829, mult_x_18_n825, mult_x_18_n823,
         mult_x_18_n821, mult_x_18_n819, mult_x_18_n817, mult_x_18_n815,
         mult_x_18_n814, mult_x_18_n813, mult_x_18_n812, mult_x_18_n810,
         mult_x_18_n809, mult_x_18_n808, mult_x_18_n807, mult_x_18_n806,
         mult_x_18_n805, mult_x_18_n804, mult_x_18_n803, mult_x_18_n802,
         mult_x_18_n801, mult_x_18_n800, mult_x_18_n799, mult_x_18_n798,
         mult_x_18_n797, mult_x_18_n794, mult_x_18_n793, mult_x_18_n792,
         mult_x_18_n791, mult_x_18_n790, mult_x_18_n789, mult_x_18_n788,
         mult_x_18_n787, mult_x_18_n786, mult_x_18_n785, mult_x_18_n784,
         mult_x_18_n782, mult_x_18_n781, mult_x_18_n780, mult_x_18_n778,
         mult_x_18_n777, mult_x_18_n776, mult_x_18_n774, mult_x_18_n773,
         mult_x_18_n770, mult_x_18_n769, mult_x_18_n768, mult_x_18_n767,
         mult_x_18_n766, mult_x_18_n765, mult_x_18_n764, mult_x_18_n762,
         mult_x_18_n761, mult_x_18_n760, mult_x_18_n759, mult_x_18_n758,
         mult_x_18_n757, mult_x_18_n753, mult_x_18_n752, mult_x_18_n750,
         mult_x_18_n749, mult_x_18_n744, mult_x_18_n740, mult_x_18_n738,
         mult_x_18_n736, mult_x_18_n735, mult_x_18_n734, mult_x_18_n726,
         mult_x_18_n723, mult_x_18_n722, mult_x_18_n721, mult_x_18_n720,
         mult_x_18_n719, mult_x_18_n718, mult_x_18_n717, mult_x_18_n716,
         mult_x_18_n715, mult_x_18_n714, mult_x_18_n713, mult_x_18_n712,
         mult_x_18_n711, mult_x_18_n710, mult_x_18_n709, mult_x_18_n708,
         mult_x_18_n707, mult_x_18_n706, mult_x_18_n705, mult_x_18_n704,
         mult_x_18_n703, mult_x_18_n702, mult_x_18_n701, mult_x_18_n700,
         mult_x_18_n699, mult_x_18_n698, mult_x_18_n697, mult_x_18_n696,
         mult_x_18_n695, mult_x_18_n694, mult_x_18_n693, mult_x_18_n692,
         mult_x_18_n691, mult_x_18_n690, mult_x_18_n689, mult_x_18_n688,
         mult_x_18_n687, mult_x_18_n686, mult_x_18_n685, mult_x_18_n684,
         mult_x_18_n683, mult_x_18_n682, mult_x_18_n681, mult_x_18_n680,
         mult_x_18_n679, mult_x_18_n678, mult_x_18_n677, mult_x_18_n676,
         mult_x_18_n675, mult_x_18_n674, mult_x_18_n673, mult_x_18_n672,
         mult_x_18_n671, mult_x_18_n670, mult_x_18_n669, mult_x_18_n668,
         mult_x_18_n667, mult_x_18_n666, mult_x_18_n665, mult_x_18_n664,
         mult_x_18_n663, mult_x_18_n662, mult_x_18_n661, mult_x_18_n660,
         mult_x_18_n659, mult_x_18_n658, mult_x_18_n657, mult_x_18_n656,
         mult_x_18_n655, mult_x_18_n654, mult_x_18_n653, mult_x_18_n652,
         mult_x_18_n651, mult_x_18_n650, mult_x_18_n649, mult_x_18_n648,
         mult_x_18_n647, mult_x_18_n646, mult_x_18_n645, mult_x_18_n644,
         mult_x_18_n643, mult_x_18_n642, mult_x_18_n641, mult_x_18_n640,
         mult_x_18_n639, mult_x_18_n638, mult_x_18_n637, mult_x_18_n636,
         mult_x_18_n635, mult_x_18_n634, mult_x_18_n633, mult_x_18_n632,
         mult_x_18_n631, mult_x_18_n630, mult_x_18_n629, mult_x_18_n628,
         mult_x_18_n627, mult_x_18_n626, mult_x_18_n625, mult_x_18_n624,
         mult_x_18_n623, mult_x_18_n622, mult_x_18_n621, mult_x_18_n620,
         mult_x_18_n619, mult_x_18_n618, mult_x_18_n617, mult_x_18_n616,
         mult_x_18_n615, mult_x_18_n614, mult_x_18_n613, mult_x_18_n612,
         mult_x_18_n611, mult_x_18_n610, mult_x_18_n609, mult_x_18_n608,
         mult_x_18_n607, mult_x_18_n606, mult_x_18_n605, mult_x_18_n604,
         mult_x_18_n603, mult_x_18_n602, mult_x_18_n601, mult_x_18_n600,
         mult_x_18_n599, mult_x_18_n598, mult_x_18_n597, mult_x_18_n596,
         mult_x_18_n595, mult_x_18_n594, mult_x_18_n593, mult_x_18_n592,
         mult_x_18_n591, mult_x_18_n590, mult_x_18_n589, mult_x_18_n588,
         mult_x_18_n587, mult_x_18_n586, mult_x_18_n585, mult_x_18_n584,
         mult_x_18_n583, mult_x_18_n582, mult_x_18_n581, mult_x_18_n580,
         mult_x_18_n579, mult_x_18_n578, mult_x_18_n577, mult_x_18_n576,
         mult_x_18_n575, mult_x_18_n574, mult_x_18_n573, mult_x_18_n572,
         mult_x_18_n571, mult_x_18_n570, mult_x_18_n569, mult_x_18_n568,
         mult_x_18_n567, mult_x_18_n566, mult_x_18_n565, mult_x_18_n564,
         mult_x_18_n563, mult_x_18_n562, mult_x_18_n561, mult_x_18_n560,
         mult_x_18_n559, mult_x_18_n558, mult_x_18_n557, mult_x_18_n556,
         mult_x_18_n555, mult_x_18_n554, mult_x_18_n553, mult_x_18_n552,
         mult_x_18_n551, mult_x_18_n550, mult_x_18_n549, mult_x_18_n548,
         mult_x_18_n547, mult_x_18_n546, mult_x_18_n545, mult_x_18_n544,
         mult_x_18_n543, mult_x_18_n542, mult_x_18_n541, mult_x_18_n540,
         mult_x_18_n539, mult_x_18_n538, mult_x_18_n537, mult_x_18_n536,
         mult_x_18_n535, mult_x_18_n534, mult_x_18_n533, mult_x_18_n532,
         mult_x_18_n531, mult_x_18_n530, mult_x_18_n529, mult_x_18_n528,
         mult_x_18_n527, mult_x_18_n526, mult_x_18_n525, mult_x_18_n524,
         mult_x_18_n523, mult_x_18_n522, mult_x_18_n521, mult_x_18_n520,
         mult_x_18_n519, mult_x_18_n518, mult_x_18_n517, mult_x_18_n516,
         mult_x_18_n515, mult_x_18_n514, mult_x_18_n513, mult_x_18_n512,
         mult_x_18_n511, mult_x_18_n510, mult_x_18_n509, mult_x_18_n508,
         mult_x_18_n507, mult_x_18_n506, mult_x_18_n505, mult_x_18_n504,
         mult_x_18_n503, mult_x_18_n502, mult_x_18_n501, mult_x_18_n500,
         mult_x_18_n499, mult_x_18_n498, mult_x_18_n497, mult_x_18_n496,
         mult_x_18_n495, mult_x_18_n494, mult_x_18_n493, mult_x_18_n492,
         mult_x_18_n491, mult_x_18_n490, mult_x_18_n489, mult_x_18_n488,
         mult_x_18_n487, mult_x_18_n486, mult_x_18_n485, mult_x_18_n484,
         mult_x_18_n483, mult_x_18_n482, mult_x_18_n481, mult_x_18_n480,
         mult_x_18_n479, mult_x_18_n478, mult_x_18_n477, mult_x_18_n476,
         mult_x_18_n475, mult_x_18_n474, mult_x_18_n473, mult_x_18_n472,
         mult_x_18_n471, mult_x_18_n470, mult_x_18_n469, mult_x_18_n468,
         mult_x_18_n467, mult_x_18_n466, mult_x_18_n465, mult_x_18_n464,
         mult_x_18_n463, mult_x_18_n462, mult_x_18_n461, mult_x_18_n460,
         mult_x_18_n459, mult_x_18_n458, mult_x_18_n457, mult_x_18_n456,
         mult_x_18_n455, mult_x_18_n454, mult_x_18_n453, mult_x_18_n452,
         mult_x_18_n451, mult_x_18_n450, mult_x_18_n449, mult_x_18_n448,
         mult_x_18_n447, mult_x_18_n446, mult_x_18_n445, mult_x_18_n444,
         mult_x_18_n443, mult_x_18_n442, mult_x_18_n441, mult_x_18_n440,
         mult_x_18_n439, mult_x_18_n438, mult_x_18_n437, mult_x_18_n436,
         mult_x_18_n435, mult_x_18_n434, mult_x_18_n433, mult_x_18_n432,
         mult_x_18_n431, mult_x_18_n430, mult_x_18_n429, mult_x_18_n428,
         mult_x_18_n427, mult_x_18_n426, mult_x_18_n425, mult_x_18_n424,
         mult_x_18_n423, mult_x_18_n422, mult_x_18_n421, mult_x_18_n420,
         mult_x_18_n419, mult_x_18_n418, mult_x_18_n417, mult_x_18_n416,
         mult_x_18_n415, mult_x_18_n414, mult_x_18_n413, mult_x_18_n412,
         mult_x_18_n411, mult_x_18_n410, mult_x_18_n409, mult_x_18_n408,
         mult_x_18_n407, mult_x_18_n406, mult_x_18_n405, mult_x_18_n404,
         mult_x_18_n403, mult_x_18_n402, mult_x_18_n400, mult_x_18_n399,
         mult_x_18_n398, mult_x_18_n397, mult_x_18_n396, mult_x_18_n395,
         mult_x_18_n394, mult_x_18_n393, mult_x_18_n392, mult_x_18_n391,
         mult_x_18_n390, mult_x_18_n389, mult_x_18_n388, mult_x_18_n387,
         mult_x_18_n386, mult_x_18_n385, mult_x_18_n384, mult_x_18_n383,
         mult_x_18_n382, mult_x_18_n381, mult_x_18_n380, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118;

  CMPE42D2BWP12T mult_x_18_U502 ( .A(mult_x_18_n710), .B(mult_x_18_n939), .C(
        mult_x_18_n714), .CIX(mult_x_18_n711), .D(mult_x_18_n708), .CO(
        mult_x_18_n705), .COX(mult_x_18_n704), .S(mult_x_18_n706) );
  CMPE42D2BWP12T mult_x_18_U495 ( .A(mult_x_18_n911), .B(mult_x_18_n888), .C(
        mult_x_18_n936), .CIX(mult_x_18_n693), .D(mult_x_18_n696), .CO(
        mult_x_18_n686), .COX(mult_x_18_n685), .S(mult_x_18_n687) );
  CMPE42D2BWP12T mult_x_18_U485 ( .A(mult_x_18_n933), .B(mult_x_18_n960), .C(
        mult_x_18_n989), .CIX(mult_x_18_n666), .D(mult_x_18_n662), .CO(
        mult_x_18_n659), .COX(mult_x_18_n658), .S(mult_x_18_n660) );
  CMPE42D1BWP12T mult_x_18_U509 ( .A(mult_x_18_n1029), .B(mult_x_18_n942), .C(
        mult_x_18_n969), .CIX(mult_x_18_n726), .D(mult_x_18_n998), .CO(
        mult_x_18_n722), .COX(mult_x_18_n721), .S(mult_x_18_n723) );
  CMPE42D1BWP12T U3 ( .A(mult_x_18_n671), .B(mult_x_18_n961), .C(
        mult_x_18_n668), .CIX(mult_x_18_n672), .D(mult_x_18_n676), .CO(
        mult_x_18_n664), .COX(mult_x_18_n663), .S(mult_x_18_n665) );
  OR2XD1BWP12T U4 ( .A1(mult_x_18_n692), .A2(mult_x_18_n699), .Z(n1491) );
  XNR2D1BWP12T U5 ( .A1(n2466), .A2(b[27]), .ZN(n2468) );
  XNR2D1BWP12T U6 ( .A1(n2516), .A2(b[27]), .ZN(n725) );
  INVD1BWP12T U7 ( .I(n2764), .ZN(n650) );
  OR2XD1BWP12T U8 ( .A1(mult_x_18_n674), .A2(mult_x_18_n683), .Z(n1487) );
  OAI21D1BWP12T U9 ( .A1(n786), .A2(n1280), .B(n785), .ZN(n1488) );
  ND2D1BWP12T U10 ( .A1(mult_x_18_n673), .A2(mult_x_18_n665), .ZN(n1325) );
  OR2XD1BWP12T U11 ( .A1(mult_x_18_n673), .A2(mult_x_18_n665), .Z(n1525) );
  OAI21D1BWP12T U12 ( .A1(n1459), .A2(n797), .B(n796), .ZN(n1464) );
  OAI21D1BWP12T U13 ( .A1(n782), .A2(n1497), .B(n781), .ZN(n1495) );
  OAI21D1BWP12T U14 ( .A1(n1240), .A2(n1239), .B(n1238), .ZN(n1241) );
  MUX2ND0BWP12T U15 ( .I0(n3102), .I1(n3101), .S(n2350), .ZN(n1122) );
  XOR2D2BWP12T U16 ( .A1(n991), .A2(n990), .Z(n1564) );
  XOR2D1BWP12T U17 ( .A1(n1529), .A2(n1528), .Z(n2703) );
  XOR2D1BWP12T U18 ( .A1(n1532), .A2(n1485), .Z(n2913) );
  AOI21D1BWP12T U19 ( .A1(n1492), .A2(n1491), .B(n1281), .ZN(n1285) );
  AOI21D1BWP12T U20 ( .A1(n1219), .A2(n2393), .B(n1248), .ZN(n2395) );
  OAI21D1BWP12T U21 ( .A1(n833), .A2(n832), .B(n831), .ZN(n1630) );
  NR2D1BWP12T U22 ( .A1(mult_x_18_n505), .A2(mult_x_18_n488), .ZN(n985) );
  OAI21D1BWP12T U23 ( .A1(n1558), .A2(n1552), .B(n1559), .ZN(n804) );
  HA1D0BWP12T U24 ( .A(n555), .B(n554), .CO(mult_x_18_n484), .S(mult_x_18_n485) );
  CMPE42D1BWP12T U25 ( .A(mult_x_18_n1013), .B(mult_x_18_n782), .C(
        mult_x_18_n901), .CIX(mult_x_18_n584), .D(mult_x_18_n586), .CO(
        mult_x_18_n570), .COX(mult_x_18_n569), .S(mult_x_18_n571) );
  OAI211D1BWP12T U26 ( .A1(n2975), .A2(n439), .B(n438), .C(n437), .ZN(
        result[5]) );
  AOI211D1BWP12T U27 ( .A1(n3076), .A2(n1425), .B(n436), .C(n435), .ZN(n437)
         );
  FA1D0BWP12T U28 ( .A(n2979), .B(b[31]), .CI(n2978), .CO(n2980), .S(n1645) );
  INVD2BWP12T U29 ( .I(n2169), .ZN(n2792) );
  BUFFD2BWP12T U30 ( .I(n2740), .Z(n2499) );
  XNR2D2BWP12T U31 ( .A1(n2870), .A2(n3100), .ZN(n2457) );
  CMPE42D1BWP12T U32 ( .A(mult_x_18_n575), .B(mult_x_18_n579), .C(
        mult_x_18_n562), .CIX(mult_x_18_n572), .D(mult_x_18_n576), .CO(
        mult_x_18_n558), .COX(mult_x_18_n557), .S(mult_x_18_n559) );
  CMPE42D1BWP12T U33 ( .A(mult_x_18_n548), .B(mult_x_18_n554), .C(
        mult_x_18_n561), .CIX(mult_x_18_n557), .D(mult_x_18_n545), .CO(
        mult_x_18_n541), .COX(mult_x_18_n540), .S(mult_x_18_n542) );
  INVD1BWP12T U34 ( .I(b[14]), .ZN(n2157) );
  INVD1BWP12T U35 ( .I(b[16]), .ZN(n2151) );
  INVD1BWP12T U36 ( .I(b[17]), .ZN(n2156) );
  INVD1BWP12T U37 ( .I(b[18]), .ZN(n2149) );
  INVD1BWP12T U38 ( .I(b[19]), .ZN(n2150) );
  INVD1BWP12T U39 ( .I(b[20]), .ZN(n2148) );
  INVD2BWP12T U40 ( .I(n2168), .ZN(n2876) );
  INVD1BWP12T U41 ( .I(a[12]), .ZN(n2193) );
  INVD1BWP12T U42 ( .I(a[14]), .ZN(n2192) );
  INVD1BWP12T U43 ( .I(n2738), .ZN(n2739) );
  INVD1BWP12T U44 ( .I(b[26]), .ZN(n2178) );
  INVD1BWP12T U45 ( .I(n2353), .ZN(n1104) );
  OR2XD1BWP12T U46 ( .A1(mult_x_18_n559), .A2(mult_x_18_n573), .Z(n1539) );
  NR2D1BWP12T U47 ( .A1(n985), .A2(n987), .ZN(n1549) );
  INVD1BWP12T U48 ( .I(n2353), .ZN(n2207) );
  INVD2BWP12T U49 ( .I(n358), .ZN(n2740) );
  INVD1BWP12T U50 ( .I(n2541), .ZN(n2544) );
  INVD1BWP12T U51 ( .I(n2652), .ZN(n2650) );
  CKBD1BWP12T U52 ( .I(a[16]), .Z(n2915) );
  INR2D1BWP12T U53 ( .A1(n916), .B1(n402), .ZN(n3020) );
  AOI22D1BWP12T U54 ( .A1(n382), .A2(n1725), .B1(n1645), .B2(n3082), .ZN(n930)
         );
  ND2D1BWP12T U55 ( .A1(n1918), .A2(n2353), .ZN(n1020) );
  OAI21D1BWP12T U56 ( .A1(n2110), .A2(n1050), .B(n1049), .ZN(n1247) );
  XNR2D1BWP12T U57 ( .A1(n2352), .A2(n2349), .ZN(n303) );
  NR2D1BWP12T U58 ( .A1(n1020), .A2(n2099), .ZN(n2109) );
  XNR2D1BWP12T U59 ( .A1(n2349), .A2(b[27]), .ZN(n550) );
  OAI22D1BWP12T U60 ( .A1(n2520), .A2(n655), .B1(n2518), .B2(n491), .ZN(n492)
         );
  XNR2D1BWP12T U61 ( .A1(n2350), .A2(a[13]), .ZN(n767) );
  INVD1BWP12T U62 ( .I(n2571), .ZN(n1820) );
  XNR2D1BWP12T U63 ( .A1(n2503), .A2(a[13]), .ZN(n766) );
  XNR2D1BWP12T U64 ( .A1(n2350), .A2(n2621), .ZN(n710) );
  OAI22D1BWP12T U65 ( .A1(n2459), .A2(n761), .B1(n760), .B2(n2457), .ZN(
        mult_x_18_n886) );
  OR2XD1BWP12T U66 ( .A1(n2157), .A2(a[14]), .Z(n1344) );
  OR2XD1BWP12T U67 ( .A1(n2151), .A2(n2915), .Z(n1446) );
  OAI21D1BWP12T U68 ( .A1(n1790), .A2(n872), .B(n871), .ZN(n1348) );
  MUX2ND0BWP12T U69 ( .I0(n2571), .I1(a[22]), .S(n1277), .ZN(n2233) );
  MUX2ND0BWP12T U70 ( .I0(n2898), .I1(n3100), .S(n1277), .ZN(n2237) );
  AOI21D1BWP12T U71 ( .A1(n2412), .A2(n3093), .B(n927), .ZN(n928) );
  MUX2ND0BWP12T U72 ( .I0(n3100), .I1(n2870), .S(n1277), .ZN(n2266) );
  OAI21D1BWP12T U73 ( .A1(n2350), .A2(n1262), .B(n1047), .ZN(n1897) );
  AOI21D1BWP12T U74 ( .A1(n1540), .A2(n1539), .B(n1466), .ZN(n1469) );
  XOR2D1BWP12T U75 ( .A1(n1546), .A2(n1545), .Z(n2537) );
  FA1D0BWP12T U76 ( .A(b[24]), .B(n2541), .CI(n1640), .CO(n1184), .S(n2538) );
  HA1D0BWP12T U77 ( .A(n2428), .B(n1817), .CO(n1816), .S(n2436) );
  HA1D0BWP12T U78 ( .A(n2544), .B(n1818), .CO(n1158), .S(n2556) );
  CMPE42D1BWP12T U79 ( .A(mult_x_18_n551), .B(mult_x_18_n570), .C(
        mult_x_18_n567), .CIX(mult_x_18_n560), .D(mult_x_18_n564), .CO(
        mult_x_18_n544), .COX(mult_x_18_n543), .S(mult_x_18_n545) );
  OAI21D1BWP12T U80 ( .A1(n1605), .A2(n1603), .B(n1782), .ZN(n1638) );
  OAI21D1BWP12T U81 ( .A1(n1577), .A2(n1575), .B(n1730), .ZN(n1574) );
  AOI21D1BWP12T U82 ( .A1(n1638), .A2(n1743), .B(n874), .ZN(n1592) );
  AOI21D1BWP12T U83 ( .A1(n1579), .A2(n1735), .B(n875), .ZN(n1577) );
  AOI21D1BWP12T U84 ( .A1(n1669), .A2(n1667), .B(n826), .ZN(n1665) );
  OAI21D1BWP12T U85 ( .A1(n1785), .A2(n1603), .B(n1782), .ZN(n1745) );
  AOI21D1BWP12T U86 ( .A1(n1448), .A2(n1446), .B(n826), .ZN(n1444) );
  OAI21D1BWP12T U87 ( .A1(n1592), .A2(n1590), .B(n1738), .ZN(n1579) );
  OAI21D1BWP12T U88 ( .A1(n1741), .A2(n1590), .B(n1738), .ZN(n1737) );
  OAI21D1BWP12T U89 ( .A1(n1410), .A2(n1406), .B(n1407), .ZN(n1448) );
  OAI21D1BWP12T U90 ( .A1(n1678), .A2(n1676), .B(n1677), .ZN(n1669) );
  OAI21D1BWP12T U91 ( .A1(n1665), .A2(n1661), .B(n1662), .ZN(n1660) );
  OAI21D1BWP12T U92 ( .A1(n1444), .A2(n1441), .B(n1442), .ZN(n1393) );
  AOI21D1BWP12T U93 ( .A1(n1346), .A2(n1344), .B(n856), .ZN(n1410) );
  CMPE42D1BWP12T U94 ( .A(mult_x_18_n474), .B(mult_x_18_n480), .C(
        mult_x_18_n471), .CIX(mult_x_18_n486), .D(mult_x_18_n490), .CO(
        mult_x_18_n467), .COX(mult_x_18_n466), .S(mult_x_18_n468) );
  CMPE42D1BWP12T U95 ( .A(mult_x_18_n660), .B(mult_x_18_n670), .C(
        mult_x_18_n657), .CIX(mult_x_18_n663), .D(mult_x_18_n667), .CO(
        mult_x_18_n653), .COX(mult_x_18_n652), .S(mult_x_18_n654) );
  HA1D0BWP12T U96 ( .A(n645), .B(n644), .CO(mult_x_18_n661), .S(mult_x_18_n662) );
  CMPE42D1BWP12T U97 ( .A(mult_x_18_n906), .B(mult_x_18_n958), .C(
        mult_x_18_n931), .CIX(mult_x_18_n644), .D(mult_x_18_n640), .CO(
        mult_x_18_n635), .COX(mult_x_18_n634), .S(mult_x_18_n636) );
  CMPE42D1BWP12T U98 ( .A(mult_x_18_n1021), .B(mult_x_18_n846), .C(
        mult_x_18_n990), .CIX(mult_x_18_n678), .D(mult_x_18_n680), .CO(
        mult_x_18_n670), .COX(mult_x_18_n669), .S(mult_x_18_n671) );
  CMPE42D1BWP12T U99 ( .A(mult_x_18_n837), .B(mult_x_18_n781), .C(
        mult_x_18_n856), .CIX(mult_x_18_n566), .D(mult_x_18_n900), .CO(
        mult_x_18_n550), .COX(mult_x_18_n549), .S(mult_x_18_n551) );
  CMPE42D1BWP12T U100 ( .A(mult_x_18_n679), .B(mult_x_18_n688), .C(
        mult_x_18_n682), .CIX(mult_x_18_n677), .D(mult_x_18_n686), .CO(
        mult_x_18_n673), .COX(mult_x_18_n672), .S(mult_x_18_n674) );
  CMPE42D1BWP12T U101 ( .A(mult_x_18_n689), .B(mult_x_18_n963), .C(
        mult_x_18_n690), .CIX(mult_x_18_n694), .D(mult_x_18_n687), .CO(
        mult_x_18_n683), .COX(mult_x_18_n682), .S(mult_x_18_n684) );
  CMPE42D1BWP12T U102 ( .A(mult_x_18_n635), .B(mult_x_18_n624), .C(
        mult_x_18_n632), .CIX(mult_x_18_n628), .D(mult_x_18_n621), .CO(
        mult_x_18_n617), .COX(mult_x_18_n616), .S(mult_x_18_n618) );
  CMPE42D1BWP12T U103 ( .A(mult_x_18_n648), .B(mult_x_18_n636), .C(
        mult_x_18_n645), .CIX(mult_x_18_n641), .D(mult_x_18_n633), .CO(
        mult_x_18_n629), .COX(mult_x_18_n628), .S(mult_x_18_n630) );
  CMPE42D1BWP12T U104 ( .A(mult_x_18_n940), .B(mult_x_18_n967), .C(
        mult_x_18_n719), .CIX(mult_x_18_n716), .D(mult_x_18_n715), .CO(
        mult_x_18_n712), .COX(mult_x_18_n711), .S(mult_x_18_n713) );
  CMPE42D1BWP12T U105 ( .A(mult_x_18_n938), .B(mult_x_18_n965), .C(
        mult_x_18_n994), .CIX(mult_x_18_n703), .D(mult_x_18_n704), .CO(
        mult_x_18_n699), .COX(mult_x_18_n698), .S(mult_x_18_n700) );
  HA1D0BWP12T U106 ( .A(n520), .B(n519), .CO(mult_x_18_n709), .S(
        mult_x_18_n710) );
  HA1D0BWP12T U107 ( .A(n585), .B(n584), .CO(mult_x_18_n521), .S(
        mult_x_18_n522) );
  INVD1BWP12T U108 ( .I(n1476), .ZN(n1532) );
  CMPE42D1BWP12T U109 ( .A(mult_x_18_n865), .B(mult_x_18_n886), .C(
        mult_x_18_n909), .CIX(mult_x_18_n675), .D(mult_x_18_n934), .CO(
        mult_x_18_n667), .COX(mult_x_18_n666), .S(mult_x_18_n668) );
  CMPE42D1BWP12T U110 ( .A(mult_x_18_n659), .B(mult_x_18_n649), .C(
        mult_x_18_n656), .CIX(mult_x_18_n652), .D(mult_x_18_n646), .CO(
        mult_x_18_n642), .COX(mult_x_18_n641), .S(mult_x_18_n643) );
  INVD1BWP12T U111 ( .I(n1282), .ZN(n784) );
  ND2D1BWP12T U112 ( .A1(mult_x_18_n654), .A2(mult_x_18_n664), .ZN(n1527) );
  HA1D0BWP12T U113 ( .A(n537), .B(n536), .CO(mult_x_18_n719), .S(
        mult_x_18_n720) );
  INVD1BWP12T U114 ( .I(n1563), .ZN(n984) );
  OA32D0BWP12T U115 ( .A1(n1307), .A2(n2029), .A3(n2080), .B1(n2740), .B2(
        n1307), .Z(n2391) );
  CKND0BWP12T U116 ( .I(n1790), .ZN(n1) );
  AOI21D0BWP12T U117 ( .A1(n1776), .A2(n1), .B(n1779), .ZN(n2) );
  CKND2D0BWP12T U118 ( .A1(n1777), .A2(n1778), .ZN(n3) );
  MAOI22D0BWP12T U119 ( .A1(n2), .A2(n3), .B1(n2), .B2(n3), .ZN(n3094) );
  INR3D0BWP12T U120 ( .A1(n3091), .B1(n2144), .B2(n2083), .ZN(n4) );
  OR4D0BWP12T U121 ( .A1(n2089), .A2(n2086), .A3(n2088), .A4(n2087), .Z(n5) );
  AOI211D0BWP12T U122 ( .A1(n2085), .A2(n2084), .B(n2403), .C(n5), .ZN(n6) );
  ND4D0BWP12T U123 ( .A1(n2767), .A2(n2985), .A3(n4), .A4(n6), .ZN(n7) );
  OR4D0BWP12T U124 ( .A1(n2950), .A2(n3036), .A3(n2435), .A4(n2986), .Z(n8) );
  ND4D0BWP12T U125 ( .A1(n3098), .A2(n2893), .A3(n2632), .A4(n2569), .ZN(n9)
         );
  ND4D0BWP12T U126 ( .A1(n2840), .A2(n2691), .A3(n2607), .A4(n2540), .ZN(n10)
         );
  NR4D0BWP12T U127 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n11) );
  ND4D0BWP12T U128 ( .A1(n2146), .A2(n2147), .A3(n2145), .A4(n11), .ZN(n2406)
         );
  CKND0BWP12T U129 ( .I(n1419), .ZN(n12) );
  CKND2D0BWP12T U130 ( .A1(n1418), .A2(n1430), .ZN(n13) );
  AOI32D0BWP12T U131 ( .A1(n12), .A2(n1420), .A3(n13), .B1(n1421), .B2(n1420), 
        .ZN(n14) );
  CKND2D0BWP12T U132 ( .A1(n1423), .A2(n1424), .ZN(n15) );
  MOAI22D0BWP12T U133 ( .A1(n14), .A2(n15), .B1(n14), .B2(n15), .ZN(n2800) );
  CKND2D0BWP12T U134 ( .A1(n1274), .A2(n1275), .ZN(n16) );
  MOAI22D0BWP12T U135 ( .A1(n1277), .A2(n16), .B1(n1277), .B2(n16), .ZN(n1612)
         );
  CKND0BWP12T U136 ( .I(n1711), .ZN(n17) );
  AN3D0BWP12T U137 ( .A1(n17), .A2(n1709), .A3(n1713), .Z(n18) );
  AOI211D0BWP12T U138 ( .A1(n1713), .A2(n1710), .B(n18), .C(n1295), .ZN(n19)
         );
  CKND2D0BWP12T U139 ( .A1(n286), .A2(n1296), .ZN(n20) );
  MAOI22D0BWP12T U140 ( .A1(n19), .A2(n20), .B1(n19), .B2(n20), .ZN(n1674) );
  CKND2D0BWP12T U141 ( .A1(n1490), .A2(n1491), .ZN(n21) );
  MOAI22D0BWP12T U142 ( .A1(n1492), .A2(n21), .B1(n1492), .B2(n21), .ZN(n2912)
         );
  CKND2D0BWP12T U143 ( .A1(n1113), .A2(n1109), .ZN(n22) );
  MAOI22D0BWP12T U144 ( .A1(n1114), .A2(n22), .B1(n1114), .B2(n22), .ZN(n1698)
         );
  IND3D0BWP12T U145 ( .A1(n2709), .B1(n2774), .B2(n2895), .ZN(n2379) );
  IND2D0BWP12T U146 ( .A1(n2550), .B1(n2740), .ZN(n23) );
  AOI222D0BWP12T U147 ( .A1(n23), .A2(n2118), .B1(n2932), .B2(n2929), .C1(
        n2933), .C2(n2930), .ZN(n2840) );
  OAI21D0BWP12T U148 ( .A1(n1711), .A2(n1671), .B(n1670), .ZN(n24) );
  CKND2D0BWP12T U149 ( .A1(n1439), .A2(n1673), .ZN(n25) );
  MOAI22D0BWP12T U150 ( .A1(n24), .A2(n25), .B1(n24), .B2(n25), .ZN(n3055) );
  CKND2D0BWP12T U151 ( .A1(n1776), .A2(n1778), .ZN(n26) );
  CKND2D0BWP12T U152 ( .A1(n1779), .A2(n1778), .ZN(n27) );
  OAI211D0BWP12T U153 ( .A1(n1790), .A2(n26), .B(n1777), .C(n27), .ZN(n28) );
  CKND2D0BWP12T U154 ( .A1(n1780), .A2(n1781), .ZN(n29) );
  MOAI22D0BWP12T U155 ( .A1(n28), .A2(n29), .B1(n28), .B2(n29), .ZN(n2897) );
  CKND0BWP12T U156 ( .I(n3105), .ZN(n30) );
  CKND0BWP12T U157 ( .I(n3106), .ZN(n31) );
  AOI221D0BWP12T U158 ( .A1(n3102), .A2(n31), .B1(n3101), .B2(n3106), .C(n3104), .ZN(n32) );
  AOI22D0BWP12T U159 ( .A1(n3104), .A2(n30), .B1(n3103), .B2(n32), .ZN(n33) );
  OAI21D0BWP12T U160 ( .A1(n3100), .A2(n3099), .B(n3103), .ZN(n34) );
  MOAI22D0BWP12T U161 ( .A1(n3097), .A2(n3098), .B1(n3106), .B2(n34), .ZN(n35)
         );
  AOI211D0BWP12T U162 ( .A1(n3107), .A2(n3108), .B(n33), .C(n35), .ZN(n3109)
         );
  NR4D0BWP12T U163 ( .A1(n2864), .A2(n3083), .A3(n2911), .A4(n1589), .ZN(n36)
         );
  NR4D0BWP12T U164 ( .A1(n1610), .A2(n1611), .A3(n2967), .A4(n1612), .ZN(n37)
         );
  NR4D0BWP12T U165 ( .A1(n2731), .A2(n2781), .A3(n2837), .A4(n2814), .ZN(n38)
         );
  NR4D0BWP12T U166 ( .A1(n2754), .A2(n1609), .A3(n2705), .A4(n1636), .ZN(n39)
         );
  NR3D0BWP12T U167 ( .A1(n2676), .A2(n3053), .A3(n2646), .ZN(n40) );
  ND4D0BWP12T U168 ( .A1(n37), .A2(n38), .A3(n39), .A4(n40), .ZN(n41) );
  NR4D0BWP12T U169 ( .A1(n2619), .A2(n2948), .A3(n2610), .A4(n41), .ZN(n42) );
  NR3D0BWP12T U170 ( .A1(n2538), .A2(n3043), .A3(n2567), .ZN(n43) );
  ND4D0BWP12T U171 ( .A1(n290), .A2(n36), .A3(n42), .A4(n43), .ZN(n44) );
  OR4D0BWP12T U172 ( .A1(n1643), .A2(n1641), .A3(n1642), .A4(n44), .Z(n45) );
  NR4D0BWP12T U173 ( .A1(n3008), .A2(n2423), .A3(n1644), .A4(n45), .ZN(n2417)
         );
  OAI22D0BWP12T U174 ( .A1(n1990), .A2(n1989), .B1(n1988), .B2(n2029), .ZN(n46) );
  AOI211D0BWP12T U175 ( .A1(n1985), .A2(n1984), .B(n2740), .C(n46), .ZN(n47)
         );
  OA21D0BWP12T U176 ( .A1(n1987), .A2(n1986), .B(n47), .Z(n2797) );
  OAI21D0BWP12T U177 ( .A1(n1687), .A2(n1686), .B(n1685), .ZN(n48) );
  CKND2D0BWP12T U178 ( .A1(n1690), .A2(n1689), .ZN(n49) );
  MOAI22D0BWP12T U179 ( .A1(n48), .A2(n49), .B1(n48), .B2(n49), .ZN(n2770) );
  CKND2D0BWP12T U180 ( .A1(n1413), .A2(n1414), .ZN(n50) );
  MAOI22D0BWP12T U181 ( .A1(n1437), .A2(n50), .B1(n1437), .B2(n50), .ZN(n2812)
         );
  OA21D0BWP12T U182 ( .A1(n1270), .A2(n2172), .B(n1271), .Z(n1763) );
  IOA21D0BWP12T U183 ( .A1(n2157), .A2(a[14]), .B(n1327), .ZN(n51) );
  MOAI22D0BWP12T U184 ( .A1(n1328), .A2(n51), .B1(n1328), .B2(n51), .ZN(n1675)
         );
  INR3D0BWP12T U185 ( .A1(n1848), .B1(n3100), .B2(n1846), .ZN(n52) );
  MOAI22D0BWP12T U186 ( .A1(n2898), .A2(n52), .B1(n2898), .B2(n52), .ZN(n2910)
         );
  NR4D0BWP12T U187 ( .A1(n2737), .A2(n2308), .A3(n2793), .A4(n2827), .ZN(n53)
         );
  AN4D0BWP12T U188 ( .A1(n2291), .A2(n2880), .A3(n2221), .A4(n53), .Z(n54) );
  CKND2D0BWP12T U189 ( .A1(n2292), .A2(n54), .ZN(n55) );
  OAI31D0BWP12T U190 ( .A1(n3107), .A2(n2905), .A3(n55), .B(n2402), .ZN(n56)
         );
  IND4D0BWP12T U191 ( .A1(n2718), .B1(n2426), .B2(n2245), .B3(n56), .ZN(n2299)
         );
  MOAI22D0BWP12T U192 ( .A1(n2679), .A2(b[16]), .B1(n2679), .B2(b[16]), .ZN(
        n57) );
  OAI22D0BWP12T U193 ( .A1(n2513), .A2(n2512), .B1(n2511), .B2(n57), .ZN(n2514) );
  CKND2D0BWP12T U194 ( .A1(n1761), .A2(n1629), .ZN(n58) );
  CKND0BWP12T U195 ( .I(n1757), .ZN(n59) );
  IND3D0BWP12T U196 ( .A1(n1759), .B1(n1756), .B2(n1768), .ZN(n60) );
  OAI211D0BWP12T U197 ( .A1(n1759), .A2(n59), .B(n1758), .C(n60), .ZN(n61) );
  MOAI22D0BWP12T U198 ( .A1(n58), .A2(n61), .B1(n58), .B2(n61), .ZN(n2828) );
  AN4D0BWP12T U199 ( .A1(n2684), .A2(n2797), .A3(n2922), .A4(n2401), .Z(n62)
         );
  ND4D0BWP12T U200 ( .A1(n2741), .A2(n2010), .A3(n2631), .A4(n62), .ZN(n63) );
  NR3D0BWP12T U201 ( .A1(n2810), .A2(n2399), .A3(n63), .ZN(n64) );
  NR4D0BWP12T U202 ( .A1(n2883), .A2(n2648), .A3(n2042), .A4(n2041), .ZN(n65)
         );
  IAO21D0BWP12T U203 ( .A1(n2740), .A2(n3112), .B(n2706), .ZN(n66) );
  ND4D0BWP12T U204 ( .A1(n2734), .A2(n2016), .A3(n2017), .A4(n66), .ZN(n67) );
  NR4D0BWP12T U205 ( .A1(n3052), .A2(n2031), .A3(n2379), .A4(n67), .ZN(n68) );
  OAI211D0BWP12T U206 ( .A1(n2740), .A2(n64), .B(n65), .C(n68), .ZN(n2407) );
  CKND2D0BWP12T U207 ( .A1(n1432), .A2(n1701), .ZN(n69) );
  IOA21D0BWP12T U208 ( .A1(n1430), .A2(n1690), .B(n1429), .ZN(n70) );
  MOAI22D0BWP12T U209 ( .A1(n69), .A2(n70), .B1(n69), .B2(n70), .ZN(n2729) );
  IND2D0BWP12T U210 ( .A1(op[0]), .B1(n415), .ZN(n392) );
  CKND2D0BWP12T U211 ( .A1(n1773), .A2(n1583), .ZN(n71) );
  IOA21D0BWP12T U212 ( .A1(n1771), .A2(n1633), .B(n1770), .ZN(n72) );
  MOAI22D0BWP12T U213 ( .A1(n71), .A2(n72), .B1(n71), .B2(n72), .ZN(n2869) );
  CKND2D0BWP12T U214 ( .A1(n1685), .A2(n1225), .ZN(n73) );
  MAOI22D0BWP12T U215 ( .A1(n1687), .A2(n73), .B1(n1687), .B2(n73), .ZN(n1699)
         );
  OR4D0BWP12T U216 ( .A1(n2868), .A2(n2783), .A3(n2384), .A4(n2856), .Z(n74)
         );
  CKND2D0BWP12T U217 ( .A1(n2386), .A2(n2387), .ZN(n75) );
  OAI211D0BWP12T U218 ( .A1(n2390), .A2(n2389), .B(n2855), .C(n75), .ZN(n76)
         );
  NR4D0BWP12T U219 ( .A1(n2835), .A2(n3081), .A3(n74), .A4(n76), .ZN(n77) );
  CKND2D0BWP12T U220 ( .A1(n3064), .A2(n2391), .ZN(n78) );
  AOI211D0BWP12T U221 ( .A1(n2396), .A2(n78), .B(n2736), .C(n2395), .ZN(n79)
         );
  OAI31D0BWP12T U222 ( .A1(n2708), .A2(n2380), .A3(n2379), .B(n2396), .ZN(n80)
         );
  IND4D0BWP12T U223 ( .A1(n2399), .B1(n2400), .B2(n2659), .B3(n2401), .ZN(n81)
         );
  IND4D0BWP12T U224 ( .A1(n2397), .B1(n2631), .B2(n2684), .B3(n2922), .ZN(n82)
         );
  OAI31D0BWP12T U225 ( .A1(n2403), .A2(n81), .A3(n82), .B(n2402), .ZN(n83) );
  ND4D0BWP12T U226 ( .A1(n77), .A2(n79), .A3(n80), .A4(n83), .ZN(n2404) );
  AOI21D0BWP12T U227 ( .A1(n1616), .A2(n1624), .B(n1618), .ZN(n84) );
  CKND2D0BWP12T U228 ( .A1(n1619), .A2(n414), .ZN(n85) );
  MAOI22D0BWP12T U229 ( .A1(n84), .A2(n85), .B1(n84), .B2(n85), .ZN(n1609) );
  CKND2D0BWP12T U230 ( .A1(n1279), .A2(n1275), .ZN(n86) );
  MOAI22D0BWP12T U231 ( .A1(n1269), .A2(n86), .B1(n1269), .B2(n86), .ZN(n1426)
         );
  CKND0BWP12T U232 ( .I(n1711), .ZN(n87) );
  AOI21D0BWP12T U233 ( .A1(n1709), .A2(n87), .B(n1710), .ZN(n88) );
  CKND2D0BWP12T U234 ( .A1(n1712), .A2(n1713), .ZN(n89) );
  MAOI22D0BWP12T U235 ( .A1(n88), .A2(n89), .B1(n88), .B2(n89), .ZN(n2890) );
  INR3D0BWP12T U236 ( .A1(n2787), .B1(n1849), .B2(n1850), .ZN(n90) );
  MOAI22D0BWP12T U237 ( .A1(n2815), .A2(n90), .B1(n2815), .B2(n90), .ZN(n2834)
         );
  OAI22D0BWP12T U238 ( .A1(n2449), .A2(n2448), .B1(n2450), .B2(n719), .ZN(n91)
         );
  IND2D0BWP12T U239 ( .A1(n1277), .B1(n2979), .ZN(n92) );
  OAI22D0BWP12T U240 ( .A1(n2504), .A2(n92), .B1(n2216), .B2(n2506), .ZN(n93)
         );
  MAOI22D0BWP12T U241 ( .A1(n91), .A2(n93), .B1(n91), .B2(n93), .ZN(
        mult_x_18_n402) );
  AN2D0BWP12T U242 ( .A1(n91), .A2(n93), .Z(n2486) );
  CKND2D0BWP12T U243 ( .A1(n858), .A2(n414), .ZN(n94) );
  IOA21D0BWP12T U244 ( .A1(n1768), .A2(n1767), .B(n1766), .ZN(n95) );
  MOAI22D0BWP12T U245 ( .A1(n94), .A2(n95), .B1(n94), .B2(n95), .ZN(n1774) );
  OAI22D0BWP12T U246 ( .A1(n1884), .A2(n2029), .B1(n1955), .B2(n1989), .ZN(n96) );
  AOI211D0BWP12T U247 ( .A1(n1984), .A2(n1952), .B(n2740), .C(n96), .ZN(n97)
         );
  OAI21D0BWP12T U248 ( .A1(n1956), .A2(n1986), .B(n97), .ZN(n2015) );
  CKND2D0BWP12T U249 ( .A1(n1581), .A2(n1583), .ZN(n98) );
  CKND2D0BWP12T U250 ( .A1(n1584), .A2(n1583), .ZN(n99) );
  OAI211D0BWP12T U251 ( .A1(n1607), .A2(n98), .B(n1582), .C(n99), .ZN(n100) );
  CKND2D0BWP12T U252 ( .A1(n1586), .A2(n1778), .ZN(n101) );
  MOAI22D0BWP12T U253 ( .A1(n100), .A2(n101), .B1(n100), .B2(n101), .ZN(n3083)
         );
  IND2D0BWP12T U254 ( .A1(n1650), .B1(n1651), .ZN(n102) );
  MAOI22D0BWP12T U255 ( .A1(n1652), .A2(n102), .B1(n1652), .B2(n102), .ZN(
        n2592) );
  OAI21D0BWP12T U256 ( .A1(n1437), .A2(n1403), .B(n1402), .ZN(n103) );
  CKND2D0BWP12T U257 ( .A1(n1713), .A2(n1404), .ZN(n104) );
  MOAI22D0BWP12T U258 ( .A1(n103), .A2(n104), .B1(n103), .B2(n104), .ZN(n2891)
         );
  AOI21D0BWP12T U259 ( .A1(n1521), .A2(n1520), .B(n1498), .ZN(n105) );
  CKND2D0BWP12T U260 ( .A1(n288), .A2(n1496), .ZN(n106) );
  MAOI22D0BWP12T U261 ( .A1(n105), .A2(n106), .B1(n105), .B2(n106), .ZN(n2889)
         );
  CKND2D0BWP12T U262 ( .A1(n1696), .A2(n1414), .ZN(n107) );
  AOI21D0BWP12T U263 ( .A1(n1691), .A2(n1703), .B(n1692), .ZN(n108) );
  OAI21D0BWP12T U264 ( .A1(n1694), .A2(n108), .B(n1693), .ZN(n109) );
  MOAI22D0BWP12T U265 ( .A1(n107), .A2(n109), .B1(n107), .B2(n109), .ZN(n2811)
         );
  NR2D0BWP12T U266 ( .A1(n2879), .A2(n2221), .ZN(n110) );
  AOI22D0BWP12T U267 ( .A1(n2087), .A2(n3090), .B1(n3076), .B2(n1426), .ZN(
        n111) );
  MUX2ND0BWP12T U268 ( .I0(n3102), .I1(n3101), .S(n1277), .ZN(n112) );
  AOI31D0BWP12T U269 ( .A1(n3103), .A2(n112), .A3(n3040), .B(n2449), .ZN(n113)
         );
  OAI22D0BWP12T U270 ( .A1(n2172), .A2(n3023), .B1(n2368), .B2(n3103), .ZN(
        n114) );
  AOI211D0BWP12T U271 ( .A1(n1272), .A2(n2208), .B(n113), .C(n114), .ZN(n115)
         );
  CKND0BWP12T U272 ( .I(n2975), .ZN(n116) );
  AOI22D0BWP12T U273 ( .A1(n3093), .A2(n1763), .B1(n1515), .B2(n116), .ZN(n117) );
  CKND0BWP12T U274 ( .I(n3004), .ZN(n118) );
  AOI22D0BWP12T U275 ( .A1(n1697), .A2(n382), .B1(n2088), .B2(n118), .ZN(n119)
         );
  ND4D0BWP12T U276 ( .A1(n111), .A2(n115), .A3(n117), .A4(n119), .ZN(n120) );
  AOI211D0BWP12T U277 ( .A1(n3082), .A2(n1612), .B(n110), .C(n120), .ZN(n121)
         );
  OAI21D0BWP12T U278 ( .A1(n1976), .A2(n2384), .B(n3084), .ZN(n122) );
  OAI211D0BWP12T U279 ( .A1(n1979), .A2(n2856), .B(n121), .C(n122), .ZN(
        result[0]) );
  MOAI22D0BWP12T U280 ( .A1(n2815), .A2(b[26]), .B1(n2815), .B2(b[26]), .ZN(
        n123) );
  OAI22D0BWP12T U281 ( .A1(n2510), .A2(n2509), .B1(n2508), .B2(n123), .ZN(
        n2515) );
  IAO21D0BWP12T U282 ( .A1(n650), .A2(n380), .B(n1431), .ZN(n1418) );
  OAI21D0BWP12T U283 ( .A1(n1222), .A2(n1221), .B(n1220), .ZN(n124) );
  CKND2D0BWP12T U284 ( .A1(n1225), .A2(n1224), .ZN(n125) );
  MOAI22D0BWP12T U285 ( .A1(n124), .A2(n125), .B1(n124), .B2(n125), .ZN(n1428)
         );
  OAI21D0BWP12T U286 ( .A1(n1790), .A2(n1786), .B(n1787), .ZN(n126) );
  AOI21D0BWP12T U287 ( .A1(n1789), .A2(n126), .B(n1788), .ZN(n127) );
  IOA21D0BWP12T U288 ( .A1(a[13]), .A2(b[13]), .B(n1791), .ZN(n128) );
  MAOI22D0BWP12T U289 ( .A1(n127), .A2(n128), .B1(n127), .B2(n128), .ZN(n3056)
         );
  CKND2D0BWP12T U290 ( .A1(n1838), .A2(n1848), .ZN(n129) );
  MAOI22D0BWP12T U291 ( .A1(a[12]), .A2(n129), .B1(a[12]), .B2(n129), .ZN(
        n1847) );
  OAI21D0BWP12T U292 ( .A1(n1607), .A2(n1588), .B(n1587), .ZN(n130) );
  CKND2D0BWP12T U293 ( .A1(n1781), .A2(n1780), .ZN(n131) );
  MOAI22D0BWP12T U294 ( .A1(n130), .A2(n131), .B1(n130), .B2(n131), .ZN(n2911)
         );
  CKND2D0BWP12T U295 ( .A1(n1493), .A2(n1494), .ZN(n132) );
  MOAI22D0BWP12T U296 ( .A1(n1495), .A2(n132), .B1(n1495), .B2(n132), .ZN(
        n3118) );
  OAI21D0BWP12T U297 ( .A1(n1970), .A2(n1949), .B(n2377), .ZN(n133) );
  IAO21D0BWP12T U298 ( .A1(n2029), .A2(n1950), .B(n133), .ZN(n134) );
  OAI21D0BWP12T U299 ( .A1(n1964), .A2(n2314), .B(n134), .ZN(n2810) );
  OR4D0BWP12T U300 ( .A1(n1675), .A2(n1674), .A3(n3115), .A4(n2890), .Z(n135)
         );
  NR4D0BWP12T U301 ( .A1(n3055), .A2(n2725), .A3(n1714), .A4(n135), .ZN(n136)
         );
  NR3D0BWP12T U302 ( .A1(n2699), .A2(n2943), .A3(n2671), .ZN(n137) );
  NR3D0BWP12T U303 ( .A1(n2641), .A2(n2592), .A3(n2971), .ZN(n138) );
  NR4D0BWP12T U304 ( .A1(n2587), .A2(n1721), .A3(n2561), .A4(n3016), .ZN(n139)
         );
  ND4D0BWP12T U305 ( .A1(n136), .A2(n137), .A3(n138), .A4(n139), .ZN(n140) );
  OR4D0BWP12T U306 ( .A1(n1723), .A2(n1722), .A3(n1724), .A4(n140), .Z(n141)
         );
  NR4D0BWP12T U307 ( .A1(n2984), .A2(n1725), .A3(n2442), .A4(n141), .ZN(n2415)
         );
  MOAI22D0BWP12T U308 ( .A1(n2870), .A2(b[24]), .B1(n2870), .B2(b[24]), .ZN(
        n142) );
  OAI22D0BWP12T U309 ( .A1(n2489), .A2(n2488), .B1(n2487), .B2(n142), .ZN(n143) );
  MOAI22D0BWP12T U310 ( .A1(n2571), .A2(n3106), .B1(n2571), .B2(n3106), .ZN(
        n144) );
  OAI22D0BWP12T U311 ( .A1(n2492), .A2(n2491), .B1(n2490), .B2(n144), .ZN(n145) );
  MAOI22D0BWP12T U312 ( .A1(n143), .A2(n145), .B1(n143), .B2(n145), .ZN(n2497)
         );
  CKND2D0BWP12T U313 ( .A1(n1770), .A2(n1633), .ZN(n146) );
  MAOI22D0BWP12T U314 ( .A1(n1790), .A2(n146), .B1(n1790), .B2(n146), .ZN(
        n2838) );
  CKND2D0BWP12T U315 ( .A1(n1766), .A2(n1767), .ZN(n147) );
  IOA21D0BWP12T U316 ( .A1(n1624), .A2(n1614), .B(n1613), .ZN(n148) );
  MOAI22D0BWP12T U317 ( .A1(n147), .A2(n148), .B1(n147), .B2(n148), .ZN(n2731)
         );
  MAOI22D0BWP12T U318 ( .A1(n2465), .A2(n2464), .B1(n2465), .B2(n2464), .ZN(
        n149) );
  MAOI22D0BWP12T U319 ( .A1(n2451), .A2(n149), .B1(n2451), .B2(n149), .ZN(n150) );
  MAOI22D0BWP12T U320 ( .A1(mult_x_18_n398), .A2(n150), .B1(mult_x_18_n398), 
        .B2(n150), .ZN(n151) );
  MAOI22D0BWP12T U321 ( .A1(mult_x_18_n393), .A2(mult_x_18_n396), .B1(
        mult_x_18_n393), .B2(mult_x_18_n396), .ZN(n152) );
  OAI22D0BWP12T U322 ( .A1(n2482), .A2(n2481), .B1(n2484), .B2(n2483), .ZN(
        n153) );
  MAOI22D0BWP12T U323 ( .A1(n2485), .A2(n153), .B1(n2485), .B2(n153), .ZN(n154) );
  MAOI22D0BWP12T U324 ( .A1(n2470), .A2(n154), .B1(n2470), .B2(n154), .ZN(n155) );
  MAOI22D0BWP12T U325 ( .A1(mult_x_18_n395), .A2(n155), .B1(mult_x_18_n395), 
        .B2(n155), .ZN(n156) );
  MAOI22D0BWP12T U326 ( .A1(n152), .A2(n156), .B1(n152), .B2(n156), .ZN(n157)
         );
  MAOI22D0BWP12T U327 ( .A1(n151), .A2(n157), .B1(n151), .B2(n157), .ZN(n158)
         );
  MAOI22D0BWP12T U328 ( .A1(mult_x_18_n386), .A2(n158), .B1(mult_x_18_n386), 
        .B2(n158), .ZN(n159) );
  MAOI22D0BWP12T U329 ( .A1(mult_x_18_n380), .A2(n159), .B1(mult_x_18_n380), 
        .B2(n159), .ZN(n2522) );
  INR2D0BWP12T U330 ( .A1(n1433), .B1(n1437), .ZN(n160) );
  OAI32D0BWP12T U331 ( .A1(n1434), .A2(n160), .A3(n1436), .B1(n1435), .B2(
        n1434), .ZN(n161) );
  CKND2D0BWP12T U332 ( .A1(n1439), .A2(n1438), .ZN(n162) );
  MAOI22D0BWP12T U333 ( .A1(n161), .A2(n162), .B1(n161), .B2(n162), .ZN(n3075)
         );
  IAO21D0BWP12T U334 ( .A1(n2432), .A2(n1989), .B(n419), .ZN(n2600) );
  OAI21D0BWP12T U335 ( .A1(n1711), .A2(n1706), .B(n1705), .ZN(n163) );
  CKND2D0BWP12T U336 ( .A1(n1401), .A2(n1708), .ZN(n164) );
  MOAI22D0BWP12T U337 ( .A1(n163), .A2(n164), .B1(n163), .B2(n164), .ZN(n3115)
         );
  CKND2D0BWP12T U338 ( .A1(n2848), .A2(n1848), .ZN(n165) );
  MAOI22D0BWP12T U339 ( .A1(n2870), .A2(n165), .B1(n2870), .B2(n165), .ZN(
        n2863) );
  IND2D0BWP12T U340 ( .A1(n776), .B1(n775), .ZN(n166) );
  MAOI22D0BWP12T U341 ( .A1(n777), .A2(n166), .B1(n777), .B2(n166), .ZN(n1517)
         );
  CKND0BWP12T U342 ( .I(n3076), .ZN(n167) );
  CKND0BWP12T U343 ( .I(n382), .ZN(n168) );
  OAI22D0BWP12T U344 ( .A1(n2526), .A2(n167), .B1(n2528), .B2(n168), .ZN(n2981) );
  AO222D0BWP12T U345 ( .A1(n2911), .A2(n3082), .B1(n3076), .B2(n2891), .C1(
        n2890), .C2(n382), .Z(n169) );
  AO211D0BWP12T U346 ( .A1(n2910), .A2(n3096), .B(n2909), .C(n169), .Z(n170)
         );
  AOI211D0BWP12T U347 ( .A1(n3093), .A2(n2897), .B(n2896), .C(n170), .ZN(n171)
         );
  IOA21D0BWP12T U348 ( .A1(n2912), .A2(n3117), .B(n171), .ZN(result[11]) );
  MOAI22D0BWP12T U349 ( .A1(n2134), .A2(n2014), .B1(n2134), .B2(n2053), .ZN(
        n172) );
  OAI21D0BWP12T U350 ( .A1(n2130), .A2(n172), .B(n2391), .ZN(n2031) );
  AOI222D0BWP12T U351 ( .A1(a[3]), .A2(n1923), .B1(n1925), .B2(n2349), .C1(
        n2352), .C2(n1924), .ZN(n173) );
  OAI22D0BWP12T U352 ( .A1(n1955), .A2(n1986), .B1(n1884), .B2(n1970), .ZN(
        n174) );
  AOI211D0BWP12T U353 ( .A1(n2076), .A2(n1952), .B(n1276), .C(n174), .ZN(n175)
         );
  OAI21D0BWP12T U354 ( .A1(n2764), .A2(n173), .B(n175), .ZN(n2087) );
  CKND0BWP12T U355 ( .I(n1437), .ZN(n176) );
  AOI21D0BWP12T U356 ( .A1(n1395), .A2(n176), .B(n1398), .ZN(n177) );
  CKND2D0BWP12T U357 ( .A1(n1396), .A2(n1397), .ZN(n178) );
  MAOI22D0BWP12T U358 ( .A1(n177), .A2(n178), .B1(n177), .B2(n178), .ZN(n2867)
         );
  AOI21D0BWP12T U359 ( .A1(n1691), .A2(n1703), .B(n1692), .ZN(n179) );
  CKND2D0BWP12T U360 ( .A1(n1693), .A2(n1424), .ZN(n180) );
  MAOI22D0BWP12T U361 ( .A1(n179), .A2(n180), .B1(n179), .B2(n180), .ZN(n2778)
         );
  NR2D0BWP12T U362 ( .A1(n2738), .A2(n1850), .ZN(n181) );
  MOAI22D0BWP12T U363 ( .A1(n2466), .A2(n181), .B1(n2466), .B2(n181), .ZN(
        n1852) );
  CKND2D0BWP12T U364 ( .A1(n1509), .A2(n1508), .ZN(n182) );
  MOAI22D0BWP12T U365 ( .A1(n1510), .A2(n182), .B1(n1510), .B2(n182), .ZN(
        n2749) );
  MAOI22D0BWP12T U366 ( .A1(n2522), .A2(n2521), .B1(n2522), .B2(n2521), .ZN(
        n183) );
  MAOI22D0BWP12T U367 ( .A1(n183), .A2(mult_x_18_n381), .B1(n183), .B2(
        mult_x_18_n381), .ZN(n184) );
  MAOI22D1BWP12T U368 ( .A1(n2523), .A2(n184), .B1(n2523), .B2(n184), .ZN(
        n2983) );
  AOI22D0BWP12T U369 ( .A1(n2809), .A2(n2810), .B1(n382), .B2(n2811), .ZN(n185) );
  AOI211D0BWP12T U370 ( .A1(n2834), .A2(n3096), .B(n2833), .C(n2832), .ZN(n186) );
  AOI22D0BWP12T U371 ( .A1(n3117), .A2(n2806), .B1(n3080), .B2(n2835), .ZN(
        n187) );
  ND3D0BWP12T U372 ( .A1(n185), .A2(n186), .A3(n187), .ZN(result[7]) );
  OA32D0BWP12T U373 ( .A1(n2028), .A2(n2029), .A3(n2432), .B1(n2740), .B2(
        n2028), .Z(n3064) );
  CKND2D0BWP12T U374 ( .A1(n1766), .A2(n1767), .ZN(n188) );
  MOAI22D0BWP12T U375 ( .A1(n1768), .A2(n188), .B1(n1768), .B2(n188), .ZN(
        n2730) );
  IAO21D0BWP12T U376 ( .A1(n1103), .A2(n1102), .B(n1213), .ZN(n1516) );
  NR4D0BWP12T U377 ( .A1(n1699), .A2(n1698), .A3(n1697), .A4(n3047), .ZN(n189)
         );
  NR3D0BWP12T U378 ( .A1(n2770), .A2(n2811), .A3(n2778), .ZN(n190) );
  NR3D0BWP12T U379 ( .A1(n1704), .A2(n2859), .A3(n2882), .ZN(n191) );
  ND4D0BWP12T U380 ( .A1(n292), .A2(n189), .A3(n190), .A4(n191), .ZN(n1714) );
  CKND2D0BWP12T U381 ( .A1(n1395), .A2(n1397), .ZN(n192) );
  CKND2D0BWP12T U382 ( .A1(n1398), .A2(n1397), .ZN(n193) );
  OAI211D0BWP12T U383 ( .A1(n1437), .A2(n192), .B(n1396), .C(n193), .ZN(n194)
         );
  CKND2D0BWP12T U384 ( .A1(n1400), .A2(n1401), .ZN(n195) );
  MOAI22D0BWP12T U385 ( .A1(n194), .A2(n195), .B1(n194), .B2(n195), .ZN(n3079)
         );
  OAI22D0BWP12T U386 ( .A1(n1918), .A2(n2544), .B1(n1919), .B2(n2202), .ZN(
        n196) );
  AOI21D0BWP12T U387 ( .A1(n2350), .A2(n1262), .B(n196), .ZN(n1941) );
  IND2D0BWP12T U388 ( .A1(n416), .B1(n400), .ZN(n3040) );
  MOAI22D0BWP12T U389 ( .A1(n2594), .A2(n2452), .B1(n2594), .B2(n2452), .ZN(
        n197) );
  OAI22D0BWP12T U390 ( .A1(n2455), .A2(n2454), .B1(n2453), .B2(n197), .ZN(n198) );
  MOAI22D0BWP12T U391 ( .A1(n2456), .A2(b[22]), .B1(n2456), .B2(b[22]), .ZN(
        n199) );
  OAI22D0BWP12T U392 ( .A1(n2459), .A2(n2458), .B1(n2457), .B2(n199), .ZN(n200) );
  MAOI22D0BWP12T U393 ( .A1(n198), .A2(n200), .B1(n198), .B2(n200), .ZN(n2465)
         );
  OA222D0BWP12T U394 ( .A1(n1972), .A2(n1986), .B1(n1971), .B2(n1970), .C1(
        n1973), .C2(n1989), .Z(n201) );
  OA211D0BWP12T U395 ( .A1(n1974), .A2(n2029), .B(n2377), .C(n201), .Z(n2028)
         );
  NR4D0BWP12T U396 ( .A1(n3056), .A2(n1792), .A3(n1793), .A4(n2704), .ZN(n202)
         );
  NR4D0BWP12T U397 ( .A1(n1765), .A2(n1764), .A3(n1763), .A4(n1762), .ZN(n203)
         );
  NR4D0BWP12T U398 ( .A1(n2730), .A2(n2758), .A3(n2780), .A4(n2828), .ZN(n204)
         );
  CKND2D0BWP12T U399 ( .A1(n203), .A2(n204), .ZN(n205) );
  NR4D0BWP12T U400 ( .A1(n1774), .A2(n2869), .A3(n2838), .A4(n205), .ZN(n206)
         );
  NR4D0BWP12T U401 ( .A1(n3094), .A2(n2677), .A3(n2897), .A4(n2914), .ZN(n207)
         );
  NR3D0BWP12T U402 ( .A1(n2620), .A2(n2949), .A3(n2647), .ZN(n208) );
  ND4D0BWP12T U403 ( .A1(n202), .A2(n206), .A3(n207), .A4(n208), .ZN(n1799) );
  CKND2D0BWP12T U404 ( .A1(n1417), .A2(n1681), .ZN(n209) );
  IOA21D0BWP12T U405 ( .A1(n1415), .A2(n1414), .B(n1413), .ZN(n210) );
  MOAI22D0BWP12T U406 ( .A1(n209), .A2(n210), .B1(n209), .B2(n210), .ZN(n2843)
         );
  MAOI22D0BWP12T U407 ( .A1(n2497), .A2(n2496), .B1(n2497), .B2(n2496), .ZN(
        n211) );
  MAOI22D0BWP12T U408 ( .A1(n2486), .A2(n211), .B1(n2486), .B2(n211), .ZN(n212) );
  MAOI22D0BWP12T U409 ( .A1(mult_x_18_n392), .A2(n212), .B1(mult_x_18_n392), 
        .B2(n212), .ZN(n213) );
  MAOI22D0BWP12T U410 ( .A1(mult_x_18_n383), .A2(n213), .B1(mult_x_18_n383), 
        .B2(n213), .ZN(n214) );
  MAOI22D0BWP12T U411 ( .A1(mult_x_18_n389), .A2(n2507), .B1(mult_x_18_n389), 
        .B2(n2507), .ZN(n215) );
  MAOI22D0BWP12T U412 ( .A1(n2515), .A2(n2514), .B1(n2515), .B2(n2514), .ZN(
        n216) );
  OAI22D0BWP12T U413 ( .A1(n2518), .A2(n2517), .B1(n2520), .B2(n2519), .ZN(
        n217) );
  MAOI22D0BWP12T U414 ( .A1(n216), .A2(n217), .B1(n216), .B2(n217), .ZN(n218)
         );
  MAOI22D0BWP12T U415 ( .A1(n215), .A2(n218), .B1(n215), .B2(n218), .ZN(n219)
         );
  MAOI22D0BWP12T U416 ( .A1(mult_x_18_n399), .A2(n219), .B1(mult_x_18_n399), 
        .B2(n219), .ZN(n220) );
  MAOI22D0BWP12T U417 ( .A1(mult_x_18_n390), .A2(n220), .B1(mult_x_18_n390), 
        .B2(n220), .ZN(n221) );
  MAOI22D0BWP12T U418 ( .A1(n214), .A2(n221), .B1(n214), .B2(n221), .ZN(n222)
         );
  MAOI22D0BWP12T U419 ( .A1(mult_x_18_n387), .A2(n222), .B1(mult_x_18_n387), 
        .B2(n222), .ZN(n223) );
  MAOI22D0BWP12T U420 ( .A1(mult_x_18_n384), .A2(n223), .B1(mult_x_18_n384), 
        .B2(n223), .ZN(n2521) );
  CKND0BWP12T U421 ( .I(n2810), .ZN(n224) );
  CKND0BWP12T U422 ( .I(n2396), .ZN(n225) );
  OAI32D0BWP12T U423 ( .A1(n224), .A2(n2808), .A3(n225), .B1(n2393), .B2(n224), 
        .ZN(n2835) );
  IND2D0BWP12T U424 ( .A1(n1511), .B1(n1512), .ZN(n226) );
  MAOI22D0BWP12T U425 ( .A1(n1513), .A2(n226), .B1(n1513), .B2(n226), .ZN(
        n2776) );
  INVD1BWP12T U426 ( .I(a[11]), .ZN(n2900) );
  INR3D0BWP12T U427 ( .A1(op[0]), .B1(op[1]), .B2(n433), .ZN(n3082) );
  CKND2D0BWP12T U428 ( .A1(n1519), .A2(n1520), .ZN(n227) );
  MOAI22D0BWP12T U429 ( .A1(n1521), .A2(n227), .B1(n1521), .B2(n227), .ZN(
        n2836) );
  CKND2D0BWP12T U430 ( .A1(n1684), .A2(n1397), .ZN(n228) );
  IOA21D0BWP12T U431 ( .A1(n1682), .A2(n1681), .B(n1680), .ZN(n229) );
  MOAI22D0BWP12T U432 ( .A1(n228), .A2(n229), .B1(n228), .B2(n229), .ZN(n2882)
         );
  AOI21D0BWP12T U433 ( .A1(n1418), .A2(n1430), .B(n1419), .ZN(n230) );
  CKND2D0BWP12T U434 ( .A1(n1420), .A2(n389), .ZN(n231) );
  MAOI22D0BWP12T U435 ( .A1(n230), .A2(n231), .B1(n230), .B2(n231), .ZN(n1425)
         );
  AOI21D0BWP12T U436 ( .A1(n2740), .A2(n3101), .B(n3020), .ZN(n232) );
  OAI21D0BWP12T U437 ( .A1(n3019), .A2(n2740), .B(n232), .ZN(n233) );
  MOAI22D0BWP12T U438 ( .A1(n2739), .A2(n233), .B1(n2739), .B2(n3023), .ZN(
        n234) );
  OAI21D0BWP12T U439 ( .A1(n2738), .A2(n3099), .B(n3103), .ZN(n235) );
  AOI22D0BWP12T U440 ( .A1(n2826), .A2(n2737), .B1(n2740), .B2(n235), .ZN(n236) );
  OAI211D0BWP12T U441 ( .A1(n2807), .A2(n2741), .B(n234), .C(n236), .ZN(n2742)
         );
  INR3D0BWP12T U442 ( .A1(n1838), .B1(n1364), .B2(n1363), .ZN(n1851) );
  NR2D0BWP12T U443 ( .A1(n2982), .A2(n2533), .ZN(n237) );
  AOI211D0BWP12T U444 ( .A1(n2982), .A2(n2533), .B(n3040), .C(n237), .ZN(n2534) );
  IAO21D0BWP12T U445 ( .A1(n1277), .A2(n2349), .B(n2208), .ZN(n1111) );
  OA21D0BWP12T U446 ( .A1(n2074), .A2(n2073), .B(n2072), .Z(n2808) );
  MOAI22D0BWP12T U447 ( .A1(n2460), .A2(n2852), .B1(n2460), .B2(n2852), .ZN(
        n238) );
  OAI22D0BWP12T U448 ( .A1(n2463), .A2(n2462), .B1(n2461), .B2(n238), .ZN(
        n2464) );
  MOAI22D0BWP12T U449 ( .A1(n2498), .A2(n2499), .B1(n2498), .B2(n2499), .ZN(
        n239) );
  OAI22D0BWP12T U450 ( .A1(n2502), .A2(n2501), .B1(n2500), .B2(n239), .ZN(n240) );
  MOAI22D0BWP12T U451 ( .A1(n2979), .A2(n2503), .B1(n2979), .B2(n2503), .ZN(
        n241) );
  OAI22D0BWP12T U452 ( .A1(n2506), .A2(n2505), .B1(n2504), .B2(n241), .ZN(n242) );
  MOAI22D0BWP12T U453 ( .A1(n240), .A2(n242), .B1(n240), .B2(n242), .ZN(n2507)
         );
  NR4D0BWP12T U454 ( .A1(b[19]), .A2(b[18]), .A3(b[21]), .A4(b[20]), .ZN(n243)
         );
  ND3D1BWP12T U455 ( .A1(n364), .A2(n365), .A3(n243), .ZN(n372) );
  CKND2D0BWP12T U456 ( .A1(n1627), .A2(n1629), .ZN(n244) );
  MAOI22D0BWP12T U457 ( .A1(n1607), .A2(n244), .B1(n1607), .B2(n244), .ZN(
        n2814) );
  AOI22D0BWP12T U458 ( .A1(n3093), .A2(n1792), .B1(n3076), .B2(n1440), .ZN(
        n245) );
  IND2D0BWP12T U459 ( .A1(n3065), .B1(n2380), .ZN(n246) );
  OAI211D0BWP12T U460 ( .A1(n2017), .A2(n3004), .B(n245), .C(n246), .ZN(n1373)
         );
  OAI21D0BWP12T U461 ( .A1(n1790), .A2(n1786), .B(n1787), .ZN(n247) );
  CKND2D0BWP12T U462 ( .A1(n1789), .A2(n1310), .ZN(n248) );
  MOAI22D0BWP12T U463 ( .A1(n247), .A2(n248), .B1(n247), .B2(n248), .ZN(n1793)
         );
  CKND2D0BWP12T U464 ( .A1(n1680), .A2(n1681), .ZN(n249) );
  MAOI22D0BWP12T U465 ( .A1(n1711), .A2(n249), .B1(n1711), .B2(n249), .ZN(
        n2859) );
  NR2D0BWP12T U466 ( .A1(n1849), .A2(n1850), .ZN(n250) );
  MOAI22D0BWP12T U467 ( .A1(n2785), .A2(n250), .B1(n2785), .B2(n250), .ZN(
        n2779) );
  MUX2ND0BWP12T U468 ( .I0(n1953), .I1(n1941), .S(n2353), .ZN(n1883) );
  NR4D0BWP12T U469 ( .A1(n2836), .A2(n2777), .A3(n2806), .A4(n1522), .ZN(n251)
         );
  NR3D0BWP12T U470 ( .A1(n1523), .A2(n3118), .A3(n2889), .ZN(n252) );
  NR3D0BWP12T U471 ( .A1(n2703), .A2(n3078), .A3(n2912), .ZN(n253) );
  NR2D0BWP12T U472 ( .A1(n2913), .A2(n1537), .ZN(n254) );
  ND4D0BWP12T U473 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(n255) );
  OR4D0BWP12T U474 ( .A1(n2675), .A2(n2947), .A3(n2645), .A4(n255), .Z(n256)
         );
  OR4D0BWP12T U475 ( .A1(n2618), .A2(n2566), .A3(n2617), .A4(n256), .Z(n257)
         );
  NR4D0BWP12T U476 ( .A1(n1547), .A2(n2537), .A3(n3051), .A4(n257), .ZN(n1566)
         );
  AOI21D0BWP12T U477 ( .A1(n1972), .A2(n1104), .B(n2263), .ZN(n258) );
  INVD1BWP12T U478 ( .I(n2432), .ZN(n259) );
  OAI22D1BWP12T U479 ( .A1(n1105), .A2(n258), .B1(n1986), .B2(n259), .ZN(n2684) );
  IND2D0BWP12T U480 ( .A1(op[2]), .B1(n916), .ZN(n3018) );
  CKND0BWP12T U481 ( .I(n3093), .ZN(n260) );
  AOI22D0BWP12T U482 ( .A1(n3082), .A2(n2980), .B1(n2982), .B2(n3096), .ZN(
        n261) );
  OAI21D0BWP12T U483 ( .A1(n2977), .A2(n260), .B(n261), .ZN(n262) );
  AO211D0BWP12T U484 ( .A1(n2983), .A2(n3117), .B(n2981), .C(n262), .Z(c_out)
         );
  CKND2D0BWP12T U485 ( .A1(n1832), .A2(n1833), .ZN(n263) );
  MAOI22D0BWP12T U486 ( .A1(n1834), .A2(n263), .B1(n1834), .B2(n263), .ZN(
        n2753) );
  MOAI22D0BWP12T U487 ( .A1(n2466), .A2(b[28]), .B1(n2466), .B2(b[28]), .ZN(
        n264) );
  OAI22D0BWP12T U488 ( .A1(n2469), .A2(n2468), .B1(n2467), .B2(n264), .ZN(
        n2470) );
  MOAI22D0BWP12T U489 ( .A1(a[13]), .A2(b[20]), .B1(a[13]), .B2(b[20]), .ZN(
        n265) );
  OAI22D0BWP12T U490 ( .A1(n2495), .A2(n2494), .B1(n2493), .B2(n265), .ZN(
        n2496) );
  OR4D0BWP12T U491 ( .A1(n2852), .A2(n2817), .A3(n2792), .A4(n2876), .Z(n370)
         );
  CKND2D0BWP12T U492 ( .A1(n1462), .A2(n1463), .ZN(n266) );
  MOAI22D0BWP12T U493 ( .A1(n1464), .A2(n266), .B1(n1464), .B2(n266), .ZN(
        n2617) );
  CKND0BWP12T U494 ( .I(n1607), .ZN(n267) );
  AOI21D0BWP12T U495 ( .A1(n1581), .A2(n267), .B(n1584), .ZN(n268) );
  CKND2D0BWP12T U496 ( .A1(n1582), .A2(n1583), .ZN(n269) );
  MAOI22D0BWP12T U497 ( .A1(n268), .A2(n269), .B1(n268), .B2(n269), .ZN(n2864)
         );
  CKND2D0BWP12T U498 ( .A1(n1212), .A2(n1211), .ZN(n270) );
  MOAI22D0BWP12T U499 ( .A1(n1213), .A2(n270), .B1(n1213), .B2(n270), .ZN(
        n1514) );
  IND2D0BWP12T U500 ( .A1(n416), .B1(n415), .ZN(n1762) );
  NR4D0BWP12T U501 ( .A1(n2867), .A2(n3079), .A3(n2891), .A4(n1405), .ZN(n271)
         );
  NR4D0BWP12T U502 ( .A1(n2751), .A2(n2843), .A3(n1425), .A4(n2800), .ZN(n272)
         );
  NR4D0BWP12T U503 ( .A1(n1428), .A2(n1427), .A3(n1426), .A4(n3089), .ZN(n273)
         );
  NR2D0BWP12T U504 ( .A1(n2729), .A2(n2812), .ZN(n274) );
  NR3D0BWP12T U505 ( .A1(n1440), .A2(n2724), .A3(n3075), .ZN(n275) );
  ND4D0BWP12T U506 ( .A1(n272), .A2(n273), .A3(n274), .A4(n275), .ZN(n276) );
  NR4D0BWP12T U507 ( .A1(n2698), .A2(n2942), .A3(n2670), .A4(n276), .ZN(n277)
         );
  NR3D0BWP12T U508 ( .A1(n2615), .A2(n2970), .A3(n2640), .ZN(n278) );
  NR3D0BWP12T U509 ( .A1(n2562), .A2(n2588), .A3(n3049), .ZN(n279) );
  ND4D0BWP12T U510 ( .A1(n271), .A2(n277), .A3(n278), .A4(n279), .ZN(n280) );
  OR4D0BWP12T U511 ( .A1(n1453), .A2(n1455), .A3(n1454), .A4(n280), .Z(n1457)
         );
  MAOI22D0BWP12T U512 ( .A1(n2201), .A2(a[28]), .B1(n2201), .B2(a[28]), .ZN(
        n2500) );
  MOAI22D0BWP12T U513 ( .A1(b[31]), .A2(n2216), .B1(b[31]), .B2(n2216), .ZN(
        n281) );
  MAOI22D0BWP12T U514 ( .A1(n2976), .A2(n281), .B1(n2976), .B2(n281), .ZN(
        n2412) );
  MAOI222D0BWP12T U515 ( .A(b[31]), .B(n282), .C(n283), .ZN(n2977) );
  CKND0BWP12T U516 ( .I(n2976), .ZN(n282) );
  CKND0BWP12T U517 ( .I(n2216), .ZN(n283) );
  AO222D0BWP12T U518 ( .A1(n896), .A2(n1160), .B1(n1111), .B2(n2320), .C1(
        n1161), .C2(n2324), .Z(n2308) );
  CKND2D0BWP12T U519 ( .A1(n2192), .A2(n1851), .ZN(n284) );
  MAOI22D0BWP12T U520 ( .A1(n2710), .A2(n284), .B1(n2710), .B2(n284), .ZN(
        n2707) );
  CKND2D0BWP12T U521 ( .A1(n1677), .A2(n1408), .ZN(n285) );
  MAOI22D0BWP12T U522 ( .A1(n1678), .A2(n285), .B1(n1678), .B2(n285), .ZN(
        n2725) );
  MAOI22D0BWP12T U523 ( .A1(n2263), .A2(n1883), .B1(n2080), .B2(n1989), .ZN(
        n2960) );
  INVD1BWP12T U524 ( .I(n374), .ZN(n2383) );
  TPOAI22D2BWP12T U525 ( .A1(n2684), .A2(n2377), .B1(n2123), .B2(n2120), .ZN(
        n2089) );
  XOR2D2BWP12T U526 ( .A1(n1926), .A2(n2764), .Z(n2134) );
  FA1D2BWP12T U527 ( .A(n2498), .B(n1377), .CI(n1647), .CO(n1646), .S(n2442)
         );
  TPNR2D1BWP12T U528 ( .A1(n1926), .A2(n902), .ZN(n2101) );
  INVD2BWP12T U529 ( .I(n1150), .ZN(n2110) );
  INVD1BWP12T U530 ( .I(n1020), .ZN(n902) );
  OAI21D1BWP12T U531 ( .A1(n790), .A2(n1324), .B(n789), .ZN(n1476) );
  FA1D2BWP12T U532 ( .A(n2571), .B(b[23]), .CI(n1798), .CO(n1727), .S(n2568)
         );
  INVD2BWP12T U533 ( .I(a[19]), .ZN(n2623) );
  TPAOI21D2BWP12T U534 ( .A1(n1495), .A2(n1494), .B(n783), .ZN(n1280) );
  BUFFXD8BWP12T U535 ( .I(n303), .Z(n2518) );
  IOA21D2BWP12T U536 ( .A1(n3078), .A2(n3117), .B(n3077), .ZN(result[13]) );
  OAI211D2BWP12T U537 ( .A1(n2975), .A2(n2702), .B(n2701), .C(n2700), .ZN(
        result[17]) );
  DCCKND16BWP12T U538 ( .I(n2368), .ZN(n1277) );
  OAI211D2BWP12T U539 ( .A1(n2975), .A2(n2946), .B(n2945), .C(n2944), .ZN(
        result[16]) );
  OAI222D0BWP12T U540 ( .A1(n2121), .A2(n2053), .B1(n2119), .B2(n2052), .C1(
        n2123), .C2(n2051), .ZN(n2950) );
  INVD3BWP12T U541 ( .I(n2052), .ZN(n2014) );
  FA1D2BWP12T U542 ( .A(b[30]), .B(a[30]), .CI(n1569), .CO(n2978), .S(n3008)
         );
  FA1D2BWP12T U543 ( .A(n2571), .B(b[23]), .CI(n1571), .CO(n1640), .S(n2567)
         );
  AOI21D1BWP12T U544 ( .A1(n1362), .A2(n1360), .B(n873), .ZN(n1605) );
  BUFFXD8BWP12T U545 ( .I(n2350), .Z(n429) );
  INVD9BWP12T U546 ( .I(n2179), .ZN(n2350) );
  INVD4BWP12T U547 ( .I(b[1]), .ZN(n2179) );
  AOI222XD4BWP12T U548 ( .A1(n2074), .A2(n2106), .B1(n2103), .B2(n2098), .C1(
        n1048), .C2(n2109), .ZN(n2052) );
  ND4D2BWP12T U549 ( .A1(n1131), .A2(n1130), .A3(n1129), .A4(n1128), .ZN(n1132) );
  TPAOI22D1BWP12T U550 ( .A1(n1107), .A2(n2387), .B1(n3091), .B2(n2089), .ZN(
        n1131) );
  AO21D4BWP12T U551 ( .A1(n2776), .A2(n3117), .B(n2775), .Z(result[3]) );
  OAI211D2BWP12T U552 ( .A1(n2894), .A2(n2774), .B(n2773), .C(n2772), .ZN(
        n2775) );
  TPND2D1BWP12T U553 ( .A1(n2933), .A2(n3091), .ZN(n2824) );
  INVD3BWP12T U554 ( .I(n1926), .ZN(n2074) );
  INR2D2BWP12T U555 ( .A1(n2207), .B1(n1918), .ZN(n1926) );
  CKND2D0BWP12T U556 ( .A1(n2110), .A2(n2233), .ZN(n905) );
  CKND2D0BWP12T U557 ( .A1(n2110), .A2(n2224), .ZN(n996) );
  CKND2D2BWP12T U558 ( .A1(n2110), .A2(n1111), .ZN(n2120) );
  OAI22D0BWP12T U559 ( .A1(n1918), .A2(n2900), .B1(n1917), .B2(n2192), .ZN(
        n1914) );
  OAI22D0BWP12T U560 ( .A1(n1918), .A2(n2819), .B1(n1917), .B2(n3104), .ZN(
        n1922) );
  OAI22D0BWP12T U561 ( .A1(n1918), .A2(n2712), .B1(n1917), .B2(n2650), .ZN(
        n1916) );
  OAI22D0BWP12T U562 ( .A1(n1918), .A2(n2917), .B1(n1919), .B2(n2682), .ZN(
        n1266) );
  OAI22D0BWP12T U563 ( .A1(n1918), .A2(n2846), .B1(n2898), .B2(n1917), .ZN(
        n1261) );
  OAI22D0BWP12T U564 ( .A1(n1918), .A2(n2739), .B1(n1917), .B2(n2819), .ZN(
        n1259) );
  OAI22D0BWP12T U565 ( .A1(n1918), .A2(n2193), .B1(n1917), .B2(n2712), .ZN(
        n1257) );
  OAI22D0BWP12T U566 ( .A1(n1918), .A2(n2952), .B1(n1920), .B2(n3022), .ZN(
        n1264) );
  TPNR2D2BWP12T U567 ( .A1(n2101), .A2(n394), .ZN(n395) );
  OAI22D0BWP12T U568 ( .A1(n1918), .A2(n3059), .B1(n1917), .B2(n2917), .ZN(
        n357) );
  OAI22D0BWP12T U569 ( .A1(n1918), .A2(n2596), .B1(n1917), .B2(n2544), .ZN(
        n338) );
  OAI22D0BWP12T U570 ( .A1(n1918), .A2(n3100), .B1(a[13]), .B2(n1917), .ZN(
        n1198) );
  OAI22D0BWP12T U571 ( .A1(n1918), .A2(n2623), .B1(n1917), .B2(n3022), .ZN(
        n1891) );
  OAI22D0BWP12T U572 ( .A1(n1918), .A2(n2574), .B1(n1917), .B2(n2200), .ZN(
        n1881) );
  OAI22D0BWP12T U573 ( .A1(n1918), .A2(n2650), .B1(n1917), .B2(n2596), .ZN(
        n1191) );
  OAI22D0BWP12T U574 ( .A1(n1918), .A2(n2787), .B1(n1917), .B2(n2872), .ZN(
        n1203) );
  OAI22D0BWP12T U575 ( .A1(n1918), .A2(n3022), .B1(n1917), .B2(n2202), .ZN(
        n1193) );
  OAI22D0BWP12T U576 ( .A1(n1918), .A2(n2192), .B1(n1917), .B2(n2682), .ZN(
        n1200) );
  TPND2D2BWP12T U577 ( .A1(n1918), .A2(n1917), .ZN(n2099) );
  INVD2BWP12T U578 ( .I(n347), .ZN(n1917) );
  DEL025D1BWP12T U579 ( .I(n1277), .Z(n306) );
  OR2D2BWP12T U580 ( .A1(n2159), .A2(a[12]), .Z(n286) );
  NR2D1BWP12T U581 ( .A1(n2350), .A2(n1277), .ZN(n291) );
  INVD1BWP12T U582 ( .I(n291), .ZN(n1918) );
  CKND0BWP12T U583 ( .I(n1277), .ZN(n1269) );
  NR2D0BWP12T U584 ( .A1(n2163), .A2(n2898), .ZN(n1286) );
  INVD2BWP12T U585 ( .I(n2171), .ZN(n2351) );
  INVD1BWP12T U586 ( .I(n2594), .ZN(n475) );
  INVD2BWP12T U587 ( .I(n2596), .ZN(n2594) );
  INVD1BWP12T U588 ( .I(n2201), .ZN(n2358) );
  INVD2BWP12T U589 ( .I(n2202), .ZN(n2460) );
  INVD2BWP12T U590 ( .I(n2623), .ZN(n2621) );
  OR2D2BWP12T U591 ( .A1(mult_x_18_n558), .A2(mult_x_18_n542), .Z(n287) );
  INVD2BWP12T U592 ( .I(n2162), .ZN(n2852) );
  OR2XD1BWP12T U593 ( .A1(mult_x_18_n706), .A2(mult_x_18_n712), .Z(n288) );
  OR2XD1BWP12T U594 ( .A1(mult_x_18_n590), .A2(mult_x_18_n603), .Z(n289) );
  INVD3BWP12T U595 ( .I(n2712), .ZN(n2710) );
  OR2XD1BWP12T U596 ( .A1(n2160), .A2(a[13]), .Z(n1439) );
  NR4D1BWP12T U597 ( .A1(n373), .A2(n372), .A3(n371), .A4(n370), .ZN(n374) );
  INVD6BWP12T U598 ( .I(n2206), .ZN(n2466) );
  NR2D1BWP12T U599 ( .A1(n860), .A2(n2817), .ZN(n1760) );
  CKBD1BWP12T U600 ( .I(n2815), .Z(n811) );
  XOR2D1BWP12T U601 ( .A1(n1638), .A2(n1637), .Z(n290) );
  INVD6BWP12T U602 ( .I(n2819), .ZN(n2815) );
  XOR2D1BWP12T U603 ( .A1(n1703), .A2(n1702), .Z(n292) );
  NR2D1BWP12T U604 ( .A1(n2170), .A2(n811), .ZN(n1695) );
  OR2D2BWP12T U605 ( .A1(mult_x_18_n654), .A2(mult_x_18_n664), .Z(n293) );
  NR2D1BWP12T U606 ( .A1(n2870), .A2(n2876), .ZN(n1772) );
  INVD2BWP12T U607 ( .I(a[1]), .ZN(n2210) );
  DCCKND12BWP12T U608 ( .I(n2210), .ZN(n2349) );
  BUFFD2BWP12T U609 ( .I(a[0]), .Z(n2172) );
  INVD2BWP12T U610 ( .I(n2172), .ZN(n2449) );
  TPND2D4BWP12T U611 ( .A1(n2349), .A2(n2449), .ZN(n2450) );
  XNR2D1BWP12T U612 ( .A1(n2349), .A2(b[22]), .ZN(n521) );
  XNR2D1BWP12T U613 ( .A1(n2349), .A2(b[23]), .ZN(n462) );
  OAI22D1BWP12T U614 ( .A1(n2450), .A2(n521), .B1(n462), .B2(n2449), .ZN(n296)
         );
  INVD2BWP12T U615 ( .I(a[15]), .ZN(n2712) );
  XNR2D2BWP12T U616 ( .A1(n2710), .A2(n2915), .ZN(n2511) );
  INVD2BWP12T U617 ( .I(a[17]), .ZN(n2682) );
  INVD4BWP12T U618 ( .I(n2682), .ZN(n2679) );
  XOR2XD1BWP12T U619 ( .A1(n2679), .A2(n2915), .Z(n294) );
  TPND2D2BWP12T U620 ( .A1(n2511), .A2(n294), .ZN(n2513) );
  INVD1BWP12T U621 ( .I(b[6]), .ZN(n2169) );
  XNR2XD1BWP12T U622 ( .A1(n2679), .A2(n2792), .ZN(n543) );
  INVD1BWP12T U623 ( .I(b[7]), .ZN(n2170) );
  INVD2BWP12T U624 ( .I(n2170), .ZN(n2817) );
  XNR2D1BWP12T U625 ( .A1(n2679), .A2(n2817), .ZN(n568) );
  OAI22D1BWP12T U626 ( .A1(n2513), .A2(n543), .B1(n568), .B2(n2511), .ZN(n295)
         );
  HA1D0BWP12T U627 ( .A(n296), .B(n295), .CO(mult_x_18_n555), .S(
        mult_x_18_n556) );
  XNR2D1BWP12T U628 ( .A1(n2349), .A2(b[18]), .ZN(n525) );
  XNR2D1BWP12T U629 ( .A1(n2349), .A2(b[19]), .ZN(n506) );
  OAI22D1BWP12T U630 ( .A1(n2450), .A2(n525), .B1(n506), .B2(n2449), .ZN(n298)
         );
  BUFFD3BWP12T U631 ( .I(b[2]), .Z(n2353) );
  XNR2D1BWP12T U632 ( .A1(n2679), .A2(n2353), .ZN(n624) );
  BUFFD12BWP12T U633 ( .I(b[3]), .Z(n2764) );
  XNR2XD1BWP12T U634 ( .A1(n2679), .A2(n2764), .ZN(n631) );
  OAI22D1BWP12T U635 ( .A1(n2513), .A2(n624), .B1(n631), .B2(n2511), .ZN(n297)
         );
  HA1D0BWP12T U636 ( .A(n298), .B(n297), .CO(mult_x_18_n614), .S(
        mult_x_18_n615) );
  BUFFD2BWP12T U637 ( .I(a[8]), .Z(n2846) );
  INVD2BWP12T U638 ( .I(a[7]), .ZN(n2819) );
  XNR2XD8BWP12T U639 ( .A1(n2846), .A2(n2815), .ZN(n2487) );
  INVD3BWP12T U640 ( .I(a[9]), .ZN(n2872) );
  INVD9BWP12T U641 ( .I(n2872), .ZN(n2870) );
  XOR2D1BWP12T U642 ( .A1(n2846), .A2(n2870), .Z(n299) );
  ND2D3BWP12T U643 ( .A1(n2487), .A2(n299), .ZN(n2489) );
  XNR2D1BWP12T U644 ( .A1(n2870), .A2(b[21]), .ZN(n626) );
  XNR2D1BWP12T U645 ( .A1(n2870), .A2(b[22]), .ZN(n748) );
  TPOAI22D0BWP12T U646 ( .A1(n2489), .A2(n626), .B1(n2487), .B2(n748), .ZN(
        mult_x_18_n893) );
  BUFFD1BWP12T U647 ( .I(a[18]), .Z(n2652) );
  XNR2D2BWP12T U648 ( .A1(n2679), .A2(n2652), .ZN(n2482) );
  XOR2XD1BWP12T U649 ( .A1(n2652), .A2(n2621), .Z(n300) );
  CKND2D2BWP12T U650 ( .A1(n2482), .A2(n300), .ZN(n2484) );
  BUFFD2BWP12T U651 ( .I(b[11]), .Z(n2904) );
  XNR2XD1BWP12T U652 ( .A1(n2621), .A2(n2904), .ZN(n679) );
  BUFFD2BWP12T U653 ( .I(b[12]), .Z(n2452) );
  XNR2XD0BWP12T U654 ( .A1(n2621), .A2(n2452), .ZN(n302) );
  OAI22D0BWP12T U655 ( .A1(n2484), .A2(n679), .B1(n2482), .B2(n302), .ZN(
        mult_x_18_n798) );
  INVD1BWP12T U656 ( .I(a[25]), .ZN(n2202) );
  XNR2D2BWP12T U657 ( .A1(a[26]), .A2(n2460), .ZN(n2476) );
  INVD1BWP12T U658 ( .I(a[27]), .ZN(n2201) );
  XNR2XD1BWP12T U659 ( .A1(n2201), .A2(a[26]), .ZN(n301) );
  TPND2D2BWP12T U660 ( .A1(n2476), .A2(n301), .ZN(n2478) );
  INVD1BWP12T U661 ( .I(b[4]), .ZN(n358) );
  XNR2XD0BWP12T U662 ( .A1(n2499), .A2(n2358), .ZN(n756) );
  INVD1BWP12T U663 ( .I(b[5]), .ZN(n2171) );
  XOR2XD0BWP12T U664 ( .A1(n2201), .A2(n2351), .Z(n2477) );
  OAI22D0BWP12T U665 ( .A1(n2478), .A2(n756), .B1(n2476), .B2(n2477), .ZN(
        mult_x_18_n757) );
  XNR2XD0BWP12T U666 ( .A1(n2621), .A2(b[13]), .ZN(n2483) );
  OAI22D0BWP12T U667 ( .A1(n2484), .A2(n302), .B1(n2482), .B2(n2483), .ZN(
        mult_x_18_n797) );
  ND2D1BWP12T U668 ( .A1(op[3]), .A2(op[0]), .ZN(n416) );
  INR3D0BWP12T U669 ( .A1(op[2]), .B1(op[1]), .B2(n416), .ZN(n3117) );
  INVD1BWP12T U670 ( .I(n3117), .ZN(n2975) );
  BUFFD2BWP12T U671 ( .I(a[2]), .Z(n2352) );
  INVD2BWP12T U672 ( .I(a[3]), .ZN(n322) );
  INVD6BWP12T U673 ( .I(n322), .ZN(n2516) );
  XOR2D1BWP12T U674 ( .A1(n2352), .A2(n2516), .Z(n304) );
  ND2D4BWP12T U675 ( .A1(n2518), .A2(n304), .ZN(n2520) );
  CKBD1BWP12T U676 ( .I(n2353), .Z(n2503) );
  XNR2D1BWP12T U677 ( .A1(n2503), .A2(n2516), .ZN(n310) );
  XNR2D1BWP12T U678 ( .A1(n2764), .A2(n2516), .ZN(n664) );
  OAI22D1BWP12T U679 ( .A1(n2520), .A2(n310), .B1(n2518), .B2(n664), .ZN(n774)
         );
  INVD3BWP12T U680 ( .I(a[5]), .ZN(n2206) );
  BUFFD2BWP12T U681 ( .I(a[4]), .Z(n2738) );
  XOR2XD2BWP12T U682 ( .A1(n2466), .A2(n2738), .Z(n305) );
  XNR2XD8BWP12T U683 ( .A1(n2738), .A2(n2516), .ZN(n2467) );
  ND2D8BWP12T U684 ( .A1(n305), .A2(n2467), .ZN(n2469) );
  INVD4BWP12T U685 ( .I(b[0]), .ZN(n2368) );
  XNR2D1BWP12T U686 ( .A1(n2466), .A2(n306), .ZN(n307) );
  XNR2D1BWP12T U687 ( .A1(n2466), .A2(n429), .ZN(n529) );
  OAI22D1BWP12T U688 ( .A1(n2469), .A2(n307), .B1(n529), .B2(n2467), .ZN(n773)
         );
  XNR2D1BWP12T U689 ( .A1(n2499), .A2(n2349), .ZN(n309) );
  XNR2D1BWP12T U690 ( .A1(n2351), .A2(n2349), .ZN(n564) );
  OAI22D1BWP12T U691 ( .A1(n2450), .A2(n309), .B1(n564), .B2(n2449), .ZN(n458)
         );
  INVD6BWP12T U692 ( .I(n2466), .ZN(n883) );
  IND2D1BWP12T U693 ( .A1(n1277), .B1(n2466), .ZN(n308) );
  OAI22D1BWP12T U694 ( .A1(n2469), .A2(n883), .B1(n2467), .B2(n308), .ZN(n457)
         );
  XNR2D1BWP12T U695 ( .A1(n2764), .A2(n2349), .ZN(n316) );
  OAI22D1BWP12T U696 ( .A1(n2450), .A2(n316), .B1(n309), .B2(n2449), .ZN(n315)
         );
  INR2D1BWP12T U697 ( .A1(n306), .B1(n2467), .ZN(n314) );
  XNR2D1BWP12T U698 ( .A1(n2350), .A2(n2516), .ZN(n317) );
  OAI22D1BWP12T U699 ( .A1(n2520), .A2(n317), .B1(n2518), .B2(n310), .ZN(n313)
         );
  NR2D1BWP12T U700 ( .A1(n312), .A2(n311), .ZN(n776) );
  ND2D1BWP12T U701 ( .A1(n312), .A2(n311), .ZN(n775) );
  FA1D0BWP12T U702 ( .A(n315), .B(n314), .CI(n313), .CO(n311), .S(n334) );
  XNR2D1BWP12T U703 ( .A1(n2503), .A2(n2349), .ZN(n323) );
  OAI22D1BWP12T U704 ( .A1(n2450), .A2(n323), .B1(n316), .B2(n2449), .ZN(n320)
         );
  XNR2D1BWP12T U705 ( .A1(n1277), .A2(n2516), .ZN(n318) );
  OAI22D1BWP12T U706 ( .A1(n2520), .A2(n318), .B1(n2518), .B2(n317), .ZN(n319)
         );
  OR2XD1BWP12T U707 ( .A1(n334), .A2(n333), .Z(n1509) );
  HA1D0BWP12T U708 ( .A(n320), .B(n319), .CO(n333), .S(n332) );
  IND2D1BWP12T U709 ( .A1(n1277), .B1(n2516), .ZN(n321) );
  OAI22D1BWP12T U710 ( .A1(n2520), .A2(n322), .B1(n2518), .B2(n321), .ZN(n331)
         );
  NR2D1BWP12T U711 ( .A1(n332), .A2(n331), .ZN(n1511) );
  XNR2D1BWP12T U712 ( .A1(n2350), .A2(n2349), .ZN(n324) );
  OAI22D1BWP12T U713 ( .A1(n2450), .A2(n324), .B1(n323), .B2(n2449), .ZN(n329)
         );
  INR2D1BWP12T U714 ( .A1(n1277), .B1(n2518), .ZN(n328) );
  OR2XD1BWP12T U715 ( .A1(n329), .A2(n328), .Z(n1212) );
  OAI22D1BWP12T U716 ( .A1(n2450), .A2(n1270), .B1(n324), .B2(n2449), .ZN(
        n1103) );
  INVD1BWP12T U717 ( .I(n1103), .ZN(n327) );
  IND2D1BWP12T U718 ( .A1(n1277), .B1(n2349), .ZN(n325) );
  ND2D1BWP12T U719 ( .A1(n2450), .A2(n325), .ZN(n1102) );
  INVD1BWP12T U720 ( .I(n1102), .ZN(n326) );
  NR2D1BWP12T U721 ( .A1(n327), .A2(n326), .ZN(n1213) );
  ND2D1BWP12T U722 ( .A1(n329), .A2(n328), .ZN(n1211) );
  INVD1BWP12T U723 ( .I(n1211), .ZN(n330) );
  AOI21D1BWP12T U724 ( .A1(n1212), .A2(n1213), .B(n330), .ZN(n1513) );
  ND2D1BWP12T U725 ( .A1(n332), .A2(n331), .ZN(n1512) );
  OAI21D1BWP12T U726 ( .A1(n1511), .A2(n1513), .B(n1512), .ZN(n1510) );
  ND2D1BWP12T U727 ( .A1(n334), .A2(n333), .ZN(n1508) );
  INVD1BWP12T U728 ( .I(n1508), .ZN(n335) );
  AOI21D1BWP12T U729 ( .A1(n1509), .A2(n1510), .B(n335), .ZN(n777) );
  INVD1BWP12T U730 ( .I(n1517), .ZN(n439) );
  CKBD1BWP12T U731 ( .I(a[3]), .Z(n1834) );
  INVD1BWP12T U732 ( .I(n2352), .ZN(n1832) );
  ND2D1BWP12T U733 ( .A1(n2760), .A2(n1832), .ZN(n336) );
  CKBD1BWP12T U734 ( .I(n2349), .Z(n1121) );
  ND2D1BWP12T U735 ( .A1(n2210), .A2(n2449), .ZN(n1243) );
  NR2D1BWP12T U736 ( .A1(n336), .A2(n1243), .ZN(n886) );
  INVD1BWP12T U737 ( .I(n886), .ZN(n1850) );
  NR2D0BWP12T U738 ( .A1(op[1]), .A2(op[2]), .ZN(n400) );
  INVD2BWP12T U739 ( .I(n3040), .ZN(n3096) );
  OR2XD1BWP12T U740 ( .A1(n2353), .A2(n2350), .Z(n1352) );
  INVD1BWP12T U741 ( .I(n1352), .ZN(n896) );
  INVD1BWP12T U742 ( .I(a[31]), .ZN(n2216) );
  INVD1BWP12T U743 ( .I(a[29]), .ZN(n2428) );
  IND2D1BWP12T U744 ( .A1(n2350), .B1(n1277), .ZN(n1919) );
  INVD1BWP12T U745 ( .I(a[30]), .ZN(n2996) );
  OAI22D1BWP12T U746 ( .A1(n1918), .A2(n2428), .B1(n1919), .B2(n2996), .ZN(
        n1092) );
  MOAI22D0BWP12T U747 ( .A1(n896), .A2(n2216), .B1(n1092), .B2(n2207), .ZN(
        n1877) );
  DCCKND4BWP12T U748 ( .I(a[21]), .ZN(n2596) );
  AN2D1BWP12T U749 ( .A1(n2350), .A2(n1277), .Z(n347) );
  CKBD1BWP12T U750 ( .I(a[24]), .Z(n2541) );
  IND2D1BWP12T U751 ( .A1(n1277), .B1(n2350), .ZN(n1920) );
  DCCKND4BWP12T U752 ( .I(a[23]), .ZN(n2574) );
  CKND1BWP12T U753 ( .I(a[22]), .ZN(n3022) );
  OAI22D1BWP12T U754 ( .A1(n1920), .A2(n2574), .B1(n1919), .B2(n3022), .ZN(
        n337) );
  NR2D1BWP12T U755 ( .A1(n338), .A2(n337), .ZN(n1973) );
  OR2XD1BWP12T U756 ( .A1(n2353), .A2(n2764), .Z(n2029) );
  INR2D1BWP12T U757 ( .A1(n2460), .B1(n1918), .ZN(n340) );
  CKND1BWP12T U758 ( .I(a[26]), .ZN(n2200) );
  NR2D1BWP12T U759 ( .A1(n1919), .A2(n2200), .ZN(n339) );
  NR2D1BWP12T U760 ( .A1(n340), .A2(n339), .ZN(n344) );
  NR2D1BWP12T U761 ( .A1(n1920), .A2(n2201), .ZN(n342) );
  CKND1BWP12T U762 ( .I(a[28]), .ZN(n2198) );
  NR2D1BWP12T U763 ( .A1(n1917), .A2(n2198), .ZN(n341) );
  NR2D1BWP12T U764 ( .A1(n342), .A2(n341), .ZN(n343) );
  ND2D1BWP12T U765 ( .A1(n344), .A2(n343), .ZN(n1093) );
  INVD1BWP12T U766 ( .I(n1093), .ZN(n1972) );
  IND2D1BWP12T U767 ( .A1(n2764), .B1(n2353), .ZN(n1970) );
  OAI22D1BWP12T U768 ( .A1(n1973), .A2(n2029), .B1(n1972), .B2(n1970), .ZN(
        n419) );
  AOI21D1BWP12T U769 ( .A1(n1877), .A2(n2764), .B(n419), .ZN(n2601) );
  ND2XD0BWP12T U770 ( .A1(n2601), .A2(n2740), .ZN(n375) );
  INVD1BWP12T U771 ( .I(n2029), .ZN(n1903) );
  AOI22D1BWP12T U772 ( .A1(n291), .A2(n2466), .B1(n347), .B2(n2846), .ZN(n346)
         );
  INVD1BWP12T U773 ( .I(n1920), .ZN(n351) );
  INVD1BWP12T U774 ( .I(n1919), .ZN(n350) );
  BUFFD2BWP12T U775 ( .I(a[6]), .Z(n2785) );
  AOI22D1BWP12T U776 ( .A1(n351), .A2(n2815), .B1(n350), .B2(n2785), .ZN(n345)
         );
  ND2D1BWP12T U777 ( .A1(n346), .A2(n345), .ZN(n1100) );
  OAI22D1BWP12T U778 ( .A1(n1918), .A2(n2682), .B1(n1919), .B2(n2650), .ZN(
        n349) );
  INVD1BWP12T U779 ( .I(a[20]), .ZN(n2952) );
  OAI22D1BWP12T U780 ( .A1(n1920), .A2(n2623), .B1(n1917), .B2(n2952), .ZN(
        n348) );
  NR2D1BWP12T U781 ( .A1(n349), .A2(n348), .ZN(n1971) );
  ND2D1BWP12T U782 ( .A1(n2764), .A2(n2353), .ZN(n1986) );
  INVD3BWP12T U783 ( .I(n2900), .ZN(n2898) );
  INVD1P75BWP12T U784 ( .I(a[10]), .ZN(n3104) );
  INVD3BWP12T U785 ( .I(n3104), .ZN(n3100) );
  AOI22D1BWP12T U786 ( .A1(n351), .A2(n2898), .B1(n350), .B2(n3100), .ZN(n355)
         );
  INR2D1BWP12T U787 ( .A1(n2870), .B1(n1918), .ZN(n353) );
  NR2D1BWP12T U788 ( .A1(n1917), .A2(n2193), .ZN(n352) );
  NR2D1BWP12T U789 ( .A1(n353), .A2(n352), .ZN(n354) );
  ND2D1BWP12T U790 ( .A1(n355), .A2(n354), .ZN(n1874) );
  INVD1BWP12T U791 ( .I(n1874), .ZN(n1095) );
  OAI22D1BWP12T U792 ( .A1(n1971), .A2(n1986), .B1(n1095), .B2(n1970), .ZN(
        n360) );
  INVD1BWP12T U793 ( .I(a[13]), .ZN(n3059) );
  CKND1BWP12T U794 ( .I(n2915), .ZN(n2917) );
  OAI22D1BWP12T U795 ( .A1(n1920), .A2(n2712), .B1(n1919), .B2(n2192), .ZN(
        n356) );
  NR2D1BWP12T U796 ( .A1(n357), .A2(n356), .ZN(n1974) );
  INVD1BWP12T U797 ( .I(n2764), .ZN(n2263) );
  NR2D1BWP12T U798 ( .A1(n2263), .A2(n2353), .ZN(n2076) );
  INVD1BWP12T U799 ( .I(n2076), .ZN(n1989) );
  BUFFD1BWP12T U800 ( .I(n358), .Z(n2377) );
  OAI21D0BWP12T U801 ( .A1(n1974), .A2(n1989), .B(n2377), .ZN(n359) );
  AOI211D1BWP12T U802 ( .A1(n1903), .A2(n1100), .B(n360), .C(n359), .ZN(n417)
         );
  NR2XD0BWP12T U803 ( .A1(b[31]), .A2(b[30]), .ZN(n363) );
  NR2D1BWP12T U804 ( .A1(b[29]), .A2(b[28]), .ZN(n362) );
  NR2D1BWP12T U805 ( .A1(b[27]), .A2(b[26]), .ZN(n361) );
  ND4D1BWP12T U806 ( .A1(n363), .A2(n362), .A3(n361), .A4(n2171), .ZN(n373) );
  NR2XD0BWP12T U807 ( .A1(b[25]), .A2(b[24]), .ZN(n365) );
  NR2XD0BWP12T U808 ( .A1(b[23]), .A2(b[22]), .ZN(n364) );
  NR2D1BWP12T U809 ( .A1(b[17]), .A2(b[16]), .ZN(n369) );
  NR2D1BWP12T U810 ( .A1(b[15]), .A2(b[14]), .ZN(n368) );
  NR2D1BWP12T U811 ( .A1(b[13]), .A2(n2452), .ZN(n367) );
  INVD1BWP12T U812 ( .I(b[10]), .ZN(n2161) );
  INVD3BWP12T U813 ( .I(n2161), .ZN(n3106) );
  NR2D1BWP12T U814 ( .A1(n2904), .A2(n3106), .ZN(n366) );
  ND4D1BWP12T U815 ( .A1(n369), .A2(n368), .A3(n367), .A4(n366), .ZN(n371) );
  INVD1BWP12T U816 ( .I(b[9]), .ZN(n2168) );
  INVD1BWP12T U817 ( .I(b[8]), .ZN(n2162) );
  NR2D1BWP12T U818 ( .A1(n417), .A2(n2383), .ZN(n424) );
  INVD2BWP12T U819 ( .I(n2383), .ZN(n2396) );
  OR2D2BWP12T U820 ( .A1(n2396), .A2(n2216), .Z(n1991) );
  INVD1BWP12T U821 ( .I(n1991), .ZN(n1976) );
  AOI21D1BWP12T U822 ( .A1(n375), .A2(n424), .B(n1976), .ZN(n1978) );
  NR2D1BWP12T U823 ( .A1(op[0]), .A2(op[1]), .ZN(n916) );
  IND2XD1BWP12T U824 ( .A1(op[3]), .B1(op[2]), .ZN(n433) );
  INR2D1BWP12T U825 ( .A1(n916), .B1(n433), .ZN(n3084) );
  INVD1BWP12T U826 ( .I(n3084), .ZN(n3071) );
  MAOI22D0BWP12T U827 ( .A1(n1852), .A2(n3096), .B1(n1978), .B2(n3071), .ZN(
        n438) );
  IND2XD1BWP12T U828 ( .A1(op[0]), .B1(op[1]), .ZN(n403) );
  NR2D1BWP12T U829 ( .A1(n433), .A2(n403), .ZN(n3076) );
  NR2D1BWP12T U830 ( .A1(n1104), .A2(n2352), .ZN(n1223) );
  INVD1BWP12T U831 ( .I(n2350), .ZN(n377) );
  CKBD1BWP12T U832 ( .I(n2349), .Z(n376) );
  NR2D1BWP12T U833 ( .A1(n377), .A2(n376), .ZN(n1221) );
  NR2D1BWP12T U834 ( .A1(n1223), .A2(n1221), .ZN(n379) );
  NR2D1BWP12T U835 ( .A1(n2172), .A2(c_in), .ZN(n1278) );
  CKND2D1BWP12T U836 ( .A1(n2172), .A2(c_in), .ZN(n1279) );
  OAI21D1BWP12T U837 ( .A1(n1277), .A2(n1278), .B(n1279), .ZN(n1108) );
  ND2D1BWP12T U838 ( .A1(n377), .A2(n376), .ZN(n1220) );
  ND2D1BWP12T U839 ( .A1(n1104), .A2(n2352), .ZN(n1224) );
  OAI21D1BWP12T U840 ( .A1(n1223), .A2(n1220), .B(n1224), .ZN(n378) );
  AOI21D1BWP12T U841 ( .A1(n379), .A2(n1108), .B(n378), .ZN(n846) );
  INVD1BWP12T U842 ( .I(n846), .ZN(n1430) );
  CKBD1BWP12T U843 ( .I(a[3]), .Z(n380) );
  INVD1BWP12T U844 ( .I(n2740), .ZN(n381) );
  NR2D1BWP12T U845 ( .A1(n381), .A2(n2738), .ZN(n1431) );
  ND2D1BWP12T U846 ( .A1(n650), .A2(n380), .ZN(n1429) );
  CKND2D1BWP12T U847 ( .A1(n381), .A2(n2738), .ZN(n1432) );
  OAI21D1BWP12T U848 ( .A1(n1431), .A2(n1429), .B(n1432), .ZN(n1419) );
  NR2D1BWP12T U849 ( .A1(n2171), .A2(n2466), .ZN(n1421) );
  ND2D1BWP12T U850 ( .A1(n2171), .A2(n2466), .ZN(n1420) );
  INR2D1BWP12T U851 ( .A1(op[1]), .B1(op[2]), .ZN(n415) );
  INR2D1BWP12T U852 ( .A1(op[3]), .B1(n392), .ZN(n382) );
  INVD1BWP12T U853 ( .I(n382), .ZN(n3047) );
  NR2D1BWP12T U854 ( .A1(n1269), .A2(n2172), .ZN(n1114) );
  CKBD1BWP12T U855 ( .I(n2349), .Z(n383) );
  NR2D1BWP12T U856 ( .A1(n377), .A2(n383), .ZN(n1112) );
  ND2D1BWP12T U857 ( .A1(n377), .A2(n383), .ZN(n1113) );
  OAI21D1BWP12T U858 ( .A1(n1114), .A2(n1112), .B(n1113), .ZN(n1242) );
  CKBD1BWP12T U859 ( .I(a[3]), .Z(n384) );
  NR2D1BWP12T U860 ( .A1(n650), .A2(n384), .ZN(n1688) );
  NR2D1BWP12T U861 ( .A1(n1104), .A2(n2352), .ZN(n1686) );
  NR2D1BWP12T U862 ( .A1(n1688), .A2(n1686), .ZN(n386) );
  CKND2D1BWP12T U863 ( .A1(n1104), .A2(n2352), .ZN(n1685) );
  ND2D1BWP12T U864 ( .A1(n650), .A2(n384), .ZN(n1689) );
  OAI21D1BWP12T U865 ( .A1(n1688), .A2(n1685), .B(n1689), .ZN(n385) );
  AOI21D1BWP12T U866 ( .A1(n1242), .A2(n386), .B(n385), .ZN(n816) );
  INVD1BWP12T U867 ( .I(n816), .ZN(n1703) );
  CKND1BWP12T U868 ( .I(n2740), .ZN(n387) );
  NR2D1BWP12T U869 ( .A1(n387), .A2(n2738), .ZN(n808) );
  INVD1BWP12T U870 ( .I(n808), .ZN(n1701) );
  CKND2D1BWP12T U871 ( .A1(n387), .A2(n2738), .ZN(n1700) );
  CKND0BWP12T U872 ( .I(n1700), .ZN(n388) );
  TPAOI21D0BWP12T U873 ( .A1(n1703), .A2(n1701), .B(n388), .ZN(n391) );
  NR2D1BWP12T U874 ( .A1(n2171), .A2(n2466), .ZN(n810) );
  CKND0BWP12T U875 ( .I(n810), .ZN(n389) );
  ND2D1BWP12T U876 ( .A1(n2171), .A2(n2466), .ZN(n809) );
  ND2XD0BWP12T U877 ( .A1(n389), .A2(n809), .ZN(n390) );
  XOR2XD1BWP12T U878 ( .A1(n391), .A2(n390), .Z(n1704) );
  INVD1BWP12T U879 ( .I(n1704), .ZN(n423) );
  TPND2D4BWP12T U880 ( .A1(n374), .A2(n2377), .ZN(n2393) );
  CKND0BWP12T U881 ( .I(op[3]), .ZN(n399) );
  INR2D1BWP12T U882 ( .A1(n399), .B1(n392), .ZN(n3067) );
  INVD1BWP12T U883 ( .I(n3067), .ZN(n2928) );
  NR2XD3BWP12T U884 ( .A1(n2393), .A2(n2928), .ZN(n3108) );
  INVD2BWP12T U885 ( .I(n3108), .ZN(n2879) );
  NR2XD3BWP12T U886 ( .A1(n2879), .A2(n2764), .ZN(n2826) );
  MUX2D1BWP12T U887 ( .I0(n2466), .I1(n2738), .S(n1277), .Z(n1160) );
  NR2D1BWP12T U888 ( .A1(n2368), .A2(n2172), .ZN(n2208) );
  IND2D1BWP12T U889 ( .A1(n2350), .B1(n2353), .ZN(n1159) );
  INVD1BWP12T U890 ( .I(n1159), .ZN(n2320) );
  MUX2ND0BWP12T U891 ( .I0(a[3]), .I1(n2352), .S(n1277), .ZN(n1144) );
  INVD1BWP12T U892 ( .I(n1144), .ZN(n1161) );
  IND2D1BWP12T U893 ( .A1(n2353), .B1(n2350), .ZN(n1353) );
  INVD1BWP12T U894 ( .I(n1353), .ZN(n2324) );
  ND2D1BWP12T U895 ( .A1(n2074), .A2(n2740), .ZN(n393) );
  ND2D1BWP12T U896 ( .A1(n2764), .A2(n2740), .ZN(n2258) );
  ND2D1BWP12T U897 ( .A1(n393), .A2(n2258), .ZN(n2892) );
  ND2XD3BWP12T U898 ( .A1(n2134), .A2(n2892), .ZN(n2123) );
  INVD1BWP12T U899 ( .I(n2123), .ZN(n2933) );
  TPND2D0BWP12T U900 ( .A1(op[0]), .A2(op[1]), .ZN(n425) );
  NR2D1BWP12T U901 ( .A1(n433), .A2(n425), .ZN(n3091) );
  ND2D1BWP12T U902 ( .A1(n2101), .A2(n2099), .ZN(n2095) );
  CKND0BWP12T U903 ( .I(n1111), .ZN(n398) );
  INVD1BWP12T U904 ( .I(n2099), .ZN(n394) );
  CKND2BWP12T U905 ( .I(n395), .ZN(n1150) );
  CKND2D1BWP12T U906 ( .A1(n2110), .A2(n1160), .ZN(n397) );
  CKND2D1BWP12T U907 ( .A1(n2109), .A2(n1161), .ZN(n396) );
  OAI211D1BWP12T U908 ( .A1(n2095), .A2(n398), .B(n397), .C(n396), .ZN(n2083)
         );
  INVD1BWP12T U909 ( .I(n2083), .ZN(n2129) );
  AN3D1BWP12T U910 ( .A1(n400), .A2(op[0]), .A3(n399), .Z(n1272) );
  INVD1BWP12T U911 ( .I(n1272), .ZN(n3099) );
  CKND2D0BWP12T U912 ( .A1(op[3]), .A2(op[2]), .ZN(n402) );
  INVD1BWP12T U913 ( .I(n3020), .ZN(n3103) );
  OAI21D1BWP12T U914 ( .A1(n2466), .A2(n3099), .B(n3103), .ZN(n401) );
  CKND2D1BWP12T U915 ( .A1(n401), .A2(n2351), .ZN(n408) );
  NR2D0BWP12T U916 ( .A1(n403), .A2(n402), .ZN(n2215) );
  NR2D1BWP12T U917 ( .A1(n1272), .A2(n2215), .ZN(n3019) );
  INVD1BWP12T U918 ( .I(n3019), .ZN(n3102) );
  INVD1BWP12T U919 ( .I(n3018), .ZN(n3101) );
  MUX2ND0BWP12T U920 ( .I0(n3102), .I1(n3101), .S(n2351), .ZN(n404) );
  CKND2D0BWP12T U921 ( .A1(n404), .A2(n3103), .ZN(n406) );
  CKND2D0BWP12T U922 ( .A1(op[2]), .A2(op[1]), .ZN(n405) );
  NR2D1BWP12T U923 ( .A1(n416), .A2(n405), .ZN(n3105) );
  MUX2ND0BWP12T U924 ( .I0(n406), .I1(n3105), .S(n2206), .ZN(n407) );
  OAI211D1BWP12T U925 ( .A1(n2824), .A2(n2129), .B(n408), .C(n407), .ZN(n409)
         );
  AOI21D1BWP12T U926 ( .A1(n2826), .A2(n2308), .B(n409), .ZN(n422) );
  CKBD1BWP12T U927 ( .I(n1277), .Z(n1270) );
  CKND2D1BWP12T U928 ( .A1(n1270), .A2(n2172), .ZN(n1271) );
  CKBD1BWP12T U929 ( .I(n2349), .Z(n410) );
  NR2D1BWP12T U930 ( .A1(n2350), .A2(n410), .ZN(n1118) );
  ND2D1BWP12T U931 ( .A1(n2350), .A2(n410), .ZN(n1119) );
  OAI21D1BWP12T U932 ( .A1(n1271), .A2(n1118), .B(n1119), .ZN(n1231) );
  CKBD1BWP12T U933 ( .I(a[3]), .Z(n411) );
  NR2D1BWP12T U934 ( .A1(n2764), .A2(n411), .ZN(n1749) );
  NR2D1BWP12T U935 ( .A1(n2353), .A2(n2352), .ZN(n1747) );
  NR2D1BWP12T U936 ( .A1(n1749), .A2(n1747), .ZN(n413) );
  ND2D1BWP12T U937 ( .A1(n2353), .A2(n2352), .ZN(n1746) );
  CKND2D1BWP12T U938 ( .A1(n2764), .A2(n411), .ZN(n1750) );
  OAI21D1BWP12T U939 ( .A1(n1749), .A2(n1746), .B(n1750), .ZN(n412) );
  AOI21D1BWP12T U940 ( .A1(n1231), .A2(n413), .B(n412), .ZN(n865) );
  INVD1BWP12T U941 ( .I(n865), .ZN(n1768) );
  NR2D1BWP12T U942 ( .A1(n2740), .A2(n2738), .ZN(n857) );
  INVD1BWP12T U943 ( .I(n857), .ZN(n1767) );
  ND2D1BWP12T U944 ( .A1(n2740), .A2(n2738), .ZN(n1766) );
  NR2D1BWP12T U945 ( .A1(n2466), .A2(n2351), .ZN(n859) );
  INVD0BWP12T U946 ( .I(n859), .ZN(n414) );
  ND2D1BWP12T U947 ( .A1(n2466), .A2(n2351), .ZN(n858) );
  INVD1BWP12T U948 ( .I(n1762), .ZN(n3093) );
  INVD1BWP12T U949 ( .I(n417), .ZN(n2085) );
  NR2D1BWP12T U950 ( .A1(n1920), .A2(n2216), .ZN(n418) );
  NR2D1BWP12T U951 ( .A1(n1092), .A2(n418), .ZN(n2432) );
  INVD1BWP12T U952 ( .I(n3091), .ZN(n3004) );
  NR2D1BWP12T U953 ( .A1(n2740), .A2(n3004), .ZN(n3090) );
  INVD1BWP12T U954 ( .I(n3090), .ZN(n2807) );
  OAI21D0BWP12T U955 ( .A1(n2600), .A2(n3004), .B(n2807), .ZN(n420) );
  AOI22D0BWP12T U956 ( .A1(n1774), .A2(n3093), .B1(n2085), .B2(n420), .ZN(n421) );
  OAI211D1BWP12T U957 ( .A1(n3047), .A2(n423), .B(n422), .C(n421), .ZN(n436)
         );
  ND2D0BWP12T U958 ( .A1(n2600), .A2(n2740), .ZN(n2084) );
  INVD1BWP12T U959 ( .I(n2084), .ZN(n2390) );
  INVD1BWP12T U960 ( .I(n424), .ZN(n2389) );
  CKND0BWP12T U961 ( .I(n425), .ZN(n427) );
  NR2D0BWP12T U962 ( .A1(op[3]), .A2(op[2]), .ZN(n426) );
  ND2D1BWP12T U963 ( .A1(n427), .A2(n426), .ZN(n2856) );
  CKBD1BWP12T U964 ( .I(n2349), .Z(n428) );
  NR2D1BWP12T U965 ( .A1(n429), .A2(n428), .ZN(n1227) );
  NR2D1BWP12T U966 ( .A1(n1747), .A2(n1227), .ZN(n431) );
  NR2D1BWP12T U967 ( .A1(n2172), .A2(c_in), .ZN(n1273) );
  CKND2D1BWP12T U968 ( .A1(n2172), .A2(c_in), .ZN(n1274) );
  OAI21D1BWP12T U969 ( .A1(n1269), .A2(n1273), .B(n1274), .ZN(n1115) );
  ND2D1BWP12T U970 ( .A1(n429), .A2(n428), .ZN(n1226) );
  OAI21D1BWP12T U971 ( .A1(n1747), .A2(n1226), .B(n1746), .ZN(n430) );
  AOI21D1BWP12T U972 ( .A1(n431), .A2(n1115), .B(n430), .ZN(n833) );
  INVD1BWP12T U973 ( .I(n833), .ZN(n1624) );
  CKBD1BWP12T U974 ( .I(a[3]), .Z(n432) );
  NR2D1BWP12T U975 ( .A1(n2764), .A2(n432), .ZN(n1608) );
  NR2D1BWP12T U976 ( .A1(n1608), .A2(n857), .ZN(n1616) );
  CKND2D1BWP12T U977 ( .A1(n2764), .A2(n432), .ZN(n1613) );
  OAI21D1BWP12T U978 ( .A1(n857), .A2(n1613), .B(n1766), .ZN(n1618) );
  NR2D1BWP12T U979 ( .A1(n2466), .A2(n2351), .ZN(n1620) );
  ND2D1BWP12T U980 ( .A1(n2466), .A2(n2351), .ZN(n1619) );
  CKND2D0BWP12T U981 ( .A1(n1609), .A2(n3082), .ZN(n434) );
  OAI31D1BWP12T U982 ( .A1(n2390), .A2(n2389), .A3(n2856), .B(n434), .ZN(n435)
         );
  XOR2D1BWP12T U983 ( .A1(n2815), .A2(n2785), .Z(n440) );
  XNR2D1BWP12T U984 ( .A1(n883), .A2(n2785), .ZN(n442) );
  INR2D1BWP12T U985 ( .A1(n440), .B1(n442), .ZN(n441) );
  INVD3BWP12T U986 ( .I(n441), .ZN(n2510) );
  XNR2D1BWP12T U987 ( .A1(n2815), .A2(b[13]), .ZN(n569) );
  INVD2BWP12T U988 ( .I(n442), .ZN(n2508) );
  XNR2D1BWP12T U989 ( .A1(n2815), .A2(b[14]), .ZN(n443) );
  OAI22D1BWP12T U990 ( .A1(n2510), .A2(n569), .B1(n2508), .B2(n443), .ZN(
        mult_x_18_n928) );
  XNR2D1BWP12T U991 ( .A1(n2815), .A2(n2876), .ZN(n448) );
  XNR2D1BWP12T U992 ( .A1(n2815), .A2(n3106), .ZN(n445) );
  OAI22D1BWP12T U993 ( .A1(n2510), .A2(n448), .B1(n2508), .B2(n445), .ZN(
        mult_x_18_n932) );
  XNR2D1BWP12T U994 ( .A1(n2815), .A2(n2792), .ZN(n447) );
  XNR2D1BWP12T U995 ( .A1(n2815), .A2(n2817), .ZN(n675) );
  OAI22D1BWP12T U996 ( .A1(n2510), .A2(n447), .B1(n2508), .B2(n675), .ZN(
        mult_x_18_n935) );
  XNR2D1BWP12T U997 ( .A1(n2815), .A2(b[21]), .ZN(n516) );
  XNR2D1BWP12T U998 ( .A1(n2815), .A2(b[22]), .ZN(n450) );
  TPOAI22D0BWP12T U999 ( .A1(n2510), .A2(n516), .B1(n2508), .B2(n450), .ZN(
        mult_x_18_n920) );
  XNR2D1BWP12T U1000 ( .A1(n2815), .A2(b[15]), .ZN(n444) );
  OAI22D1BWP12T U1001 ( .A1(n2510), .A2(n443), .B1(n2508), .B2(n444), .ZN(
        mult_x_18_n927) );
  XNR2D1BWP12T U1002 ( .A1(n2815), .A2(b[16]), .ZN(n607) );
  OAI22D1BWP12T U1003 ( .A1(n2510), .A2(n444), .B1(n2508), .B2(n607), .ZN(
        mult_x_18_n926) );
  XNR2D1BWP12T U1004 ( .A1(n2815), .A2(n2904), .ZN(n446) );
  OAI22D1BWP12T U1005 ( .A1(n2510), .A2(n445), .B1(n2508), .B2(n446), .ZN(
        mult_x_18_n931) );
  XNR2D1BWP12T U1006 ( .A1(n2815), .A2(n2452), .ZN(n570) );
  OAI22D1BWP12T U1007 ( .A1(n2510), .A2(n446), .B1(n2508), .B2(n570), .ZN(
        mult_x_18_n930) );
  XNR2D1BWP12T U1008 ( .A1(n2815), .A2(n2351), .ZN(n549) );
  OAI22D1BWP12T U1009 ( .A1(n2510), .A2(n549), .B1(n2508), .B2(n447), .ZN(
        mult_x_18_n936) );
  XNR2D1BWP12T U1010 ( .A1(n2815), .A2(n2852), .ZN(n674) );
  OAI22D1BWP12T U1011 ( .A1(n2510), .A2(n674), .B1(n2508), .B2(n448), .ZN(
        mult_x_18_n933) );
  INVD4BWP12T U1012 ( .I(n2898), .ZN(n879) );
  INVD8BWP12T U1013 ( .I(n879), .ZN(n2456) );
  XNR2XD4BWP12T U1014 ( .A1(n2456), .A2(a[12]), .ZN(n2493) );
  CKXOR2D1BWP12T U1015 ( .A1(a[13]), .A2(a[12]), .Z(n449) );
  TPND2D3BWP12T U1016 ( .A1(n2493), .A2(n449), .ZN(n2495) );
  XNR2XD1BWP12T U1017 ( .A1(a[13]), .A2(b[18]), .ZN(n722) );
  XNR2D0BWP12T U1018 ( .A1(a[13]), .A2(b[19]), .ZN(n2494) );
  OAI22D0BWP12T U1019 ( .A1(n2495), .A2(n722), .B1(n2493), .B2(n2494), .ZN(
        mult_x_18_n848) );
  XNR2D1BWP12T U1020 ( .A1(n2815), .A2(b[17]), .ZN(n606) );
  XNR2D1BWP12T U1021 ( .A1(n2815), .A2(b[18]), .ZN(n452) );
  OAI22D1BWP12T U1022 ( .A1(n2510), .A2(n606), .B1(n2508), .B2(n452), .ZN(
        mult_x_18_n924) );
  XNR2D1BWP12T U1023 ( .A1(n2815), .A2(b[23]), .ZN(n451) );
  TPOAI22D0BWP12T U1024 ( .A1(n2510), .A2(n450), .B1(n2508), .B2(n451), .ZN(
        mult_x_18_n919) );
  XNR2D1BWP12T U1025 ( .A1(n2815), .A2(b[24]), .ZN(n759) );
  TPOAI22D0BWP12T U1026 ( .A1(n2510), .A2(n451), .B1(n2508), .B2(n759), .ZN(
        mult_x_18_n918) );
  XNR2D1BWP12T U1027 ( .A1(n2815), .A2(b[19]), .ZN(n611) );
  OAI22D1BWP12T U1028 ( .A1(n2510), .A2(n452), .B1(n2508), .B2(n611), .ZN(
        mult_x_18_n923) );
  XNR2D1BWP12T U1029 ( .A1(n2349), .A2(b[28]), .ZN(n470) );
  XNR2D1BWP12T U1030 ( .A1(n2349), .A2(b[29]), .ZN(n720) );
  OAI22D1BWP12T U1031 ( .A1(n2450), .A2(n470), .B1(n720), .B2(n2449), .ZN(n456) );
  INVD1BWP12T U1032 ( .I(n2428), .ZN(n2498) );
  XOR2XD1BWP12T U1033 ( .A1(n2498), .A2(a[28]), .Z(n453) );
  ND2D1BWP12T U1034 ( .A1(n453), .A2(n2500), .ZN(n2502) );
  IND2D0BWP12T U1035 ( .A1(n1277), .B1(n2498), .ZN(n454) );
  OAI22D1BWP12T U1036 ( .A1(n2502), .A2(n2428), .B1(n2500), .B2(n454), .ZN(
        n455) );
  HA1D0BWP12T U1037 ( .A(n456), .B(n455), .CO(mult_x_18_n444), .S(
        mult_x_18_n445) );
  HA1D0BWP12T U1038 ( .A(n458), .B(n457), .CO(mult_x_18_n726), .S(n772) );
  XNR2D2BWP12T U1039 ( .A1(a[20]), .A2(n2621), .ZN(n2453) );
  XOR2D1BWP12T U1040 ( .A1(a[20]), .A2(n2594), .Z(n459) );
  ND2D3BWP12T U1041 ( .A1(n2453), .A2(n459), .ZN(n2455) );
  XNR2D1BWP12T U1042 ( .A1(n2594), .A2(n2876), .ZN(n639) );
  XNR2D1BWP12T U1043 ( .A1(n2594), .A2(n3106), .ZN(n750) );
  TPOAI22D0BWP12T U1044 ( .A1(n2455), .A2(n639), .B1(n2453), .B2(n750), .ZN(
        mult_x_18_n785) );
  XNR2D1BWP12T U1045 ( .A1(n2349), .A2(b[30]), .ZN(n719) );
  XNR2D1BWP12T U1046 ( .A1(n2349), .A2(b[31]), .ZN(n2448) );
  XNR2XD1BWP12T U1047 ( .A1(n2498), .A2(a[30]), .ZN(n2504) );
  INVD1BWP12T U1048 ( .I(n2216), .ZN(n2979) );
  CKXOR2D0BWP12T U1049 ( .A1(n2979), .A2(a[30]), .Z(n460) );
  CKND2D1BWP12T U1050 ( .A1(n2504), .A2(n460), .ZN(n2506) );
  XNR2D2BWP12T U1051 ( .A1(a[14]), .A2(a[13]), .ZN(n2472) );
  XOR2XD1BWP12T U1052 ( .A1(a[14]), .A2(n2710), .Z(n461) );
  TPND2D3BWP12T U1053 ( .A1(n2472), .A2(n461), .ZN(n2474) );
  XNR2D0BWP12T U1054 ( .A1(n2710), .A2(b[15]), .ZN(n714) );
  XNR2XD0BWP12T U1055 ( .A1(n2710), .A2(b[16]), .ZN(n753) );
  TPOAI22D0BWP12T U1056 ( .A1(n2474), .A2(n714), .B1(n2472), .B2(n753), .ZN(
        mult_x_18_n830) );
  XNR2D1BWP12T U1057 ( .A1(n2349), .A2(b[24]), .ZN(n581) );
  OAI22D1BWP12T U1058 ( .A1(n2450), .A2(n462), .B1(n581), .B2(n2449), .ZN(n465) );
  INVD2BWP12T U1059 ( .I(n2574), .ZN(n2571) );
  XNR2D1BWP12T U1060 ( .A1(n2571), .A2(n2541), .ZN(n2461) );
  INR2D1BWP12T U1061 ( .A1(n306), .B1(n2461), .ZN(n464) );
  XNR2D1BWP12T U1062 ( .A1(n2516), .A2(b[21]), .ZN(n706) );
  XNR2D1BWP12T U1063 ( .A1(n2516), .A2(b[22]), .ZN(n484) );
  OAI22D1BWP12T U1064 ( .A1(n2520), .A2(n706), .B1(n2518), .B2(n484), .ZN(n463) );
  FA1D0BWP12T U1065 ( .A(n465), .B(n464), .CI(n463), .CO(mult_x_18_n538), .S(
        mult_x_18_n539) );
  INR2D1BWP12T U1066 ( .A1(n1277), .B1(n2508), .ZN(mult_x_18_n942) );
  XNR2XD4BWP12T U1067 ( .A1(a[22]), .A2(n2594), .ZN(n2490) );
  INR2D1BWP12T U1068 ( .A1(n306), .B1(n2490), .ZN(mult_x_18_n782) );
  IND2D0BWP12T U1069 ( .A1(n306), .B1(a[13]), .ZN(n466) );
  OAI22D1BWP12T U1070 ( .A1(n2495), .A2(n3059), .B1(n2493), .B2(n466), .ZN(
        n469) );
  XNR2D1BWP12T U1071 ( .A1(n2466), .A2(n2852), .ZN(n671) );
  XNR2D1BWP12T U1072 ( .A1(n2466), .A2(n2876), .ZN(n724) );
  OAI22D1BWP12T U1073 ( .A1(n2469), .A2(n671), .B1(n724), .B2(n2467), .ZN(n468) );
  XNR2D1BWP12T U1074 ( .A1(n2516), .A2(n3106), .ZN(n491) );
  XNR2D1BWP12T U1075 ( .A1(n2516), .A2(n2904), .ZN(n587) );
  OAI22D1BWP12T U1076 ( .A1(n2520), .A2(n491), .B1(n2518), .B2(n587), .ZN(n467) );
  FA1D0BWP12T U1077 ( .A(n469), .B(n468), .CI(n467), .CO(mult_x_18_n678), .S(
        mult_x_18_n679) );
  OAI22D1BWP12T U1078 ( .A1(n2450), .A2(n550), .B1(n470), .B2(n2449), .ZN(n473) );
  INR2D1BWP12T U1079 ( .A1(n1277), .B1(n2500), .ZN(n472) );
  XNR2D1BWP12T U1080 ( .A1(n2516), .A2(b[25]), .ZN(n548) );
  XNR2D1BWP12T U1081 ( .A1(n2516), .A2(b[26]), .ZN(n512) );
  OAI22D1BWP12T U1082 ( .A1(n2520), .A2(n548), .B1(n2518), .B2(n512), .ZN(n471) );
  FA1D0BWP12T U1083 ( .A(n473), .B(n472), .CI(n471), .CO(mult_x_18_n464), .S(
        mult_x_18_n465) );
  INR2D1BWP12T U1084 ( .A1(n306), .B1(n2457), .ZN(mult_x_18_n890) );
  IND2D1BWP12T U1085 ( .A1(n306), .B1(n2594), .ZN(n474) );
  TPOAI22D1BWP12T U1086 ( .A1(n2455), .A2(n475), .B1(n2453), .B2(n474), .ZN(
        n479) );
  XOR2D1BWP12T U1087 ( .A1(n2456), .A2(n3100), .Z(n476) );
  TPND2D8BWP12T U1088 ( .A1(n476), .A2(n2457), .ZN(n2459) );
  XNR2D1BWP12T U1089 ( .A1(n2456), .A2(n3106), .ZN(n667) );
  XNR2D1BWP12T U1090 ( .A1(n2456), .A2(n2904), .ZN(n633) );
  OAI22D1BWP12T U1091 ( .A1(n2459), .A2(n667), .B1(n633), .B2(n2457), .ZN(n478) );
  XNR2D1BWP12T U1092 ( .A1(n2516), .A2(b[18]), .ZN(n507) );
  XNR2D1BWP12T U1093 ( .A1(n2516), .A2(b[19]), .ZN(n688) );
  OAI22D1BWP12T U1094 ( .A1(n2520), .A2(n507), .B1(n2518), .B2(n688), .ZN(n477) );
  FA1D0BWP12T U1095 ( .A(n479), .B(n478), .CI(n477), .CO(mult_x_18_n584), .S(
        mult_x_18_n585) );
  XNR2D1BWP12T U1096 ( .A1(n2349), .A2(b[15]), .ZN(n642) );
  XNR2D1BWP12T U1097 ( .A1(n2349), .A2(b[16]), .ZN(n593) );
  OAI22D1BWP12T U1098 ( .A1(n2450), .A2(n642), .B1(n593), .B2(n2449), .ZN(n482) );
  INR2D1BWP12T U1099 ( .A1(n1277), .B1(n2511), .ZN(n481) );
  XNR2D1BWP12T U1100 ( .A1(n2516), .A2(b[13]), .ZN(n652) );
  XNR2D1BWP12T U1101 ( .A1(n2516), .A2(b[14]), .ZN(n496) );
  OAI22D1BWP12T U1102 ( .A1(n2520), .A2(n652), .B1(n2518), .B2(n496), .ZN(n480) );
  FA1D0BWP12T U1103 ( .A(n482), .B(n481), .CI(n480), .CO(mult_x_18_n650), .S(
        mult_x_18_n651) );
  INR2D1BWP12T U1104 ( .A1(n1277), .B1(n2476), .ZN(mult_x_18_n762) );
  XNR2D1BWP12T U1105 ( .A1(n2456), .A2(b[14]), .ZN(n546) );
  XNR2D1BWP12T U1106 ( .A1(n2456), .A2(b[15]), .ZN(n542) );
  OAI22D1BWP12T U1107 ( .A1(n2459), .A2(n546), .B1(n542), .B2(n2457), .ZN(n487) );
  XOR2D1BWP12T U1108 ( .A1(n2571), .A2(a[22]), .Z(n483) );
  ND2D1BWP12T U1109 ( .A1(n2490), .A2(n483), .ZN(n2492) );
  XNR2D1BWP12T U1110 ( .A1(n2571), .A2(n2353), .ZN(n522) );
  XNR2D1BWP12T U1111 ( .A1(n2764), .A2(n2571), .ZN(n613) );
  OAI22D1BWP12T U1112 ( .A1(n2492), .A2(n522), .B1(n613), .B2(n2490), .ZN(n486) );
  XNR2D1BWP12T U1113 ( .A1(n2516), .A2(b[23]), .ZN(n558) );
  OAI22D1BWP12T U1114 ( .A1(n2520), .A2(n484), .B1(n2518), .B2(n558), .ZN(n485) );
  FA1D0BWP12T U1115 ( .A(n487), .B(n486), .CI(n485), .CO(mult_x_18_n519), .S(
        mult_x_18_n520) );
  XNR2D1BWP12T U1116 ( .A1(n2817), .A2(n2349), .ZN(n533) );
  XNR2D1BWP12T U1117 ( .A1(n2349), .A2(n2852), .ZN(n518) );
  OAI22D1BWP12T U1118 ( .A1(n2450), .A2(n533), .B1(n518), .B2(n2449), .ZN(n490) );
  INR2D1BWP12T U1119 ( .A1(n306), .B1(n2487), .ZN(n489) );
  XNR2D1BWP12T U1120 ( .A1(n2516), .A2(n2351), .ZN(n634) );
  XNR2D1BWP12T U1121 ( .A1(n2516), .A2(n2792), .ZN(n502) );
  OAI22D1BWP12T U1122 ( .A1(n2520), .A2(n634), .B1(n2518), .B2(n502), .ZN(n488) );
  FA1D0BWP12T U1123 ( .A(n490), .B(n489), .CI(n488), .CO(mult_x_18_n714), .S(
        mult_x_18_n715) );
  INR2D1BWP12T U1124 ( .A1(n306), .B1(n2482), .ZN(mult_x_18_n810) );
  XNR2D1BWP12T U1125 ( .A1(n2349), .A2(n2904), .ZN(n614) );
  XNR2D1BWP12T U1126 ( .A1(n2349), .A2(n2452), .ZN(n589) );
  OAI22D1BWP12T U1127 ( .A1(n2450), .A2(n614), .B1(n589), .B2(n2449), .ZN(n494) );
  INR2D1BWP12T U1128 ( .A1(n1277), .B1(n2493), .ZN(n493) );
  XNR2D1BWP12T U1129 ( .A1(n2516), .A2(n2876), .ZN(n655) );
  FA1D0BWP12T U1130 ( .A(n494), .B(n493), .CI(n492), .CO(mult_x_18_n688), .S(
        mult_x_18_n689) );
  XNR2D1BWP12T U1131 ( .A1(n2456), .A2(n2792), .ZN(n762) );
  XNR2D1BWP12T U1132 ( .A1(n2456), .A2(n2817), .ZN(n636) );
  OAI22D1BWP12T U1133 ( .A1(n2459), .A2(n762), .B1(n636), .B2(n2457), .ZN(n499) );
  XNR2D1BWP12T U1134 ( .A1(n2679), .A2(n306), .ZN(n495) );
  XNR2D1BWP12T U1135 ( .A1(n2679), .A2(n429), .ZN(n625) );
  OAI22D1BWP12T U1136 ( .A1(n2513), .A2(n495), .B1(n625), .B2(n2511), .ZN(n498) );
  XNR2D1BWP12T U1137 ( .A1(n2516), .A2(b[15]), .ZN(n545) );
  OAI22D1BWP12T U1138 ( .A1(n2520), .A2(n496), .B1(n2518), .B2(n545), .ZN(n497) );
  FA1D0BWP12T U1139 ( .A(n499), .B(n498), .CI(n497), .CO(mult_x_18_n637), .S(
        mult_x_18_n638) );
  INVD1BWP12T U1140 ( .I(n2870), .ZN(n877) );
  IND2D1BWP12T U1141 ( .A1(n306), .B1(n2870), .ZN(n500) );
  OAI22D1BWP12T U1142 ( .A1(n2489), .A2(n877), .B1(n2487), .B2(n500), .ZN(n505) );
  XNR2D1BWP12T U1143 ( .A1(n1277), .A2(n2870), .ZN(n501) );
  XNR2D1BWP12T U1144 ( .A1(n429), .A2(n2870), .ZN(n566) );
  OAI22D1BWP12T U1145 ( .A1(n2489), .A2(n501), .B1(n2487), .B2(n566), .ZN(n504) );
  XNR2D1BWP12T U1146 ( .A1(n2516), .A2(n2817), .ZN(n705) );
  OAI22D1BWP12T U1147 ( .A1(n2520), .A2(n502), .B1(n2518), .B2(n705), .ZN(n503) );
  FA1D0BWP12T U1148 ( .A(n505), .B(n504), .CI(n503), .CO(mult_x_18_n707), .S(
        mult_x_18_n708) );
  XNR2D1BWP12T U1149 ( .A1(n2349), .A2(b[20]), .ZN(n576) );
  OAI22D1BWP12T U1150 ( .A1(n2450), .A2(n506), .B1(n576), .B2(n2449), .ZN(n510) );
  INR2D1BWP12T U1151 ( .A1(n1270), .B1(n2453), .ZN(n509) );
  XNR2D1BWP12T U1152 ( .A1(n2516), .A2(b[17]), .ZN(n659) );
  OAI22D1BWP12T U1153 ( .A1(n2520), .A2(n659), .B1(n2518), .B2(n507), .ZN(n508) );
  FA1D0BWP12T U1154 ( .A(n510), .B(n509), .CI(n508), .CO(mult_x_18_n600), .S(
        mult_x_18_n601) );
  XNR2D1BWP12T U1155 ( .A1(n2571), .A2(n2792), .ZN(n599) );
  XNR2D1BWP12T U1156 ( .A1(n2571), .A2(n2817), .ZN(n742) );
  OAI22D1BWP12T U1157 ( .A1(n2492), .A2(n599), .B1(n742), .B2(n2490), .ZN(n515) );
  XNR2XD1BWP12T U1158 ( .A1(n306), .A2(n2498), .ZN(n511) );
  XNR2XD1BWP12T U1159 ( .A1(n2498), .A2(b[1]), .ZN(n713) );
  OAI22D1BWP12T U1160 ( .A1(n2502), .A2(n511), .B1(n713), .B2(n2500), .ZN(n514) );
  OAI22D1BWP12T U1161 ( .A1(n2520), .A2(n512), .B1(n2518), .B2(n725), .ZN(n513) );
  FA1D0BWP12T U1162 ( .A(n515), .B(n514), .CI(n513), .CO(mult_x_18_n442), .S(
        mult_x_18_n443) );
  INR2D1BWP12T U1163 ( .A1(n306), .B1(n2504), .ZN(mult_x_18_n750) );
  INR2D1BWP12T U1164 ( .A1(n1277), .B1(n2472), .ZN(mult_x_18_n846) );
  XNR2D1BWP12T U1165 ( .A1(n2815), .A2(b[20]), .ZN(n610) );
  OAI22D1BWP12T U1166 ( .A1(n2510), .A2(n610), .B1(n2508), .B2(n516), .ZN(
        mult_x_18_n921) );
  XNR2D1BWP12T U1167 ( .A1(n2571), .A2(n2499), .ZN(n612) );
  XNR2D1BWP12T U1168 ( .A1(n2571), .A2(n2351), .ZN(n600) );
  OAI22D1BWP12T U1169 ( .A1(n2492), .A2(n612), .B1(n600), .B2(n2490), .ZN(
        mult_x_18_n777) );
  XNR2D1BWP12T U1170 ( .A1(n1277), .A2(n2571), .ZN(n517) );
  XNR2D1BWP12T U1171 ( .A1(n2571), .A2(n429), .ZN(n523) );
  OAI22D1BWP12T U1172 ( .A1(n2492), .A2(n517), .B1(n523), .B2(n2490), .ZN(
        mult_x_18_n781) );
  XNR2D1BWP12T U1173 ( .A1(n2349), .A2(n2876), .ZN(n524) );
  OAI22D1BWP12T U1174 ( .A1(n2450), .A2(n518), .B1(n524), .B2(n2449), .ZN(n520) );
  XNR2D1BWP12T U1175 ( .A1(n2466), .A2(n2499), .ZN(n527) );
  XNR2D1BWP12T U1176 ( .A1(n2466), .A2(n2351), .ZN(n539) );
  OAI22D1BWP12T U1177 ( .A1(n2469), .A2(n527), .B1(n539), .B2(n2467), .ZN(n519) );
  XNR2XD1BWP12T U1178 ( .A1(n429), .A2(n2358), .ZN(n622) );
  XNR2D1BWP12T U1179 ( .A1(n2503), .A2(n2358), .ZN(n651) );
  OAI22D1BWP12T U1180 ( .A1(n2478), .A2(n622), .B1(n651), .B2(n2476), .ZN(
        mult_x_18_n760) );
  XNR2D1BWP12T U1181 ( .A1(n2466), .A2(b[16]), .ZN(n702) );
  XNR2D1BWP12T U1182 ( .A1(n2466), .A2(b[17]), .ZN(n565) );
  OAI22D1BWP12T U1183 ( .A1(n2469), .A2(n702), .B1(n565), .B2(n2467), .ZN(
        mult_x_18_n954) );
  XNR2D1BWP12T U1184 ( .A1(n2349), .A2(b[21]), .ZN(n575) );
  OAI22D1BWP12T U1185 ( .A1(n2450), .A2(n575), .B1(n521), .B2(n2449), .ZN(
        mult_x_18_n1013) );
  OAI22D1BWP12T U1186 ( .A1(n2492), .A2(n523), .B1(n522), .B2(n2490), .ZN(
        mult_x_18_n780) );
  XNR2D1BWP12T U1187 ( .A1(n2349), .A2(n3106), .ZN(n615) );
  OAI22D1BWP12T U1188 ( .A1(n2450), .A2(n524), .B1(n615), .B2(n2449), .ZN(
        mult_x_18_n1025) );
  XNR2D1BWP12T U1189 ( .A1(n2466), .A2(b[14]), .ZN(n571) );
  XNR2D1BWP12T U1190 ( .A1(n2466), .A2(b[15]), .ZN(n703) );
  OAI22D1BWP12T U1191 ( .A1(n2469), .A2(n571), .B1(n703), .B2(n2467), .ZN(
        mult_x_18_n956) );
  XNR2D1BWP12T U1192 ( .A1(n2349), .A2(b[17]), .ZN(n592) );
  OAI22D1BWP12T U1193 ( .A1(n2450), .A2(n592), .B1(n525), .B2(n2449), .ZN(
        mult_x_18_n1017) );
  OR2D0BWP12T U1194 ( .A1(n1277), .A2(n2201), .Z(n526) );
  OAI22D1BWP12T U1195 ( .A1(n2478), .A2(n2201), .B1(n2476), .B2(n526), .ZN(
        mult_x_18_n734) );
  XNR2D1BWP12T U1196 ( .A1(n2349), .A2(b[25]), .ZN(n580) );
  XNR2D1BWP12T U1197 ( .A1(n2349), .A2(b[26]), .ZN(n551) );
  OAI22D1BWP12T U1198 ( .A1(n2450), .A2(n580), .B1(n551), .B2(n2449), .ZN(
        mult_x_18_n1009) );
  XNR2XD1BWP12T U1199 ( .A1(n2679), .A2(n2904), .ZN(n552) );
  XNR2XD1BWP12T U1200 ( .A1(n2679), .A2(n2452), .ZN(n605) );
  OAI22D1BWP12T U1201 ( .A1(n2513), .A2(n552), .B1(n605), .B2(n2511), .ZN(
        mult_x_18_n815) );
  XNR2D1BWP12T U1202 ( .A1(n2466), .A2(n2764), .ZN(n534) );
  OAI22D1BWP12T U1203 ( .A1(n2469), .A2(n534), .B1(n527), .B2(n2467), .ZN(
        mult_x_18_n967) );
  XNR2D1BWP12T U1204 ( .A1(n306), .A2(n2815), .ZN(n528) );
  XNR2D1BWP12T U1205 ( .A1(n429), .A2(n2815), .ZN(n603) );
  OAI22D1BWP12T U1206 ( .A1(n2510), .A2(n528), .B1(n2508), .B2(n603), .ZN(
        mult_x_18_n941) );
  XNR2XD1BWP12T U1207 ( .A1(a[13]), .A2(b[13]), .ZN(n648) );
  XNR2XD1BWP12T U1208 ( .A1(a[13]), .A2(b[14]), .ZN(n654) );
  OAI22D1BWP12T U1209 ( .A1(n2495), .A2(n648), .B1(n2493), .B2(n654), .ZN(
        mult_x_18_n853) );
  XNR2D1BWP12T U1210 ( .A1(n2466), .A2(n2353), .ZN(n535) );
  OAI22D1BWP12T U1211 ( .A1(n2469), .A2(n529), .B1(n535), .B2(n2467), .ZN(
        mult_x_18_n969) );
  XNR2XD1BWP12T U1212 ( .A1(a[13]), .A2(n2876), .ZN(n740) );
  XNR2D1BWP12T U1213 ( .A1(a[13]), .A2(n3106), .ZN(n530) );
  OAI22D1BWP12T U1214 ( .A1(n2495), .A2(n740), .B1(n2493), .B2(n530), .ZN(
        mult_x_18_n857) );
  XNR2D1BWP12T U1215 ( .A1(n2466), .A2(b[22]), .ZN(n531) );
  XNR2D1BWP12T U1216 ( .A1(n2466), .A2(b[23]), .ZN(n541) );
  OAI22D1BWP12T U1217 ( .A1(n2469), .A2(n531), .B1(n541), .B2(n2467), .ZN(
        mult_x_18_n948) );
  XNR2D1BWP12T U1218 ( .A1(n2466), .A2(b[20]), .ZN(n544) );
  XNR2D1BWP12T U1219 ( .A1(n2466), .A2(b[21]), .ZN(n532) );
  OAI22D1BWP12T U1220 ( .A1(n2469), .A2(n544), .B1(n532), .B2(n2467), .ZN(
        mult_x_18_n950) );
  XNR2D1BWP12T U1221 ( .A1(n2466), .A2(n2452), .ZN(n556) );
  XNR2D1BWP12T U1222 ( .A1(n2466), .A2(b[13]), .ZN(n572) );
  OAI22D1BWP12T U1223 ( .A1(n2469), .A2(n556), .B1(n572), .B2(n2467), .ZN(
        mult_x_18_n958) );
  XNR2D1BWP12T U1224 ( .A1(a[13]), .A2(n2904), .ZN(n670) );
  OAI22D1BWP12T U1225 ( .A1(n2495), .A2(n530), .B1(n2493), .B2(n670), .ZN(
        mult_x_18_n856) );
  OAI22D1BWP12T U1226 ( .A1(n2469), .A2(n532), .B1(n531), .B2(n2467), .ZN(
        mult_x_18_n949) );
  XNR2D1BWP12T U1227 ( .A1(n2792), .A2(n2349), .ZN(n563) );
  OAI22D1BWP12T U1228 ( .A1(n2450), .A2(n563), .B1(n533), .B2(n2449), .ZN(n537) );
  OAI22D1BWP12T U1229 ( .A1(n2469), .A2(n535), .B1(n534), .B2(n2467), .ZN(n536) );
  IND2D1BWP12T U1230 ( .A1(n306), .B1(n2815), .ZN(n538) );
  OAI22D1BWP12T U1231 ( .A1(n2510), .A2(n884), .B1(n2508), .B2(n538), .ZN(
        mult_x_18_n744) );
  XNR2D1BWP12T U1232 ( .A1(n2870), .A2(b[19]), .ZN(n728) );
  XNR2D1BWP12T U1233 ( .A1(n2870), .A2(b[20]), .ZN(n627) );
  OAI22D1BWP12T U1234 ( .A1(n2489), .A2(n728), .B1(n2487), .B2(n627), .ZN(
        mult_x_18_n895) );
  XNR2D1BWP12T U1235 ( .A1(n2466), .A2(n2792), .ZN(n567) );
  OAI22D1BWP12T U1236 ( .A1(n2469), .A2(n539), .B1(n567), .B2(n2467), .ZN(
        mult_x_18_n965) );
  XOR2D1BWP12T U1237 ( .A1(n2460), .A2(n2541), .Z(n540) );
  TPND2D2BWP12T U1238 ( .A1(n2461), .A2(n540), .ZN(n2463) );
  XNR2XD1BWP12T U1239 ( .A1(n2764), .A2(n2460), .ZN(n656) );
  XNR2XD1BWP12T U1240 ( .A1(n2499), .A2(n2460), .ZN(n629) );
  OAI22D1BWP12T U1241 ( .A1(n2463), .A2(n656), .B1(n2461), .B2(n629), .ZN(
        mult_x_18_n767) );
  XNR2D1BWP12T U1242 ( .A1(n2466), .A2(b[24]), .ZN(n609) );
  OAI22D1BWP12T U1243 ( .A1(n2469), .A2(n541), .B1(n609), .B2(n2467), .ZN(
        mult_x_18_n947) );
  XNR2D1BWP12T U1244 ( .A1(n2456), .A2(b[16]), .ZN(n547) );
  OAI22D1BWP12T U1245 ( .A1(n2459), .A2(n542), .B1(n547), .B2(n2457), .ZN(
        mult_x_18_n874) );
  XNR2XD1BWP12T U1246 ( .A1(n2679), .A2(n2876), .ZN(n582) );
  XNR2XD1BWP12T U1247 ( .A1(n2679), .A2(n3106), .ZN(n553) );
  OAI22D1BWP12T U1248 ( .A1(n2513), .A2(n582), .B1(n553), .B2(n2511), .ZN(
        mult_x_18_n817) );
  XNR2XD1BWP12T U1249 ( .A1(n2679), .A2(n2351), .ZN(n577) );
  OAI22D1BWP12T U1250 ( .A1(n2513), .A2(n577), .B1(n543), .B2(n2511), .ZN(
        mult_x_18_n821) );
  XNR2D1BWP12T U1251 ( .A1(n2456), .A2(b[18]), .ZN(n692) );
  XNR2D1BWP12T U1252 ( .A1(n2456), .A2(b[19]), .ZN(n745) );
  OAI22D1BWP12T U1253 ( .A1(n2459), .A2(n692), .B1(n745), .B2(n2457), .ZN(
        mult_x_18_n871) );
  XNR2D1BWP12T U1254 ( .A1(n2466), .A2(b[19]), .ZN(n573) );
  OAI22D1BWP12T U1255 ( .A1(n2469), .A2(n573), .B1(n544), .B2(n2467), .ZN(
        mult_x_18_n951) );
  XNR2D1BWP12T U1256 ( .A1(n2516), .A2(b[16]), .ZN(n660) );
  OAI22D1BWP12T U1257 ( .A1(n2520), .A2(n545), .B1(n2518), .B2(n660), .ZN(
        mult_x_18_n986) );
  XNR2D1BWP12T U1258 ( .A1(n2456), .A2(b[13]), .ZN(n561) );
  OAI22D1BWP12T U1259 ( .A1(n2459), .A2(n561), .B1(n546), .B2(n2457), .ZN(
        mult_x_18_n876) );
  XNR2D1BWP12T U1260 ( .A1(n2456), .A2(b[17]), .ZN(n693) );
  OAI22D1BWP12T U1261 ( .A1(n2459), .A2(n547), .B1(n693), .B2(n2457), .ZN(
        mult_x_18_n873) );
  XNR2D1BWP12T U1262 ( .A1(n2594), .A2(n2792), .ZN(n676) );
  XNR2D1BWP12T U1263 ( .A1(n2594), .A2(n2817), .ZN(n560) );
  OAI22D1BWP12T U1264 ( .A1(n2455), .A2(n676), .B1(n2453), .B2(n560), .ZN(
        mult_x_18_n788) );
  XNR2D1BWP12T U1265 ( .A1(n2516), .A2(b[24]), .ZN(n557) );
  OAI22D1BWP12T U1266 ( .A1(n2520), .A2(n557), .B1(n2518), .B2(n548), .ZN(
        mult_x_18_n977) );
  XNR2D1BWP12T U1267 ( .A1(n2499), .A2(n2815), .ZN(n598) );
  OAI22D1BWP12T U1268 ( .A1(n2510), .A2(n598), .B1(n2508), .B2(n549), .ZN(
        mult_x_18_n937) );
  OAI22D1BWP12T U1269 ( .A1(n2450), .A2(n551), .B1(n550), .B2(n2449), .ZN(n555) );
  OAI22D1BWP12T U1270 ( .A1(n2513), .A2(n553), .B1(n552), .B2(n2511), .ZN(n554) );
  XNR2D1BWP12T U1271 ( .A1(n2466), .A2(n2904), .ZN(n768) );
  OAI22D1BWP12T U1272 ( .A1(n2469), .A2(n768), .B1(n556), .B2(n2467), .ZN(
        mult_x_18_n959) );
  XNR2XD1BWP12T U1273 ( .A1(n2621), .A2(n2792), .ZN(n559) );
  XNR2D1BWP12T U1274 ( .A1(n2621), .A2(n2817), .ZN(n689) );
  OAI22D1BWP12T U1275 ( .A1(n2484), .A2(n559), .B1(n2482), .B2(n689), .ZN(
        mult_x_18_n803) );
  OAI22D1BWP12T U1276 ( .A1(n2520), .A2(n558), .B1(n2518), .B2(n557), .ZN(
        mult_x_18_n978) );
  XNR2D1BWP12T U1277 ( .A1(n2349), .A2(b[13]), .ZN(n588) );
  XNR2D1BWP12T U1278 ( .A1(n2349), .A2(b[14]), .ZN(n643) );
  OAI22D1BWP12T U1279 ( .A1(n2450), .A2(n588), .B1(n643), .B2(n2449), .ZN(
        mult_x_18_n1021) );
  XNR2XD1BWP12T U1280 ( .A1(n2621), .A2(n2351), .ZN(n738) );
  OAI22D1BWP12T U1281 ( .A1(n2484), .A2(n738), .B1(n2482), .B2(n559), .ZN(
        mult_x_18_n804) );
  XNR2D1BWP12T U1282 ( .A1(n2710), .A2(n2852), .ZN(n736) );
  XNR2XD1BWP12T U1283 ( .A1(n2710), .A2(n2876), .ZN(n638) );
  OAI22D1BWP12T U1284 ( .A1(n2474), .A2(n736), .B1(n2472), .B2(n638), .ZN(
        mult_x_18_n837) );
  XNR2D1BWP12T U1285 ( .A1(n2870), .A2(b[13]), .ZN(n682) );
  XNR2D1BWP12T U1286 ( .A1(n2870), .A2(b[14]), .ZN(n666) );
  OAI22D1BWP12T U1287 ( .A1(n2489), .A2(n682), .B1(n2487), .B2(n666), .ZN(
        mult_x_18_n901) );
  XNR2D1BWP12T U1288 ( .A1(n2594), .A2(n2852), .ZN(n640) );
  OAI22D1BWP12T U1289 ( .A1(n2455), .A2(n560), .B1(n2453), .B2(n640), .ZN(
        mult_x_18_n787) );
  XNR2D1BWP12T U1290 ( .A1(n2456), .A2(n2452), .ZN(n632) );
  OAI22D1BWP12T U1291 ( .A1(n2459), .A2(n632), .B1(n561), .B2(n2457), .ZN(
        mult_x_18_n877) );
  XNR2D1BWP12T U1292 ( .A1(n2456), .A2(n306), .ZN(n562) );
  XNR2D1BWP12T U1293 ( .A1(n2456), .A2(n429), .ZN(n765) );
  OAI22D1BWP12T U1294 ( .A1(n2459), .A2(n562), .B1(n765), .B2(n2457), .ZN(
        mult_x_18_n889) );
  OAI22D1BWP12T U1295 ( .A1(n2450), .A2(n564), .B1(n563), .B2(n2449), .ZN(
        mult_x_18_n1029) );
  XNR2D1BWP12T U1296 ( .A1(n2466), .A2(b[18]), .ZN(n574) );
  OAI22D1BWP12T U1297 ( .A1(n2469), .A2(n565), .B1(n574), .B2(n2467), .ZN(
        mult_x_18_n953) );
  XNR2D1BWP12T U1298 ( .A1(n2503), .A2(n2870), .ZN(n687) );
  OAI22D1BWP12T U1299 ( .A1(n2489), .A2(n566), .B1(n2487), .B2(n687), .ZN(
        mult_x_18_n913) );
  XNR2D1BWP12T U1300 ( .A1(n2466), .A2(n2817), .ZN(n672) );
  OAI22D1BWP12T U1301 ( .A1(n2469), .A2(n567), .B1(n672), .B2(n2467), .ZN(
        mult_x_18_n964) );
  XNR2XD1BWP12T U1302 ( .A1(n2679), .A2(n2852), .ZN(n583) );
  OAI22D1BWP12T U1303 ( .A1(n2513), .A2(n568), .B1(n583), .B2(n2511), .ZN(
        mult_x_18_n819) );
  OAI22D1BWP12T U1304 ( .A1(n2510), .A2(n570), .B1(n2508), .B2(n569), .ZN(
        mult_x_18_n929) );
  OAI22D1BWP12T U1305 ( .A1(n2469), .A2(n572), .B1(n571), .B2(n2467), .ZN(
        mult_x_18_n957) );
  XNR2D1BWP12T U1306 ( .A1(n2764), .A2(n2870), .ZN(n686) );
  XNR2D1BWP12T U1307 ( .A1(n2499), .A2(n2870), .ZN(n647) );
  OAI22D1BWP12T U1308 ( .A1(n2489), .A2(n686), .B1(n2487), .B2(n647), .ZN(
        mult_x_18_n911) );
  OAI22D1BWP12T U1309 ( .A1(n2469), .A2(n574), .B1(n573), .B2(n2467), .ZN(
        mult_x_18_n952) );
  OAI22D1BWP12T U1310 ( .A1(n2450), .A2(n576), .B1(n575), .B2(n2449), .ZN(n579) );
  XNR2D1BWP12T U1311 ( .A1(n2679), .A2(n2499), .ZN(n630) );
  TPOAI22D1BWP12T U1312 ( .A1(n2513), .A2(n630), .B1(n577), .B2(n2511), .ZN(
        n578) );
  HA1D1BWP12T U1313 ( .A(n579), .B(n578), .CO(mult_x_18_n586), .S(
        mult_x_18_n587) );
  OAI22D1BWP12T U1314 ( .A1(n2450), .A2(n581), .B1(n580), .B2(n2449), .ZN(n585) );
  OAI22D1BWP12T U1315 ( .A1(n2513), .A2(n583), .B1(n582), .B2(n2511), .ZN(n584) );
  XNR2XD1BWP12T U1316 ( .A1(n306), .A2(a[13]), .ZN(n586) );
  OAI22D1BWP12T U1317 ( .A1(n2495), .A2(n586), .B1(n2493), .B2(n767), .ZN(
        mult_x_18_n866) );
  XNR2D1BWP12T U1318 ( .A1(n2764), .A2(n2594), .ZN(n608) );
  XNR2D1BWP12T U1319 ( .A1(n2499), .A2(n2594), .ZN(n619) );
  OAI22D1BWP12T U1320 ( .A1(n2455), .A2(n608), .B1(n2453), .B2(n619), .ZN(
        mult_x_18_n791) );
  XNR2D1BWP12T U1321 ( .A1(n2870), .A2(b[15]), .ZN(n665) );
  XNR2D1BWP12T U1322 ( .A1(n2870), .A2(b[16]), .ZN(n602) );
  OAI22D1BWP12T U1323 ( .A1(n2489), .A2(n665), .B1(n2487), .B2(n602), .ZN(
        mult_x_18_n899) );
  XNR2D1BWP12T U1324 ( .A1(n2516), .A2(n2452), .ZN(n653) );
  OAI22D1BWP12T U1325 ( .A1(n2520), .A2(n587), .B1(n2518), .B2(n653), .ZN(
        mult_x_18_n990) );
  OAI22D1BWP12T U1326 ( .A1(n2450), .A2(n589), .B1(n588), .B2(n2449), .ZN(n591) );
  XNR2D1BWP12T U1327 ( .A1(n2456), .A2(n2353), .ZN(n764) );
  XNR2D1BWP12T U1328 ( .A1(n2456), .A2(n2764), .ZN(n761) );
  OAI22D1BWP12T U1329 ( .A1(n2459), .A2(n764), .B1(n761), .B2(n2457), .ZN(n590) );
  HA1D1BWP12T U1330 ( .A(n591), .B(n590), .CO(mult_x_18_n680), .S(
        mult_x_18_n681) );
  XNR2XD1BWP12T U1331 ( .A1(a[13]), .A2(n2351), .ZN(n641) );
  XNR2D1BWP12T U1332 ( .A1(a[13]), .A2(n2792), .ZN(n646) );
  OAI22D1BWP12T U1333 ( .A1(n2495), .A2(n641), .B1(n2493), .B2(n646), .ZN(
        mult_x_18_n861) );
  OAI22D1BWP12T U1334 ( .A1(n2450), .A2(n593), .B1(n592), .B2(n2449), .ZN(n597) );
  CKND0BWP12T U1335 ( .I(n2679), .ZN(n595) );
  IND2D0BWP12T U1336 ( .A1(n1277), .B1(n2679), .ZN(n594) );
  OAI22D1BWP12T U1337 ( .A1(n2513), .A2(n595), .B1(n2511), .B2(n594), .ZN(n596) );
  HA1D1BWP12T U1338 ( .A(n597), .B(n596), .CO(mult_x_18_n639), .S(
        mult_x_18_n640) );
  XNR2D1BWP12T U1339 ( .A1(n2764), .A2(n2815), .ZN(n620) );
  OAI22D1BWP12T U1340 ( .A1(n2510), .A2(n620), .B1(n2508), .B2(n598), .ZN(
        mult_x_18_n938) );
  OAI22D1BWP12T U1341 ( .A1(n2492), .A2(n600), .B1(n599), .B2(n2490), .ZN(
        mult_x_18_n776) );
  XNR2XD1BWP12T U1342 ( .A1(n306), .A2(n2460), .ZN(n601) );
  XNR2XD1BWP12T U1343 ( .A1(n2350), .A2(n2460), .ZN(n649) );
  OAI22D1BWP12T U1344 ( .A1(n2463), .A2(n601), .B1(n2461), .B2(n649), .ZN(
        mult_x_18_n770) );
  XNR2D1BWP12T U1345 ( .A1(n2870), .A2(b[17]), .ZN(n604) );
  OAI22D1BWP12T U1346 ( .A1(n2489), .A2(n602), .B1(n2487), .B2(n604), .ZN(
        mult_x_18_n898) );
  XNR2D1BWP12T U1347 ( .A1(n2503), .A2(n2815), .ZN(n621) );
  OAI22D1BWP12T U1348 ( .A1(n2510), .A2(n603), .B1(n2508), .B2(n621), .ZN(
        mult_x_18_n940) );
  XNR2D1BWP12T U1349 ( .A1(n2870), .A2(b[18]), .ZN(n729) );
  OAI22D1BWP12T U1350 ( .A1(n2489), .A2(n604), .B1(n2487), .B2(n729), .ZN(
        mult_x_18_n897) );
  XNR2XD1BWP12T U1351 ( .A1(n2679), .A2(b[13]), .ZN(n747) );
  OAI22D1BWP12T U1352 ( .A1(n2513), .A2(n605), .B1(n747), .B2(n2511), .ZN(
        mult_x_18_n814) );
  OAI22D1BWP12T U1353 ( .A1(n2510), .A2(n607), .B1(n2508), .B2(n606), .ZN(
        mult_x_18_n925) );
  XNR2D1BWP12T U1354 ( .A1(n2456), .A2(n2852), .ZN(n635) );
  XNR2D1BWP12T U1355 ( .A1(n2456), .A2(n2876), .ZN(n668) );
  OAI22D1BWP12T U1356 ( .A1(n2459), .A2(n635), .B1(n668), .B2(n2457), .ZN(
        mult_x_18_n881) );
  XNR2D1BWP12T U1357 ( .A1(n2503), .A2(n2594), .ZN(n743) );
  OAI22D1BWP12T U1358 ( .A1(n2455), .A2(n743), .B1(n2453), .B2(n608), .ZN(
        mult_x_18_n792) );
  XNR2D1BWP12T U1359 ( .A1(n2466), .A2(b[25]), .ZN(n721) );
  OAI22D1BWP12T U1360 ( .A1(n2469), .A2(n609), .B1(n721), .B2(n2467), .ZN(
        mult_x_18_n946) );
  OAI22D1BWP12T U1361 ( .A1(n2510), .A2(n611), .B1(n2508), .B2(n610), .ZN(
        mult_x_18_n922) );
  OAI22D1BWP12T U1362 ( .A1(n2492), .A2(n613), .B1(n612), .B2(n2490), .ZN(
        mult_x_18_n778) );
  OAI22D1BWP12T U1363 ( .A1(n2450), .A2(n615), .B1(n614), .B2(n2449), .ZN(n618) );
  IND2D1BWP12T U1364 ( .A1(n306), .B1(n2456), .ZN(n616) );
  OAI22D1BWP12T U1365 ( .A1(n2459), .A2(n879), .B1(n2457), .B2(n616), .ZN(n617) );
  HA1D1BWP12T U1366 ( .A(n618), .B(n617), .CO(mult_x_18_n696), .S(
        mult_x_18_n697) );
  XNR2D1BWP12T U1367 ( .A1(n2594), .A2(n2351), .ZN(n677) );
  OAI22D1BWP12T U1368 ( .A1(n2455), .A2(n619), .B1(n2453), .B2(n677), .ZN(
        mult_x_18_n790) );
  OAI22D1BWP12T U1369 ( .A1(n2510), .A2(n621), .B1(n2508), .B2(n620), .ZN(
        mult_x_18_n939) );
  XNR2D0BWP12T U1370 ( .A1(n306), .A2(n2358), .ZN(n623) );
  OAI22D1BWP12T U1371 ( .A1(n2478), .A2(n623), .B1(n2476), .B2(n622), .ZN(
        mult_x_18_n761) );
  OAI22D1BWP12T U1372 ( .A1(n2513), .A2(n625), .B1(n624), .B2(n2511), .ZN(
        mult_x_18_n825) );
  OAI22D1BWP12T U1373 ( .A1(n2489), .A2(n627), .B1(n2487), .B2(n626), .ZN(
        mult_x_18_n894) );
  IND2D1BWP12T U1374 ( .A1(n1270), .B1(n2571), .ZN(n628) );
  OAI22D1BWP12T U1375 ( .A1(n2492), .A2(n1820), .B1(n2490), .B2(n628), .ZN(
        mult_x_18_n736) );
  XNR2XD1BWP12T U1376 ( .A1(n2460), .A2(n2351), .ZN(n755) );
  OAI22D1BWP12T U1377 ( .A1(n2463), .A2(n629), .B1(n2461), .B2(n755), .ZN(
        mult_x_18_n766) );
  OAI22D1BWP12T U1378 ( .A1(n2513), .A2(n631), .B1(n630), .B2(n2511), .ZN(
        mult_x_18_n823) );
  OAI22D1BWP12T U1379 ( .A1(n2459), .A2(n633), .B1(n632), .B2(n2457), .ZN(
        mult_x_18_n878) );
  XNR2D1BWP12T U1380 ( .A1(n2499), .A2(n2516), .ZN(n663) );
  OAI22D1BWP12T U1381 ( .A1(n2520), .A2(n663), .B1(n2518), .B2(n634), .ZN(
        mult_x_18_n997) );
  OAI22D1BWP12T U1382 ( .A1(n2459), .A2(n636), .B1(n635), .B2(n2457), .ZN(
        mult_x_18_n882) );
  XNR2D1BWP12T U1383 ( .A1(n2710), .A2(n3106), .ZN(n637) );
  XNR2D1BWP12T U1384 ( .A1(n2710), .A2(n2904), .ZN(n734) );
  OAI22D1BWP12T U1385 ( .A1(n2474), .A2(n637), .B1(n2472), .B2(n734), .ZN(
        mult_x_18_n835) );
  OAI22D1BWP12T U1386 ( .A1(n2474), .A2(n638), .B1(n2472), .B2(n637), .ZN(
        mult_x_18_n836) );
  OAI22D1BWP12T U1387 ( .A1(n2455), .A2(n640), .B1(n2453), .B2(n639), .ZN(
        mult_x_18_n786) );
  XNR2XD1BWP12T U1388 ( .A1(n2499), .A2(a[13]), .ZN(n684) );
  OAI22D1BWP12T U1389 ( .A1(n2495), .A2(n684), .B1(n2493), .B2(n641), .ZN(
        mult_x_18_n862) );
  OAI22D1BWP12T U1390 ( .A1(n2450), .A2(n643), .B1(n642), .B2(n2449), .ZN(n645) );
  XNR2D1BWP12T U1391 ( .A1(n2456), .A2(n2499), .ZN(n760) );
  XNR2D1BWP12T U1392 ( .A1(n2456), .A2(n2351), .ZN(n763) );
  OAI22D1BWP12T U1393 ( .A1(n2459), .A2(n760), .B1(n763), .B2(n2457), .ZN(n644) );
  XNR2D1BWP12T U1394 ( .A1(a[13]), .A2(n2817), .ZN(n732) );
  OAI22D1BWP12T U1395 ( .A1(n2495), .A2(n646), .B1(n2493), .B2(n732), .ZN(
        mult_x_18_n860) );
  XNR2D1BWP12T U1396 ( .A1(n2870), .A2(n2351), .ZN(n662) );
  OAI22D1BWP12T U1397 ( .A1(n2489), .A2(n647), .B1(n2487), .B2(n662), .ZN(
        mult_x_18_n910) );
  XNR2XD1BWP12T U1398 ( .A1(a[13]), .A2(n2452), .ZN(n669) );
  OAI22D1BWP12T U1399 ( .A1(n2495), .A2(n669), .B1(n2493), .B2(n648), .ZN(
        mult_x_18_n854) );
  XNR2D1BWP12T U1400 ( .A1(n2503), .A2(n2460), .ZN(n657) );
  OAI22D1BWP12T U1401 ( .A1(n2463), .A2(n649), .B1(n2461), .B2(n657), .ZN(
        mult_x_18_n769) );
  XNR2D1BWP12T U1402 ( .A1(n2201), .A2(n650), .ZN(n757) );
  OAI22D1BWP12T U1403 ( .A1(n2478), .A2(n651), .B1(n757), .B2(n2476), .ZN(
        mult_x_18_n759) );
  OAI22D1BWP12T U1404 ( .A1(n2520), .A2(n653), .B1(n2518), .B2(n652), .ZN(
        mult_x_18_n989) );
  XNR2D1BWP12T U1405 ( .A1(n2503), .A2(n2621), .ZN(n709) );
  XNR2D1BWP12T U1406 ( .A1(n2764), .A2(n2621), .ZN(n708) );
  OAI22D1BWP12T U1407 ( .A1(n2484), .A2(n709), .B1(n2482), .B2(n708), .ZN(
        mult_x_18_n807) );
  XNR2XD0BWP12T U1408 ( .A1(a[13]), .A2(b[15]), .ZN(n696) );
  OAI22D1BWP12T U1409 ( .A1(n2495), .A2(n654), .B1(n2493), .B2(n696), .ZN(
        mult_x_18_n852) );
  XNR2XD1BWP12T U1410 ( .A1(n2621), .A2(n2876), .ZN(n697) );
  XNR2XD1BWP12T U1411 ( .A1(n2621), .A2(n3106), .ZN(n680) );
  OAI22D1BWP12T U1412 ( .A1(n2484), .A2(n697), .B1(n2482), .B2(n680), .ZN(
        mult_x_18_n800) );
  XNR2D1BWP12T U1413 ( .A1(n2870), .A2(n2817), .ZN(n726) );
  XNR2D1BWP12T U1414 ( .A1(n2870), .A2(n2852), .ZN(n661) );
  OAI22D1BWP12T U1415 ( .A1(n2489), .A2(n726), .B1(n2487), .B2(n661), .ZN(
        mult_x_18_n907) );
  XNR2D1BWP12T U1416 ( .A1(n2516), .A2(n2852), .ZN(n704) );
  OAI22D1BWP12T U1417 ( .A1(n2520), .A2(n704), .B1(n2518), .B2(n655), .ZN(
        mult_x_18_n993) );
  OAI22D1BWP12T U1418 ( .A1(n2463), .A2(n657), .B1(n656), .B2(n2461), .ZN(
        mult_x_18_n768) );
  XNR2D1BWP12T U1419 ( .A1(n2870), .A2(n2904), .ZN(n717) );
  XNR2D1BWP12T U1420 ( .A1(n2870), .A2(n2452), .ZN(n683) );
  OAI22D1BWP12T U1421 ( .A1(n2489), .A2(n717), .B1(n2487), .B2(n683), .ZN(
        mult_x_18_n903) );
  XNR2D1BWP12T U1422 ( .A1(n1270), .A2(n2594), .ZN(n658) );
  XNR2D1BWP12T U1423 ( .A1(n429), .A2(n2594), .ZN(n744) );
  OAI22D1BWP12T U1424 ( .A1(n2455), .A2(n658), .B1(n2453), .B2(n744), .ZN(
        mult_x_18_n794) );
  XNR2XD1BWP12T U1425 ( .A1(n2499), .A2(n2710), .ZN(n711) );
  XNR2D1BWP12T U1426 ( .A1(n2710), .A2(n2351), .ZN(n731) );
  OAI22D1BWP12T U1427 ( .A1(n2474), .A2(n711), .B1(n2472), .B2(n731), .ZN(
        mult_x_18_n841) );
  OAI22D1BWP12T U1428 ( .A1(n2520), .A2(n660), .B1(n2518), .B2(n659), .ZN(
        mult_x_18_n985) );
  XNR2D1BWP12T U1429 ( .A1(n2870), .A2(n2876), .ZN(n673) );
  OAI22D1BWP12T U1430 ( .A1(n2489), .A2(n661), .B1(n2487), .B2(n673), .ZN(
        mult_x_18_n906) );
  XNR2D1BWP12T U1431 ( .A1(n2870), .A2(n2792), .ZN(n727) );
  OAI22D1BWP12T U1432 ( .A1(n2489), .A2(n662), .B1(n2487), .B2(n727), .ZN(
        mult_x_18_n909) );
  OAI22D1BWP12T U1433 ( .A1(n2520), .A2(n664), .B1(n2518), .B2(n663), .ZN(
        mult_x_18_n998) );
  OAI22D1BWP12T U1434 ( .A1(n2489), .A2(n666), .B1(n2487), .B2(n665), .ZN(
        mult_x_18_n900) );
  OAI22D1BWP12T U1435 ( .A1(n2459), .A2(n668), .B1(n667), .B2(n2457), .ZN(
        mult_x_18_n880) );
  OAI22D1BWP12T U1436 ( .A1(n2495), .A2(n670), .B1(n2493), .B2(n669), .ZN(
        mult_x_18_n855) );
  XNR2D1BWP12T U1437 ( .A1(n2764), .A2(a[13]), .ZN(n685) );
  OAI22D1BWP12T U1438 ( .A1(n2495), .A2(n766), .B1(n2493), .B2(n685), .ZN(
        mult_x_18_n864) );
  OAI22D1BWP12T U1439 ( .A1(n2469), .A2(n672), .B1(n671), .B2(n2467), .ZN(
        mult_x_18_n963) );
  XNR2XD1BWP12T U1440 ( .A1(n2710), .A2(n2452), .ZN(n733) );
  XNR2XD1BWP12T U1441 ( .A1(n2710), .A2(b[13]), .ZN(n694) );
  OAI22D1BWP12T U1442 ( .A1(n2474), .A2(n733), .B1(n2472), .B2(n694), .ZN(
        mult_x_18_n833) );
  XNR2D1BWP12T U1443 ( .A1(n2870), .A2(n3106), .ZN(n718) );
  OAI22D1BWP12T U1444 ( .A1(n2489), .A2(n673), .B1(n2487), .B2(n718), .ZN(
        mult_x_18_n905) );
  OAI22D1BWP12T U1445 ( .A1(n2510), .A2(n675), .B1(n2508), .B2(n674), .ZN(
        mult_x_18_n934) );
  OAI22D1BWP12T U1446 ( .A1(n2455), .A2(n677), .B1(n2453), .B2(n676), .ZN(
        mult_x_18_n789) );
  XNR2D1BWP12T U1447 ( .A1(n2503), .A2(n2710), .ZN(n699) );
  XNR2XD1BWP12T U1448 ( .A1(n2764), .A2(n2710), .ZN(n712) );
  OAI22D1BWP12T U1449 ( .A1(n2474), .A2(n699), .B1(n2472), .B2(n712), .ZN(
        mult_x_18_n843) );
  XNR2XD1BWP12T U1450 ( .A1(n306), .A2(n2710), .ZN(n678) );
  XNR2XD1BWP12T U1451 ( .A1(n429), .A2(n2710), .ZN(n700) );
  OAI22D1BWP12T U1452 ( .A1(n2474), .A2(n678), .B1(n2472), .B2(n700), .ZN(
        mult_x_18_n845) );
  OAI22D1BWP12T U1453 ( .A1(n2484), .A2(n680), .B1(n2482), .B2(n679), .ZN(
        mult_x_18_n799) );
  XNR2XD1BWP12T U1454 ( .A1(n306), .A2(n2621), .ZN(n681) );
  OAI22D1BWP12T U1455 ( .A1(n2484), .A2(n681), .B1(n2482), .B2(n710), .ZN(
        mult_x_18_n809) );
  OAI22D1BWP12T U1456 ( .A1(n2489), .A2(n683), .B1(n2487), .B2(n682), .ZN(
        mult_x_18_n902) );
  OAI22D1BWP12T U1457 ( .A1(n2495), .A2(n685), .B1(n2493), .B2(n684), .ZN(
        mult_x_18_n863) );
  OAI22D1BWP12T U1458 ( .A1(n2489), .A2(n687), .B1(n2487), .B2(n686), .ZN(
        mult_x_18_n912) );
  XNR2D1BWP12T U1459 ( .A1(n2516), .A2(b[20]), .ZN(n707) );
  OAI22D1BWP12T U1460 ( .A1(n2520), .A2(n688), .B1(n2518), .B2(n707), .ZN(
        mult_x_18_n982) );
  XNR2XD1BWP12T U1461 ( .A1(n2621), .A2(n2852), .ZN(n698) );
  OAI22D1BWP12T U1462 ( .A1(n2484), .A2(n689), .B1(n2482), .B2(n698), .ZN(
        mult_x_18_n802) );
  CKND0BWP12T U1463 ( .I(n2710), .ZN(n691) );
  IND2D0BWP12T U1464 ( .A1(n1277), .B1(n2710), .ZN(n690) );
  OAI22D1BWP12T U1465 ( .A1(n2474), .A2(n691), .B1(n2472), .B2(n690), .ZN(
        mult_x_18_n740) );
  OAI22D1BWP12T U1466 ( .A1(n2459), .A2(n693), .B1(n692), .B2(n2457), .ZN(
        mult_x_18_n872) );
  XNR2D0BWP12T U1467 ( .A1(n2710), .A2(b[14]), .ZN(n715) );
  OAI22D1BWP12T U1468 ( .A1(n2474), .A2(n694), .B1(n2472), .B2(n715), .ZN(
        mult_x_18_n832) );
  IND2D0BWP12T U1469 ( .A1(n1270), .B1(n2621), .ZN(n695) );
  OAI22D1BWP12T U1470 ( .A1(n2484), .A2(n2623), .B1(n2482), .B2(n695), .ZN(
        mult_x_18_n738) );
  XNR2XD0BWP12T U1471 ( .A1(a[13]), .A2(b[16]), .ZN(n716) );
  OAI22D1BWP12T U1472 ( .A1(n2495), .A2(n696), .B1(n2493), .B2(n716), .ZN(
        mult_x_18_n851) );
  OAI22D1BWP12T U1473 ( .A1(n2484), .A2(n698), .B1(n2482), .B2(n697), .ZN(
        mult_x_18_n801) );
  OAI22D1BWP12T U1474 ( .A1(n2474), .A2(n700), .B1(n2472), .B2(n699), .ZN(
        mult_x_18_n844) );
  XNR2XD1BWP12T U1475 ( .A1(n1270), .A2(n2979), .ZN(n701) );
  XNR2XD1BWP12T U1476 ( .A1(n2979), .A2(b[1]), .ZN(n2505) );
  OAI22D1BWP12T U1477 ( .A1(n2506), .A2(n701), .B1(n2505), .B2(n2504), .ZN(
        mult_x_18_n749) );
  OAI22D1BWP12T U1478 ( .A1(n2469), .A2(n703), .B1(n702), .B2(n2467), .ZN(
        mult_x_18_n955) );
  OAI22D1BWP12T U1479 ( .A1(n2520), .A2(n705), .B1(n2518), .B2(n704), .ZN(
        mult_x_18_n994) );
  OAI22D1BWP12T U1480 ( .A1(n2520), .A2(n707), .B1(n2518), .B2(n706), .ZN(
        mult_x_18_n981) );
  XNR2XD1BWP12T U1481 ( .A1(n2499), .A2(n2621), .ZN(n739) );
  OAI22D1BWP12T U1482 ( .A1(n2484), .A2(n708), .B1(n2482), .B2(n739), .ZN(
        mult_x_18_n806) );
  OAI22D1BWP12T U1483 ( .A1(n2484), .A2(n710), .B1(n2482), .B2(n709), .ZN(
        mult_x_18_n808) );
  OAI22D1BWP12T U1484 ( .A1(n2474), .A2(n712), .B1(n2472), .B2(n711), .ZN(
        mult_x_18_n842) );
  XNR2D1BWP12T U1485 ( .A1(n2503), .A2(n2498), .ZN(n735) );
  OAI22D1BWP12T U1486 ( .A1(n2502), .A2(n713), .B1(n735), .B2(n2500), .ZN(
        mult_x_18_n753) );
  XNR2XD1BWP12T U1487 ( .A1(n2710), .A2(n2792), .ZN(n730) );
  XNR2D1BWP12T U1488 ( .A1(n2710), .A2(n2817), .ZN(n737) );
  OAI22D1BWP12T U1489 ( .A1(n2474), .A2(n730), .B1(n2472), .B2(n737), .ZN(
        mult_x_18_n839) );
  OAI22D1BWP12T U1490 ( .A1(n2474), .A2(n715), .B1(n2472), .B2(n714), .ZN(
        mult_x_18_n831) );
  XNR2XD1BWP12T U1491 ( .A1(a[13]), .A2(b[17]), .ZN(n723) );
  OAI22D1BWP12T U1492 ( .A1(n2495), .A2(n716), .B1(n2493), .B2(n723), .ZN(
        mult_x_18_n850) );
  OAI22D1BWP12T U1493 ( .A1(n2489), .A2(n718), .B1(n2487), .B2(n717), .ZN(
        mult_x_18_n904) );
  OAI22D1BWP12T U1494 ( .A1(n2450), .A2(n720), .B1(n719), .B2(n2449), .ZN(
        mult_x_18_n1005) );
  XNR2D1BWP12T U1495 ( .A1(n2466), .A2(b[26]), .ZN(n746) );
  OAI22D1BWP12T U1496 ( .A1(n2469), .A2(n721), .B1(n746), .B2(n2467), .ZN(
        mult_x_18_n945) );
  OAI22D1BWP12T U1497 ( .A1(n2495), .A2(n723), .B1(n2493), .B2(n722), .ZN(
        mult_x_18_n849) );
  XNR2D1BWP12T U1498 ( .A1(n2466), .A2(n3106), .ZN(n769) );
  OAI22D1BWP12T U1499 ( .A1(n2469), .A2(n724), .B1(n769), .B2(n2467), .ZN(
        mult_x_18_n961) );
  XNR2D1BWP12T U1500 ( .A1(n2516), .A2(b[28]), .ZN(n749) );
  OAI22D1BWP12T U1501 ( .A1(n2520), .A2(n725), .B1(n2518), .B2(n749), .ZN(
        mult_x_18_n974) );
  OAI22D1BWP12T U1502 ( .A1(n2489), .A2(n727), .B1(n2487), .B2(n726), .ZN(
        mult_x_18_n908) );
  OAI22D1BWP12T U1503 ( .A1(n2489), .A2(n729), .B1(n2487), .B2(n728), .ZN(
        mult_x_18_n896) );
  OAI22D1BWP12T U1504 ( .A1(n2474), .A2(n731), .B1(n2472), .B2(n730), .ZN(
        mult_x_18_n840) );
  XNR2XD1BWP12T U1505 ( .A1(a[13]), .A2(n2852), .ZN(n741) );
  OAI22D1BWP12T U1506 ( .A1(n2495), .A2(n732), .B1(n2493), .B2(n741), .ZN(
        mult_x_18_n859) );
  OAI22D1BWP12T U1507 ( .A1(n2474), .A2(n734), .B1(n2472), .B2(n733), .ZN(
        mult_x_18_n834) );
  XNR2XD1BWP12T U1508 ( .A1(n2764), .A2(n2498), .ZN(n2501) );
  OAI22D1BWP12T U1509 ( .A1(n2502), .A2(n735), .B1(n2501), .B2(n2500), .ZN(
        mult_x_18_n752) );
  OAI22D1BWP12T U1510 ( .A1(n2474), .A2(n737), .B1(n2472), .B2(n736), .ZN(
        mult_x_18_n838) );
  OAI22D1BWP12T U1511 ( .A1(n2484), .A2(n739), .B1(n2482), .B2(n738), .ZN(
        mult_x_18_n805) );
  OAI22D1BWP12T U1512 ( .A1(n2495), .A2(n741), .B1(n2493), .B2(n740), .ZN(
        mult_x_18_n858) );
  XNR2D1BWP12T U1513 ( .A1(n2571), .A2(n2852), .ZN(n752) );
  OAI22D1BWP12T U1514 ( .A1(n2492), .A2(n742), .B1(n752), .B2(n2490), .ZN(
        mult_x_18_n774) );
  OAI22D1BWP12T U1515 ( .A1(n2455), .A2(n744), .B1(n2453), .B2(n743), .ZN(
        mult_x_18_n793) );
  XNR2D1BWP12T U1516 ( .A1(n2456), .A2(b[20]), .ZN(n754) );
  OAI22D1BWP12T U1517 ( .A1(n2459), .A2(n745), .B1(n754), .B2(n2457), .ZN(
        mult_x_18_n870) );
  OAI22D1BWP12T U1518 ( .A1(n2469), .A2(n746), .B1(n2468), .B2(n2467), .ZN(
        mult_x_18_n944) );
  XNR2XD0BWP12T U1519 ( .A1(n2679), .A2(b[14]), .ZN(n751) );
  OAI22D1BWP12T U1520 ( .A1(n2513), .A2(n747), .B1(n751), .B2(n2511), .ZN(
        mult_x_18_n813) );
  XNR2D1BWP12T U1521 ( .A1(n2870), .A2(b[23]), .ZN(n2488) );
  OAI22D1BWP12T U1522 ( .A1(n2489), .A2(n748), .B1(n2487), .B2(n2488), .ZN(
        mult_x_18_n892) );
  XNR2D1BWP12T U1523 ( .A1(n2516), .A2(b[29]), .ZN(n2519) );
  OAI22D1BWP12T U1524 ( .A1(n2520), .A2(n749), .B1(n2518), .B2(n2519), .ZN(
        mult_x_18_n973) );
  XNR2D1BWP12T U1525 ( .A1(n2594), .A2(n2904), .ZN(n2454) );
  OAI22D1BWP12T U1526 ( .A1(n2455), .A2(n750), .B1(n2453), .B2(n2454), .ZN(
        mult_x_18_n784) );
  XNR2XD0BWP12T U1527 ( .A1(n2679), .A2(b[15]), .ZN(n2512) );
  OAI22D1BWP12T U1528 ( .A1(n2513), .A2(n751), .B1(n2512), .B2(n2511), .ZN(
        mult_x_18_n812) );
  XNR2D1BWP12T U1529 ( .A1(n2571), .A2(n2876), .ZN(n2491) );
  OAI22D1BWP12T U1530 ( .A1(n2492), .A2(n752), .B1(n2491), .B2(n2490), .ZN(
        mult_x_18_n773) );
  XNR2XD1BWP12T U1531 ( .A1(n2710), .A2(b[17]), .ZN(n2473) );
  OAI22D1BWP12T U1532 ( .A1(n2474), .A2(n753), .B1(n2472), .B2(n2473), .ZN(
        mult_x_18_n829) );
  XNR2D1BWP12T U1533 ( .A1(n2456), .A2(b[21]), .ZN(n2458) );
  OAI22D1BWP12T U1534 ( .A1(n2459), .A2(n754), .B1(n2458), .B2(n2457), .ZN(
        mult_x_18_n869) );
  XNR2XD1BWP12T U1535 ( .A1(n2460), .A2(n2792), .ZN(n758) );
  OAI22D1BWP12T U1536 ( .A1(n2463), .A2(n755), .B1(n2461), .B2(n758), .ZN(
        mult_x_18_n765) );
  OAI22D1BWP12T U1537 ( .A1(n2478), .A2(n757), .B1(n756), .B2(n2476), .ZN(
        mult_x_18_n758) );
  XNR2D1BWP12T U1538 ( .A1(n2460), .A2(n2817), .ZN(n2462) );
  OAI22D1BWP12T U1539 ( .A1(n2463), .A2(n758), .B1(n2461), .B2(n2462), .ZN(
        mult_x_18_n764) );
  XNR2D1BWP12T U1540 ( .A1(n2815), .A2(b[25]), .ZN(n2509) );
  OAI22D0BWP12T U1541 ( .A1(n2510), .A2(n759), .B1(n2508), .B2(n2509), .ZN(
        mult_x_18_n917) );
  TPOAI22D2BWP12T U1542 ( .A1(n2459), .A2(n763), .B1(n762), .B2(n2457), .ZN(
        mult_x_18_n884) );
  TPOAI22D2BWP12T U1543 ( .A1(n2459), .A2(n765), .B1(n764), .B2(n2457), .ZN(
        mult_x_18_n888) );
  TPOAI22D1BWP12T U1544 ( .A1(n2495), .A2(n767), .B1(n2493), .B2(n766), .ZN(
        mult_x_18_n865) );
  TPOAI22D1BWP12T U1545 ( .A1(n2469), .A2(n769), .B1(n768), .B2(n2467), .ZN(
        mult_x_18_n960) );
  IND2D0BWP12T U1546 ( .A1(n1277), .B1(n2460), .ZN(n770) );
  TPOAI22D1BWP12T U1547 ( .A1(n2463), .A2(n2202), .B1(n2461), .B2(n770), .ZN(
        mult_x_18_n735) );
  ND2D1BWP12T U1548 ( .A1(n287), .A2(n1539), .ZN(n801) );
  NR2D1BWP12T U1549 ( .A1(mult_x_18_n642), .A2(mult_x_18_n630), .ZN(n771) );
  INVD1BWP12T U1550 ( .I(n771), .ZN(n1534) );
  NR2D1BWP12T U1551 ( .A1(mult_x_18_n643), .A2(mult_x_18_n653), .ZN(n1531) );
  INVD1BWP12T U1552 ( .I(n1531), .ZN(n1484) );
  ND2D1BWP12T U1553 ( .A1(n1534), .A2(n1484), .ZN(n1478) );
  NR2D1BWP12T U1554 ( .A1(mult_x_18_n618), .A2(mult_x_18_n629), .ZN(n1479) );
  NR2D1BWP12T U1555 ( .A1(n1478), .A2(n1479), .ZN(n794) );
  CKND2D1BWP12T U1556 ( .A1(n293), .A2(n1525), .ZN(n790) );
  OR2D2BWP12T U1557 ( .A1(mult_x_18_n684), .A2(mult_x_18_n691), .Z(n1283) );
  ND2D1BWP12T U1558 ( .A1(n1283), .A2(n1491), .ZN(n786) );
  OR2XD1BWP12T U1559 ( .A1(mult_x_18_n717), .A2(mult_x_18_n713), .Z(n1520) );
  CKND2D1BWP12T U1560 ( .A1(n288), .A2(n1520), .ZN(n782) );
  FA1D0BWP12T U1561 ( .A(n774), .B(n773), .CI(n772), .CO(n778), .S(n312) );
  NR2D1BWP12T U1562 ( .A1(mult_x_18_n723), .A2(n778), .ZN(n1503) );
  OA21D1BWP12T U1563 ( .A1(n777), .A2(n776), .B(n775), .Z(n1506) );
  ND2D1BWP12T U1564 ( .A1(mult_x_18_n723), .A2(n778), .ZN(n1504) );
  OAI21D1BWP12T U1565 ( .A1(n1503), .A2(n1506), .B(n1504), .ZN(n1501) );
  OR2XD1BWP12T U1566 ( .A1(mult_x_18_n718), .A2(mult_x_18_n722), .Z(n1500) );
  ND2D1BWP12T U1567 ( .A1(mult_x_18_n718), .A2(mult_x_18_n722), .ZN(n1499) );
  INVD1BWP12T U1568 ( .I(n1499), .ZN(n779) );
  AOI21D1BWP12T U1569 ( .A1(n1501), .A2(n1500), .B(n779), .ZN(n1497) );
  ND2D1BWP12T U1570 ( .A1(mult_x_18_n717), .A2(mult_x_18_n713), .ZN(n1519) );
  INVD1BWP12T U1571 ( .I(n1519), .ZN(n1498) );
  ND2D1BWP12T U1572 ( .A1(mult_x_18_n706), .A2(mult_x_18_n712), .ZN(n1496) );
  INVD1BWP12T U1573 ( .I(n1496), .ZN(n780) );
  AOI21D1BWP12T U1574 ( .A1(n288), .A2(n1498), .B(n780), .ZN(n781) );
  OR2XD1BWP12T U1575 ( .A1(mult_x_18_n700), .A2(mult_x_18_n705), .Z(n1494) );
  ND2D1BWP12T U1576 ( .A1(mult_x_18_n700), .A2(mult_x_18_n705), .ZN(n1493) );
  INVD1BWP12T U1577 ( .I(n1493), .ZN(n783) );
  ND2D1BWP12T U1578 ( .A1(mult_x_18_n692), .A2(mult_x_18_n699), .ZN(n1490) );
  INVD1BWP12T U1579 ( .I(n1490), .ZN(n1281) );
  ND2D1BWP12T U1580 ( .A1(mult_x_18_n684), .A2(mult_x_18_n691), .ZN(n1282) );
  TPAOI21D2BWP12T U1581 ( .A1(n1283), .A2(n1281), .B(n784), .ZN(n785) );
  ND2D1BWP12T U1582 ( .A1(mult_x_18_n674), .A2(mult_x_18_n683), .ZN(n1486) );
  INVD1BWP12T U1583 ( .I(n1486), .ZN(n787) );
  TPAOI21D1BWP12T U1584 ( .A1(n1488), .A2(n1487), .B(n787), .ZN(n1324) );
  INVD1BWP12T U1585 ( .I(n1325), .ZN(n1524) );
  INVD1BWP12T U1586 ( .I(n1527), .ZN(n788) );
  AOI21D1BWP12T U1587 ( .A1(n293), .A2(n1524), .B(n788), .ZN(n789) );
  ND2D1BWP12T U1588 ( .A1(mult_x_18_n643), .A2(mult_x_18_n653), .ZN(n1530) );
  INVD1BWP12T U1589 ( .I(n1530), .ZN(n792) );
  ND2D1BWP12T U1590 ( .A1(mult_x_18_n642), .A2(mult_x_18_n630), .ZN(n1533) );
  INVD1BWP12T U1591 ( .I(n1533), .ZN(n791) );
  AOI21D1BWP12T U1592 ( .A1(n1534), .A2(n792), .B(n791), .ZN(n1477) );
  ND2D1BWP12T U1593 ( .A1(mult_x_18_n618), .A2(mult_x_18_n629), .ZN(n1480) );
  OAI21D1BWP12T U1594 ( .A1(n1477), .A2(n1479), .B(n1480), .ZN(n793) );
  TPAOI21D1BWP12T U1595 ( .A1(n794), .A2(n1476), .B(n793), .ZN(n1459) );
  OR2XD1BWP12T U1596 ( .A1(mult_x_18_n604), .A2(mult_x_18_n617), .Z(n1471) );
  CKND2D1BWP12T U1597 ( .A1(n289), .A2(n1471), .ZN(n797) );
  ND2D1BWP12T U1598 ( .A1(mult_x_18_n604), .A2(mult_x_18_n617), .ZN(n1460) );
  INVD1BWP12T U1599 ( .I(n1460), .ZN(n1470) );
  ND2D1BWP12T U1600 ( .A1(mult_x_18_n590), .A2(mult_x_18_n603), .ZN(n1473) );
  INVD1BWP12T U1601 ( .I(n1473), .ZN(n795) );
  AOI21D1BWP12T U1602 ( .A1(n289), .A2(n1470), .B(n795), .ZN(n796) );
  OR2XD1BWP12T U1603 ( .A1(mult_x_18_n574), .A2(mult_x_18_n589), .Z(n1463) );
  ND2D1BWP12T U1604 ( .A1(mult_x_18_n574), .A2(mult_x_18_n589), .ZN(n1462) );
  INVD1BWP12T U1605 ( .I(n1462), .ZN(n798) );
  TPAOI21D1BWP12T U1606 ( .A1(n1464), .A2(n1463), .B(n798), .ZN(n1465) );
  ND2D1BWP12T U1607 ( .A1(mult_x_18_n559), .A2(mult_x_18_n573), .ZN(n1538) );
  INVD1BWP12T U1608 ( .I(n1538), .ZN(n1466) );
  ND2D1BWP12T U1609 ( .A1(mult_x_18_n558), .A2(mult_x_18_n542), .ZN(n1467) );
  INVD1BWP12T U1610 ( .I(n1467), .ZN(n799) );
  TPAOI21D1BWP12T U1611 ( .A1(n287), .A2(n1466), .B(n799), .ZN(n800) );
  TPOAI21D1BWP12T U1612 ( .A1(n801), .A2(n1465), .B(n800), .ZN(n1134) );
  TPNR2D1BWP12T U1613 ( .A1(mult_x_18_n506), .A2(mult_x_18_n524), .ZN(n1135)
         );
  TPNR2D1BWP12T U1614 ( .A1(mult_x_18_n525), .A2(mult_x_18_n541), .ZN(n1542)
         );
  NR2D1BWP12T U1615 ( .A1(n1135), .A2(n1542), .ZN(n803) );
  ND2D1BWP12T U1616 ( .A1(mult_x_18_n525), .A2(mult_x_18_n541), .ZN(n1543) );
  ND2D1BWP12T U1617 ( .A1(mult_x_18_n506), .A2(mult_x_18_n524), .ZN(n1136) );
  TPOAI21D1BWP12T U1618 ( .A1(n1135), .A2(n1543), .B(n1136), .ZN(n802) );
  TPAOI21D1BWP12T U1619 ( .A1(n1134), .A2(n803), .B(n802), .ZN(n932) );
  NR2D1BWP12T U1620 ( .A1(mult_x_18_n447), .A2(mult_x_18_n426), .ZN(n1558) );
  NR2D1BWP12T U1621 ( .A1(mult_x_18_n467), .A2(mult_x_18_n448), .ZN(n1553) );
  NR2D1BWP12T U1622 ( .A1(n1558), .A2(n1553), .ZN(n805) );
  TPNR2D2BWP12T U1623 ( .A1(mult_x_18_n487), .A2(mult_x_18_n468), .ZN(n987) );
  ND2D1BWP12T U1624 ( .A1(n805), .A2(n1549), .ZN(n807) );
  ND2D1BWP12T U1625 ( .A1(mult_x_18_n505), .A2(mult_x_18_n488), .ZN(n1039) );
  ND2D1BWP12T U1626 ( .A1(mult_x_18_n487), .A2(mult_x_18_n468), .ZN(n988) );
  OAI21D1BWP12T U1627 ( .A1(n987), .A2(n1039), .B(n988), .ZN(n1551) );
  ND2D1BWP12T U1628 ( .A1(mult_x_18_n467), .A2(mult_x_18_n448), .ZN(n1552) );
  ND2D1BWP12T U1629 ( .A1(mult_x_18_n447), .A2(mult_x_18_n426), .ZN(n1559) );
  AOI21D1BWP12T U1630 ( .A1(n805), .A2(n1551), .B(n804), .ZN(n806) );
  OAI21D1BWP12T U1631 ( .A1(n932), .A2(n807), .B(n806), .ZN(n1548) );
  CKND0BWP12T U1632 ( .I(b[28]), .ZN(n937) );
  INVD1BWP12T U1633 ( .I(b[22]), .ZN(n1720) );
  NR2D1BWP12T U1634 ( .A1(n808), .A2(n810), .ZN(n1691) );
  INVD1P75BWP12T U1635 ( .I(n2792), .ZN(n841) );
  NR2D1BWP12T U1636 ( .A1(n841), .A2(n2785), .ZN(n1694) );
  NR2D1BWP12T U1637 ( .A1(n1695), .A2(n1694), .ZN(n813) );
  CKND2D1BWP12T U1638 ( .A1(n1691), .A2(n813), .ZN(n815) );
  OAI21D1BWP12T U1639 ( .A1(n1700), .A2(n810), .B(n809), .ZN(n1692) );
  CKND2D1BWP12T U1640 ( .A1(n841), .A2(n2785), .ZN(n1693) );
  ND2D1BWP12T U1641 ( .A1(n2170), .A2(n811), .ZN(n1696) );
  OAI21D1BWP12T U1642 ( .A1(n1695), .A2(n1693), .B(n1696), .ZN(n812) );
  TPAOI21D0BWP12T U1643 ( .A1(n1692), .A2(n813), .B(n812), .ZN(n814) );
  OAI21D1BWP12T U1644 ( .A1(n816), .A2(n815), .B(n814), .ZN(n1682) );
  INVD1P75BWP12T U1645 ( .I(n1682), .ZN(n1711) );
  INVD1P75BWP12T U1646 ( .I(n2904), .ZN(n2163) );
  OR2D2BWP12T U1647 ( .A1(n2163), .A2(n2898), .Z(n1713) );
  INVD1P75BWP12T U1648 ( .I(n2452), .ZN(n2159) );
  ND2D1BWP12T U1649 ( .A1(n1713), .A2(n286), .ZN(n821) );
  INVD1BWP12T U1650 ( .I(n3106), .ZN(n818) );
  NR2D1BWP12T U1651 ( .A1(n818), .A2(n3100), .ZN(n1707) );
  NR2D1BWP12T U1652 ( .A1(n821), .A2(n1707), .ZN(n823) );
  INVD1BWP12T U1653 ( .I(n2876), .ZN(n817) );
  NR2D1BWP12T U1654 ( .A1(n817), .A2(n2870), .ZN(n1683) );
  NR2D1BWP12T U1655 ( .A1(n2162), .A2(n2846), .ZN(n1679) );
  NR2D1BWP12T U1656 ( .A1(n1683), .A2(n1679), .ZN(n1293) );
  ND2D1BWP12T U1657 ( .A1(n823), .A2(n1293), .ZN(n1671) );
  INVD1P75BWP12T U1658 ( .I(b[13]), .ZN(n2160) );
  NR2D1BWP12T U1659 ( .A1(n2160), .A2(a[13]), .ZN(n1672) );
  OR2D0BWP12T U1660 ( .A1(n1671), .A2(n1672), .Z(n825) );
  CKND2D1BWP12T U1661 ( .A1(n2162), .A2(n2846), .ZN(n1680) );
  ND2D1BWP12T U1662 ( .A1(n817), .A2(n2870), .ZN(n1684) );
  OAI21D1BWP12T U1663 ( .A1(n1683), .A2(n1680), .B(n1684), .ZN(n1294) );
  ND2D1BWP12T U1664 ( .A1(n818), .A2(n3100), .ZN(n1708) );
  ND2D1BWP12T U1665 ( .A1(n2163), .A2(n2898), .ZN(n1712) );
  INVD1BWP12T U1666 ( .I(n1712), .ZN(n1295) );
  ND2D1BWP12T U1667 ( .A1(n2159), .A2(a[12]), .ZN(n1296) );
  INVD1BWP12T U1668 ( .I(n1296), .ZN(n819) );
  AOI21D1BWP12T U1669 ( .A1(n286), .A2(n1295), .B(n819), .ZN(n820) );
  OAI21D1BWP12T U1670 ( .A1(n821), .A2(n1708), .B(n820), .ZN(n822) );
  AOI21D1BWP12T U1671 ( .A1(n823), .A2(n1294), .B(n822), .ZN(n1670) );
  ND2D1BWP12T U1672 ( .A1(n2160), .A2(a[13]), .ZN(n1673) );
  OA21D1BWP12T U1673 ( .A1(n1670), .A2(n1672), .B(n1673), .Z(n824) );
  TPOAI21D1BWP12T U1674 ( .A1(n1711), .A2(n825), .B(n824), .ZN(n1328) );
  OR2XD1BWP12T U1675 ( .A1(n2157), .A2(a[14]), .Z(n1327) );
  TPAOI21D1BWP12T U1676 ( .A1(n1328), .A2(n1327), .B(n856), .ZN(n1678) );
  INVD1P75BWP12T U1677 ( .I(b[15]), .ZN(n2158) );
  NR2D1BWP12T U1678 ( .A1(n2158), .A2(n2710), .ZN(n1676) );
  ND2D1BWP12T U1679 ( .A1(n2158), .A2(n2710), .ZN(n1677) );
  OR2XD1BWP12T U1680 ( .A1(n2151), .A2(n2915), .Z(n1667) );
  ND2D1BWP12T U1681 ( .A1(n2151), .A2(n2915), .ZN(n1666) );
  INVD1BWP12T U1682 ( .I(n1666), .ZN(n826) );
  NR2D1BWP12T U1683 ( .A1(n2156), .A2(n2679), .ZN(n1661) );
  ND2D1BWP12T U1684 ( .A1(n2156), .A2(n2679), .ZN(n1662) );
  OR2XD1BWP12T U1685 ( .A1(n2149), .A2(n2652), .Z(n1658) );
  ND2D1BWP12T U1686 ( .A1(n2149), .A2(n2652), .ZN(n1657) );
  INVD1BWP12T U1687 ( .I(n1657), .ZN(n827) );
  TPAOI21D1BWP12T U1688 ( .A1(n1660), .A2(n1658), .B(n827), .ZN(n1718) );
  NR2D1BWP12T U1689 ( .A1(n2150), .A2(n2621), .ZN(n1715) );
  ND2D1BWP12T U1690 ( .A1(n2150), .A2(n2621), .ZN(n1716) );
  TPOAI21D1BWP12T U1691 ( .A1(n1718), .A2(n1715), .B(n1716), .ZN(n1656) );
  OR2XD1BWP12T U1692 ( .A1(n2148), .A2(a[20]), .Z(n1654) );
  ND2D1BWP12T U1693 ( .A1(n2148), .A2(a[20]), .ZN(n1653) );
  INVD1BWP12T U1694 ( .I(n1653), .ZN(n828) );
  TPAOI21D1BWP12T U1695 ( .A1(n1656), .A2(n1654), .B(n828), .ZN(n1652) );
  NR2D1BWP12T U1696 ( .A1(n1450), .A2(n2594), .ZN(n1650) );
  ND2D1BWP12T U1697 ( .A1(n1450), .A2(n2594), .ZN(n1651) );
  OAI21D1BWP12T U1698 ( .A1(n1652), .A2(n1650), .B(n1651), .ZN(n1719) );
  NR2D1BWP12T U1699 ( .A1(n2792), .A2(n2785), .ZN(n1759) );
  NR2D1BWP12T U1700 ( .A1(n1620), .A2(n1759), .ZN(n830) );
  ND2D1BWP12T U1701 ( .A1(n1616), .A2(n830), .ZN(n832) );
  ND2D1BWP12T U1702 ( .A1(n2792), .A2(n2785), .ZN(n1758) );
  OAI21D1BWP12T U1703 ( .A1(n1759), .A2(n1619), .B(n1758), .ZN(n829) );
  AOI21D1BWP12T U1704 ( .A1(n1618), .A2(n830), .B(n829), .ZN(n831) );
  INVD2BWP12T U1705 ( .I(n1630), .ZN(n1607) );
  NR2D1BWP12T U1706 ( .A1(n811), .A2(n2817), .ZN(n1606) );
  NR2D1BWP12T U1707 ( .A1(n2852), .A2(n2846), .ZN(n1631) );
  NR2D1BWP12T U1708 ( .A1(n1606), .A2(n1631), .ZN(n1581) );
  NR2D1BWP12T U1709 ( .A1(n2870), .A2(n2876), .ZN(n1580) );
  NR2D1BWP12T U1710 ( .A1(n3106), .A2(n3100), .ZN(n1585) );
  NR2D1BWP12T U1711 ( .A1(n1580), .A2(n1585), .ZN(n835) );
  ND2D1BWP12T U1712 ( .A1(n1581), .A2(n835), .ZN(n1588) );
  NR2D1BWP12T U1713 ( .A1(n2898), .A2(n2904), .ZN(n1297) );
  NR2D1BWP12T U1714 ( .A1(n2452), .A2(a[12]), .ZN(n866) );
  NR2D1BWP12T U1715 ( .A1(n1297), .A2(n866), .ZN(n1595) );
  OR2XD1BWP12T U1716 ( .A1(a[13]), .A2(b[13]), .Z(n1600) );
  CKND2D1BWP12T U1717 ( .A1(n1595), .A2(n1600), .ZN(n838) );
  OR2XD1BWP12T U1718 ( .A1(n1588), .A2(n838), .Z(n840) );
  ND2D1BWP12T U1719 ( .A1(n811), .A2(n2817), .ZN(n1627) );
  CKND2D1BWP12T U1720 ( .A1(n2852), .A2(n2846), .ZN(n1632) );
  OAI21D1BWP12T U1721 ( .A1(n1631), .A2(n1627), .B(n1632), .ZN(n1584) );
  ND2D1BWP12T U1722 ( .A1(n2870), .A2(n2876), .ZN(n1582) );
  ND2D1BWP12T U1723 ( .A1(n3106), .A2(n3100), .ZN(n1586) );
  OAI21D1BWP12T U1724 ( .A1(n1585), .A2(n1582), .B(n1586), .ZN(n834) );
  AOI21D1BWP12T U1725 ( .A1(n835), .A2(n1584), .B(n834), .ZN(n1587) );
  ND2D1BWP12T U1726 ( .A1(n2898), .A2(n2904), .ZN(n1780) );
  ND2D1BWP12T U1727 ( .A1(n2452), .A2(a[12]), .ZN(n1310) );
  OAI21D1BWP12T U1728 ( .A1(n866), .A2(n1780), .B(n1310), .ZN(n1594) );
  CKND2D1BWP12T U1729 ( .A1(a[13]), .A2(b[13]), .ZN(n1599) );
  INVD1BWP12T U1730 ( .I(n1599), .ZN(n836) );
  AOI21D1BWP12T U1731 ( .A1(n1594), .A2(n1600), .B(n836), .ZN(n837) );
  OA21D1BWP12T U1732 ( .A1(n1587), .A2(n838), .B(n837), .Z(n839) );
  TPOAI21D1BWP12T U1733 ( .A1(n1607), .A2(n840), .B(n839), .ZN(n1362) );
  OR2XD1BWP12T U1734 ( .A1(b[14]), .A2(a[14]), .Z(n1360) );
  ND2D1BWP12T U1735 ( .A1(b[14]), .A2(a[14]), .ZN(n1359) );
  INVD1BWP12T U1736 ( .I(n1359), .ZN(n873) );
  NR2D1BWP12T U1737 ( .A1(n2710), .A2(b[15]), .ZN(n1603) );
  ND2D1BWP12T U1738 ( .A1(n2710), .A2(b[15]), .ZN(n1782) );
  OR2XD1BWP12T U1739 ( .A1(b[16]), .A2(n2915), .Z(n1743) );
  ND2D1BWP12T U1740 ( .A1(b[16]), .A2(n2915), .ZN(n1742) );
  INVD1BWP12T U1741 ( .I(n1742), .ZN(n874) );
  NR2D1BWP12T U1742 ( .A1(n2679), .A2(b[17]), .ZN(n1590) );
  ND2D1BWP12T U1743 ( .A1(n2679), .A2(b[17]), .ZN(n1738) );
  OR2XD1BWP12T U1744 ( .A1(b[18]), .A2(n2652), .Z(n1735) );
  ND2D1BWP12T U1745 ( .A1(b[18]), .A2(n2652), .ZN(n1734) );
  INVD1BWP12T U1746 ( .I(n1734), .ZN(n875) );
  NR2D1BWP12T U1747 ( .A1(n2621), .A2(b[19]), .ZN(n1575) );
  ND2D1BWP12T U1748 ( .A1(n2621), .A2(b[19]), .ZN(n1730) );
  OR2XD1BWP12T U1749 ( .A1(b[20]), .A2(a[20]), .Z(n1795) );
  ND2D1BWP12T U1750 ( .A1(b[20]), .A2(a[20]), .ZN(n1794) );
  INVD1BWP12T U1751 ( .I(n1794), .ZN(n876) );
  AO21D1BWP12T U1752 ( .A1(n1574), .A2(n1795), .B(n876), .Z(n1639) );
  INVD1BWP12T U1753 ( .I(b[29]), .ZN(n1377) );
  INVD1BWP12T U1754 ( .I(b[27]), .ZN(n993) );
  INVD1BWP12T U1755 ( .I(b[25]), .ZN(n1141) );
  INVD1BWP12T U1756 ( .I(b[24]), .ZN(n1452) );
  INVD1BWP12T U1757 ( .I(b[23]), .ZN(n1379) );
  INVD1BWP12T U1758 ( .I(b[21]), .ZN(n1450) );
  NR2D1BWP12T U1759 ( .A1(n841), .A2(n2785), .ZN(n1422) );
  NR2D1BWP12T U1760 ( .A1(n1421), .A2(n1422), .ZN(n843) );
  CKND2D1BWP12T U1761 ( .A1(n1418), .A2(n843), .ZN(n845) );
  CKND2D1BWP12T U1762 ( .A1(n841), .A2(n2785), .ZN(n1423) );
  OAI21D1BWP12T U1763 ( .A1(n1422), .A2(n1420), .B(n1423), .ZN(n842) );
  AOI21D1BWP12T U1764 ( .A1(n1419), .A2(n843), .B(n842), .ZN(n844) );
  OAI21D1BWP12T U1765 ( .A1(n846), .A2(n845), .B(n844), .ZN(n1415) );
  INVD2BWP12T U1766 ( .I(n1415), .ZN(n1437) );
  NR2D1BWP12T U1767 ( .A1(n2170), .A2(n2815), .ZN(n1411) );
  NR2D1BWP12T U1768 ( .A1(n2162), .A2(n2846), .ZN(n1416) );
  NR2D1BWP12T U1769 ( .A1(n1411), .A2(n1416), .ZN(n1395) );
  INVD1BWP12T U1770 ( .I(n2876), .ZN(n847) );
  NR2D1BWP12T U1771 ( .A1(n847), .A2(n2870), .ZN(n1394) );
  INVD1BWP12T U1772 ( .I(n3106), .ZN(n848) );
  NR2D1BWP12T U1773 ( .A1(n848), .A2(n3100), .ZN(n1399) );
  NR2D1BWP12T U1774 ( .A1(n1394), .A2(n1399), .ZN(n850) );
  ND2D1BWP12T U1775 ( .A1(n1395), .A2(n850), .ZN(n1403) );
  NR2D1BWP12T U1776 ( .A1(n2159), .A2(a[12]), .ZN(n1289) );
  NR2D1BWP12T U1777 ( .A1(n1286), .A2(n1289), .ZN(n1435) );
  CKND2D1BWP12T U1778 ( .A1(n1435), .A2(n1439), .ZN(n853) );
  OR2XD1BWP12T U1779 ( .A1(n1403), .A2(n853), .Z(n855) );
  ND2D1BWP12T U1780 ( .A1(n2170), .A2(n2815), .ZN(n1413) );
  CKND2D1BWP12T U1781 ( .A1(n2162), .A2(n2846), .ZN(n1417) );
  OAI21D1BWP12T U1782 ( .A1(n1416), .A2(n1413), .B(n1417), .ZN(n1398) );
  ND2D1BWP12T U1783 ( .A1(n847), .A2(n2870), .ZN(n1396) );
  ND2D1BWP12T U1784 ( .A1(n848), .A2(n3100), .ZN(n1400) );
  OAI21D1BWP12T U1785 ( .A1(n1399), .A2(n1396), .B(n1400), .ZN(n849) );
  AOI21D1BWP12T U1786 ( .A1(n850), .A2(n1398), .B(n849), .ZN(n1402) );
  ND2D1BWP12T U1787 ( .A1(n2163), .A2(n2898), .ZN(n1404) );
  CKND2D1BWP12T U1788 ( .A1(n2159), .A2(a[12]), .ZN(n1290) );
  OAI21D1BWP12T U1789 ( .A1(n1289), .A2(n1404), .B(n1290), .ZN(n1434) );
  ND2D1BWP12T U1790 ( .A1(n2160), .A2(a[13]), .ZN(n1438) );
  INVD1BWP12T U1791 ( .I(n1438), .ZN(n851) );
  AOI21D1BWP12T U1792 ( .A1(n1434), .A2(n1439), .B(n851), .ZN(n852) );
  OA21D1BWP12T U1793 ( .A1(n1402), .A2(n853), .B(n852), .Z(n854) );
  TPOAI21D2BWP12T U1794 ( .A1(n1437), .A2(n855), .B(n854), .ZN(n1346) );
  ND2D1BWP12T U1795 ( .A1(n2157), .A2(a[14]), .ZN(n1343) );
  INVD1BWP12T U1796 ( .I(n1343), .ZN(n856) );
  NR2D1BWP12T U1797 ( .A1(n2158), .A2(n2710), .ZN(n1406) );
  ND2D1BWP12T U1798 ( .A1(n2158), .A2(n2710), .ZN(n1407) );
  ND2D1BWP12T U1799 ( .A1(n2151), .A2(n2915), .ZN(n1445) );
  NR2D1BWP12T U1800 ( .A1(n2156), .A2(n2679), .ZN(n1441) );
  ND2D1BWP12T U1801 ( .A1(n2156), .A2(n2679), .ZN(n1442) );
  OR2XD1BWP12T U1802 ( .A1(n2149), .A2(n2652), .Z(n1391) );
  ND2D1BWP12T U1803 ( .A1(n2149), .A2(n2652), .ZN(n1390) );
  TPAOI21D1BWP12T U1804 ( .A1(n1393), .A2(n1391), .B(n827), .ZN(n1389) );
  NR2D1BWP12T U1805 ( .A1(n2150), .A2(n2621), .ZN(n1385) );
  ND2D1BWP12T U1806 ( .A1(n2150), .A2(n2621), .ZN(n1386) );
  TPOAI21D1BWP12T U1807 ( .A1(n1389), .A2(n1385), .B(n1386), .ZN(n1384) );
  OR2XD1BWP12T U1808 ( .A1(n2148), .A2(a[20]), .Z(n1382) );
  ND2D1BWP12T U1809 ( .A1(n2148), .A2(a[20]), .ZN(n1381) );
  AO21D1BWP12T U1810 ( .A1(n1384), .A2(n1382), .B(n828), .Z(n1449) );
  TPND2D2BWP12T U1811 ( .A1(n2421), .A2(n3076), .ZN(n929) );
  NR2D1BWP12T U1812 ( .A1(n857), .A2(n859), .ZN(n1756) );
  CKBD1BWP12T U1813 ( .I(n2815), .Z(n860) );
  TPNR2D2BWP12T U1814 ( .A1(n1760), .A2(n1759), .ZN(n862) );
  ND2D1BWP12T U1815 ( .A1(n1756), .A2(n862), .ZN(n864) );
  OAI21D1BWP12T U1816 ( .A1(n1766), .A2(n859), .B(n858), .ZN(n1757) );
  ND2D1BWP12T U1817 ( .A1(n860), .A2(n2817), .ZN(n1761) );
  TPOAI21D1BWP12T U1818 ( .A1(n1760), .A2(n1758), .B(n1761), .ZN(n861) );
  TPAOI21D1BWP12T U1819 ( .A1(n1757), .A2(n862), .B(n861), .ZN(n863) );
  TPOAI21D1BWP12T U1820 ( .A1(n865), .A2(n864), .B(n863), .ZN(n1771) );
  INVD2BWP12T U1821 ( .I(n1771), .ZN(n1790) );
  NR2D1BWP12T U1822 ( .A1(n2852), .A2(n2846), .ZN(n1769) );
  NR2D1BWP12T U1823 ( .A1(n1772), .A2(n1769), .ZN(n1776) );
  NR2D1BWP12T U1824 ( .A1(n3106), .A2(n3100), .ZN(n1775) );
  NR2D1BWP12T U1825 ( .A1(n1297), .A2(n1775), .ZN(n868) );
  ND2D1BWP12T U1826 ( .A1(n1776), .A2(n868), .ZN(n1786) );
  OR2XD1BWP12T U1827 ( .A1(a[13]), .A2(b[13]), .Z(n1791) );
  INVD1BWP12T U1828 ( .I(n866), .ZN(n1789) );
  CKND2D1BWP12T U1829 ( .A1(n1791), .A2(n1789), .ZN(n870) );
  OR2D0BWP12T U1830 ( .A1(n1786), .A2(n870), .Z(n872) );
  CKND2D1BWP12T U1831 ( .A1(n2852), .A2(n2846), .ZN(n1770) );
  ND2D1BWP12T U1832 ( .A1(n2870), .A2(n2876), .ZN(n1773) );
  OAI21D1BWP12T U1833 ( .A1(n1772), .A2(n1770), .B(n1773), .ZN(n1779) );
  ND2D1BWP12T U1834 ( .A1(n3106), .A2(n3100), .ZN(n1777) );
  TPOAI21D0BWP12T U1835 ( .A1(n1297), .A2(n1777), .B(n1780), .ZN(n867) );
  AOI21D1BWP12T U1836 ( .A1(n868), .A2(n1779), .B(n867), .ZN(n1787) );
  CKND1BWP12T U1837 ( .I(n1310), .ZN(n1788) );
  AOI21D1BWP12T U1838 ( .A1(n1791), .A2(n1788), .B(n836), .ZN(n869) );
  OA21D1BWP12T U1839 ( .A1(n1787), .A2(n870), .B(n869), .Z(n871) );
  TPAOI21D1BWP12T U1840 ( .A1(n1348), .A2(n1360), .B(n873), .ZN(n1785) );
  TPAOI21D1BWP12T U1841 ( .A1(n1745), .A2(n1743), .B(n874), .ZN(n1741) );
  TPAOI21D1BWP12T U1842 ( .A1(n1737), .A2(n1735), .B(n875), .ZN(n1733) );
  TPOAI21D1BWP12T U1843 ( .A1(n1733), .A2(n1575), .B(n1730), .ZN(n1797) );
  AO21D1BWP12T U1844 ( .A1(n1797), .A2(n1795), .B(n876), .Z(n1729) );
  INVD1BWP12T U1845 ( .I(n2594), .ZN(n1830) );
  INVD1BWP12T U1846 ( .I(n2846), .ZN(n2848) );
  ND2D1BWP12T U1847 ( .A1(n877), .A2(n2848), .ZN(n1846) );
  INVD1BWP12T U1848 ( .I(n3100), .ZN(n878) );
  ND2D1BWP12T U1849 ( .A1(n879), .A2(n878), .ZN(n880) );
  NR2D1BWP12T U1850 ( .A1(n1846), .A2(n880), .ZN(n1838) );
  ND2D1BWP12T U1851 ( .A1(n3059), .A2(n2193), .ZN(n1363) );
  CKND2D1BWP12T U1852 ( .A1(n691), .A2(n2192), .ZN(n881) );
  NR2D1BWP12T U1853 ( .A1(n1363), .A2(n881), .ZN(n882) );
  CKND2D1BWP12T U1854 ( .A1(n1838), .A2(n882), .ZN(n888) );
  ND2D1BWP12T U1855 ( .A1(n883), .A2(n2739), .ZN(n1849) );
  INVD1BWP12T U1856 ( .I(n2815), .ZN(n884) );
  INVD1BWP12T U1857 ( .I(n2785), .ZN(n2787) );
  ND2D1BWP12T U1858 ( .A1(n884), .A2(n2787), .ZN(n885) );
  NR2D1BWP12T U1859 ( .A1(n1849), .A2(n885), .ZN(n887) );
  ND2D1BWP12T U1860 ( .A1(n887), .A2(n886), .ZN(n1364) );
  NR2D1BWP12T U1861 ( .A1(n888), .A2(n1364), .ZN(n1822) );
  NR2XD0BWP12T U1862 ( .A1(n2679), .A2(n2915), .ZN(n1824) );
  ND2D1BWP12T U1863 ( .A1(n1824), .A2(n2650), .ZN(n1827) );
  NR2XD0BWP12T U1864 ( .A1(n1827), .A2(n2621), .ZN(n889) );
  ND2D1BWP12T U1865 ( .A1(n1822), .A2(n889), .ZN(n1831) );
  XNR2D1BWP12T U1866 ( .A1(n2532), .A2(n2979), .ZN(n2533) );
  INVD1BWP12T U1867 ( .I(n2533), .ZN(n926) );
  NR2D1BWP12T U1868 ( .A1(n2263), .A2(n2740), .ZN(n2333) );
  MUX2ND0BWP12T U1869 ( .I0(n2594), .I1(a[20]), .S(n1277), .ZN(n2223) );
  AOI22D0BWP12T U1870 ( .A1(n896), .A2(n2233), .B1(n2223), .B2(n2324), .ZN(
        n891) );
  ND2D1BWP12T U1871 ( .A1(n2350), .A2(n2353), .ZN(n2228) );
  INVD1BWP12T U1872 ( .I(n2228), .ZN(n2323) );
  MUX2ND0BWP12T U1873 ( .I0(n2679), .I1(n2915), .S(n1277), .ZN(n2225) );
  MUX2D1BWP12T U1874 ( .I0(n2621), .I1(n2652), .S(n1277), .Z(n1149) );
  INVD1BWP12T U1875 ( .I(n1149), .ZN(n2224) );
  AOI22D0BWP12T U1876 ( .A1(n2323), .A2(n2225), .B1(n2224), .B2(n2320), .ZN(
        n890) );
  CKND2D1BWP12T U1877 ( .A1(n891), .A2(n890), .ZN(n2317) );
  OAI22D0BWP12T U1878 ( .A1(n1111), .A2(n2228), .B1(n1160), .B2(n1353), .ZN(
        n893) );
  MUX2D1BWP12T U1879 ( .I0(n2815), .I1(n2785), .S(n1277), .Z(n2022) );
  OAI22D0BWP12T U1880 ( .A1(n1161), .A2(n1159), .B1(n2022), .B2(n1352), .ZN(
        n892) );
  NR2D1BWP12T U1881 ( .A1(n893), .A2(n892), .ZN(n2827) );
  MUX2D1BWP12T U1882 ( .I0(n2710), .I1(a[14]), .S(n1277), .Z(n2229) );
  MUX2ND0BWP12T U1883 ( .I0(a[13]), .I1(a[12]), .S(n1277), .ZN(n2238) );
  INVD0BWP12T U1884 ( .I(n2238), .ZN(n2024) );
  OAI22D0BWP12T U1885 ( .A1(n2229), .A2(n1352), .B1(n2024), .B2(n1353), .ZN(
        n895) );
  INVD1BWP12T U1886 ( .I(n2237), .ZN(n2023) );
  MUX2ND0BWP12T U1887 ( .I0(n2870), .I1(n2846), .S(n1277), .ZN(n2239) );
  INVD0BWP12T U1888 ( .I(n2239), .ZN(n2021) );
  OAI22D0BWP12T U1889 ( .A1(n2023), .A2(n1159), .B1(n2021), .B2(n2228), .ZN(
        n894) );
  NR2D1BWP12T U1890 ( .A1(n895), .A2(n894), .ZN(n2315) );
  IND2XD1BWP12T U1891 ( .A1(n2764), .B1(n2740), .ZN(n2337) );
  OAI22D0BWP12T U1892 ( .A1(n2827), .A2(n2258), .B1(n2315), .B2(n2337), .ZN(
        n901) );
  OR2XD1BWP12T U1893 ( .A1(n2764), .A2(n2740), .Z(n2327) );
  NR2D1BWP12T U1894 ( .A1(n2074), .A2(n2327), .ZN(n2114) );
  CKND0BWP12T U1895 ( .I(n2114), .ZN(n1811) );
  MUX2ND0BWP12T U1896 ( .I0(n2460), .I1(n2541), .S(n1277), .ZN(n2232) );
  INVD0BWP12T U1897 ( .I(n2232), .ZN(n2062) );
  MUX2ND0BWP12T U1898 ( .I0(n2498), .I1(a[28]), .S(n1277), .ZN(n2231) );
  CKND0BWP12T U1899 ( .I(n2231), .ZN(n2065) );
  OAI22D0BWP12T U1900 ( .A1(n2062), .A2(n2228), .B1(n2065), .B2(n1353), .ZN(
        n898) );
  MUX2ND0BWP12T U1901 ( .I0(n2358), .I1(a[26]), .S(n1277), .ZN(n2230) );
  CKND0BWP12T U1902 ( .I(n2230), .ZN(n2064) );
  ND2D1BWP12T U1903 ( .A1(n896), .A2(n1277), .ZN(n2250) );
  OAI22D0BWP12T U1904 ( .A1(n2064), .A2(n1159), .B1(n2250), .B2(a[30]), .ZN(
        n897) );
  INVD1BWP12T U1905 ( .I(n2327), .ZN(n2316) );
  OAI21D0BWP12T U1906 ( .A1(n898), .A2(n897), .B(n2316), .ZN(n899) );
  OAI211D0BWP12T U1907 ( .A1(n2979), .A2(n1811), .B(n899), .C(n2396), .ZN(n900) );
  AOI211D1BWP12T U1908 ( .A1(n2333), .A2(n2317), .B(n901), .C(n900), .ZN(n2279) );
  NR2D1BWP12T U1909 ( .A1(n2134), .A2(n2892), .ZN(n2988) );
  NR2D1BWP12T U1910 ( .A1(n2099), .A2(n902), .ZN(n2108) );
  AOI22D1BWP12T U1911 ( .A1(n1160), .A2(n2109), .B1(n2108), .B2(n1111), .ZN(
        n904) );
  CKND2D1BWP12T U1912 ( .A1(n2110), .A2(n2022), .ZN(n903) );
  OAI211D1BWP12T U1913 ( .A1(n2095), .A2(n1144), .B(n904), .C(n903), .ZN(n2144) );
  INVD1BWP12T U1914 ( .I(n2134), .ZN(n2139) );
  ND2D1BWP12T U1915 ( .A1(n2139), .A2(n2892), .ZN(n2121) );
  AOI22D0BWP12T U1916 ( .A1(n2109), .A2(n2223), .B1(n2108), .B2(n2225), .ZN(
        n906) );
  OAI211D0BWP12T U1917 ( .A1(n1149), .A2(n2095), .B(n906), .C(n905), .ZN(n2141) );
  NR2D0BWP12T U1918 ( .A1(n2892), .A2(n2114), .ZN(n907) );
  ND2D1BWP12T U1919 ( .A1(n907), .A2(n2134), .ZN(n2119) );
  INVD3BWP12T U1920 ( .I(n1150), .ZN(n2103) );
  TPNR2D0BWP12T U1921 ( .A1(n2095), .A2(n2237), .ZN(n909) );
  INVD1BWP12T U1922 ( .I(n2108), .ZN(n2046) );
  INVD1BWP12T U1923 ( .I(n2109), .ZN(n2047) );
  OAI22D1BWP12T U1924 ( .A1(n2046), .A2(n2239), .B1(n2047), .B2(n2238), .ZN(
        n908) );
  AOI211D1BWP12T U1925 ( .A1(n2229), .A2(n2103), .B(n909), .C(n908), .ZN(n2140) );
  TPNR2D0BWP12T U1926 ( .A1(n2095), .A2(n2230), .ZN(n911) );
  TPOAI22D0BWP12T U1927 ( .A1(n2046), .A2(n2232), .B1(n2047), .B2(n2231), .ZN(
        n910) );
  AOI211D1BWP12T U1928 ( .A1(n2103), .A2(a[30]), .B(n911), .C(n910), .ZN(n912)
         );
  OAI222D1BWP12T U1929 ( .A1(n2121), .A2(n2141), .B1(n2119), .B2(n2140), .C1(
        n2123), .C2(n912), .ZN(n2041) );
  AOI21D1BWP12T U1930 ( .A1(n2988), .A2(n2144), .B(n2041), .ZN(n913) );
  NR2D1BWP12T U1931 ( .A1(n913), .A2(n3004), .ZN(n924) );
  NR2D0BWP12T U1932 ( .A1(n2216), .A2(n2764), .ZN(n914) );
  TPND2D0BWP12T U1933 ( .A1(n1926), .A2(n914), .ZN(n2378) );
  NR2D1BWP12T U1934 ( .A1(n2393), .A2(n2856), .ZN(n1176) );
  NR2D1BWP12T U1935 ( .A1(n1176), .A2(n3090), .ZN(n3029) );
  XNR2D1BWP12T U1936 ( .A1(b[31]), .A2(n2979), .ZN(n2530) );
  INVD1BWP12T U1937 ( .I(n2530), .ZN(n915) );
  AOI22D1BWP12T U1938 ( .A1(n915), .A2(n1272), .B1(b[31]), .B2(n3020), .ZN(
        n922) );
  NR2D1BWP12T U1939 ( .A1(b[31]), .A2(op[2]), .ZN(n919) );
  CKND0BWP12T U1940 ( .I(n916), .ZN(n918) );
  CKND0BWP12T U1941 ( .I(n2215), .ZN(n917) );
  OAI22D1BWP12T U1942 ( .A1(n919), .A2(n918), .B1(b[31]), .B2(n917), .ZN(n920)
         );
  MUX2NXD0BWP12T U1943 ( .I0(n3105), .I1(n920), .S(n2979), .ZN(n921) );
  OAI211D1BWP12T U1944 ( .A1(n2378), .A2(n3029), .B(n922), .C(n921), .ZN(n923)
         );
  AOI211D1BWP12T U1945 ( .A1(n3067), .A2(n2279), .B(n924), .C(n923), .ZN(n925)
         );
  OAI21D1BWP12T U1946 ( .A1(n926), .A2(n3040), .B(n925), .ZN(n927) );
  ND3D1BWP12T U1947 ( .A1(n930), .A2(n929), .A3(n928), .ZN(n931) );
  AO21D1BWP12T U1948 ( .A1(n2524), .A2(n3117), .B(n931), .Z(result[31]) );
  INVD1P75BWP12T U1949 ( .I(n932), .ZN(n1557) );
  AOI21D1BWP12T U1950 ( .A1(n1557), .A2(n1549), .B(n1551), .ZN(n935) );
  INVD1BWP12T U1951 ( .I(n1553), .ZN(n933) );
  ND2D1BWP12T U1952 ( .A1(n933), .A2(n1552), .ZN(n934) );
  XOR2XD2BWP12T U1953 ( .A1(n935), .A2(n934), .Z(n1563) );
  FA1D0BWP12T U1954 ( .A(n937), .B(a[28]), .CI(n936), .CO(n1647), .S(n1722) );
  FA1D2BWP12T U1955 ( .A(b[28]), .B(a[28]), .CI(n938), .CO(n1570), .S(n1644)
         );
  CKND2D1BWP12T U1956 ( .A1(n1644), .A2(n3082), .ZN(n979) );
  FA1D0BWP12T U1957 ( .A(b[28]), .B(a[28]), .CI(n939), .CO(n1803), .S(n1806)
         );
  CKND2D1BWP12T U1958 ( .A1(n1806), .A2(n3093), .ZN(n978) );
  INR2D1BWP12T U1959 ( .A1(n2172), .B1(n1918), .ZN(n2106) );
  MUX2ND0BWP12T U1960 ( .I0(n2738), .I1(a[3]), .S(n1277), .ZN(n2271) );
  INVD1BWP12T U1961 ( .I(n2271), .ZN(n2098) );
  MUX2ND0BWP12T U1962 ( .I0(n2352), .I1(n2349), .S(n1277), .ZN(n2272) );
  INVD1BWP12T U1963 ( .I(n2272), .ZN(n1048) );
  MUX2ND0BWP12T U1964 ( .I0(a[12]), .I1(n2898), .S(n1277), .ZN(n2265) );
  CKND0BWP12T U1965 ( .I(n2265), .ZN(n942) );
  MUX2ND0BWP12T U1966 ( .I0(n2785), .I1(n2466), .S(n1277), .ZN(n2273) );
  OAI22D0BWP12T U1967 ( .A1(n2046), .A2(n2273), .B1(n2047), .B2(n2266), .ZN(
        n941) );
  MUX2ND0BWP12T U1968 ( .I0(n2846), .I1(n2815), .S(n1277), .ZN(n2274) );
  NR2D0BWP12T U1969 ( .A1(n2095), .A2(n2274), .ZN(n940) );
  AOI211D1BWP12T U1970 ( .A1(n942), .A2(n2103), .B(n941), .C(n940), .ZN(n2053)
         );
  MUX2ND0BWP12T U1971 ( .I0(a[20]), .I1(n2621), .S(n1277), .ZN(n2321) );
  CKND0BWP12T U1972 ( .I(n2321), .ZN(n945) );
  MUX2ND0BWP12T U1973 ( .I0(n2652), .I1(n2679), .S(n1277), .ZN(n2322) );
  MUX2ND0BWP12T U1974 ( .I0(a[14]), .I1(a[13]), .S(n1277), .ZN(n2267) );
  OAI22D0BWP12T U1975 ( .A1(n2047), .A2(n2322), .B1(n2046), .B2(n2267), .ZN(
        n944) );
  MUX2ND0BWP12T U1976 ( .I0(n2915), .I1(n2710), .S(n1277), .ZN(n2268) );
  NR2D0BWP12T U1977 ( .A1(n2095), .A2(n2268), .ZN(n943) );
  AOI211D1BWP12T U1978 ( .A1(n945), .A2(n2103), .B(n944), .C(n943), .ZN(n2051)
         );
  OAI22D0BWP12T U1979 ( .A1(n2053), .A2(n2119), .B1(n2051), .B2(n2121), .ZN(
        n951) );
  MUX2ND0BWP12T U1980 ( .I0(n2541), .I1(n2571), .S(n1277), .ZN(n2326) );
  CKND0BWP12T U1981 ( .I(n2326), .ZN(n948) );
  INVD1BWP12T U1982 ( .I(n2095), .ZN(n2107) );
  MUX2ND0BWP12T U1983 ( .I0(a[26]), .I1(n2460), .S(n1277), .ZN(n2246) );
  MUX2NXD1BWP12T U1984 ( .I0(a[22]), .I1(n2594), .S(n1277), .ZN(n2325) );
  OAI22D0BWP12T U1985 ( .A1(n2047), .A2(n2246), .B1(n2046), .B2(n2325), .ZN(
        n947) );
  MUX2ND0BWP12T U1986 ( .I0(a[28]), .I1(n2358), .S(n1277), .ZN(n2247) );
  NR2D1BWP12T U1987 ( .A1(n1150), .A2(n2247), .ZN(n946) );
  AOI211D0BWP12T U1988 ( .A1(n948), .A2(n2107), .B(n947), .C(n946), .ZN(n949)
         );
  NR2D0BWP12T U1989 ( .A1(n949), .A2(n2123), .ZN(n950) );
  AO211D1BWP12T U1990 ( .A1(n2988), .A2(n2014), .B(n951), .C(n950), .Z(n2042)
         );
  AOI21D0BWP12T U1991 ( .A1(n2198), .A2(n1272), .B(n3020), .ZN(n960) );
  ND2D1BWP12T U1992 ( .A1(n2393), .A2(n2979), .ZN(n1908) );
  OAI22D1BWP12T U1993 ( .A1(n1918), .A2(n2198), .B1(n2216), .B2(n1917), .ZN(
        n953) );
  OAI22D1BWP12T U1994 ( .A1(n1920), .A2(n2996), .B1(n1919), .B2(n2428), .ZN(
        n952) );
  NR2D1BWP12T U1995 ( .A1(n953), .A2(n952), .ZN(n2080) );
  CKND0BWP12T U1996 ( .I(n2080), .ZN(n954) );
  MUX2NXD0BWP12T U1997 ( .I0(n2979), .I1(n954), .S(n1903), .ZN(n1308) );
  IND2D0BWP12T U1998 ( .A1(n2979), .B1(n2740), .ZN(n955) );
  ND2D1BWP12T U1999 ( .A1(n2396), .A2(n955), .ZN(n2549) );
  INVD1BWP12T U2000 ( .I(n2549), .ZN(n1945) );
  NR2D1BWP12T U2001 ( .A1(n1945), .A2(n1976), .ZN(n1878) );
  AOI21D0BWP12T U2002 ( .A1(n1908), .A2(n1308), .B(n1878), .ZN(n1944) );
  CKND2D0BWP12T U2003 ( .A1(n1944), .A2(n3084), .ZN(n959) );
  MUX2ND0BWP12T U2004 ( .I0(n3102), .I1(n3101), .S(b[28]), .ZN(n956) );
  CKND2D0BWP12T U2005 ( .A1(n956), .A2(n3103), .ZN(n957) );
  MUX2ND0BWP12T U2006 ( .I0(n957), .I1(n3105), .S(n2198), .ZN(n958) );
  OAI211D1BWP12T U2007 ( .A1(n960), .A2(n937), .B(n959), .C(n958), .ZN(n974)
         );
  INVD0BWP12T U2008 ( .I(n3029), .ZN(n961) );
  ND2D1BWP12T U2009 ( .A1(n961), .A2(n1903), .ZN(n2991) );
  OAI22D0BWP12T U2010 ( .A1(n1048), .A2(n1353), .B1(n2106), .B2(n2207), .ZN(
        n963) );
  NR2XD0BWP12T U2011 ( .A1(n2098), .A2(n1352), .ZN(n962) );
  NR2D1BWP12T U2012 ( .A1(n963), .A2(n962), .ZN(n2737) );
  AOI22D0BWP12T U2013 ( .A1(n896), .A2(n2321), .B1(n2322), .B2(n2324), .ZN(
        n965) );
  AOI22D0BWP12T U2014 ( .A1(n2323), .A2(n2267), .B1(n2268), .B2(n2320), .ZN(
        n964) );
  ND2D1BWP12T U2015 ( .A1(n965), .A2(n964), .ZN(n2284) );
  AOI22D0BWP12T U2016 ( .A1(n896), .A2(n2247), .B1(n2325), .B2(n2323), .ZN(
        n967) );
  AOI22D0BWP12T U2017 ( .A1(n2324), .A2(n2246), .B1(n2326), .B2(n2320), .ZN(
        n966) );
  AOI21D0BWP12T U2018 ( .A1(n967), .A2(n966), .B(n2327), .ZN(n968) );
  AOI211D0BWP12T U2019 ( .A1(n2333), .A2(n2284), .B(n968), .C(n2383), .ZN(n972) );
  AOI22D0BWP12T U2020 ( .A1(n896), .A2(n2265), .B1(n2273), .B2(n2323), .ZN(
        n970) );
  AOI22D0BWP12T U2021 ( .A1(n2324), .A2(n2266), .B1(n2274), .B2(n2320), .ZN(
        n969) );
  ND2D1BWP12T U2022 ( .A1(n970), .A2(n969), .ZN(n2283) );
  INVD1BWP12T U2023 ( .I(n2337), .ZN(n2255) );
  TPND2D0BWP12T U2024 ( .A1(n2283), .A2(n2255), .ZN(n971) );
  OAI211D0BWP12T U2025 ( .A1(n2737), .A2(n2258), .B(n972), .C(n971), .ZN(n2245) );
  OAI22D1BWP12T U2026 ( .A1(n2991), .A2(n2080), .B1(n2245), .B2(n2928), .ZN(
        n973) );
  RCAOI211D0BWP12T U2027 ( .A1(n2042), .A2(n3091), .B(n974), .C(n973), .ZN(
        n977) );
  HA1D1BWP12T U2028 ( .A(n2198), .B(n975), .CO(n1817), .S(n1861) );
  ND2D1BWP12T U2029 ( .A1(n1861), .A2(n3096), .ZN(n976) );
  ND4D1BWP12T U2030 ( .A1(n979), .A2(n978), .A3(n977), .A4(n976), .ZN(n980) );
  AOI21D1BWP12T U2031 ( .A1(n382), .A2(n1722), .B(n980), .ZN(n983) );
  FA1D0BWP12T U2032 ( .A(n937), .B(a[28]), .CI(n981), .CO(n1376), .S(n1458) );
  CKND2D1BWP12T U2033 ( .A1(n1458), .A2(n3076), .ZN(n982) );
  OAI211D2BWP12T U2034 ( .A1(n2975), .A2(n984), .B(n983), .C(n982), .ZN(
        result[28]) );
  INVD1BWP12T U2035 ( .I(n985), .ZN(n1040) );
  INVD1BWP12T U2036 ( .I(n1039), .ZN(n986) );
  AOI21D1BWP12T U2037 ( .A1(n1557), .A2(n1040), .B(n986), .ZN(n991) );
  INVD1BWP12T U2038 ( .I(n987), .ZN(n989) );
  ND2D1BWP12T U2039 ( .A1(n989), .A2(n988), .ZN(n990) );
  FA1D0BWP12T U2040 ( .A(n993), .B(n2358), .CI(n992), .CO(n981), .S(n1453) );
  FA1D0BWP12T U2041 ( .A(n993), .B(n2358), .CI(n994), .CO(n936), .S(n1724) );
  INVD1BWP12T U2042 ( .I(n1724), .ZN(n1036) );
  FA1D0BWP12T U2043 ( .A(n2358), .B(b[27]), .CI(n995), .CO(n939), .S(n1805) );
  AOI22D0BWP12T U2044 ( .A1(n2109), .A2(n2225), .B1(n2108), .B2(n2238), .ZN(
        n997) );
  OAI211D0BWP12T U2045 ( .A1(n2229), .A2(n2095), .B(n997), .C(n996), .ZN(n2136) );
  INVD0BWP12T U2046 ( .I(n2136), .ZN(n1007) );
  NR2D1BWP12T U2047 ( .A1(n2101), .A2(n2099), .ZN(n2096) );
  CKND2D1BWP12T U2048 ( .A1(n2096), .A2(n1111), .ZN(n999) );
  CKND2D1BWP12T U2049 ( .A1(n2110), .A2(n1161), .ZN(n998) );
  ND2D1BWP12T U2050 ( .A1(n999), .A2(n998), .ZN(n2138) );
  INVD1BWP12T U2051 ( .I(n2138), .ZN(n2767) );
  INVD1BWP12T U2052 ( .I(n2022), .ZN(n2240) );
  TPAOI22D0BWP12T U2053 ( .A1(n2107), .A2(n2240), .B1(n2096), .B2(n2239), .ZN(
        n1001) );
  INVD1BWP12T U2054 ( .I(n1160), .ZN(n1145) );
  AOI22D1BWP12T U2055 ( .A1(n2103), .A2(n2237), .B1(n2108), .B2(n1145), .ZN(
        n1000) );
  ND2D1BWP12T U2056 ( .A1(n1001), .A2(n1000), .ZN(n2135) );
  MUX2D1BWP12T U2057 ( .I0(n2767), .I1(n2135), .S(n2134), .Z(n2893) );
  INVD1BWP12T U2058 ( .I(n2892), .ZN(n2130) );
  ND2XD0BWP12T U2059 ( .A1(n2893), .A2(n2130), .ZN(n1006) );
  CKND2D0BWP12T U2060 ( .A1(n2107), .A2(n2233), .ZN(n1003) );
  AOI22D0BWP12T U2061 ( .A1(n2109), .A2(n2232), .B1(n2108), .B2(n2223), .ZN(
        n1002) );
  OAI211D1BWP12T U2062 ( .A1(n2064), .A2(n1150), .B(n1003), .C(n1002), .ZN(
        n1004) );
  AOI21D0BWP12T U2063 ( .A1(n1004), .A2(n2933), .B(n2114), .ZN(n1005) );
  OAI211D1BWP12T U2064 ( .A1(n1007), .A2(n2121), .B(n1006), .C(n1005), .ZN(
        n2145) );
  HA1D1BWP12T U2065 ( .A(n2201), .B(n1008), .CO(n975), .S(n1864) );
  ND2D1BWP12T U2066 ( .A1(n1864), .A2(n3096), .ZN(n1031) );
  OA22XD1BWP12T U2067 ( .A1(n2022), .A2(n1159), .B1(n1160), .B2(n2228), .Z(
        n1010) );
  AOI22D0BWP12T U2068 ( .A1(n896), .A2(n2237), .B1(n2239), .B2(n2324), .ZN(
        n1009) );
  ND2D1BWP12T U2069 ( .A1(n1010), .A2(n1009), .ZN(n2294) );
  AOI22D1BWP12T U2070 ( .A1(n1161), .A2(n896), .B1(n2324), .B2(n1111), .ZN(
        n2292) );
  MUX2NXD0BWP12T U2071 ( .I0(n2294), .I1(n2292), .S(n2764), .ZN(n2905) );
  AOI22D0BWP12T U2072 ( .A1(n2224), .A2(n896), .B1(n2324), .B2(n2225), .ZN(
        n1012) );
  TPND2D0BWP12T U2073 ( .A1(n2238), .A2(n2323), .ZN(n1011) );
  OAI211D1BWP12T U2074 ( .A1(n2229), .A2(n1159), .B(n1012), .C(n1011), .ZN(
        n2293) );
  AOI22D0BWP12T U2075 ( .A1(n896), .A2(n2230), .B1(n2232), .B2(n2324), .ZN(
        n1014) );
  AOI22D0BWP12T U2076 ( .A1(n2323), .A2(n2223), .B1(n2233), .B2(n2320), .ZN(
        n1013) );
  AOI21D0BWP12T U2077 ( .A1(n1014), .A2(n1013), .B(n2327), .ZN(n1015) );
  AOI211D0BWP12T U2078 ( .A1(n2293), .A2(n2333), .B(n1015), .C(n2383), .ZN(
        n1016) );
  OA21XD0BWP12T U2079 ( .A1(n2905), .A2(n2377), .B(n1016), .Z(n2341) );
  OAI22D0BWP12T U2080 ( .A1(n1918), .A2(n2201), .B1(n1917), .B2(n2996), .ZN(
        n1018) );
  OAI22D1BWP12T U2081 ( .A1(n1920), .A2(n2428), .B1(n1919), .B2(n2198), .ZN(
        n1017) );
  NR2D1BWP12T U2082 ( .A1(n1018), .A2(n1017), .ZN(n1894) );
  MUX2D1BWP12T U2083 ( .I0(n2216), .I1(n1894), .S(n2207), .Z(n1019) );
  INR2D1BWP12T U2084 ( .A1(n1020), .B1(n1019), .ZN(n2013) );
  INVD1BWP12T U2085 ( .I(n2013), .ZN(n1021) );
  NR2D1BWP12T U2086 ( .A1(n1021), .A2(n2764), .ZN(n2020) );
  INVD1BWP12T U2087 ( .I(n2020), .ZN(n2401) );
  NR2XD0BWP12T U2088 ( .A1(n2401), .A2(n3029), .ZN(n1029) );
  INVD1BWP12T U2089 ( .I(n1970), .ZN(n1984) );
  ND2D1BWP12T U2090 ( .A1(n2764), .A2(n2979), .ZN(n2073) );
  INVD1BWP12T U2091 ( .I(n2073), .ZN(n1968) );
  AOI21D0BWP12T U2092 ( .A1(n1984), .A2(n2979), .B(n1968), .ZN(n1022) );
  OAI21D0BWP12T U2093 ( .A1(n1894), .A2(n2029), .B(n1022), .ZN(n1938) );
  TPND2D0BWP12T U2094 ( .A1(n1945), .A2(n1938), .ZN(n1942) );
  INVD1BWP12T U2095 ( .I(n1908), .ZN(n1966) );
  ND2D1BWP12T U2096 ( .A1(n1966), .A2(n3084), .ZN(n3028) );
  OAI21D0BWP12T U2097 ( .A1(n2358), .A2(n3099), .B(n3103), .ZN(n1026) );
  MUX2ND0BWP12T U2098 ( .I0(n3019), .I1(n3018), .S(b[27]), .ZN(n1023) );
  NR2D0BWP12T U2099 ( .A1(n1023), .A2(n3020), .ZN(n1024) );
  INVD1BWP12T U2100 ( .I(n3105), .ZN(n3023) );
  MUX2ND0BWP12T U2101 ( .I0(n1024), .I1(n3023), .S(n2201), .ZN(n1025) );
  AOI21D0BWP12T U2102 ( .A1(b[27]), .A2(n1026), .B(n1025), .ZN(n1027) );
  OAI211D0BWP12T U2103 ( .A1(n1942), .A2(n3071), .B(n3028), .C(n1027), .ZN(
        n1028) );
  RCAOI211D0BWP12T U2104 ( .A1(n3067), .A2(n2341), .B(n1029), .C(n1028), .ZN(
        n1030) );
  OAI211D1BWP12T U2105 ( .A1(n2145), .A2(n3004), .B(n1031), .C(n1030), .ZN(
        n1032) );
  AOI21D1BWP12T U2106 ( .A1(n1805), .A2(n3093), .B(n1032), .ZN(n1035) );
  FA1D2BWP12T U2107 ( .A(n2358), .B(b[27]), .CI(n1033), .CO(n938), .S(n1641)
         );
  CKND2D1BWP12T U2108 ( .A1(n1641), .A2(n3082), .ZN(n1034) );
  OAI211D1BWP12T U2109 ( .A1(n3047), .A2(n1036), .B(n1035), .C(n1034), .ZN(
        n1037) );
  AOI21D1BWP12T U2110 ( .A1(n3076), .A2(n1453), .B(n1037), .ZN(n1038) );
  IOA21D2BWP12T U2111 ( .A1(n1564), .A2(n3117), .B(n1038), .ZN(result[27]) );
  ND2D1BWP12T U2112 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XNR2XD2BWP12T U2113 ( .A1(n1557), .A2(n1041), .ZN(n1568) );
  INVD1P75BWP12T U2114 ( .I(n1568), .ZN(n1091) );
  FA1D0BWP12T U2115 ( .A(n2178), .B(a[26]), .CI(n1042), .CO(n992), .S(n1455)
         );
  FA1D0BWP12T U2116 ( .A(n2178), .B(a[26]), .CI(n1043), .CO(n994), .S(n1723)
         );
  INVD1BWP12T U2117 ( .I(n1723), .ZN(n1088) );
  FA1D0BWP12T U2118 ( .A(b[26]), .B(a[26]), .CI(n1044), .CO(n995), .S(n1800)
         );
  OAI22D1BWP12T U2119 ( .A1(n1918), .A2(n2996), .B1(n1919), .B2(n2216), .ZN(
        n2077) );
  MUX2D1BWP12T U2120 ( .I0(a[26]), .I1(n2358), .S(n1277), .Z(n1262) );
  NR2D1BWP12T U2121 ( .A1(n1920), .A2(a[28]), .ZN(n1046) );
  NR2D1BWP12T U2122 ( .A1(n1917), .A2(n2498), .ZN(n1045) );
  NR2D1BWP12T U2123 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  INVD1BWP12T U2124 ( .I(n1897), .ZN(n1194) );
  MUX2D1BWP12T U2125 ( .I0(n2077), .I1(n1194), .S(n2207), .Z(n2086) );
  INVD1BWP12T U2126 ( .I(n2086), .ZN(n1250) );
  INR2D1BWP12T U2127 ( .A1(n2172), .B1(n1920), .ZN(n1351) );
  CKND1BWP12T U2128 ( .I(n1351), .ZN(n1334) );
  NR2D0BWP12T U2129 ( .A1(n2101), .A2(n1334), .ZN(n1050) );
  NR2D1BWP12T U2130 ( .A1(n1048), .A2(n1351), .ZN(n1356) );
  INVD1BWP12T U2131 ( .I(n1356), .ZN(n1049) );
  TPAOI22D0BWP12T U2132 ( .A1(n2107), .A2(n2273), .B1(n2108), .B2(n2271), .ZN(
        n1052) );
  AOI22D1BWP12T U2133 ( .A1(n2103), .A2(n2266), .B1(n2096), .B2(n2274), .ZN(
        n1051) );
  ND2D1BWP12T U2134 ( .A1(n1052), .A2(n1051), .ZN(n2034) );
  MUX2D1BWP12T U2135 ( .I0(n1247), .I1(n2034), .S(n2134), .Z(n3098) );
  INVD0BWP12T U2136 ( .I(n3098), .ZN(n1061) );
  CKND2D0BWP12T U2137 ( .A1(n2107), .A2(n2267), .ZN(n1055) );
  AOI22D0BWP12T U2138 ( .A1(n2109), .A2(n2268), .B1(n2108), .B2(n2265), .ZN(
        n1054) );
  CKND2D0BWP12T U2139 ( .A1(n2110), .A2(n2322), .ZN(n1053) );
  ND3D1BWP12T U2140 ( .A1(n1055), .A2(n1054), .A3(n1053), .ZN(n2035) );
  INVD1BWP12T U2141 ( .I(n2121), .ZN(n2929) );
  CKND2D0BWP12T U2142 ( .A1(n2107), .A2(n2325), .ZN(n1058) );
  AOI22D0BWP12T U2143 ( .A1(n2109), .A2(n2326), .B1(n2108), .B2(n2321), .ZN(
        n1057) );
  CKND2D0BWP12T U2144 ( .A1(n2110), .A2(n2246), .ZN(n1056) );
  AOI31D0BWP12T U2145 ( .A1(n1058), .A2(n1057), .A3(n1056), .B(n2123), .ZN(
        n1059) );
  AOI211D0BWP12T U2146 ( .A1(n2035), .A2(n2929), .B(n2114), .C(n1059), .ZN(
        n1060) );
  OAI21D0BWP12T U2147 ( .A1(n1061), .A2(n2892), .B(n1060), .ZN(n2146) );
  OA21D1BWP12T U2148 ( .A1(n1250), .A2(n2327), .B(n2146), .Z(n1083) );
  HA1D1BWP12T U2149 ( .A(n2200), .B(n1062), .CO(n1008), .S(n1863) );
  ND2D1BWP12T U2150 ( .A1(n1863), .A2(n3096), .ZN(n1082) );
  AOI22D0BWP12T U2151 ( .A1(n2323), .A2(n2271), .B1(n2273), .B2(n2320), .ZN(
        n1064) );
  AOI22D0BWP12T U2152 ( .A1(n896), .A2(n2266), .B1(n2274), .B2(n2324), .ZN(
        n1063) );
  ND2D1BWP12T U2153 ( .A1(n1064), .A2(n1063), .ZN(n2306) );
  AOI21D1BWP12T U2154 ( .A1(n1351), .A2(n1104), .B(n896), .ZN(n1065) );
  NR2D1BWP12T U2155 ( .A1(n1356), .A2(n1065), .ZN(n2264) );
  INVD1BWP12T U2156 ( .I(n2264), .ZN(n1239) );
  MUX2ND0BWP12T U2157 ( .I0(n2306), .I1(n1239), .S(n2764), .ZN(n3107) );
  NR2D0BWP12T U2158 ( .A1(n3107), .A2(n2377), .ZN(n1070) );
  OAI22D0BWP12T U2159 ( .A1(n1352), .A2(n2322), .B1(n2268), .B2(n1353), .ZN(
        n2303) );
  OAI22D0BWP12T U2160 ( .A1(n2228), .A2(n2265), .B1(n2267), .B2(n1159), .ZN(
        n2302) );
  INVD1BWP12T U2161 ( .I(n2333), .ZN(n2287) );
  TPNR3D0BWP12T U2162 ( .A1(n2303), .A2(n2302), .A3(n2287), .ZN(n1069) );
  AOI22D0BWP12T U2163 ( .A1(n2323), .A2(n2321), .B1(n2325), .B2(n2320), .ZN(
        n1067) );
  AOI22D0BWP12T U2164 ( .A1(n896), .A2(n2246), .B1(n2326), .B2(n2324), .ZN(
        n1066) );
  AOI21D0BWP12T U2165 ( .A1(n1067), .A2(n1066), .B(n2327), .ZN(n1068) );
  NR4D0BWP12T U2166 ( .A1(n1070), .A2(n1069), .A3(n1068), .A4(n2383), .ZN(
        n2342) );
  ND2D1BWP12T U2167 ( .A1(n1918), .A2(n2979), .ZN(n1071) );
  INR2D1BWP12T U2168 ( .A1(n1071), .B1(n2077), .ZN(n1332) );
  CKND0BWP12T U2169 ( .I(n1332), .ZN(n1072) );
  MUX2ND0BWP12T U2170 ( .I0(n1072), .I1(n1194), .S(n2207), .ZN(n1073) );
  OA21XD1BWP12T U2171 ( .A1(n1073), .A2(n2764), .B(n2073), .Z(n1901) );
  INVD1BWP12T U2172 ( .I(n1878), .ZN(n1886) );
  ND2D0BWP12T U2173 ( .A1(n1886), .A2(n3084), .ZN(n1179) );
  AOI21D0BWP12T U2174 ( .A1(n1901), .A2(n1908), .B(n1179), .ZN(n1080) );
  CKND0BWP12T U2175 ( .I(n1176), .ZN(n2660) );
  INVD1BWP12T U2176 ( .I(n2764), .ZN(n2314) );
  INR2D1BWP12T U2177 ( .A1(n2314), .B1(n1250), .ZN(n3092) );
  INVD1BWP12T U2178 ( .I(n3092), .ZN(n2400) );
  MUX2ND0BWP12T U2179 ( .I0(n3102), .I1(n3101), .S(b[26]), .ZN(n1074) );
  CKND2D0BWP12T U2180 ( .A1(n1074), .A2(n3103), .ZN(n1075) );
  MUX2ND0BWP12T U2181 ( .I0(n1075), .I1(n3105), .S(n2200), .ZN(n1078) );
  OAI21D0BWP12T U2182 ( .A1(a[26]), .A2(n3099), .B(n3103), .ZN(n1076) );
  CKND2D0BWP12T U2183 ( .A1(n1076), .A2(b[26]), .ZN(n1077) );
  OAI211D1BWP12T U2184 ( .A1(n2660), .A2(n2400), .B(n1078), .C(n1077), .ZN(
        n1079) );
  AOI211XD0BWP12T U2185 ( .A1(n3067), .A2(n2342), .B(n1080), .C(n1079), .ZN(
        n1081) );
  OAI211D1BWP12T U2186 ( .A1(n1083), .A2(n3004), .B(n1082), .C(n1081), .ZN(
        n1084) );
  AOI21D1BWP12T U2187 ( .A1(n1800), .A2(n3093), .B(n1084), .ZN(n1087) );
  FA1D2BWP12T U2188 ( .A(b[26]), .B(a[26]), .CI(n1085), .CO(n1033), .S(n1643)
         );
  CKND2D1BWP12T U2189 ( .A1(n1643), .A2(n3082), .ZN(n1086) );
  OAI211D1BWP12T U2190 ( .A1(n3047), .A2(n1088), .B(n1087), .C(n1086), .ZN(
        n1089) );
  AOI21D1BWP12T U2191 ( .A1(n3076), .A2(n1455), .B(n1089), .ZN(n1090) );
  RCOAI21D2BWP12T U2192 ( .A1(n1091), .A2(n2975), .B(n1090), .ZN(result[26])
         );
  MUX2ND0BWP12T U2193 ( .I0(n1093), .I1(n1092), .S(n2353), .ZN(n1094) );
  OAI21D0BWP12T U2194 ( .A1(n2216), .A2(n2228), .B(n1094), .ZN(n1869) );
  OAI22D1BWP12T U2195 ( .A1(n1973), .A2(n1970), .B1(n1971), .B2(n2029), .ZN(
        n1105) );
  AOI21D1BWP12T U2196 ( .A1(n1869), .A2(n2764), .B(n1105), .ZN(n1895) );
  INVD1BWP12T U2197 ( .I(n1895), .ZN(n2688) );
  OAI22D1BWP12T U2198 ( .A1(n1974), .A2(n1986), .B1(n1095), .B2(n1989), .ZN(
        n1099) );
  INVD1BWP12T U2199 ( .I(n2250), .ZN(n1925) );
  AOI22D1BWP12T U2200 ( .A1(n1925), .A2(n2352), .B1(n1926), .B2(n2349), .ZN(
        n1097) );
  INR2D1BWP12T U2201 ( .A1(n1277), .B1(n1353), .ZN(n1923) );
  NR2D1BWP12T U2202 ( .A1(n1353), .A2(n1277), .ZN(n1924) );
  AOI22D1BWP12T U2203 ( .A1(n2738), .A2(n1923), .B1(n1924), .B2(a[3]), .ZN(
        n1096) );
  AOI21D0BWP12T U2204 ( .A1(n1097), .A2(n1096), .B(n2764), .ZN(n1098) );
  AOI211D1BWP12T U2205 ( .A1(n1984), .A2(n1100), .B(n1099), .C(n1098), .ZN(
        n2010) );
  AOI21D1BWP12T U2206 ( .A1(n2010), .A2(n2377), .B(n2383), .ZN(n2387) );
  OAI21D1BWP12T U2207 ( .A1(n2688), .A2(n2377), .B(n2387), .ZN(n1101) );
  CKND2D1BWP12T U2208 ( .A1(n1101), .A2(n1991), .ZN(n1981) );
  ND2D1BWP12T U2209 ( .A1(n2684), .A2(n2740), .ZN(n2386) );
  INVD1BWP12T U2210 ( .I(n2386), .ZN(n1106) );
  NR2D1BWP12T U2211 ( .A1(n1106), .A2(n2856), .ZN(n1107) );
  INVD1BWP12T U2212 ( .I(n1108), .ZN(n1222) );
  INVD1BWP12T U2213 ( .I(n1221), .ZN(n1109) );
  ND2D1BWP12T U2214 ( .A1(n1109), .A2(n1220), .ZN(n1110) );
  CKXOR2D1BWP12T U2215 ( .A1(n1222), .A2(n1110), .Z(n1427) );
  ND2D1BWP12T U2216 ( .A1(n1111), .A2(n896), .ZN(n2291) );
  INVD1BWP12T U2217 ( .I(n2291), .ZN(n1164) );
  AOI22D1BWP12T U2218 ( .A1(n1427), .A2(n3076), .B1(n2826), .B2(n1164), .ZN(
        n1130) );
  INVD1BWP12T U2219 ( .I(n1115), .ZN(n1228) );
  INVD1BWP12T U2220 ( .I(n1227), .ZN(n1116) );
  CKND2D1BWP12T U2221 ( .A1(n1116), .A2(n1226), .ZN(n1117) );
  CKXOR2D1BWP12T U2222 ( .A1(n1228), .A2(n1117), .Z(n1611) );
  AOI22D0BWP12T U2223 ( .A1(n1698), .A2(n382), .B1(n3082), .B2(n1611), .ZN(
        n1129) );
  ND2D1BWP12T U2224 ( .A1(n1116), .A2(n1119), .ZN(n1120) );
  XOR2XD1BWP12T U2225 ( .A1(n1120), .A2(n1271), .Z(n1764) );
  NR2D1BWP12T U2226 ( .A1(n2010), .A2(n2807), .ZN(n1127) );
  XNR2XD0BWP12T U2227 ( .A1(n1121), .A2(n2449), .ZN(n1836) );
  AOI21D1BWP12T U2228 ( .A1(n1122), .A2(n3103), .B(n2210), .ZN(n1125) );
  AOI21D1BWP12T U2229 ( .A1(n2210), .A2(n1272), .B(n3020), .ZN(n1123) );
  OAI22D1BWP12T U2230 ( .A1(n1123), .A2(n2179), .B1(n2349), .B2(n3023), .ZN(
        n1124) );
  AO211D0BWP12T U2231 ( .A1(n1836), .A2(n3096), .B(n1125), .C(n1124), .Z(n1126) );
  AOI211D1BWP12T U2232 ( .A1(n1764), .A2(n3093), .B(n1127), .C(n1126), .ZN(
        n1128) );
  AOI21D1BWP12T U2233 ( .A1(n1516), .A2(n3117), .B(n1132), .ZN(n1133) );
  IOA21D2BWP12T U2234 ( .A1(n3084), .A2(n1981), .B(n1133), .ZN(result[1]) );
  INVD1P75BWP12T U2235 ( .I(n1134), .ZN(n1546) );
  TPOAI21D1BWP12T U2236 ( .A1(n1546), .A2(n1542), .B(n1543), .ZN(n1139) );
  INVD1BWP12T U2237 ( .I(n1135), .ZN(n1137) );
  ND2D1BWP12T U2238 ( .A1(n1137), .A2(n1136), .ZN(n1138) );
  XNR2XD2BWP12T U2239 ( .A1(n1139), .A2(n1138), .ZN(n1547) );
  FA1D0BWP12T U2240 ( .A(n1141), .B(n2460), .CI(n1140), .CO(n1042), .S(n1454)
         );
  FA1D0BWP12T U2241 ( .A(n1141), .B(n2460), .CI(n1142), .CO(n1043), .S(n1721)
         );
  INVD1BWP12T U2242 ( .I(n1721), .ZN(n1187) );
  FA1D2BWP12T U2243 ( .A(n2460), .B(b[25]), .CI(n1143), .CO(n1044), .S(n1802)
         );
  TPAOI22D0BWP12T U2244 ( .A1(n2107), .A2(n1145), .B1(n2108), .B2(n1144), .ZN(
        n1147) );
  AOI22D1BWP12T U2245 ( .A1(n2103), .A2(n2239), .B1(n2096), .B2(n2240), .ZN(
        n1146) );
  ND2D1BWP12T U2246 ( .A1(n1147), .A2(n1146), .ZN(n2122) );
  MUX2D1BWP12T U2247 ( .I0(n2120), .I1(n2122), .S(n2134), .Z(n2033) );
  CKND2D0BWP12T U2248 ( .A1(n2033), .A2(n2130), .ZN(n1157) );
  INVD0BWP12T U2249 ( .I(n2225), .ZN(n2059) );
  AOI22D1BWP12T U2250 ( .A1(n2103), .A2(n2059), .B1(n2108), .B2(n2023), .ZN(
        n2124) );
  CKND2D0BWP12T U2251 ( .A1(n2109), .A2(n2229), .ZN(n1148) );
  OA21XD0BWP12T U2252 ( .A1(n2095), .A2(n2238), .B(n1148), .Z(n2125) );
  CKND0BWP12T U2253 ( .I(n2233), .ZN(n2063) );
  OAI22D0BWP12T U2254 ( .A1(n2047), .A2(n2063), .B1(n2046), .B2(n1149), .ZN(
        n1152) );
  NR2D1BWP12T U2255 ( .A1(n1150), .A2(n2062), .ZN(n1151) );
  AOI211D0BWP12T U2256 ( .A1(n2107), .A2(n2223), .B(n1152), .C(n1151), .ZN(
        n1153) );
  OAI21D0BWP12T U2257 ( .A1(n1153), .A2(n2123), .B(n1811), .ZN(n1154) );
  AOI31D0BWP12T U2258 ( .A1(n2929), .A2(n2124), .A3(n2125), .B(n1154), .ZN(
        n1156) );
  MUX2NXD0BWP12T U2259 ( .I0(n2432), .I1(n1972), .S(n2207), .ZN(n1155) );
  AOI22D1BWP12T U2260 ( .A1(n1157), .A2(n1156), .B1(n2316), .B2(n1155), .ZN(
        n2147) );
  HA1D1BWP12T U2261 ( .A(n2202), .B(n1158), .CO(n1062), .S(n1859) );
  CKND2D1BWP12T U2262 ( .A1(n1859), .A2(n3096), .ZN(n1182) );
  OAI22D0BWP12T U2263 ( .A1(n2021), .A2(n1352), .B1(n2022), .B2(n1353), .ZN(
        n1163) );
  OAI22D0BWP12T U2264 ( .A1(n1161), .A2(n2228), .B1(n1160), .B2(n1159), .ZN(
        n1162) );
  NR2D1BWP12T U2265 ( .A1(n1163), .A2(n1162), .ZN(n2288) );
  MUX2NXD0BWP12T U2266 ( .I0(n2288), .I1(n1164), .S(n2764), .ZN(n2880) );
  CKND0BWP12T U2267 ( .I(n2880), .ZN(n1171) );
  CKND0BWP12T U2268 ( .I(n2229), .ZN(n2056) );
  AOI22D0BWP12T U2269 ( .A1(n2324), .A2(n2056), .B1(n896), .B2(n2225), .ZN(
        n1166) );
  AOI22D0BWP12T U2270 ( .A1(n2323), .A2(n2237), .B1(n2238), .B2(n2320), .ZN(
        n1165) );
  ND2D1BWP12T U2271 ( .A1(n1166), .A2(n1165), .ZN(n2286) );
  AOI22D0BWP12T U2272 ( .A1(n896), .A2(n2232), .B1(n2233), .B2(n2324), .ZN(
        n1168) );
  AOI22D0BWP12T U2273 ( .A1(n2224), .A2(n2323), .B1(n2223), .B2(n2320), .ZN(
        n1167) );
  AOI21D0BWP12T U2274 ( .A1(n1168), .A2(n1167), .B(n2327), .ZN(n1169) );
  AOI211D0BWP12T U2275 ( .A1(n2286), .A2(n2333), .B(n1169), .C(n2383), .ZN(
        n1170) );
  OAI21D0BWP12T U2276 ( .A1(n1171), .A2(n2377), .B(n1170), .ZN(n2296) );
  CKND2D1BWP12T U2277 ( .A1(n1908), .A2(n2073), .ZN(n1876) );
  AOI21D0BWP12T U2278 ( .A1(n1869), .A2(n2263), .B(n1876), .ZN(n1879) );
  OAI21D0BWP12T U2279 ( .A1(n2460), .A2(n3099), .B(n3103), .ZN(n1175) );
  MUX2ND0BWP12T U2280 ( .I0(n3019), .I1(n3018), .S(b[25]), .ZN(n1172) );
  NR2D0BWP12T U2281 ( .A1(n1172), .A2(n3020), .ZN(n1173) );
  MUX2ND0BWP12T U2282 ( .I0(n1173), .I1(n3023), .S(n2202), .ZN(n1174) );
  AOI21D0BWP12T U2283 ( .A1(b[25]), .A2(n1175), .B(n1174), .ZN(n1178) );
  OAI22D1BWP12T U2284 ( .A1(n2432), .A2(n1970), .B1(n1972), .B2(n2029), .ZN(
        n2397) );
  TPND2D0BWP12T U2285 ( .A1(n1176), .A2(n2397), .ZN(n1177) );
  OAI211D1BWP12T U2286 ( .A1(n1179), .A2(n1879), .B(n1178), .C(n1177), .ZN(
        n1180) );
  IAO21D1BWP12T U2287 ( .A1(n2296), .A2(n2928), .B(n1180), .ZN(n1181) );
  OAI211D1BWP12T U2288 ( .A1(n2147), .A2(n3004), .B(n1182), .C(n1181), .ZN(
        n1183) );
  AOI21D1BWP12T U2289 ( .A1(n1802), .A2(n3093), .B(n1183), .ZN(n1186) );
  FA1D2BWP12T U2290 ( .A(n2460), .B(b[25]), .CI(n1184), .CO(n1085), .S(n1642)
         );
  CKND2D1BWP12T U2291 ( .A1(n1642), .A2(n3082), .ZN(n1185) );
  OAI211D1BWP12T U2292 ( .A1(n3047), .A2(n1187), .B(n1186), .C(n1185), .ZN(
        n1188) );
  AOI21D1BWP12T U2293 ( .A1(n3076), .A2(n1454), .B(n1188), .ZN(n1189) );
  IOA21D2BWP12T U2294 ( .A1(n1547), .A2(n3117), .B(n1189), .ZN(result[25]) );
  OAI22D1BWP12T U2295 ( .A1(n1920), .A2(n2952), .B1(n1919), .B2(n2623), .ZN(
        n1190) );
  NR2D1BWP12T U2296 ( .A1(n1191), .A2(n1190), .ZN(n1987) );
  OAI22D1BWP12T U2297 ( .A1(n1920), .A2(n2544), .B1(n1919), .B2(n2574), .ZN(
        n1192) );
  NR2D1BWP12T U2298 ( .A1(n1193), .A2(n1192), .ZN(n1896) );
  MUX2ND0BWP12T U2299 ( .I0(n1987), .I1(n1896), .S(n2353), .ZN(n1906) );
  NR2D1BWP12T U2300 ( .A1(n1906), .A2(n2764), .ZN(n2040) );
  NR2D1BWP12T U2301 ( .A1(n1194), .A2(n1989), .ZN(n1195) );
  TPNR2D1BWP12T U2302 ( .A1(n2040), .A2(n1195), .ZN(n1215) );
  CKND0BWP12T U2303 ( .I(n1986), .ZN(n1214) );
  CKND2D1BWP12T U2304 ( .A1(n1332), .A2(n1214), .ZN(n1196) );
  ND2D1BWP12T U2305 ( .A1(n1215), .A2(n1196), .ZN(n1909) );
  OAI21D0BWP12T U2306 ( .A1(n1909), .A2(n2383), .B(n2393), .ZN(n1210) );
  OAI22D1BWP12T U2307 ( .A1(a[12]), .A2(n1920), .B1(n1919), .B2(n2898), .ZN(
        n1197) );
  NR2D1BWP12T U2308 ( .A1(n1198), .A2(n1197), .ZN(n1985) );
  OAI22D1BWP12T U2309 ( .A1(n1920), .A2(n2917), .B1(n1919), .B2(n2712), .ZN(
        n1199) );
  NR2D1BWP12T U2310 ( .A1(n1200), .A2(n1199), .ZN(n1990) );
  NR2D1BWP12T U2311 ( .A1(n1990), .A2(n1986), .ZN(n1201) );
  AOI211D1BWP12T U2312 ( .A1(n1985), .A2(n2076), .B(n1201), .C(n2740), .ZN(
        n1209) );
  OAI22D1BWP12T U2313 ( .A1(n1920), .A2(n2848), .B1(n1919), .B2(n2819), .ZN(
        n1202) );
  NR2D1BWP12T U2314 ( .A1(n1203), .A2(n1202), .ZN(n1988) );
  ND2D1BWP12T U2315 ( .A1(n1988), .A2(n2353), .ZN(n1207) );
  TPAOI21D0BWP12T U2316 ( .A1(n1926), .A2(n1832), .B(n2764), .ZN(n1206) );
  INVD1BWP12T U2317 ( .I(a[3]), .ZN(n2760) );
  AOI22D1BWP12T U2318 ( .A1(n1925), .A2(n2760), .B1(n1923), .B2(n2206), .ZN(
        n1205) );
  TPND2D0BWP12T U2319 ( .A1(n1924), .A2(n2739), .ZN(n1204) );
  ND4D1BWP12T U2320 ( .A1(n1207), .A2(n1206), .A3(n1205), .A4(n1204), .ZN(
        n1208) );
  ND2D1BWP12T U2321 ( .A1(n1209), .A2(n1208), .ZN(n1218) );
  AOI21D1BWP12T U2322 ( .A1(n1210), .A2(n1218), .B(n1976), .ZN(n1995) );
  ND2XD0BWP12T U2323 ( .A1(n1514), .A2(n3117), .ZN(n1255) );
  INVD1BWP12T U2324 ( .I(n2077), .ZN(n2992) );
  CKND2D1BWP12T U2325 ( .A1(n2992), .A2(n1214), .ZN(n1217) );
  INVD1BWP12T U2326 ( .I(n1215), .ZN(n1216) );
  INR2D2BWP12T U2327 ( .A1(n1217), .B1(n1216), .ZN(n2398) );
  CKND2D1BWP12T U2328 ( .A1(n2398), .A2(n2396), .ZN(n1219) );
  INVD1BWP12T U2329 ( .I(n1218), .ZN(n1248) );
  INVD1BWP12T U2330 ( .I(n2856), .ZN(n3080) );
  CKND1BWP12T U2331 ( .I(n3076), .ZN(n3089) );
  INVD0BWP12T U2332 ( .I(n1223), .ZN(n1225) );
  INVD1BWP12T U2333 ( .I(n1428), .ZN(n1246) );
  TPOAI21D0BWP12T U2334 ( .A1(n1228), .A2(n1227), .B(n1226), .ZN(n1230) );
  CKND0BWP12T U2335 ( .I(n1747), .ZN(n1232) );
  CKND2D0BWP12T U2336 ( .A1(n1232), .A2(n1746), .ZN(n1229) );
  XNR2D1BWP12T U2337 ( .A1(n1230), .A2(n1229), .ZN(n1610) );
  INVD1P75BWP12T U2338 ( .I(n2826), .ZN(n1240) );
  INVD1BWP12T U2339 ( .I(n1231), .ZN(n1748) );
  CKND2D0BWP12T U2340 ( .A1(n1232), .A2(n1746), .ZN(n1233) );
  XOR2XD1BWP12T U2341 ( .A1(n1748), .A2(n1233), .Z(n1765) );
  MUX2ND0BWP12T U2342 ( .I0(n3102), .I1(n3101), .S(n2353), .ZN(n1234) );
  AOI21D0BWP12T U2343 ( .A1(n3103), .A2(n1234), .B(n1832), .ZN(n1237) );
  AOI21D0BWP12T U2344 ( .A1(n1272), .A2(n1832), .B(n3020), .ZN(n1235) );
  OAI22D0BWP12T U2345 ( .A1(n1235), .A2(n2207), .B1(n2352), .B2(n3023), .ZN(
        n1236) );
  AOI211D1BWP12T U2346 ( .A1(n1765), .A2(n3093), .B(n1237), .C(n1236), .ZN(
        n1238) );
  AOI21D1BWP12T U2347 ( .A1(n3082), .A2(n1610), .B(n1241), .ZN(n1245) );
  INVD1BWP12T U2348 ( .I(n1242), .ZN(n1687) );
  CKND0BWP12T U2349 ( .I(n1243), .ZN(n1833) );
  XNR2D0BWP12T U2350 ( .A1(n1833), .A2(n2352), .ZN(n1835) );
  AOI22D0BWP12T U2351 ( .A1(n1699), .A2(n382), .B1(n3096), .B2(n1835), .ZN(
        n1244) );
  OAI211D1BWP12T U2352 ( .A1(n3089), .A2(n1246), .B(n1245), .C(n1244), .ZN(
        n1253) );
  INVD1BWP12T U2353 ( .I(n1247), .ZN(n2037) );
  CKND0BWP12T U2354 ( .I(n2258), .ZN(n2332) );
  NR2D1BWP12T U2355 ( .A1(n1906), .A2(n2337), .ZN(n1249) );
  AOI211D1BWP12T U2356 ( .A1(n2332), .A2(n1250), .B(n1249), .C(n1248), .ZN(
        n1251) );
  AOI21D1BWP12T U2357 ( .A1(n2037), .A2(n2933), .B(n1251), .ZN(n2016) );
  NR2D1BWP12T U2358 ( .A1(n2016), .A2(n3004), .ZN(n1252) );
  AOI211D1BWP12T U2359 ( .A1(n2395), .A2(n3080), .B(n1253), .C(n1252), .ZN(
        n1254) );
  OAI211D2BWP12T U2360 ( .A1(n1995), .A2(n3071), .B(n1255), .C(n1254), .ZN(
        result[2]) );
  OAI22D1BWP12T U2361 ( .A1(n1920), .A2(n2192), .B1(n1919), .B2(n3059), .ZN(
        n1256) );
  NR2D1BWP12T U2362 ( .A1(n1257), .A2(n1256), .ZN(n1955) );
  OAI22D1BWP12T U2363 ( .A1(n1920), .A2(n2787), .B1(n1919), .B2(n2206), .ZN(
        n1258) );
  NR2D1BWP12T U2364 ( .A1(n1259), .A2(n1258), .ZN(n1884) );
  OAI22D1BWP12T U2365 ( .A1(n3100), .A2(n1920), .B1(n1919), .B2(n2870), .ZN(
        n1260) );
  NR2D1BWP12T U2366 ( .A1(n1261), .A2(n1260), .ZN(n1952) );
  INR2D1BWP12T U2367 ( .A1(n2106), .B1(n2029), .ZN(n1276) );
  INVD1BWP12T U2368 ( .I(n2393), .ZN(n2402) );
  OAI22D1BWP12T U2369 ( .A1(n1919), .A2(n2596), .B1(n1917), .B2(n2574), .ZN(
        n1263) );
  NR2D1BWP12T U2370 ( .A1(n1264), .A2(n1263), .ZN(n1953) );
  OAI22D0BWP12T U2371 ( .A1(n1941), .A2(n1989), .B1(n1953), .B2(n1970), .ZN(
        n1268) );
  OAI22D1BWP12T U2372 ( .A1(n1920), .A2(n2650), .B1(n1917), .B2(n2623), .ZN(
        n1265) );
  NR2D1BWP12T U2373 ( .A1(n1266), .A2(n1265), .ZN(n1956) );
  OAI22D0BWP12T U2374 ( .A1(n2080), .A2(n1986), .B1(n1956), .B2(n2029), .ZN(
        n1267) );
  NR2D1BWP12T U2375 ( .A1(n1268), .A2(n1267), .ZN(n2922) );
  NR2D1BWP12T U2376 ( .A1(n2922), .A2(n2377), .ZN(n2088) );
  AOI22D1BWP12T U2377 ( .A1(n2087), .A2(n2402), .B1(n2396), .B2(n2088), .ZN(
        n1979) );
  XNR2XD0BWP12T U2378 ( .A1(n1269), .A2(n2172), .ZN(n1697) );
  INR2D0BWP12T U2379 ( .A1(n306), .B1(n2449), .ZN(n1515) );
  INVD1BWP12T U2380 ( .I(n1273), .ZN(n1275) );
  INVD1BWP12T U2381 ( .I(n1276), .ZN(n2221) );
  INVD1BWP12T U2382 ( .I(n1979), .ZN(n2384) );
  INVD1BWP12T U2383 ( .I(n1280), .ZN(n1492) );
  ND2D1BWP12T U2384 ( .A1(n1283), .A2(n1282), .ZN(n1284) );
  XOR2XD1BWP12T U2385 ( .A1(n1285), .A2(n1284), .Z(n1523) );
  INVD1BWP12T U2386 ( .I(n1403), .ZN(n1433) );
  CKND2D1BWP12T U2387 ( .A1(n1433), .A2(n1713), .ZN(n1288) );
  INVD1BWP12T U2388 ( .I(n1402), .ZN(n1436) );
  AOI21D1BWP12T U2389 ( .A1(n1436), .A2(n1713), .B(n1295), .ZN(n1287) );
  OAI21D1BWP12T U2390 ( .A1(n1437), .A2(n1288), .B(n1287), .ZN(n1292) );
  ND2D1BWP12T U2391 ( .A1(n286), .A2(n1290), .ZN(n1291) );
  XNR2XD1BWP12T U2392 ( .A1(n1292), .A2(n1291), .ZN(n1405) );
  INVD1BWP12T U2393 ( .I(n1293), .ZN(n1706) );
  NR2XD0BWP12T U2394 ( .A1(n1706), .A2(n1707), .ZN(n1709) );
  INVD1BWP12T U2395 ( .I(n1294), .ZN(n1705) );
  OAI21D1BWP12T U2396 ( .A1(n1705), .A2(n1707), .B(n1708), .ZN(n1710) );
  INVD1BWP12T U2397 ( .I(n1588), .ZN(n1593) );
  INVD1BWP12T U2398 ( .I(n1297), .ZN(n1781) );
  ND2XD0BWP12T U2399 ( .A1(n1593), .A2(n1781), .ZN(n1300) );
  INVD1BWP12T U2400 ( .I(n1587), .ZN(n1596) );
  INVD1BWP12T U2401 ( .I(n1780), .ZN(n1298) );
  AOI21D1BWP12T U2402 ( .A1(n1596), .A2(n1781), .B(n1298), .ZN(n1299) );
  OAI21D1BWP12T U2403 ( .A1(n1607), .A2(n1300), .B(n1299), .ZN(n1302) );
  CKND2D1BWP12T U2404 ( .A1(n1789), .A2(n1310), .ZN(n1301) );
  XNR2XD1BWP12T U2405 ( .A1(n1302), .A2(n1301), .ZN(n1589) );
  INVD0BWP12T U2406 ( .I(n1955), .ZN(n1303) );
  AOI21D0BWP12T U2407 ( .A1(n1303), .A2(n1903), .B(n2740), .ZN(n1304) );
  OAI21D0BWP12T U2408 ( .A1(n1956), .A2(n1970), .B(n1304), .ZN(n1305) );
  AOI21D1BWP12T U2409 ( .A1(n2764), .A2(n1883), .B(n1305), .ZN(n1307) );
  AOI22D0BWP12T U2410 ( .A1(n3082), .A2(n1589), .B1(n2031), .B2(n3091), .ZN(
        n1306) );
  IOA21D1BWP12T U2411 ( .A1(n1674), .A2(n382), .B(n1306), .ZN(n1322) );
  AOI211D0BWP12T U2412 ( .A1(n2740), .A2(n1308), .B(n1307), .C(n2383), .ZN(
        n1309) );
  NR2XD0BWP12T U2413 ( .A1(n1309), .A2(n1976), .ZN(n1888) );
  INVD1BWP12T U2414 ( .I(n1364), .ZN(n1848) );
  AOI22D0BWP12T U2415 ( .A1(n3096), .A2(n1847), .B1(n1793), .B2(n3093), .ZN(
        n1320) );
  INVD1BWP12T U2416 ( .I(n2283), .ZN(n1311) );
  MUX2NXD0BWP12T U2417 ( .I0(n1311), .I1(n2737), .S(n2764), .ZN(n1312) );
  NR2D1BWP12T U2418 ( .A1(n1312), .A2(n2393), .ZN(n2313) );
  ND2D1BWP12T U2419 ( .A1(n2396), .A2(n3080), .ZN(n3065) );
  TPNR2D0BWP12T U2420 ( .A1(n2391), .A2(n3065), .ZN(n1318) );
  OAI21D0BWP12T U2421 ( .A1(a[12]), .A2(n3099), .B(n3103), .ZN(n1316) );
  MUX2ND0BWP12T U2422 ( .I0(n3102), .I1(n3101), .S(n2452), .ZN(n1313) );
  CKND2D0BWP12T U2423 ( .A1(n1313), .A2(n3103), .ZN(n1314) );
  MUX2NXD0BWP12T U2424 ( .I0(n1314), .I1(n3105), .S(n2193), .ZN(n1315) );
  IOA21D1BWP12T U2425 ( .A1(n2452), .A2(n1316), .B(n1315), .ZN(n1317) );
  AOI211XD0BWP12T U2426 ( .A1(n3067), .A2(n2313), .B(n1318), .C(n1317), .ZN(
        n1319) );
  OAI211D1BWP12T U2427 ( .A1(n1888), .A2(n3071), .B(n1320), .C(n1319), .ZN(
        n1321) );
  AOI211D1BWP12T U2428 ( .A1(n3076), .A2(n1405), .B(n1322), .C(n1321), .ZN(
        n1323) );
  IOA21D1BWP12T U2429 ( .A1(n1523), .A2(n3117), .B(n1323), .ZN(result[12]) );
  BUFFXD0BWP12T U2430 ( .I(result[31]), .Z(n) );
  INVD1BWP12T U2431 ( .I(n1324), .ZN(n1526) );
  ND2D1BWP12T U2432 ( .A1(n1525), .A2(n1325), .ZN(n1326) );
  XNR2D1BWP12T U2433 ( .A1(n1526), .A2(n1326), .ZN(n1537) );
  MUX2D1BWP12T U2434 ( .I0(n1896), .I1(n1897), .S(n2353), .Z(n1329) );
  AOI21D0BWP12T U2435 ( .A1(n1329), .A2(n2377), .B(n2316), .ZN(n1331) );
  OAI22D1BWP12T U2436 ( .A1(n1990), .A2(n2029), .B1(n1987), .B2(n1970), .ZN(
        n1330) );
  NR2D1BWP12T U2437 ( .A1(n1331), .A2(n1330), .ZN(n1341) );
  MUX2ND0BWP12T U2438 ( .I0(n1332), .I1(n2216), .S(n2353), .ZN(n1898) );
  TPAOI21D0BWP12T U2439 ( .A1(n1898), .A2(n2263), .B(n1968), .ZN(n1899) );
  INVD1BWP12T U2440 ( .I(n1899), .ZN(n3000) );
  NR2D0BWP12T U2441 ( .A1(n3000), .A2(n2377), .ZN(n1333) );
  OAI31D0BWP12T U2442 ( .A1(n2383), .A2(n1341), .A3(n1333), .B(n1991), .ZN(
        n1993) );
  INVD1BWP12T U2443 ( .I(n2273), .ZN(n2097) );
  CKND0BWP12T U2444 ( .I(n2101), .ZN(n1335) );
  OAI22D1BWP12T U2445 ( .A1(n1335), .A2(n1334), .B1(n2047), .B2(n2271), .ZN(
        n1337) );
  NR2D1BWP12T U2446 ( .A1(n2095), .A2(n2272), .ZN(n1336) );
  AOI211D1BWP12T U2447 ( .A1(n2097), .A2(n2103), .B(n1337), .C(n1336), .ZN(
        n2985) );
  INVD1BWP12T U2448 ( .I(n2267), .ZN(n2091) );
  OAI22D0BWP12T U2449 ( .A1(n2046), .A2(n2274), .B1(n2047), .B2(n2265), .ZN(
        n1339) );
  TPNR2D0BWP12T U2450 ( .A1(n2095), .A2(n2266), .ZN(n1338) );
  AOI211D1BWP12T U2451 ( .A1(n2091), .A2(n2103), .B(n1339), .C(n1338), .ZN(
        n2055) );
  MUX2NXD0BWP12T U2452 ( .I0(n2985), .I1(n2055), .S(n2134), .ZN(n1342) );
  AOI21D0BWP12T U2453 ( .A1(n2077), .A2(n1903), .B(n2377), .ZN(n1340) );
  NR2D1BWP12T U2454 ( .A1(n1341), .A2(n1340), .ZN(n2380) );
  TPAOI21D0BWP12T U2455 ( .A1(n2892), .A2(n1342), .B(n2380), .ZN(n2017) );
  CKND2D1BWP12T U2456 ( .A1(n1344), .A2(n1343), .ZN(n1345) );
  XNR2XD0BWP12T U2457 ( .A1(n1346), .A2(n1345), .ZN(n1440) );
  CKND2D0BWP12T U2458 ( .A1(n1360), .A2(n1359), .ZN(n1347) );
  XNR2XD0BWP12T U2459 ( .A1(n1348), .A2(n1347), .ZN(n1792) );
  AOI22D0BWP12T U2460 ( .A1(n896), .A2(n2267), .B1(n2266), .B2(n2320), .ZN(
        n1350) );
  AOI22D0BWP12T U2461 ( .A1(n2323), .A2(n2274), .B1(n2265), .B2(n2324), .ZN(
        n1349) );
  ND2D1BWP12T U2462 ( .A1(n1350), .A2(n1349), .ZN(n2262) );
  OAI22D0BWP12T U2463 ( .A1(n2097), .A2(n1352), .B1(n1351), .B2(n2228), .ZN(
        n1355) );
  NR2D0BWP12T U2464 ( .A1(n2098), .A2(n1353), .ZN(n1354) );
  AOI211D1BWP12T U2465 ( .A1(n1356), .A2(n2353), .B(n1355), .C(n1354), .ZN(
        n2793) );
  INVD0BWP12T U2466 ( .I(n2793), .ZN(n1357) );
  MUX2NXD0BWP12T U2467 ( .I0(n2262), .I1(n1357), .S(n2764), .ZN(n1358) );
  CKND2D1BWP12T U2468 ( .A1(n1358), .A2(n2402), .ZN(n2339) );
  ND2XD0BWP12T U2469 ( .A1(n1360), .A2(n1359), .ZN(n1361) );
  XNR2XD0BWP12T U2470 ( .A1(n1362), .A2(n1361), .ZN(n1636) );
  CKND2D0BWP12T U2471 ( .A1(n1636), .A2(n3082), .ZN(n1371) );
  XNR2XD0BWP12T U2472 ( .A1(n1851), .A2(a[14]), .ZN(n1853) );
  MUX2ND0BWP12T U2473 ( .I0(n3019), .I1(n3018), .S(b[14]), .ZN(n1365) );
  NR2D0BWP12T U2474 ( .A1(n1365), .A2(n3020), .ZN(n1366) );
  MUX2NXD0BWP12T U2475 ( .I0(n1366), .I1(n3023), .S(n2192), .ZN(n1369) );
  NR2D0BWP12T U2476 ( .A1(a[14]), .A2(n3099), .ZN(n1367) );
  OA21D0BWP12T U2477 ( .A1(n1367), .A2(n3020), .B(b[14]), .Z(n1368) );
  AOI211D1BWP12T U2478 ( .A1(n1853), .A2(n3096), .B(n1369), .C(n1368), .ZN(
        n1370) );
  OAI211D1BWP12T U2479 ( .A1(n2928), .A2(n2339), .B(n1371), .C(n1370), .ZN(
        n1372) );
  AOI211D1BWP12T U2480 ( .A1(n3084), .A2(n1993), .B(n1373), .C(n1372), .ZN(
        n1374) );
  IOA21D1BWP12T U2481 ( .A1(n382), .A2(n1675), .B(n1374), .ZN(n1375) );
  AO21D2BWP12T U2482 ( .A1(n1537), .A2(n3117), .B(n1375), .Z(result[14]) );
  FA1D0BWP12T U2483 ( .A(n2498), .B(n1377), .CI(n1376), .CO(n1456), .S(n2443)
         );
  FA1D1BWP12T U2484 ( .A(n1379), .B(n2571), .CI(n1378), .CO(n1451), .S(n2588)
         );
  FA1D2BWP12T U2485 ( .A(n1720), .B(a[22]), .CI(n1380), .CO(n1378), .S(n3049)
         );
  ND2D0BWP12T U2486 ( .A1(n1382), .A2(n1381), .ZN(n1383) );
  XNR2XD0BWP12T U2487 ( .A1(n1384), .A2(n1383), .ZN(n2970) );
  INVD0BWP12T U2488 ( .I(n1385), .ZN(n1387) );
  ND2XD0BWP12T U2489 ( .A1(n1387), .A2(n1386), .ZN(n1388) );
  XOR2XD0BWP12T U2490 ( .A1(n1389), .A2(n1388), .Z(n2640) );
  ND2XD0BWP12T U2491 ( .A1(n1391), .A2(n1390), .ZN(n1392) );
  XNR2XD0BWP12T U2492 ( .A1(n1393), .A2(n1392), .ZN(n2670) );
  INVD1BWP12T U2493 ( .I(n1394), .ZN(n1397) );
  INVD0BWP12T U2494 ( .I(n1399), .ZN(n1401) );
  INVD0BWP12T U2495 ( .I(n1406), .ZN(n1408) );
  TPND2D0BWP12T U2496 ( .A1(n1408), .A2(n1407), .ZN(n1409) );
  XOR2XD0BWP12T U2497 ( .A1(n1410), .A2(n1409), .Z(n2724) );
  INVD1BWP12T U2498 ( .I(n1411), .ZN(n1414) );
  ND2XD0BWP12T U2499 ( .A1(n1690), .A2(n1429), .ZN(n1412) );
  XNR2D1BWP12T U2500 ( .A1(n1430), .A2(n1412), .ZN(n2751) );
  INVD0BWP12T U2501 ( .I(n1422), .ZN(n1424) );
  TPND2D0BWP12T U2502 ( .A1(n1663), .A2(n1442), .ZN(n1443) );
  XOR2XD0BWP12T U2503 ( .A1(n1444), .A2(n1443), .Z(n2698) );
  CKND2D1BWP12T U2504 ( .A1(n1446), .A2(n1445), .ZN(n1447) );
  XNR2XD0BWP12T U2505 ( .A1(n1448), .A2(n1447), .ZN(n2942) );
  FA1D2BWP12T U2506 ( .A(n1450), .B(n2594), .CI(n1449), .CO(n1380), .S(n2615)
         );
  FA1D0BWP12T U2507 ( .A(n1452), .B(n2541), .CI(n1451), .CO(n1140), .S(n2562)
         );
  FA1D0BWP12T U2508 ( .A(n2177), .B(a[30]), .CI(n1456), .CO(n2525), .S(n3013)
         );
  OR4D0BWP12T U2509 ( .A1(n2443), .A2(n1458), .A3(n1457), .A4(n3013), .Z(n2420) );
  CKND0BWP12T U2510 ( .I(n2524), .ZN(n1567) );
  INVD1BWP12T U2511 ( .I(n1459), .ZN(n1472) );
  CKND2D1BWP12T U2512 ( .A1(n1471), .A2(n1460), .ZN(n1461) );
  XNR2D1BWP12T U2513 ( .A1(n1472), .A2(n1461), .ZN(n2618) );
  INVD1BWP12T U2514 ( .I(n1465), .ZN(n1540) );
  ND2D1BWP12T U2515 ( .A1(n287), .A2(n1467), .ZN(n1468) );
  XOR2XD1BWP12T U2516 ( .A1(n1469), .A2(n1468), .Z(n2566) );
  AOI21D1BWP12T U2517 ( .A1(n1472), .A2(n1471), .B(n1470), .ZN(n1475) );
  CKND2D1BWP12T U2518 ( .A1(n289), .A2(n1473), .ZN(n1474) );
  XOR2XD1BWP12T U2519 ( .A1(n1475), .A2(n1474), .Z(n2947) );
  OAI21D1BWP12T U2520 ( .A1(n1532), .A2(n1478), .B(n1477), .ZN(n1483) );
  INVD1BWP12T U2521 ( .I(n1479), .ZN(n1481) );
  CKND2D1BWP12T U2522 ( .A1(n1481), .A2(n1480), .ZN(n1482) );
  XNR2XD1BWP12T U2523 ( .A1(n1483), .A2(n1482), .ZN(n2645) );
  ND2D1BWP12T U2524 ( .A1(n1484), .A2(n1530), .ZN(n1485) );
  ND2D1BWP12T U2525 ( .A1(n1487), .A2(n1486), .ZN(n1489) );
  XNR2D1BWP12T U2526 ( .A1(n1489), .A2(n1488), .ZN(n3078) );
  INVD1BWP12T U2527 ( .I(n1497), .ZN(n1521) );
  ND2D1BWP12T U2528 ( .A1(n1500), .A2(n1499), .ZN(n1502) );
  XNR2D1BWP12T U2529 ( .A1(n1502), .A2(n1501), .ZN(n2806) );
  INVD1BWP12T U2530 ( .I(n1503), .ZN(n1505) );
  ND2D1BWP12T U2531 ( .A1(n1505), .A2(n1504), .ZN(n1507) );
  XOR2XD1BWP12T U2532 ( .A1(n1507), .A2(n1506), .Z(n2777) );
  OR4D1BWP12T U2533 ( .A1(n1516), .A2(n1515), .A3(n2975), .A4(n1514), .Z(n1518) );
  OR4D1BWP12T U2534 ( .A1(n2749), .A2(n2776), .A3(n1518), .A4(n1517), .Z(n1522) );
  AOI21D1BWP12T U2535 ( .A1(n1526), .A2(n1525), .B(n1524), .ZN(n1529) );
  ND2D1BWP12T U2536 ( .A1(n293), .A2(n1527), .ZN(n1528) );
  OAI21D1BWP12T U2537 ( .A1(n1532), .A2(n1531), .B(n1530), .ZN(n1536) );
  ND2D1BWP12T U2538 ( .A1(n1534), .A2(n1533), .ZN(n1535) );
  XNR2XD4BWP12T U2539 ( .A1(n1536), .A2(n1535), .ZN(n2675) );
  ND2D1BWP12T U2540 ( .A1(n1539), .A2(n1538), .ZN(n1541) );
  XNR2D1BWP12T U2541 ( .A1(n1541), .A2(n1540), .ZN(n3051) );
  INVD1BWP12T U2542 ( .I(n1542), .ZN(n1544) );
  ND2D1BWP12T U2543 ( .A1(n1544), .A2(n1543), .ZN(n1545) );
  FA1D1BWP12T U2544 ( .A(mult_x_18_n425), .B(mult_x_18_n405), .CI(n1548), .CO(
        n2447), .S(n3015) );
  CKND1BWP12T U2545 ( .I(n1549), .ZN(n1550) );
  NR2D1BWP12T U2546 ( .A1(n1550), .A2(n1553), .ZN(n1556) );
  INVD1BWP12T U2547 ( .I(n1551), .ZN(n1554) );
  OAI21D1BWP12T U2548 ( .A1(n1554), .A2(n1553), .B(n1552), .ZN(n1555) );
  AOI21D1BWP12T U2549 ( .A1(n1557), .A2(n1556), .B(n1555), .ZN(n1562) );
  INVD1BWP12T U2550 ( .I(n1558), .ZN(n1560) );
  ND2D1BWP12T U2551 ( .A1(n1560), .A2(n1559), .ZN(n1561) );
  XOR2D1BWP12T U2552 ( .A1(n1562), .A2(n1561), .Z(n2422) );
  NR4D0BWP12T U2553 ( .A1(n1564), .A2(n3015), .A3(n1563), .A4(n2422), .ZN(
        n1565) );
  IND4D1BWP12T U2554 ( .A1(n1568), .B1(n1567), .B2(n1566), .B3(n1565), .ZN(
        n2419) );
  FA1D0BWP12T U2555 ( .A(n2498), .B(b[29]), .CI(n1570), .CO(n1569), .S(n2423)
         );
  FA1D1BWP12T U2556 ( .A(b[22]), .B(a[22]), .CI(n1572), .CO(n1571), .S(n3043)
         );
  CKND2D0BWP12T U2557 ( .A1(n1795), .A2(n1794), .ZN(n1573) );
  XNR2XD0BWP12T U2558 ( .A1(n1574), .A2(n1573), .ZN(n2948) );
  INVD1BWP12T U2559 ( .I(n1575), .ZN(n1731) );
  CKND2D0BWP12T U2560 ( .A1(n1731), .A2(n1730), .ZN(n1576) );
  XOR2XD0BWP12T U2561 ( .A1(n1577), .A2(n1576), .Z(n2619) );
  CKND2D0BWP12T U2562 ( .A1(n1735), .A2(n1734), .ZN(n1578) );
  XNR2XD0BWP12T U2563 ( .A1(n1579), .A2(n1578), .ZN(n2646) );
  INVD1BWP12T U2564 ( .I(n1580), .ZN(n1583) );
  INVD1BWP12T U2565 ( .I(n1590), .ZN(n1739) );
  CKND2D0BWP12T U2566 ( .A1(n1739), .A2(n1738), .ZN(n1591) );
  XOR2XD0BWP12T U2567 ( .A1(n1592), .A2(n1591), .Z(n2676) );
  CKND2D1BWP12T U2568 ( .A1(n1593), .A2(n1595), .ZN(n1598) );
  AOI21D1BWP12T U2569 ( .A1(n1596), .A2(n1595), .B(n1594), .ZN(n1597) );
  OAI21D1BWP12T U2570 ( .A1(n1607), .A2(n1598), .B(n1597), .ZN(n1602) );
  ND2D1BWP12T U2571 ( .A1(n1600), .A2(n1599), .ZN(n1601) );
  XNR2XD1BWP12T U2572 ( .A1(n1602), .A2(n1601), .ZN(n3053) );
  INVD1BWP12T U2573 ( .I(n1603), .ZN(n1783) );
  TPND2D0BWP12T U2574 ( .A1(n1783), .A2(n1782), .ZN(n1604) );
  XOR2XD0BWP12T U2575 ( .A1(n1605), .A2(n1604), .Z(n2705) );
  INVD1BWP12T U2576 ( .I(n1606), .ZN(n1629) );
  INVD1BWP12T U2577 ( .I(n1608), .ZN(n1614) );
  INVD1BWP12T U2578 ( .I(n3082), .ZN(n2967) );
  CKND2D1BWP12T U2579 ( .A1(n1614), .A2(n1613), .ZN(n1615) );
  XNR2D1BWP12T U2580 ( .A1(n1624), .A2(n1615), .ZN(n2754) );
  CKND0BWP12T U2581 ( .I(n1616), .ZN(n1617) );
  NR2D1BWP12T U2582 ( .A1(n1617), .A2(n1620), .ZN(n1623) );
  CKND0BWP12T U2583 ( .I(n1618), .ZN(n1621) );
  OAI21D1BWP12T U2584 ( .A1(n1621), .A2(n1620), .B(n1619), .ZN(n1622) );
  AOI21D1BWP12T U2585 ( .A1(n1624), .A2(n1623), .B(n1622), .ZN(n1626) );
  INVD1BWP12T U2586 ( .I(n1759), .ZN(n1753) );
  ND2XD0BWP12T U2587 ( .A1(n1753), .A2(n1758), .ZN(n1625) );
  XOR2XD1BWP12T U2588 ( .A1(n1626), .A2(n1625), .Z(n2781) );
  INVD1BWP12T U2589 ( .I(n1627), .ZN(n1628) );
  AOI21D1BWP12T U2590 ( .A1(n1630), .A2(n1629), .B(n1628), .ZN(n1635) );
  INVD0BWP12T U2591 ( .I(n1631), .ZN(n1633) );
  CKND2D1BWP12T U2592 ( .A1(n1633), .A2(n1632), .ZN(n1634) );
  XOR2XD1BWP12T U2593 ( .A1(n1635), .A2(n1634), .Z(n2837) );
  CKND2D0BWP12T U2594 ( .A1(n1743), .A2(n1742), .ZN(n1637) );
  FA1D2BWP12T U2595 ( .A(n2594), .B(b[21]), .CI(n1639), .CO(n1572), .S(n2610)
         );
  INVD1BWP12T U2596 ( .I(n1645), .ZN(n2416) );
  FA1D2BWP12T U2597 ( .A(n2177), .B(a[30]), .CI(n1646), .CO(n2527), .S(n2984)
         );
  FA1D2BWP12T U2598 ( .A(n1452), .B(n2541), .CI(n1648), .CO(n1142), .S(n2561)
         );
  FA1D0BWP12T U2599 ( .A(n1379), .B(n2571), .CI(n1649), .CO(n1648), .S(n2587)
         );
  CKND2D1BWP12T U2600 ( .A1(n1654), .A2(n1653), .ZN(n1655) );
  XNR2XD0BWP12T U2601 ( .A1(n1656), .A2(n1655), .ZN(n2971) );
  CKND2D1BWP12T U2602 ( .A1(n1658), .A2(n1657), .ZN(n1659) );
  XNR2XD0BWP12T U2603 ( .A1(n1660), .A2(n1659), .ZN(n2671) );
  INVD1BWP12T U2604 ( .I(n1661), .ZN(n1663) );
  CKND2D1BWP12T U2605 ( .A1(n1663), .A2(n1662), .ZN(n1664) );
  XOR2XD0BWP12T U2606 ( .A1(n1665), .A2(n1664), .Z(n2699) );
  CKND2D1BWP12T U2607 ( .A1(n1667), .A2(n1666), .ZN(n1668) );
  XNR2XD0BWP12T U2608 ( .A1(n1669), .A2(n1668), .ZN(n2943) );
  INVD1BWP12T U2609 ( .I(n1679), .ZN(n1681) );
  INVD0BWP12T U2610 ( .I(n1688), .ZN(n1690) );
  ND2D1BWP12T U2611 ( .A1(n1701), .A2(n1700), .ZN(n1702) );
  CKND2D1BWP12T U2612 ( .A1(n1387), .A2(n1716), .ZN(n1717) );
  XOR2XD0BWP12T U2613 ( .A1(n1718), .A2(n1717), .Z(n2641) );
  FA1D0BWP12T U2614 ( .A(n1720), .B(a[22]), .CI(n1719), .CO(n1649), .S(n3016)
         );
  FA1D2BWP12T U2615 ( .A(b[30]), .B(a[30]), .CI(n1726), .CO(n2976), .S(n3007)
         );
  FA1D2BWP12T U2616 ( .A(b[24]), .B(n2541), .CI(n1727), .CO(n1143), .S(n2539)
         );
  FA1D0BWP12T U2617 ( .A(b[22]), .B(a[22]), .CI(n1728), .CO(n1798), .S(n3042)
         );
  FA1D0BWP12T U2618 ( .A(n2594), .B(b[21]), .CI(n1729), .CO(n1728), .S(n2609)
         );
  ND2XD0BWP12T U2619 ( .A1(n1731), .A2(n1730), .ZN(n1732) );
  XOR2XD0BWP12T U2620 ( .A1(n1733), .A2(n1732), .Z(n2620) );
  ND2XD0BWP12T U2621 ( .A1(n1735), .A2(n1734), .ZN(n1736) );
  XNR2XD0BWP12T U2622 ( .A1(n1737), .A2(n1736), .ZN(n2647) );
  TPND2D0BWP12T U2623 ( .A1(n1739), .A2(n1738), .ZN(n1740) );
  XOR2XD0BWP12T U2624 ( .A1(n1741), .A2(n1740), .Z(n2677) );
  TPND2D0BWP12T U2625 ( .A1(n1743), .A2(n1742), .ZN(n1744) );
  XNR2XD0BWP12T U2626 ( .A1(n1745), .A2(n1744), .ZN(n2914) );
  OAI21D1BWP12T U2627 ( .A1(n1748), .A2(n1747), .B(n1746), .ZN(n1752) );
  CKND2D1BWP12T U2628 ( .A1(n1614), .A2(n1750), .ZN(n1751) );
  XNR2D1BWP12T U2629 ( .A1(n1752), .A2(n1751), .ZN(n2758) );
  AOI21D1BWP12T U2630 ( .A1(n1768), .A2(n1756), .B(n1757), .ZN(n1755) );
  ND2XD0BWP12T U2631 ( .A1(n1753), .A2(n1758), .ZN(n1754) );
  XOR2XD1BWP12T U2632 ( .A1(n1755), .A2(n1754), .Z(n2780) );
  INVD1BWP12T U2633 ( .I(n1775), .ZN(n1778) );
  TPND2D0BWP12T U2634 ( .A1(n1783), .A2(n1782), .ZN(n1784) );
  XOR2XD0BWP12T U2635 ( .A1(n1785), .A2(n1784), .Z(n2704) );
  CKND2D0BWP12T U2636 ( .A1(n1795), .A2(n1794), .ZN(n1796) );
  XNR2XD0BWP12T U2637 ( .A1(n1797), .A2(n1796), .ZN(n2949) );
  OR4D1BWP12T U2638 ( .A1(n3042), .A2(n2609), .A3(n1799), .A4(n2568), .Z(n1801) );
  OR4D1BWP12T U2639 ( .A1(n1802), .A2(n2539), .A3(n1801), .A4(n1800), .Z(n1804) );
  FA1D2BWP12T U2640 ( .A(n2498), .B(b[29]), .CI(n1803), .CO(n1726), .S(n2424)
         );
  OR4D1BWP12T U2641 ( .A1(n1806), .A2(n1805), .A3(n1804), .A4(n2424), .Z(n2413) );
  NR4D0BWP12T U2642 ( .A1(n2979), .A2(a[26]), .A3(n2358), .A4(n2541), .ZN(
        n1810) );
  NR4D0BWP12T U2643 ( .A1(n2498), .A2(a[28]), .A3(n2460), .A4(n3100), .ZN(
        n1809) );
  NR4D0BWP12T U2644 ( .A1(a[14]), .A2(n2870), .A3(n2846), .A4(n2898), .ZN(
        n1808) );
  NR4D0BWP12T U2645 ( .A1(n2652), .A2(n2710), .A3(a[13]), .A4(a[12]), .ZN(
        n1807) );
  ND4D1BWP12T U2646 ( .A1(n1810), .A2(n1809), .A3(n1808), .A4(n1807), .ZN(
        n1868) );
  NR2D0BWP12T U2647 ( .A1(n1811), .A2(a[30]), .ZN(n2251) );
  NR4D0BWP12T U2648 ( .A1(n2594), .A2(a[20]), .A3(n2621), .A4(a[22]), .ZN(
        n1815) );
  NR4D0BWP12T U2649 ( .A1(n2466), .A2(n2738), .A3(a[3]), .A4(n2349), .ZN(n1812) );
  AN4XD1BWP12T U2650 ( .A1(n2574), .A2(n1832), .A3(n3020), .A4(n1812), .Z(
        n1814) );
  NR4D0BWP12T U2651 ( .A1(n2679), .A2(n2915), .A3(n2785), .A4(n2815), .ZN(
        n1813) );
  ND4D0BWP12T U2652 ( .A1(n2251), .A2(n1815), .A3(n1814), .A4(n1813), .ZN(
        n1867) );
  HA1D0BWP12T U2653 ( .A(n2996), .B(n1816), .CO(n2532), .S(n2989) );
  HA1D1BWP12T U2654 ( .A(n1820), .B(n1819), .CO(n1818), .S(n2582) );
  HA1D0BWP12T U2655 ( .A(n3022), .B(n1821), .CO(n1819), .S(n3017) );
  INVD1BWP12T U2656 ( .I(n1822), .ZN(n1842) );
  NR2XD0BWP12T U2657 ( .A1(n1842), .A2(n2915), .ZN(n1823) );
  XNR2XD1BWP12T U2658 ( .A1(n1823), .A2(n2679), .ZN(n2693) );
  CKND0BWP12T U2659 ( .I(n1824), .ZN(n1825) );
  NR2D1BWP12T U2660 ( .A1(n1842), .A2(n1825), .ZN(n1826) );
  XNR2XD0BWP12T U2661 ( .A1(n1826), .A2(n2652), .ZN(n2665) );
  NR2XD0BWP12T U2662 ( .A1(n1842), .A2(n1827), .ZN(n1828) );
  XNR2XD1BWP12T U2663 ( .A1(n1828), .A2(n2621), .ZN(n2635) );
  HA1D0BWP12T U2664 ( .A(n1830), .B(n1829), .CO(n1821), .S(n2593) );
  NR4D0BWP12T U2665 ( .A1(n2693), .A2(n2665), .A3(n2635), .A4(n2593), .ZN(
        n1858) );
  HICIND1BWP12T U2666 ( .A(n2952), .CIN(n1831), .CO(n1829), .S(n2964) );
  CKXOR2D0BWP12T U2667 ( .A1(n1850), .A2(n2738), .Z(n2744) );
  OR4D0BWP12T U2668 ( .A1(n1836), .A2(n3040), .A3(n2753), .A4(n1835), .Z(n1837) );
  XNR2XD1BWP12T U2669 ( .A1(n1848), .A2(n2846), .ZN(n2842) );
  OR4D0BWP12T U2670 ( .A1(n2964), .A2(n2744), .A3(n1837), .A4(n2842), .Z(n1843) );
  CKND0BWP12T U2671 ( .I(n1838), .ZN(n1839) );
  NR2D0BWP12T U2672 ( .A1(n1839), .A2(a[12]), .ZN(n1840) );
  CKND2D1BWP12T U2673 ( .A1(n1840), .A2(n1848), .ZN(n1841) );
  XOR2XD1BWP12T U2674 ( .A1(n1841), .A2(a[13]), .Z(n3057) );
  CKXOR2D0BWP12T U2675 ( .A1(n1842), .A2(n2915), .Z(n2938) );
  NR3D0BWP12T U2676 ( .A1(n1843), .A2(n3057), .A3(n2938), .ZN(n1857) );
  CKND0BWP12T U2677 ( .I(n1846), .ZN(n1844) );
  CKND2D1BWP12T U2678 ( .A1(n1848), .A2(n1844), .ZN(n1845) );
  XOR2D1BWP12T U2679 ( .A1(n1845), .A2(n3100), .Z(n3095) );
  OR4D0BWP12T U2680 ( .A1(n2834), .A2(n3095), .A3(n2910), .A4(n1847), .Z(n1855) );
  OR3XD0BWP12T U2681 ( .A1(n1853), .A2(n2707), .A3(n1852), .Z(n1854) );
  NR4D0BWP12T U2682 ( .A1(n1855), .A2(n2863), .A3(n2779), .A4(n1854), .ZN(
        n1856) );
  IND4D1BWP12T U2683 ( .A1(n3017), .B1(n1858), .B2(n1857), .B3(n1856), .ZN(
        n1860) );
  OR4D1BWP12T U2684 ( .A1(n2556), .A2(n2582), .A3(n1860), .A4(n1859), .Z(n1862) );
  OR4D1BWP12T U2685 ( .A1(n1864), .A2(n1863), .A3(n1862), .A4(n1861), .Z(n1865) );
  OR4XD1BWP12T U2686 ( .A1(n2989), .A2(n2436), .A3(n1865), .A4(n2533), .Z(
        n1866) );
  OAI31D0BWP12T U2687 ( .A1(n1868), .A2(n2383), .A3(n1867), .B(n1866), .ZN(
        n2410) );
  CKND0BWP12T U2688 ( .I(n1869), .ZN(n1870) );
  CKND2D1BWP12T U2689 ( .A1(n2396), .A2(n2258), .ZN(n2289) );
  AOI21D0BWP12T U2690 ( .A1(n1870), .A2(n2740), .B(n2289), .ZN(n1871) );
  TPNR2D0BWP12T U2691 ( .A1(n1871), .A2(n1968), .ZN(n1875) );
  OAI22D0BWP12T U2692 ( .A1(n1973), .A2(n1986), .B1(n1974), .B2(n1970), .ZN(
        n1873) );
  OAI21D0BWP12T U2693 ( .A1(n1971), .A2(n1989), .B(n2377), .ZN(n1872) );
  AOI211D1BWP12T U2694 ( .A1(n1903), .A2(n1874), .B(n1873), .C(n1872), .ZN(
        n2381) );
  TPOAI21D0BWP12T U2695 ( .A1(n1875), .A2(n2381), .B(n1991), .ZN(n2866) );
  INVD1BWP12T U2696 ( .I(n1876), .ZN(n2542) );
  CKND2D0BWP12T U2697 ( .A1(n1877), .A2(n2263), .ZN(n1967) );
  AOI21D0BWP12T U2698 ( .A1(n2542), .A2(n1967), .B(n1878), .ZN(n2425) );
  AOI21D0BWP12T U2699 ( .A1(n1901), .A2(n1879), .B(n1878), .ZN(n1882) );
  OAI22D1BWP12T U2700 ( .A1(n1920), .A2(n2202), .B1(n1919), .B2(n2544), .ZN(
        n1880) );
  NR2D1BWP12T U2701 ( .A1(n1881), .A2(n1880), .ZN(n1934) );
  MUX2ND0BWP12T U2702 ( .I0(n1934), .I1(n1894), .S(n2353), .ZN(n1963) );
  CKND2D1BWP12T U2703 ( .A1(n1963), .A2(n2314), .ZN(n2072) );
  TPOAI21D0BWP12T U2704 ( .A1(n2549), .A2(n2072), .B(n2542), .ZN(n2570) );
  NR4D0BWP12T U2705 ( .A1(n2866), .A2(n2425), .A3(n1882), .A4(n2570), .ZN(
        n1889) );
  OAI211D0BWP12T U2706 ( .A1(n2207), .A2(n2073), .B(n2960), .C(n2740), .ZN(
        n1885) );
  TPAOI31D0BWP12T U2707 ( .A1(n1885), .A2(n2396), .A3(n2015), .B(n1976), .ZN(
        n2747) );
  AOI21D0BWP12T U2708 ( .A1(n2207), .A2(n1908), .B(n2542), .ZN(n1887) );
  INVD1BWP12T U2709 ( .I(n2960), .ZN(n2392) );
  OAI21D1BWP12T U2710 ( .A1(n1887), .A2(n2392), .B(n1886), .ZN(n2961) );
  ND4D0BWP12T U2711 ( .A1(n1889), .A2(n2747), .A3(n1888), .A4(n2961), .ZN(
        n1911) );
  OAI22D1BWP12T U2712 ( .A1(n2596), .A2(n1920), .B1(n1919), .B2(n2952), .ZN(
        n1890) );
  NR2D1BWP12T U2713 ( .A1(n1891), .A2(n1890), .ZN(n1947) );
  MUX2ND0BWP12T U2714 ( .I0(n1947), .I1(n1934), .S(n2353), .ZN(n1892) );
  NR2D1BWP12T U2715 ( .A1(n1892), .A2(n2764), .ZN(n2011) );
  NR2D1BWP12T U2716 ( .A1(n1986), .A2(n2979), .ZN(n1893) );
  AO211D1BWP12T U2717 ( .A1(n2076), .A2(n1894), .B(n2011), .C(n1893), .Z(n2630) );
  AN4D0BWP12T U2718 ( .A1(n2630), .A2(n1895), .A3(n2922), .A4(n2601), .Z(n1900) );
  OAI22D1BWP12T U2719 ( .A1(n1897), .A2(n1970), .B1(n1896), .B2(n2029), .ZN(
        n2075) );
  AOI21D1BWP12T U2720 ( .A1(n1898), .A2(n2764), .B(n2075), .ZN(n3032) );
  AOI31D0BWP12T U2721 ( .A1(n1900), .A2(n1899), .A3(n3032), .B(n2549), .ZN(
        n1910) );
  INVD0BWP12T U2722 ( .I(n1901), .ZN(n1902) );
  AOI21D0BWP12T U2723 ( .A1(n1902), .A2(n2396), .B(n2402), .ZN(n1907) );
  AOI21D0BWP12T U2724 ( .A1(n1985), .A2(n1903), .B(n2740), .ZN(n1904) );
  OAI21D1BWP12T U2725 ( .A1(n1990), .A2(n1970), .B(n1904), .ZN(n1905) );
  AOI21D1BWP12T U2726 ( .A1(n2764), .A2(n1906), .B(n1905), .ZN(n3112) );
  TPOAI21D0BWP12T U2727 ( .A1(n1907), .A2(n3112), .B(n1991), .ZN(n3085) );
  TPOAI21D0BWP12T U2728 ( .A1(n1909), .A2(n2549), .B(n1908), .ZN(n2661) );
  NR4D0BWP12T U2729 ( .A1(n1911), .A2(n1910), .A3(n3085), .A4(n2661), .ZN(
        n1997) );
  INVD1BWP12T U2730 ( .I(n2630), .ZN(n1912) );
  TPAOI21D0BWP12T U2731 ( .A1(n1912), .A2(n2396), .B(n2402), .ZN(n1933) );
  OAI22D1BWP12T U2732 ( .A1(n1920), .A2(n3059), .B1(n1919), .B2(n2193), .ZN(
        n1913) );
  NR2D1BWP12T U2733 ( .A1(n1914), .A2(n1913), .ZN(n1949) );
  OAI22D1BWP12T U2734 ( .A1(n1920), .A2(n2682), .B1(n1919), .B2(n2917), .ZN(
        n1915) );
  NR2D1BWP12T U2735 ( .A1(n1916), .A2(n1915), .ZN(n1948) );
  TPOAI22D0BWP12T U2736 ( .A1(n1949), .A2(n1989), .B1(n1948), .B2(n1986), .ZN(
        n1932) );
  OAI22D1BWP12T U2737 ( .A1(n1920), .A2(n2872), .B1(n1919), .B2(n2848), .ZN(
        n1921) );
  NR2D1BWP12T U2738 ( .A1(n1922), .A2(n1921), .ZN(n1950) );
  OAI21D0BWP12T U2739 ( .A1(n1950), .A2(n1970), .B(n2377), .ZN(n1931) );
  AOI22D1BWP12T U2740 ( .A1(n2466), .A2(n1924), .B1(n1923), .B2(n2785), .ZN(
        n1929) );
  CKND2D0BWP12T U2741 ( .A1(n1925), .A2(n2738), .ZN(n1928) );
  ND2D1BWP12T U2742 ( .A1(n1926), .A2(a[3]), .ZN(n1927) );
  TPAOI31D0BWP12T U2743 ( .A1(n1929), .A2(n1928), .A3(n1927), .B(n2764), .ZN(
        n1930) );
  NR3D1BWP12T U2744 ( .A1(n1932), .A2(n1931), .A3(n1930), .ZN(n2018) );
  OAI21D1BWP12T U2745 ( .A1(n1933), .A2(n2018), .B(n1991), .ZN(n2771) );
  CKND0BWP12T U2746 ( .I(n1948), .ZN(n1937) );
  OAI22D0BWP12T U2747 ( .A1(n1934), .A2(n1986), .B1(n1947), .B2(n1989), .ZN(
        n1936) );
  OAI21D0BWP12T U2748 ( .A1(n1949), .A2(n2029), .B(n2377), .ZN(n1935) );
  AO211D1BWP12T U2749 ( .A1(n1984), .A2(n1937), .B(n1936), .C(n1935), .Z(n2019) );
  CKND0BWP12T U2750 ( .I(n1938), .ZN(n1939) );
  OAI21D1BWP12T U2751 ( .A1(n1939), .A2(n2383), .B(n2393), .ZN(n1940) );
  RCAOI21D0BWP12T U2752 ( .A1(n2019), .A2(n1940), .B(n1976), .ZN(n2908) );
  OAI22D1BWP12T U2753 ( .A1(n1941), .A2(n2029), .B1(n2080), .B2(n1970), .ZN(
        n2550) );
  CKND2D0BWP12T U2754 ( .A1(n1942), .A2(n3084), .ZN(n1943) );
  AOI211D0BWP12T U2755 ( .A1(n1945), .A2(n2550), .B(n1944), .C(n1943), .ZN(
        n1962) );
  OAI21D0BWP12T U2756 ( .A1(n1963), .A2(n2377), .B(n2258), .ZN(n1946) );
  CKND2D0BWP12T U2757 ( .A1(n1946), .A2(n2073), .ZN(n1951) );
  MUX2D1BWP12T U2758 ( .I0(n1948), .I1(n1947), .S(n2353), .Z(n1964) );
  TPAOI31D0BWP12T U2759 ( .A1(n1951), .A2(n2396), .A3(n2810), .B(n1976), .ZN(
        n2813) );
  CKND0BWP12T U2760 ( .I(n1952), .ZN(n1954) );
  OAI22D0BWP12T U2761 ( .A1(n1954), .A2(n2029), .B1(n1953), .B2(n1986), .ZN(
        n1959) );
  OAI21D0BWP12T U2762 ( .A1(n1955), .A2(n1970), .B(n2377), .ZN(n1958) );
  NR2D0BWP12T U2763 ( .A1(n1956), .A2(n1989), .ZN(n1957) );
  NR3D1BWP12T U2764 ( .A1(n1959), .A2(n1958), .A3(n1957), .ZN(n1960) );
  INVD1BWP12T U2765 ( .I(n1960), .ZN(n2118) );
  CKND2D0BWP12T U2766 ( .A1(n2550), .A2(n2396), .ZN(n1961) );
  AOI21D1BWP12T U2767 ( .A1(n2393), .A2(n1961), .B(n1960), .ZN(n2388) );
  AOI211D1BWP12T U2768 ( .A1(n1968), .A2(n2118), .B(n2388), .C(n1976), .ZN(
        n2844) );
  ND4D0BWP12T U2769 ( .A1(n2908), .A2(n1962), .A3(n2813), .A4(n2844), .ZN(
        n1982) );
  CKND0BWP12T U2770 ( .I(n1963), .ZN(n1965) );
  OAI22D1BWP12T U2771 ( .A1(n1965), .A2(n2287), .B1(n1964), .B2(n2327), .ZN(
        n2709) );
  AOI21D0BWP12T U2772 ( .A1(n2709), .A2(n2396), .B(n1966), .ZN(n2721) );
  CKND0BWP12T U2773 ( .I(n1967), .ZN(n1969) );
  OAI21D0BWP12T U2774 ( .A1(n1969), .A2(n1968), .B(n2396), .ZN(n1975) );
  AOI21D1BWP12T U2775 ( .A1(n1975), .A2(n2393), .B(n2028), .ZN(n1977) );
  NR2XD0BWP12T U2776 ( .A1(n1977), .A2(n1976), .ZN(n3072) );
  ND4D0BWP12T U2777 ( .A1(n1979), .A2(n2721), .A3(n1978), .A4(n3072), .ZN(
        n1980) );
  NR4D0BWP12T U2778 ( .A1(n2771), .A2(n1982), .A3(n1981), .A4(n1980), .ZN(
        n1996) );
  CKND0BWP12T U2779 ( .I(n3032), .ZN(n1983) );
  AOI21D0BWP12T U2780 ( .A1(n1983), .A2(n2396), .B(n2402), .ZN(n1992) );
  TPOAI21D0BWP12T U2781 ( .A1(n1992), .A2(n2797), .B(n1991), .ZN(n2801) );
  NR2D0BWP12T U2782 ( .A1(n2801), .A2(n1993), .ZN(n1994) );
  ND4D0BWP12T U2783 ( .A1(n1997), .A2(n1996), .A3(n1995), .A4(n1994), .ZN(
        n2009) );
  ND4D1BWP12T U2784 ( .A1(n2870), .A2(n2846), .A3(n3100), .A4(n2898), .ZN(
        n2001) );
  ND4D1BWP12T U2785 ( .A1(n2498), .A2(a[28]), .A3(n2460), .A4(n2541), .ZN(
        n2000) );
  ND4D1BWP12T U2786 ( .A1(a[3]), .A2(n2352), .A3(n2349), .A4(n2172), .ZN(n1999) );
  ND4D0BWP12T U2787 ( .A1(n2571), .A2(a[22]), .A3(n2594), .A4(a[20]), .ZN(
        n1998) );
  NR4D0BWP12T U2788 ( .A1(n2001), .A2(n2000), .A3(n1999), .A4(n1998), .ZN(
        n2007) );
  AN4XD1BWP12T U2789 ( .A1(n2358), .A2(a[26]), .A3(n2738), .A4(n2466), .Z(
        n2006) );
  CKND2D0BWP12T U2790 ( .A1(n2710), .A2(n2785), .ZN(n2003) );
  ND4D0BWP12T U2791 ( .A1(n2679), .A2(n2915), .A3(a[13]), .A4(a[12]), .ZN(
        n2002) );
  NR4D0BWP12T U2792 ( .A1(n2192), .A2(n2003), .A3(n2002), .A4(n3023), .ZN(
        n2005) );
  AN4XD1BWP12T U2793 ( .A1(n2652), .A2(n2621), .A3(a[30]), .A4(n2815), .Z(
        n2004) );
  ND4D1BWP12T U2794 ( .A1(n2007), .A2(n2006), .A3(n2005), .A4(n2004), .ZN(
        n2008) );
  MUX2ND0BWP12T U2795 ( .I0(n2009), .I1(n2008), .S(n2979), .ZN(n2409) );
  INVD1BWP12T U2796 ( .I(n2015), .ZN(n2741) );
  INVD1BWP12T U2797 ( .I(n2011), .ZN(n2012) );
  OAI21D1BWP12T U2798 ( .A1(n2013), .A2(n2314), .B(n2012), .ZN(n2631) );
  CKND2D0BWP12T U2799 ( .A1(n2960), .A2(n2600), .ZN(n2399) );
  INVD1BWP12T U2800 ( .I(n2144), .ZN(n2823) );
  OAI22D1BWP12T U2801 ( .A1(n2823), .A2(n2121), .B1(n2140), .B2(n2123), .ZN(
        n2706) );
  AOI22D1BWP12T U2802 ( .A1(n2015), .A2(n2392), .B1(n2933), .B2(n2014), .ZN(
        n2734) );
  AO21D1BWP12T U2803 ( .A1(n2631), .A2(n2740), .B(n2018), .Z(n2774) );
  OAI21D1BWP12T U2804 ( .A1(n2020), .A2(n2377), .B(n2019), .ZN(n2895) );
  TPND2D0BWP12T U2805 ( .A1(n2107), .A2(n2021), .ZN(n2027) );
  AOI22D0BWP12T U2806 ( .A1(n2109), .A2(n2023), .B1(n2108), .B2(n2022), .ZN(
        n2026) );
  TPND2D0BWP12T U2807 ( .A1(n2110), .A2(n2024), .ZN(n2025) );
  ND3D1BWP12T U2808 ( .A1(n2027), .A2(n2026), .A3(n2025), .ZN(n2133) );
  MUX2ND0BWP12T U2809 ( .I0(n2133), .I1(n2083), .S(n2139), .ZN(n2030) );
  OAI21D1BWP12T U2810 ( .A1(n2030), .A2(n2130), .B(n3064), .ZN(n3052) );
  NR2D0BWP12T U2811 ( .A1(n2397), .A2(n2377), .ZN(n2032) );
  OAI22D1BWP12T U2812 ( .A1(n2033), .A2(n2130), .B1(n2381), .B2(n2032), .ZN(
        n2883) );
  AOI21D0BWP12T U2813 ( .A1(n2086), .A2(n2377), .B(n2316), .ZN(n2039) );
  AOI22D0BWP12T U2814 ( .A1(n2933), .A2(n2035), .B1(n2034), .B2(n2139), .ZN(
        n2036) );
  NR2D1BWP12T U2815 ( .A1(n2988), .A2(n2114), .ZN(n2142) );
  OAI211D0BWP12T U2816 ( .A1(n2037), .A2(n2892), .B(n2036), .C(n2142), .ZN(
        n2038) );
  OAI21D1BWP12T U2817 ( .A1(n2040), .A2(n2039), .B(n2038), .ZN(n2648) );
  INVD1BWP12T U2818 ( .I(n2325), .ZN(n2045) );
  TPOAI22D0BWP12T U2819 ( .A1(n2047), .A2(n2321), .B1(n2046), .B2(n2268), .ZN(
        n2044) );
  TPNR2D0BWP12T U2820 ( .A1(n2095), .A2(n2322), .ZN(n2043) );
  AOI211D1BWP12T U2821 ( .A1(n2045), .A2(n2103), .B(n2044), .C(n2043), .ZN(
        n2054) );
  OAI22D0BWP12T U2822 ( .A1(n2047), .A2(n2247), .B1(n2046), .B2(n2326), .ZN(
        n2049) );
  NR2D0BWP12T U2823 ( .A1(n2095), .A2(n2246), .ZN(n2048) );
  AOI211D1BWP12T U2824 ( .A1(n2103), .A2(n2498), .B(n2049), .C(n2048), .ZN(
        n2050) );
  OAI222D1BWP12T U2825 ( .A1(n2121), .A2(n2054), .B1(n2119), .B2(n2055), .C1(
        n2123), .C2(n2050), .ZN(n2986) );
  OAI222D1BWP12T U2826 ( .A1(n2119), .A2(n2985), .B1(n2121), .B2(n2055), .C1(
        n2123), .C2(n2054), .ZN(n3036) );
  AOI22D0BWP12T U2827 ( .A1(n2109), .A2(n2224), .B1(n2108), .B2(n2056), .ZN(
        n2058) );
  CKND2D0BWP12T U2828 ( .A1(n2110), .A2(n2223), .ZN(n2057) );
  CKND2D1BWP12T U2829 ( .A1(n2058), .A2(n2057), .ZN(n2061) );
  TPNR2D0BWP12T U2830 ( .A1(n2095), .A2(n2059), .ZN(n2060) );
  NR2D1BWP12T U2831 ( .A1(n2061), .A2(n2060), .ZN(n2128) );
  AOI22D0BWP12T U2832 ( .A1(n2988), .A2(n2083), .B1(n2128), .B2(n2929), .ZN(
        n2071) );
  INVD1BWP12T U2833 ( .I(n2119), .ZN(n2931) );
  CKND2D0BWP12T U2834 ( .A1(n2107), .A2(n2062), .ZN(n2068) );
  AOI22D0BWP12T U2835 ( .A1(n2109), .A2(n2064), .B1(n2108), .B2(n2063), .ZN(
        n2067) );
  CKND2D0BWP12T U2836 ( .A1(n2110), .A2(n2065), .ZN(n2066) );
  AOI31D0BWP12T U2837 ( .A1(n2068), .A2(n2067), .A3(n2066), .B(n2123), .ZN(
        n2069) );
  AOI21D0BWP12T U2838 ( .A1(n2133), .A2(n2931), .B(n2069), .ZN(n2070) );
  CKND2D1BWP12T U2839 ( .A1(n2071), .A2(n2070), .ZN(n2435) );
  INVD0BWP12T U2840 ( .I(n2075), .ZN(n2079) );
  CKND2D0BWP12T U2841 ( .A1(n2077), .A2(n2076), .ZN(n2078) );
  ND2D1BWP12T U2842 ( .A1(n2079), .A2(n2078), .ZN(n2784) );
  ND4D0BWP12T U2843 ( .A1(n2432), .A2(n2080), .A3(n2378), .A4(n2992), .ZN(
        n2081) );
  NR3D0BWP12T U2844 ( .A1(n2784), .A2(n2550), .A3(n2081), .ZN(n2082) );
  CKND2D0BWP12T U2845 ( .A1(n2808), .A2(n2082), .ZN(n2403) );
  INVD0BWP12T U2846 ( .I(n2266), .ZN(n2090) );
  TPAOI22D0BWP12T U2847 ( .A1(n2109), .A2(n2091), .B1(n2108), .B2(n2090), .ZN(
        n2094) );
  INVD0BWP12T U2848 ( .I(n2268), .ZN(n2092) );
  TPND2D0BWP12T U2849 ( .A1(n2110), .A2(n2092), .ZN(n2093) );
  OAI211D1BWP12T U2850 ( .A1(n2095), .A2(n2265), .B(n2094), .C(n2093), .ZN(
        n2934) );
  AOI22D1BWP12T U2851 ( .A1(n2107), .A2(n2098), .B1(n2097), .B2(n2096), .ZN(
        n2105) );
  INVD0BWP12T U2852 ( .I(n2274), .ZN(n2102) );
  NR2D0BWP12T U2853 ( .A1(n2099), .A2(n2272), .ZN(n2100) );
  AOI22D1BWP12T U2854 ( .A1(n2103), .A2(n2102), .B1(n2101), .B2(n2100), .ZN(
        n2104) );
  ND2D1BWP12T U2855 ( .A1(n2105), .A2(n2104), .ZN(n2930) );
  OR3D0BWP12T U2856 ( .A1(n2892), .A2(n2139), .A3(n2930), .Z(n2117) );
  INR2D1BWP12T U2857 ( .A1(n2106), .B1(n2353), .ZN(n2932) );
  CKND0BWP12T U2858 ( .I(n2932), .ZN(n2331) );
  CKND2D0BWP12T U2859 ( .A1(n2107), .A2(n2321), .ZN(n2113) );
  AOI22D0BWP12T U2860 ( .A1(n2109), .A2(n2325), .B1(n2108), .B2(n2322), .ZN(
        n2112) );
  CKND2D0BWP12T U2861 ( .A1(n2110), .A2(n2326), .ZN(n2111) );
  TPAOI31D0BWP12T U2862 ( .A1(n2113), .A2(n2112), .A3(n2111), .B(n2123), .ZN(
        n2115) );
  AOI211D0BWP12T U2863 ( .A1(n2988), .A2(n2331), .B(n2115), .C(n2114), .ZN(
        n2116) );
  OAI211D1BWP12T U2864 ( .A1(n2121), .A2(n2934), .B(n2117), .C(n2116), .ZN(
        n2540) );
  OAI22D0BWP12T U2865 ( .A1(n2122), .A2(n2121), .B1(n2120), .B2(n2119), .ZN(
        n2127) );
  AOI21D0BWP12T U2866 ( .A1(n2125), .A2(n2124), .B(n2123), .ZN(n2126) );
  NR2D1BWP12T U2867 ( .A1(n2127), .A2(n2126), .ZN(n2691) );
  INVD1BWP12T U2868 ( .I(n2128), .ZN(n2131) );
  AOI22D0BWP12T U2869 ( .A1(n2131), .A2(n2933), .B1(n2130), .B2(n2129), .ZN(
        n2132) );
  OAI211D0BWP12T U2870 ( .A1(n2134), .A2(n2133), .B(n2132), .C(n2142), .ZN(
        n2607) );
  AOI22D0BWP12T U2871 ( .A1(n2933), .A2(n2136), .B1(n2135), .B2(n2139), .ZN(
        n2137) );
  OAI211D0BWP12T U2872 ( .A1(n2892), .A2(n2138), .B(n2137), .C(n2142), .ZN(
        n2632) );
  AOI22D0BWP12T U2873 ( .A1(n2141), .A2(n2933), .B1(n2140), .B2(n2139), .ZN(
        n2143) );
  OAI211D0BWP12T U2874 ( .A1(n2892), .A2(n2144), .B(n2143), .C(n2142), .ZN(
        n2569) );
  AOI22D0BWP12T U2875 ( .A1(a[22]), .A2(n1720), .B1(n1141), .B2(n2460), .ZN(
        n2155) );
  AOI22D1BWP12T U2876 ( .A1(a[20]), .A2(n2148), .B1(n1379), .B2(n2571), .ZN(
        n2154) );
  AOI22D1BWP12T U2877 ( .A1(n2652), .A2(n2149), .B1(n1450), .B2(n2594), .ZN(
        n2153) );
  AOI22D1BWP12T U2878 ( .A1(n2915), .A2(n2151), .B1(n2150), .B2(n2621), .ZN(
        n2152) );
  ND4D1BWP12T U2879 ( .A1(n2155), .A2(n2154), .A3(n2153), .A4(n2152), .ZN(
        n2187) );
  AOI22D1BWP12T U2880 ( .A1(a[14]), .A2(n2157), .B1(n2156), .B2(n2679), .ZN(
        n2167) );
  AOI22D1BWP12T U2881 ( .A1(a[12]), .A2(n2159), .B1(n2158), .B2(n2710), .ZN(
        n2166) );
  AOI22D1BWP12T U2882 ( .A1(n3100), .A2(n2161), .B1(n2160), .B2(a[13]), .ZN(
        n2165) );
  AOI22D1BWP12T U2883 ( .A1(n2898), .A2(n2163), .B1(n2162), .B2(n2846), .ZN(
        n2164) );
  ND4D1BWP12T U2884 ( .A1(n2167), .A2(n2166), .A3(n2165), .A4(n2164), .ZN(
        n2186) );
  AOI22D1BWP12T U2885 ( .A1(n2785), .A2(n2169), .B1(n2168), .B2(n2870), .ZN(
        n2176) );
  AOI22D1BWP12T U2886 ( .A1(n2738), .A2(n2377), .B1(n2170), .B2(n2815), .ZN(
        n2175) );
  AOI22D1BWP12T U2887 ( .A1(n2352), .A2(n2207), .B1(n2171), .B2(n2466), .ZN(
        n2174) );
  AOI22D1BWP12T U2888 ( .A1(a[3]), .A2(n2263), .B1(n2368), .B2(n2172), .ZN(
        n2173) );
  ND4D1BWP12T U2889 ( .A1(n2176), .A2(n2175), .A3(n2174), .A4(n2173), .ZN(
        n2185) );
  CKND0BWP12T U2890 ( .I(b[30]), .ZN(n2177) );
  AOI22D0BWP12T U2891 ( .A1(a[28]), .A2(n937), .B1(n2177), .B2(a[30]), .ZN(
        n2183) );
  AOI22D1BWP12T U2892 ( .A1(a[26]), .A2(n2178), .B1(n1377), .B2(n2498), .ZN(
        n2182) );
  AOI22D1BWP12T U2893 ( .A1(n2541), .A2(n1452), .B1(n993), .B2(n2358), .ZN(
        n2181) );
  ND2D1BWP12T U2894 ( .A1(n2179), .A2(n2349), .ZN(n2180) );
  ND4D1BWP12T U2895 ( .A1(n2183), .A2(n2182), .A3(n2181), .A4(n2180), .ZN(
        n2184) );
  NR4D0BWP12T U2896 ( .A1(n2187), .A2(n2186), .A3(n2185), .A4(n2184), .ZN(
        n2376) );
  AOI22D1BWP12T U2897 ( .A1(b[23]), .A2(n2574), .B1(n3022), .B2(b[22]), .ZN(
        n2191) );
  AOI22D1BWP12T U2898 ( .A1(b[20]), .A2(n2952), .B1(n2596), .B2(b[21]), .ZN(
        n2190) );
  AOI22D0BWP12T U2899 ( .A1(b[18]), .A2(n2650), .B1(n2623), .B2(b[19]), .ZN(
        n2189) );
  AOI22D0BWP12T U2900 ( .A1(b[16]), .A2(n2917), .B1(n2682), .B2(b[17]), .ZN(
        n2188) );
  ND4D1BWP12T U2901 ( .A1(n2191), .A2(n2190), .A3(n2189), .A4(n2188), .ZN(
        n2220) );
  AOI22D0BWP12T U2902 ( .A1(b[15]), .A2(n2712), .B1(n2192), .B2(b[14]), .ZN(
        n2197) );
  AOI22D0BWP12T U2903 ( .A1(n2452), .A2(n2193), .B1(n3059), .B2(b[13]), .ZN(
        n2196) );
  AOI22D0BWP12T U2904 ( .A1(n2904), .A2(n2900), .B1(n3104), .B2(n3106), .ZN(
        n2195) );
  AOI22D1BWP12T U2905 ( .A1(n2852), .A2(n2848), .B1(n2872), .B2(n2876), .ZN(
        n2194) );
  ND4D1BWP12T U2906 ( .A1(n2197), .A2(n2196), .A3(n2195), .A4(n2194), .ZN(
        n2219) );
  AO22D0BWP12T U2907 ( .A1(b[28]), .A2(n2198), .B1(n2428), .B2(b[29]), .Z(
        n2199) );
  AOI211D0BWP12T U2908 ( .A1(b[30]), .A2(n2996), .B(n2199), .C(n3099), .ZN(
        n2205) );
  AOI22D0BWP12T U2909 ( .A1(b[27]), .A2(n2201), .B1(n2200), .B2(b[26]), .ZN(
        n2204) );
  AOI22D0BWP12T U2910 ( .A1(b[24]), .A2(n2544), .B1(n2202), .B2(b[25]), .ZN(
        n2203) );
  ND4D0BWP12T U2911 ( .A1(n2205), .A2(n2204), .A3(n2203), .A4(n2530), .ZN(
        n2214) );
  AOI22D1BWP12T U2912 ( .A1(n2817), .A2(n2819), .B1(n2787), .B2(n2792), .ZN(
        n2213) );
  AOI22D1BWP12T U2913 ( .A1(n2740), .A2(n2739), .B1(n2206), .B2(n2351), .ZN(
        n2212) );
  OAI22D1BWP12T U2914 ( .A1(n2352), .A2(n2207), .B1(n2314), .B2(a[3]), .ZN(
        n2209) );
  AOI211D1BWP12T U2915 ( .A1(n2350), .A2(n2210), .B(n2209), .C(n2208), .ZN(
        n2211) );
  IND4D1BWP12T U2916 ( .A1(n2214), .B1(n2213), .B2(n2212), .B3(n2211), .ZN(
        n2218) );
  OAI21D1BWP12T U2917 ( .A1(n2216), .A2(b[31]), .B(n2215), .ZN(n2217) );
  TPOAI31D0BWP12T U2918 ( .A1(n2220), .A2(n2219), .A3(n2218), .B(n2217), .ZN(
        n2375) );
  MUX2ND0BWP12T U2919 ( .I0(n2315), .I1(n2827), .S(n2764), .ZN(n2222) );
  NR2D1BWP12T U2920 ( .A1(n2222), .A2(n2393), .ZN(n2718) );
  AOI22D0BWP12T U2921 ( .A1(n2324), .A2(n2224), .B1(n896), .B2(n2223), .ZN(
        n2227) );
  CKND2D0BWP12T U2922 ( .A1(n2225), .A2(n2320), .ZN(n2226) );
  OAI211D0BWP12T U2923 ( .A1(n2229), .A2(n2228), .B(n2227), .C(n2226), .ZN(
        n2280) );
  AOI22D0BWP12T U2924 ( .A1(n896), .A2(n2231), .B1(n2230), .B2(n2324), .ZN(
        n2235) );
  AOI22D0BWP12T U2925 ( .A1(n2323), .A2(n2233), .B1(n2232), .B2(n2320), .ZN(
        n2234) );
  AOI21D0BWP12T U2926 ( .A1(n2235), .A2(n2234), .B(n2327), .ZN(n2236) );
  AOI211D0BWP12T U2927 ( .A1(n2280), .A2(n2333), .B(n2236), .C(n2383), .ZN(
        n2244) );
  AOI22D0BWP12T U2928 ( .A1(n896), .A2(n2238), .B1(n2237), .B2(n2324), .ZN(
        n2242) );
  AOI22D0BWP12T U2929 ( .A1(n2240), .A2(n2323), .B1(n2239), .B2(n2320), .ZN(
        n2241) );
  ND2D1BWP12T U2930 ( .A1(n2242), .A2(n2241), .ZN(n2307) );
  CKND2D1BWP12T U2931 ( .A1(n2307), .A2(n2255), .ZN(n2243) );
  OAI211D0BWP12T U2932 ( .A1(n2308), .A2(n2258), .B(n2244), .C(n2243), .ZN(
        n2426) );
  AOI22D0BWP12T U2933 ( .A1(n2323), .A2(n2326), .B1(n2246), .B2(n2320), .ZN(
        n2249) );
  CKND2D0BWP12T U2934 ( .A1(n2247), .A2(n2324), .ZN(n2248) );
  OAI211D0BWP12T U2935 ( .A1(n2498), .A2(n2250), .B(n2249), .C(n2248), .ZN(
        n2252) );
  AOI211D0BWP12T U2936 ( .A1(n2252), .A2(n2316), .B(n2251), .C(n2383), .ZN(
        n2257) );
  AOI22D0BWP12T U2937 ( .A1(n2324), .A2(n2321), .B1(n2322), .B2(n2320), .ZN(
        n2254) );
  AOI22D0BWP12T U2938 ( .A1(n896), .A2(n2325), .B1(n2268), .B2(n2323), .ZN(
        n2253) );
  CKND2D1BWP12T U2939 ( .A1(n2254), .A2(n2253), .ZN(n2259) );
  AOI22D0BWP12T U2940 ( .A1(n2333), .A2(n2259), .B1(n2262), .B2(n2255), .ZN(
        n2256) );
  OA211D0BWP12T U2941 ( .A1(n2793), .A2(n2258), .B(n2257), .C(n2256), .Z(n2990) );
  INVD1BWP12T U2942 ( .I(n2259), .ZN(n2260) );
  OAI22D0BWP12T U2943 ( .A1(n2793), .A2(n2377), .B1(n2260), .B2(n2327), .ZN(
        n2261) );
  AOI211XD0BWP12T U2944 ( .A1(n2764), .A2(n2262), .B(n2261), .C(n2289), .ZN(
        n3035) );
  CKND2D0BWP12T U2945 ( .A1(n2264), .A2(n2263), .ZN(n2300) );
  AOI22D0BWP12T U2946 ( .A1(n2323), .A2(n2266), .B1(n2265), .B2(n2320), .ZN(
        n2270) );
  AOI22D0BWP12T U2947 ( .A1(n896), .A2(n2268), .B1(n2267), .B2(n2324), .ZN(
        n2269) );
  ND2D1BWP12T U2948 ( .A1(n2270), .A2(n2269), .ZN(n2334) );
  AOI22D0BWP12T U2949 ( .A1(n2323), .A2(n2272), .B1(n2271), .B2(n2320), .ZN(
        n2276) );
  AOI22D0BWP12T U2950 ( .A1(n896), .A2(n2274), .B1(n2273), .B2(n2324), .ZN(
        n2275) );
  ND2D1BWP12T U2951 ( .A1(n2276), .A2(n2275), .ZN(n2311) );
  AOI22D0BWP12T U2952 ( .A1(n2316), .A2(n2334), .B1(n2311), .B2(n2764), .ZN(
        n2277) );
  INVD1BWP12T U2953 ( .I(n2289), .ZN(n2318) );
  OAI211D1BWP12T U2954 ( .A1(n2932), .A2(n2377), .B(n2277), .C(n2318), .ZN(
        n2927) );
  OAI211D1BWP12T U2955 ( .A1(n2300), .A2(n2393), .B(n2927), .C(n3067), .ZN(
        n2278) );
  NR4D0BWP12T U2956 ( .A1(n2990), .A2(n3035), .A3(n2279), .A4(n2278), .ZN(
        n2298) );
  INVD1BWP12T U2957 ( .I(n2280), .ZN(n2281) );
  OAI22D0BWP12T U2958 ( .A1(n2281), .A2(n2327), .B1(n2308), .B2(n2377), .ZN(
        n2282) );
  AOI211XD0BWP12T U2959 ( .A1(n2764), .A2(n2307), .B(n2282), .C(n2289), .ZN(
        n2604) );
  AOI22D0BWP12T U2960 ( .A1(n2316), .A2(n2284), .B1(n2283), .B2(n2764), .ZN(
        n2285) );
  OA211D0BWP12T U2961 ( .A1(n2737), .A2(n2377), .B(n2285), .C(n2318), .Z(n2957) );
  MOAI22D0BWP12T U2962 ( .A1(n2288), .A2(n2287), .B1(n2316), .B2(n2286), .ZN(
        n2290) );
  RCAOI211D0BWP12T U2963 ( .A1(n2740), .A2(n2291), .B(n2290), .C(n2289), .ZN(
        n2687) );
  INVD1BWP12T U2964 ( .I(n2292), .ZN(n2752) );
  ND3D0BWP12T U2965 ( .A1(n2752), .A2(n2396), .A3(n2314), .ZN(n2295) );
  AOI222D1BWP12T U2966 ( .A1(n2295), .A2(n2393), .B1(n2294), .B2(n2333), .C1(
        n2293), .C2(n2316), .ZN(n2627) );
  NR4D0BWP12T U2967 ( .A1(n2604), .A2(n2957), .A3(n2687), .A4(n2627), .ZN(
        n2297) );
  IND4D0BWP12T U2968 ( .A1(n2299), .B1(n2298), .B2(n2297), .B3(n2296), .ZN(
        n2344) );
  INVD1BWP12T U2969 ( .I(n2300), .ZN(n2301) );
  AOI21D0BWP12T U2970 ( .A1(n2396), .A2(n2301), .B(n2402), .ZN(n2305) );
  NR3D0BWP12T U2971 ( .A1(n2303), .A2(n2302), .A3(n2327), .ZN(n2304) );
  RCAOI211D0BWP12T U2972 ( .A1(n2333), .A2(n2306), .B(n2305), .C(n2304), .ZN(
        n2656) );
  INVD0BWP12T U2973 ( .I(n2307), .ZN(n2309) );
  MUX2NXD0BWP12T U2974 ( .I0(n2309), .I1(n2308), .S(n2764), .ZN(n2310) );
  NR2D1BWP12T U2975 ( .A1(n2310), .A2(n2393), .ZN(n3068) );
  INVD1BWP12T U2976 ( .I(n2311), .ZN(n2338) );
  MUX2NXD0BWP12T U2977 ( .I0(n2338), .I1(n2932), .S(n2764), .ZN(n2312) );
  NR2D1BWP12T U2978 ( .A1(n2312), .A2(n2393), .ZN(n2845) );
  NR4D0BWP12T U2979 ( .A1(n2656), .A2(n3068), .A3(n2845), .A4(n2313), .ZN(
        n2340) );
  MAOI22D0BWP12T U2980 ( .A1(n2317), .A2(n2316), .B1(n2315), .B2(n2314), .ZN(
        n2319) );
  OAI211D0BWP12T U2981 ( .A1(n2827), .A2(n2377), .B(n2319), .C(n2318), .ZN(
        n2572) );
  AOI22D0BWP12T U2982 ( .A1(n2323), .A2(n2322), .B1(n2321), .B2(n2320), .ZN(
        n2329) );
  AOI22D0BWP12T U2983 ( .A1(n896), .A2(n2326), .B1(n2325), .B2(n2324), .ZN(
        n2328) );
  AOI21D0BWP12T U2984 ( .A1(n2329), .A2(n2328), .B(n2327), .ZN(n2330) );
  AOI211D0BWP12T U2985 ( .A1(n2332), .A2(n2331), .B(n2330), .C(n2383), .ZN(
        n2336) );
  ND2XD0BWP12T U2986 ( .A1(n2334), .A2(n2333), .ZN(n2335) );
  OAI211D1BWP12T U2987 ( .A1(n2338), .A2(n2337), .B(n2336), .C(n2335), .ZN(
        n2553) );
  ND4D0BWP12T U2988 ( .A1(n2340), .A2(n2339), .A3(n2572), .A4(n2553), .ZN(
        n2343) );
  NR4D0BWP12T U2989 ( .A1(n2344), .A2(n2343), .A3(n2342), .A4(n2341), .ZN(
        n2374) );
  AOI22D0BWP12T U2990 ( .A1(n2852), .A2(n2846), .B1(n2792), .B2(n2785), .ZN(
        n2348) );
  AOI22D1BWP12T U2991 ( .A1(n2979), .A2(b[31]), .B1(n2817), .B2(n2815), .ZN(
        n2347) );
  AOI22D0BWP12T U2992 ( .A1(b[13]), .A2(a[13]), .B1(b[14]), .B2(a[14]), .ZN(
        n2346) );
  AOI22D1BWP12T U2993 ( .A1(n2904), .A2(n2898), .B1(n3106), .B2(n3100), .ZN(
        n2345) );
  ND4D1BWP12T U2994 ( .A1(n2348), .A2(n2347), .A3(n2346), .A4(n2345), .ZN(
        n2372) );
  AOI22D1BWP12T U2995 ( .A1(b[26]), .A2(a[26]), .B1(n2350), .B2(n2349), .ZN(
        n2357) );
  AOI22D1BWP12T U2996 ( .A1(b[24]), .A2(n2541), .B1(b[25]), .B2(n2460), .ZN(
        n2356) );
  AOI22D1BWP12T U2997 ( .A1(n2351), .A2(n2466), .B1(n2740), .B2(n2738), .ZN(
        n2355) );
  AOI22D1BWP12T U2998 ( .A1(n2764), .A2(a[3]), .B1(n2353), .B2(n2352), .ZN(
        n2354) );
  ND4D1BWP12T U2999 ( .A1(n2357), .A2(n2356), .A3(n2355), .A4(n2354), .ZN(
        n2371) );
  AOI22D1BWP12T U3000 ( .A1(b[21]), .A2(n2594), .B1(b[20]), .B2(a[20]), .ZN(
        n2362) );
  AOI22D0BWP12T U3001 ( .A1(b[22]), .A2(a[22]), .B1(b[30]), .B2(a[30]), .ZN(
        n2361) );
  AOI22D0BWP12T U3002 ( .A1(b[27]), .A2(n2358), .B1(b[29]), .B2(n2498), .ZN(
        n2360) );
  AOI22D1BWP12T U3003 ( .A1(b[28]), .A2(a[28]), .B1(b[23]), .B2(n2571), .ZN(
        n2359) );
  ND4D1BWP12T U3004 ( .A1(n2362), .A2(n2361), .A3(n2360), .A4(n2359), .ZN(
        n2370) );
  AOI22D0BWP12T U3005 ( .A1(n2452), .A2(a[12]), .B1(b[15]), .B2(n2710), .ZN(
        n2365) );
  AOI22D0BWP12T U3006 ( .A1(b[18]), .A2(n2652), .B1(b[16]), .B2(n2915), .ZN(
        n2364) );
  AOI22D0BWP12T U3007 ( .A1(b[19]), .A2(n2621), .B1(b[17]), .B2(n2679), .ZN(
        n2363) );
  ND3D1BWP12T U3008 ( .A1(n2365), .A2(n2364), .A3(n2363), .ZN(n2366) );
  AOI211D1BWP12T U3009 ( .A1(n2876), .A2(n2870), .B(n3018), .C(n2366), .ZN(
        n2367) );
  OAI21D1BWP12T U3010 ( .A1(n2368), .A2(n2449), .B(n2367), .ZN(n2369) );
  NR4D0BWP12T U3011 ( .A1(n2372), .A2(n2371), .A3(n2370), .A4(n2369), .ZN(
        n2373) );
  AOI211XD0BWP12T U3012 ( .A1(n2376), .A2(n2375), .B(n2374), .C(n2373), .ZN(
        n2405) );
  NR2D0BWP12T U3013 ( .A1(n2378), .A2(n2377), .ZN(n2708) );
  CKND2D0BWP12T U3014 ( .A1(n2397), .A2(n2396), .ZN(n2382) );
  AOI21D1BWP12T U3015 ( .A1(n2382), .A2(n2393), .B(n2381), .ZN(n2868) );
  INVD1BWP12T U3016 ( .I(n2784), .ZN(n3030) );
  AOI211D1BWP12T U3017 ( .A1(n2740), .A2(n3030), .B(n2797), .C(n2383), .ZN(
        n2783) );
  CKND2D0BWP12T U3018 ( .A1(n3092), .A2(n2396), .ZN(n2385) );
  AOI21D1BWP12T U3019 ( .A1(n2385), .A2(n2393), .B(n3112), .ZN(n3081) );
  INVD1BWP12T U3020 ( .I(n2388), .ZN(n2855) );
  CKND2D0BWP12T U3021 ( .A1(n2392), .A2(n2396), .ZN(n2394) );
  AOI21D1BWP12T U3022 ( .A1(n2394), .A2(n2393), .B(n2741), .ZN(n2736) );
  INVD1BWP12T U3023 ( .I(n2398), .ZN(n2659) );
  OAI211D1BWP12T U3024 ( .A1(n2407), .A2(n2406), .B(n2405), .C(n2404), .ZN(
        n2408) );
  AOI211D1BWP12T U3025 ( .A1(n2410), .A2(n2449), .B(n2409), .C(n2408), .ZN(
        n2411) );
  OAI31D0BWP12T U3026 ( .A1(n3007), .A2(n2413), .A3(n2412), .B(n2411), .ZN(
        n2414) );
  AOI211D1BWP12T U3027 ( .A1(n2417), .A2(n2416), .B(n2415), .C(n2414), .ZN(
        n2418) );
  OAI211D1BWP12T U3028 ( .A1(n2421), .A2(n2420), .B(n2419), .C(n2418), .ZN(z)
         );
  INVD1BWP12T U3029 ( .I(n2422), .ZN(n2446) );
  TPND2D0BWP12T U3030 ( .A1(n2423), .A2(n3082), .ZN(n2440) );
  CKND2D1BWP12T U3031 ( .A1(n2424), .A2(n3093), .ZN(n2439) );
  MOAI22D0BWP12T U3032 ( .A1(n2426), .A2(n2928), .B1(n2425), .B2(n3084), .ZN(
        n2434) );
  OAI21D0BWP12T U3033 ( .A1(n2498), .A2(n3099), .B(n3103), .ZN(n2427) );
  AOI22D0BWP12T U3034 ( .A1(n3105), .A2(n2428), .B1(n2427), .B2(b[29]), .ZN(
        n2431) );
  MUX2ND0BWP12T U3035 ( .I0(n3019), .I1(n3018), .S(b[29]), .ZN(n2429) );
  OAI21D0BWP12T U3036 ( .A1(n2429), .A2(n3020), .B(n2498), .ZN(n2430) );
  OAI211D1BWP12T U3037 ( .A1(n2432), .A2(n2991), .B(n2431), .C(n2430), .ZN(
        n2433) );
  AOI211XD0BWP12T U3038 ( .A1(n3091), .A2(n2435), .B(n2434), .C(n2433), .ZN(
        n2438) );
  ND2D1BWP12T U3039 ( .A1(n2436), .A2(n3096), .ZN(n2437) );
  ND4D1BWP12T U3040 ( .A1(n2440), .A2(n2439), .A3(n2438), .A4(n2437), .ZN(
        n2441) );
  AOI21D1BWP12T U3041 ( .A1(n382), .A2(n2442), .B(n2441), .ZN(n2445) );
  CKND2D1BWP12T U3042 ( .A1(n2443), .A2(n3076), .ZN(n2444) );
  OAI211D1BWP12T U3043 ( .A1(n2975), .A2(n2446), .B(n2445), .C(n2444), .ZN(
        result[29]) );
  FA1D1BWP12T U3044 ( .A(mult_x_18_n404), .B(mult_x_18_n382), .CI(n2447), .CO(
        n2523), .S(n2524) );
  AO21D0BWP12T U3045 ( .A1(n2450), .A2(n2449), .B(n2448), .Z(n2451) );
  XNR2XD0BWP12T U3046 ( .A1(n2710), .A2(b[18]), .ZN(n2471) );
  OAI22D0BWP12T U3047 ( .A1(n2474), .A2(n2473), .B1(n2472), .B2(n2471), .ZN(
        n2480) );
  XOR2XD0BWP12T U3048 ( .A1(n2792), .A2(n2201), .Z(n2475) );
  OAI22D0BWP12T U3049 ( .A1(n2478), .A2(n2477), .B1(n2476), .B2(n2475), .ZN(
        n2479) );
  CKXOR2D1BWP12T U3050 ( .A1(n2480), .A2(n2479), .Z(n2485) );
  XNR2XD0BWP12T U3051 ( .A1(n2621), .A2(b[14]), .ZN(n2481) );
  XNR2D1BWP12T U3052 ( .A1(n2516), .A2(b[30]), .ZN(n2517) );
  XOR2D1BWP12T U3053 ( .A1(n2983), .A2(n2524), .Z(n2536) );
  CKND2D0BWP12T U3054 ( .A1(n3047), .A2(n3089), .ZN(n2529) );
  FA1D2BWP12T U3055 ( .A(n2216), .B(b[31]), .CI(n2525), .CO(n2526), .S(n2421)
         );
  FA1D1BWP12T U3056 ( .A(n2216), .B(b[31]), .CI(n2527), .CO(n2528), .S(n1725)
         );
  MUX2NXD0BWP12T U3057 ( .I0(n2529), .I1(n2981), .S(n2979), .ZN(n2531) );
  NR2D1BWP12T U3058 ( .A1(n2531), .A2(n2530), .ZN(n2535) );
  NR2D0BWP12T U3059 ( .A1(n2532), .A2(n2979), .ZN(n2982) );
  AO211D1BWP12T U3060 ( .A1(n2536), .A2(n3117), .B(n2535), .C(n2534), .Z(v) );
  INVD1BWP12T U3061 ( .I(n2537), .ZN(n2565) );
  INVD1BWP12T U3062 ( .I(n2538), .ZN(n2559) );
  CKND2D1BWP12T U3063 ( .A1(n2539), .A2(n3093), .ZN(n2558) );
  NR2D1BWP12T U3064 ( .A1(n2540), .A2(n3004), .ZN(n2555) );
  OAI21D1BWP12T U3065 ( .A1(n2541), .A2(n3099), .B(n3103), .ZN(n2548) );
  NR2D0BWP12T U3066 ( .A1(n2542), .A2(n3071), .ZN(n2547) );
  MUX2ND0BWP12T U3067 ( .I0(n3019), .I1(n3018), .S(b[24]), .ZN(n2543) );
  NR2D0BWP12T U3068 ( .A1(n2543), .A2(n3020), .ZN(n2545) );
  MUX2ND0BWP12T U3069 ( .I0(n2545), .I1(n3023), .S(n2544), .ZN(n2546) );
  AOI211D0BWP12T U3070 ( .A1(b[24]), .A2(n2548), .B(n2547), .C(n2546), .ZN(
        n2552) );
  NR2D1BWP12T U3071 ( .A1(n2549), .A2(n3071), .ZN(n3001) );
  INVD1BWP12T U3072 ( .I(n3001), .ZN(n3031) );
  CKND2D1BWP12T U3073 ( .A1(n3029), .A2(n3031), .ZN(n2924) );
  CKND2D1BWP12T U3074 ( .A1(n2924), .A2(n2550), .ZN(n2551) );
  OAI211D1BWP12T U3075 ( .A1(n2928), .A2(n2553), .B(n2552), .C(n2551), .ZN(
        n2554) );
  RCAOI211D0BWP12T U3076 ( .A1(n2556), .A2(n3096), .B(n2555), .C(n2554), .ZN(
        n2557) );
  OAI211D1BWP12T U3077 ( .A1(n2559), .A2(n2967), .B(n2558), .C(n2557), .ZN(
        n2560) );
  AOI21D1BWP12T U3078 ( .A1(n382), .A2(n2561), .B(n2560), .ZN(n2564) );
  CKND2D1BWP12T U3079 ( .A1(n2562), .A2(n3076), .ZN(n2563) );
  OAI211D1BWP12T U3080 ( .A1(n2975), .A2(n2565), .B(n2564), .C(n2563), .ZN(
        result[24]) );
  INVD1BWP12T U3081 ( .I(n2566), .ZN(n2591) );
  INVD1BWP12T U3082 ( .I(n2567), .ZN(n2585) );
  CKND2D1BWP12T U3083 ( .A1(n2568), .A2(n3093), .ZN(n2584) );
  MAOI22D0BWP12T U3084 ( .A1(n3084), .A2(n2570), .B1(n2569), .B2(n3004), .ZN(
        n2580) );
  OAI21D1BWP12T U3085 ( .A1(n2571), .A2(n3099), .B(n3103), .ZN(n2578) );
  NR2XD0BWP12T U3086 ( .A1(n2572), .A2(n2928), .ZN(n2577) );
  MUX2ND0BWP12T U3087 ( .I0(n3019), .I1(n3018), .S(b[23]), .ZN(n2573) );
  NR2D0BWP12T U3088 ( .A1(n2573), .A2(n3020), .ZN(n2575) );
  MUX2ND0BWP12T U3089 ( .I0(n2575), .I1(n3023), .S(n2574), .ZN(n2576) );
  AOI211D0BWP12T U3090 ( .A1(b[23]), .A2(n2578), .B(n2577), .C(n2576), .ZN(
        n2579) );
  OAI211D1BWP12T U3091 ( .A1(n2808), .A2(n3029), .B(n2580), .C(n2579), .ZN(
        n2581) );
  AOI21D1BWP12T U3092 ( .A1(n2582), .A2(n3096), .B(n2581), .ZN(n2583) );
  OAI211D1BWP12T U3093 ( .A1(n2585), .A2(n2967), .B(n2584), .C(n2583), .ZN(
        n2586) );
  AOI21D1BWP12T U3094 ( .A1(n382), .A2(n2587), .B(n2586), .ZN(n2590) );
  CKND2D1BWP12T U3095 ( .A1(n2588), .A2(n3076), .ZN(n2589) );
  OAI211D1BWP12T U3096 ( .A1(n2975), .A2(n2591), .B(n2590), .C(n2589), .ZN(
        result[23]) );
  INVD1BWP12T U3097 ( .I(n2592), .ZN(n2613) );
  CKND2D1BWP12T U3098 ( .A1(n2593), .A2(n3096), .ZN(n2606) );
  OAI21D1BWP12T U3099 ( .A1(n2594), .A2(n3099), .B(n3103), .ZN(n2599) );
  INVD1BWP12T U3100 ( .I(n3028), .ZN(n2920) );
  MUX2ND0BWP12T U3101 ( .I0(n3019), .I1(n3018), .S(b[21]), .ZN(n2595) );
  NR2D0BWP12T U3102 ( .A1(n2595), .A2(n3020), .ZN(n2597) );
  MUX2ND0BWP12T U3103 ( .I0(n2597), .I1(n3023), .S(n2596), .ZN(n2598) );
  AO211D0BWP12T U3104 ( .A1(b[21]), .A2(n2599), .B(n2920), .C(n2598), .Z(n2603) );
  OAI22D0BWP12T U3105 ( .A1(n2601), .A2(n3031), .B1(n3029), .B2(n2600), .ZN(
        n2602) );
  RCAOI211D0BWP12T U3106 ( .A1(n3067), .A2(n2604), .B(n2603), .C(n2602), .ZN(
        n2605) );
  OAI211D1BWP12T U3107 ( .A1(n2607), .A2(n3004), .B(n2606), .C(n2605), .ZN(
        n2608) );
  AOI21D1BWP12T U3108 ( .A1(n2609), .A2(n3093), .B(n2608), .ZN(n2612) );
  CKND2D1BWP12T U3109 ( .A1(n2610), .A2(n3082), .ZN(n2611) );
  OAI211D1BWP12T U3110 ( .A1(n3047), .A2(n2613), .B(n2612), .C(n2611), .ZN(
        n2614) );
  AOI21D1BWP12T U3111 ( .A1(n3076), .A2(n2615), .B(n2614), .ZN(n2616) );
  IOA21D2BWP12T U3112 ( .A1(n2617), .A2(n3117), .B(n2616), .ZN(result[21]) );
  INVD1BWP12T U3113 ( .I(n2618), .ZN(n2644) );
  INVD1BWP12T U3114 ( .I(n2619), .ZN(n2638) );
  CKND2D1BWP12T U3115 ( .A1(n2620), .A2(n3093), .ZN(n2637) );
  OAI21D0BWP12T U3116 ( .A1(n2621), .A2(n3099), .B(n3103), .ZN(n2626) );
  MUX2ND0BWP12T U3117 ( .I0(n3019), .I1(n3018), .S(b[19]), .ZN(n2622) );
  NR2D0BWP12T U3118 ( .A1(n2622), .A2(n3020), .ZN(n2624) );
  MUX2ND0BWP12T U3119 ( .I0(n2624), .I1(n3023), .S(n2623), .ZN(n2625) );
  RCAOI211D0BWP12T U3120 ( .A1(b[19]), .A2(n2626), .B(n2920), .C(n2625), .ZN(
        n2629) );
  ND2XD0BWP12T U3121 ( .A1(n2627), .A2(n3067), .ZN(n2628) );
  OAI211D1BWP12T U3122 ( .A1(n3031), .A2(n2630), .B(n2629), .C(n2628), .ZN(
        n2634) );
  OAI22D1BWP12T U3123 ( .A1(n2632), .A2(n3004), .B1(n3029), .B2(n2631), .ZN(
        n2633) );
  AOI211D1BWP12T U3124 ( .A1(n2635), .A2(n3096), .B(n2634), .C(n2633), .ZN(
        n2636) );
  OAI211D1BWP12T U3125 ( .A1(n2638), .A2(n2967), .B(n2637), .C(n2636), .ZN(
        n2639) );
  AOI21D1BWP12T U3126 ( .A1(n3076), .A2(n2640), .B(n2639), .ZN(n2643) );
  CKND2D1BWP12T U3127 ( .A1(n2641), .A2(n382), .ZN(n2642) );
  OAI211D1BWP12T U3128 ( .A1(n2975), .A2(n2644), .B(n2643), .C(n2642), .ZN(
        result[19]) );
  INVD1BWP12T U3129 ( .I(n2645), .ZN(n2674) );
  INVD1BWP12T U3130 ( .I(n2646), .ZN(n2668) );
  TPND2D0BWP12T U3131 ( .A1(n2647), .A2(n3093), .ZN(n2667) );
  CKND2D0BWP12T U3132 ( .A1(n2648), .A2(n3091), .ZN(n2658) );
  MUX2ND0BWP12T U3133 ( .I0(n3019), .I1(n3018), .S(b[18]), .ZN(n2649) );
  NR2D0BWP12T U3134 ( .A1(n2649), .A2(n3020), .ZN(n2651) );
  MUX2NXD0BWP12T U3135 ( .I0(n2651), .I1(n3023), .S(n2650), .ZN(n2655) );
  NR2D0BWP12T U3136 ( .A1(n2652), .A2(n3099), .ZN(n2653) );
  OA21XD0BWP12T U3137 ( .A1(n2653), .A2(n3020), .B(b[18]), .Z(n2654) );
  RCAOI211D0BWP12T U3138 ( .A1(n2656), .A2(n3067), .B(n2655), .C(n2654), .ZN(
        n2657) );
  OAI211D1BWP12T U3139 ( .A1(n2660), .A2(n2659), .B(n2658), .C(n2657), .ZN(
        n2664) );
  INVD1BWP12T U3140 ( .I(n2661), .ZN(n2662) );
  NR2D1BWP12T U3141 ( .A1(n2662), .A2(n3071), .ZN(n2663) );
  RCAOI211D0BWP12T U3142 ( .A1(n2665), .A2(n3096), .B(n2664), .C(n2663), .ZN(
        n2666) );
  OAI211D1BWP12T U3143 ( .A1(n2967), .A2(n2668), .B(n2667), .C(n2666), .ZN(
        n2669) );
  AOI21D1BWP12T U3144 ( .A1(n3076), .A2(n2670), .B(n2669), .ZN(n2673) );
  CKND2D1BWP12T U3145 ( .A1(n2671), .A2(n382), .ZN(n2672) );
  OAI211D1BWP12T U3146 ( .A1(n2975), .A2(n2674), .B(n2673), .C(n2672), .ZN(
        result[18]) );
  INVD1BWP12T U3147 ( .I(n2675), .ZN(n2702) );
  INVD1BWP12T U3148 ( .I(n2676), .ZN(n2696) );
  TPND2D0BWP12T U3149 ( .A1(n2677), .A2(n3093), .ZN(n2695) );
  MUX2ND0BWP12T U3150 ( .I0(n3019), .I1(n3018), .S(b[17]), .ZN(n2678) );
  NR2D0BWP12T U3151 ( .A1(n2678), .A2(n3020), .ZN(n2683) );
  OAI21D0BWP12T U3152 ( .A1(n2679), .A2(n3099), .B(n3103), .ZN(n2680) );
  AOI22D0BWP12T U3153 ( .A1(n3105), .A2(n2682), .B1(n2680), .B2(b[17]), .ZN(
        n2681) );
  OAI211D0BWP12T U3154 ( .A1(n2683), .A2(n2682), .B(n3028), .C(n2681), .ZN(
        n2686) );
  TPNR2D0BWP12T U3155 ( .A1(n3029), .A2(n2684), .ZN(n2685) );
  RCAOI211D0BWP12T U3156 ( .A1(n2687), .A2(n3067), .B(n2686), .C(n2685), .ZN(
        n2690) );
  CKND2D1BWP12T U3157 ( .A1(n2688), .A2(n3001), .ZN(n2689) );
  OAI211D1BWP12T U3158 ( .A1(n2691), .A2(n3004), .B(n2690), .C(n2689), .ZN(
        n2692) );
  AOI21D1BWP12T U3159 ( .A1(n2693), .A2(n3096), .B(n2692), .ZN(n2694) );
  OAI211D1BWP12T U3160 ( .A1(n2696), .A2(n2967), .B(n2695), .C(n2694), .ZN(
        n2697) );
  AOI21D1BWP12T U3161 ( .A1(n3076), .A2(n2698), .B(n2697), .ZN(n2701) );
  CKND2D1BWP12T U3162 ( .A1(n2699), .A2(n382), .ZN(n2700) );
  INVD1BWP12T U3163 ( .I(n2703), .ZN(n2728) );
  AO22XD1BWP12T U3164 ( .A1(n2705), .A2(n3082), .B1(n2704), .B2(n3093), .Z(
        n2723) );
  AOI22D0BWP12T U3165 ( .A1(n3096), .A2(n2707), .B1(n2706), .B2(n3091), .ZN(
        n2720) );
  CKND2D1BWP12T U3166 ( .A1(n3065), .A2(n3004), .ZN(n2750) );
  OA21D1BWP12T U3167 ( .A1(n2709), .A2(n2708), .B(n2750), .Z(n2717) );
  OAI21D0BWP12T U3168 ( .A1(n2710), .A2(n3099), .B(n3103), .ZN(n2715) );
  MUX2ND0BWP12T U3169 ( .I0(n3102), .I1(n3101), .S(b[15]), .ZN(n2711) );
  CKND2D0BWP12T U3170 ( .A1(n2711), .A2(n3103), .ZN(n2713) );
  MUX2ND0BWP12T U3171 ( .I0(n2713), .I1(n3105), .S(n2712), .ZN(n2714) );
  IOA21D1BWP12T U3172 ( .A1(b[15]), .A2(n2715), .B(n2714), .ZN(n2716) );
  RCAOI211D0BWP12T U3173 ( .A1(n3067), .A2(n2718), .B(n2717), .C(n2716), .ZN(
        n2719) );
  OAI211D1BWP12T U3174 ( .A1(n2721), .A2(n3071), .B(n2720), .C(n2719), .ZN(
        n2722) );
  AOI211D1BWP12T U3175 ( .A1(n3076), .A2(n2724), .B(n2723), .C(n2722), .ZN(
        n2727) );
  CKND2D1BWP12T U3176 ( .A1(n2725), .A2(n382), .ZN(n2726) );
  OAI211D1BWP12T U3177 ( .A1(n2975), .A2(n2728), .B(n2727), .C(n2726), .ZN(
        result[15]) );
  CKND2D0BWP12T U3178 ( .A1(n2729), .A2(n3076), .ZN(n2733) );
  AOI22D0BWP12T U3179 ( .A1(n2731), .A2(n3082), .B1(n2730), .B2(n3093), .ZN(
        n2732) );
  OAI211D1BWP12T U3180 ( .A1(n2734), .A2(n3004), .B(n2733), .C(n2732), .ZN(
        n2735) );
  AOI21D1BWP12T U3181 ( .A1(n3080), .A2(n2736), .B(n2735), .ZN(n2746) );
  NR2D0BWP12T U3182 ( .A1(n292), .A2(n3047), .ZN(n2743) );
  AOI211D1BWP12T U3183 ( .A1(n2744), .A2(n3096), .B(n2743), .C(n2742), .ZN(
        n2745) );
  OAI211D1BWP12T U3184 ( .A1(n2747), .A2(n3071), .B(n2746), .C(n2745), .ZN(
        n2748) );
  AO21D1BWP12T U3185 ( .A1(n2749), .A2(n3117), .B(n2748), .Z(result[4]) );
  INVD1BWP12T U3186 ( .I(n2750), .ZN(n2894) );
  INVD1BWP12T U3187 ( .I(n2751), .ZN(n2757) );
  AOI22D1BWP12T U3188 ( .A1(n3096), .A2(n2753), .B1(n2826), .B2(n2752), .ZN(
        n2756) );
  CKND2D0BWP12T U3189 ( .A1(n2754), .A2(n3082), .ZN(n2755) );
  OAI211D1BWP12T U3190 ( .A1(n3089), .A2(n2757), .B(n2756), .C(n2755), .ZN(
        n2769) );
  CKND2D0BWP12T U3191 ( .A1(n2758), .A2(n3093), .ZN(n2766) );
  OAI21D1BWP12T U3192 ( .A1(a[3]), .A2(n3099), .B(n3103), .ZN(n2763) );
  MUX2ND0BWP12T U3193 ( .I0(n3019), .I1(n3018), .S(n2764), .ZN(n2759) );
  NR2D0BWP12T U3194 ( .A1(n2759), .A2(n3020), .ZN(n2761) );
  MUX2ND0BWP12T U3195 ( .I0(n2761), .I1(n3023), .S(n2760), .ZN(n2762) );
  RCAOI21D0BWP12T U3196 ( .A1(n2764), .A2(n2763), .B(n2762), .ZN(n2765) );
  OAI211D1BWP12T U3197 ( .A1(n2767), .A2(n2824), .B(n2766), .C(n2765), .ZN(
        n2768) );
  AOI211D1BWP12T U3198 ( .A1(n382), .A2(n2770), .B(n2769), .C(n2768), .ZN(
        n2773) );
  CKND2D1BWP12T U3199 ( .A1(n2771), .A2(n3084), .ZN(n2772) );
  ND2XD0BWP12T U3200 ( .A1(n2777), .A2(n3117), .ZN(n2805) );
  AOI22D0BWP12T U3201 ( .A1(n3096), .A2(n2779), .B1(n2778), .B2(n382), .ZN(
        n2804) );
  AOI22D0BWP12T U3202 ( .A1(n3082), .A2(n2781), .B1(n2780), .B2(n3093), .ZN(
        n2782) );
  IOA21D1BWP12T U3203 ( .A1(n2783), .A2(n3080), .B(n2782), .ZN(n2799) );
  AOI21D0BWP12T U3204 ( .A1(n2784), .A2(n3091), .B(n3090), .ZN(n2796) );
  OAI21D0BWP12T U3205 ( .A1(n2785), .A2(n3099), .B(n3103), .ZN(n2791) );
  NR2D1BWP12T U3206 ( .A1(n2985), .A2(n2824), .ZN(n2790) );
  MUX2ND0BWP12T U3207 ( .I0(n3019), .I1(n3018), .S(n2792), .ZN(n2786) );
  NR2D0BWP12T U3208 ( .A1(n2786), .A2(n3020), .ZN(n2788) );
  MUX2NXD0BWP12T U3209 ( .I0(n2788), .I1(n3023), .S(n2787), .ZN(n2789) );
  AOI211D1BWP12T U3210 ( .A1(n2792), .A2(n2791), .B(n2790), .C(n2789), .ZN(
        n2795) );
  ND2D1BWP12T U3211 ( .A1(n2826), .A2(n2793), .ZN(n2794) );
  OAI211D1BWP12T U3212 ( .A1(n2797), .A2(n2796), .B(n2795), .C(n2794), .ZN(
        n2798) );
  AOI211D1BWP12T U3213 ( .A1(n3076), .A2(n2800), .B(n2799), .C(n2798), .ZN(
        n2803) );
  TPND2D0BWP12T U3214 ( .A1(n2801), .A2(n3084), .ZN(n2802) );
  ND4D1BWP12T U3215 ( .A1(n2805), .A2(n2804), .A3(n2803), .A4(n2802), .ZN(
        result[6]) );
  OAI21D0BWP12T U3216 ( .A1(n2808), .A2(n3004), .B(n2807), .ZN(n2809) );
  MOAI22D0BWP12T U3217 ( .A1(n2813), .A2(n3071), .B1(n2812), .B2(n3076), .ZN(
        n2833) );
  INVD1BWP12T U3218 ( .I(n2814), .ZN(n2831) );
  OAI21D1BWP12T U3219 ( .A1(n2815), .A2(n3099), .B(n3103), .ZN(n2816) );
  ND2D1BWP12T U3220 ( .A1(n2816), .A2(n2817), .ZN(n2822) );
  MUX2ND0BWP12T U3221 ( .I0(n3102), .I1(n3101), .S(n2817), .ZN(n2818) );
  CKND2D0BWP12T U3222 ( .A1(n2818), .A2(n3103), .ZN(n2820) );
  MUX2ND0BWP12T U3223 ( .I0(n2820), .I1(n3105), .S(n2819), .ZN(n2821) );
  OAI211D1BWP12T U3224 ( .A1(n2824), .A2(n2823), .B(n2822), .C(n2821), .ZN(
        n2825) );
  AOI21D1BWP12T U3225 ( .A1(n2827), .A2(n2826), .B(n2825), .ZN(n2830) );
  CKND2D0BWP12T U3226 ( .A1(n2828), .A2(n3093), .ZN(n2829) );
  OAI211D1BWP12T U3227 ( .A1(n2831), .A2(n2967), .B(n2830), .C(n2829), .ZN(
        n2832) );
  INVD1BWP12T U3228 ( .I(n2836), .ZN(n2862) );
  AOI22D0BWP12T U3229 ( .A1(n3093), .A2(n2838), .B1(n2837), .B2(n3082), .ZN(
        n2839) );
  OAI21D1BWP12T U3230 ( .A1(n2840), .A2(n3004), .B(n2839), .ZN(n2841) );
  AOI21D1BWP12T U3231 ( .A1(n3096), .A2(n2842), .B(n2841), .ZN(n2861) );
  MOAI22D0BWP12T U3232 ( .A1(n2844), .A2(n3071), .B1(n2843), .B2(n3076), .ZN(
        n2858) );
  TPND2D0BWP12T U3233 ( .A1(n2845), .A2(n3067), .ZN(n2854) );
  OAI21D0BWP12T U3234 ( .A1(n2846), .A2(n3099), .B(n3103), .ZN(n2851) );
  MUX2ND0BWP12T U3235 ( .I0(n3019), .I1(n3018), .S(n2852), .ZN(n2847) );
  NR2D0BWP12T U3236 ( .A1(n2847), .A2(n3020), .ZN(n2849) );
  MUX2NXD0BWP12T U3237 ( .I0(n2849), .I1(n3023), .S(n2848), .ZN(n2850) );
  RCAOI21D0BWP12T U3238 ( .A1(n2852), .A2(n2851), .B(n2850), .ZN(n2853) );
  OAI211D1BWP12T U3239 ( .A1(n2856), .A2(n2855), .B(n2854), .C(n2853), .ZN(
        n2857) );
  AOI211XD0BWP12T U3240 ( .A1(n382), .A2(n2859), .B(n2858), .C(n2857), .ZN(
        n2860) );
  OAI211D1BWP12T U3241 ( .A1(n2975), .A2(n2862), .B(n2861), .C(n2860), .ZN(
        result[8]) );
  AOI22D0BWP12T U3242 ( .A1(n3082), .A2(n2864), .B1(n2863), .B2(n3096), .ZN(
        n2865) );
  IOA21D1BWP12T U3243 ( .A1(n3084), .A2(n2866), .B(n2865), .ZN(n2888) );
  INVD1BWP12T U3244 ( .I(n2867), .ZN(n2886) );
  AOI22D0BWP12T U3245 ( .A1(n2869), .A2(n3093), .B1(n3080), .B2(n2868), .ZN(
        n2878) );
  OAI21D1BWP12T U3246 ( .A1(n2870), .A2(n3099), .B(n3103), .ZN(n2875) );
  MUX2ND0BWP12T U3247 ( .I0(n3019), .I1(n3018), .S(n2876), .ZN(n2871) );
  NR2D0BWP12T U3248 ( .A1(n2871), .A2(n3020), .ZN(n2873) );
  MUX2ND0BWP12T U3249 ( .I0(n2873), .I1(n3023), .S(n2872), .ZN(n2874) );
  RCAOI21D0BWP12T U3250 ( .A1(n2876), .A2(n2875), .B(n2874), .ZN(n2877) );
  OAI211D1BWP12T U3251 ( .A1(n2880), .A2(n2879), .B(n2878), .C(n2877), .ZN(
        n2881) );
  RCAOI21D0BWP12T U3252 ( .A1(n382), .A2(n2882), .B(n2881), .ZN(n2885) );
  ND2XD0BWP12T U3253 ( .A1(n2883), .A2(n3091), .ZN(n2884) );
  OAI211D1BWP12T U3254 ( .A1(n2886), .A2(n3089), .B(n2885), .C(n2884), .ZN(
        n2887) );
  AO211D1BWP12T U3255 ( .A1(n2889), .A2(n3117), .B(n2888), .C(n2887), .Z(
        result[9]) );
  CKND2D0BWP12T U3256 ( .A1(n2892), .A2(n3091), .ZN(n3097) );
  OAI22D1BWP12T U3257 ( .A1(n2895), .A2(n2894), .B1(n2893), .B2(n3097), .ZN(
        n2896) );
  OAI21D1BWP12T U3258 ( .A1(n2898), .A2(n3099), .B(n3103), .ZN(n2903) );
  MUX2ND0BWP12T U3259 ( .I0(n3019), .I1(n3018), .S(n2904), .ZN(n2899) );
  NR2D0BWP12T U3260 ( .A1(n2899), .A2(n3020), .ZN(n2901) );
  MUX2ND0BWP12T U3261 ( .I0(n2901), .I1(n3023), .S(n2900), .ZN(n2902) );
  RCAOI21D0BWP12T U3262 ( .A1(n2904), .A2(n2903), .B(n2902), .ZN(n2907) );
  ND2D1BWP12T U3263 ( .A1(n2905), .A2(n3108), .ZN(n2906) );
  OAI211D1BWP12T U3264 ( .A1(n3071), .A2(n2908), .B(n2907), .C(n2906), .ZN(
        n2909) );
  INVD1BWP12T U3265 ( .I(n2913), .ZN(n2946) );
  TPND2D0BWP12T U3266 ( .A1(n2914), .A2(n3093), .ZN(n2940) );
  OAI21D0BWP12T U3267 ( .A1(n2915), .A2(n3099), .B(n3103), .ZN(n2921) );
  MUX2ND0BWP12T U3268 ( .I0(n3019), .I1(n3018), .S(b[16]), .ZN(n2916) );
  NR2D0BWP12T U3269 ( .A1(n2916), .A2(n3020), .ZN(n2918) );
  MUX2ND0BWP12T U3270 ( .I0(n2918), .I1(n3023), .S(n2917), .ZN(n2919) );
  RCAOI211D0BWP12T U3271 ( .A1(b[16]), .A2(n2921), .B(n2920), .C(n2919), .ZN(
        n2926) );
  INVD0BWP12T U3272 ( .I(n2922), .ZN(n2923) );
  ND2D1BWP12T U3273 ( .A1(n2924), .A2(n2923), .ZN(n2925) );
  OAI211D1BWP12T U3274 ( .A1(n2928), .A2(n2927), .B(n2926), .C(n2925), .ZN(
        n2937) );
  AOI222D1BWP12T U3275 ( .A1(n2934), .A2(n2933), .B1(n2932), .B2(n2931), .C1(
        n2930), .C2(n2929), .ZN(n2935) );
  NR2D1BWP12T U3276 ( .A1(n2935), .A2(n3004), .ZN(n2936) );
  RCAOI211D0BWP12T U3277 ( .A1(n2938), .A2(n3096), .B(n2937), .C(n2936), .ZN(
        n2939) );
  OAI211D1BWP12T U3278 ( .A1(n290), .A2(n2967), .B(n2940), .C(n2939), .ZN(
        n2941) );
  AOI21D1BWP12T U3279 ( .A1(n3076), .A2(n2942), .B(n2941), .ZN(n2945) );
  CKND2D1BWP12T U3280 ( .A1(n2943), .A2(n382), .ZN(n2944) );
  INVD1BWP12T U3281 ( .I(n2947), .ZN(n2974) );
  INVD1BWP12T U3282 ( .I(n2948), .ZN(n2968) );
  CKND2D1BWP12T U3283 ( .A1(n2949), .A2(n3093), .ZN(n2966) );
  CKND2D0BWP12T U3284 ( .A1(n2950), .A2(n3091), .ZN(n2959) );
  MUX2ND0BWP12T U3285 ( .I0(n3019), .I1(n3018), .S(b[20]), .ZN(n2951) );
  NR2D0BWP12T U3286 ( .A1(n2951), .A2(n3020), .ZN(n2953) );
  MUX2ND0BWP12T U3287 ( .I0(n2953), .I1(n3023), .S(n2952), .ZN(n2956) );
  NR2D0BWP12T U3288 ( .A1(a[20]), .A2(n3099), .ZN(n2954) );
  OA21XD0BWP12T U3289 ( .A1(n2954), .A2(n3020), .B(b[20]), .Z(n2955) );
  RCAOI211D0BWP12T U3290 ( .A1(n2957), .A2(n3067), .B(n2956), .C(n2955), .ZN(
        n2958) );
  OAI211D1BWP12T U3291 ( .A1(n2960), .A2(n3029), .B(n2959), .C(n2958), .ZN(
        n2963) );
  NR2D1BWP12T U3292 ( .A1(n2961), .A2(n3071), .ZN(n2962) );
  AOI211D1BWP12T U3293 ( .A1(n2964), .A2(n3096), .B(n2963), .C(n2962), .ZN(
        n2965) );
  OAI211D1BWP12T U3294 ( .A1(n2968), .A2(n2967), .B(n2966), .C(n2965), .ZN(
        n2969) );
  AOI21D1BWP12T U3295 ( .A1(n3076), .A2(n2970), .B(n2969), .ZN(n2973) );
  CKND2D1BWP12T U3296 ( .A1(n2971), .A2(n382), .ZN(n2972) );
  OAI211D1BWP12T U3297 ( .A1(n2975), .A2(n2974), .B(n2973), .C(n2972), .ZN(
        result[20]) );
  INVD1BWP12T U3298 ( .I(n2984), .ZN(n3011) );
  INVD0BWP12T U3299 ( .I(n2985), .ZN(n2987) );
  AOI21D1BWP12T U3300 ( .A1(n2988), .A2(n2987), .B(n2986), .ZN(n3005) );
  ND2D1BWP12T U3301 ( .A1(n2989), .A2(n3096), .ZN(n3003) );
  MOAI22D0BWP12T U3302 ( .A1(n2992), .A2(n2991), .B1(n2990), .B2(n3067), .ZN(
        n2999) );
  MUX2ND0BWP12T U3303 ( .I0(n3019), .I1(n3018), .S(b[30]), .ZN(n2993) );
  NR2D0BWP12T U3304 ( .A1(n2993), .A2(n3020), .ZN(n2997) );
  OAI21D0BWP12T U3305 ( .A1(a[30]), .A2(n3099), .B(n3103), .ZN(n2994) );
  AOI22D0BWP12T U3306 ( .A1(n3105), .A2(n2996), .B1(n2994), .B2(b[30]), .ZN(
        n2995) );
  OAI211D1BWP12T U3307 ( .A1(n2997), .A2(n2996), .B(n3028), .C(n2995), .ZN(
        n2998) );
  RCAOI211D0BWP12T U3308 ( .A1(n3001), .A2(n3000), .B(n2999), .C(n2998), .ZN(
        n3002) );
  OAI211D1BWP12T U3309 ( .A1(n3005), .A2(n3004), .B(n3003), .C(n3002), .ZN(
        n3006) );
  TPAOI21D1BWP12T U3310 ( .A1(n3007), .A2(n3093), .B(n3006), .ZN(n3010) );
  CKND2D1BWP12T U3311 ( .A1(n3008), .A2(n3082), .ZN(n3009) );
  OAI211D1BWP12T U3312 ( .A1(n3047), .A2(n3011), .B(n3010), .C(n3009), .ZN(
        n3012) );
  TPAOI21D1BWP12T U3313 ( .A1(n3076), .A2(n3013), .B(n3012), .ZN(n3014) );
  IOA21D1BWP12T U3314 ( .A1(n3015), .A2(n3117), .B(n3014), .ZN(result[30]) );
  INVD1BWP12T U3315 ( .I(n3016), .ZN(n3046) );
  INVD1BWP12T U3316 ( .I(n3017), .ZN(n3039) );
  OAI21D0BWP12T U3317 ( .A1(a[22]), .A2(n3099), .B(n3103), .ZN(n3026) );
  MUX2ND0BWP12T U3318 ( .I0(n3019), .I1(n3018), .S(b[22]), .ZN(n3021) );
  NR2D0BWP12T U3319 ( .A1(n3021), .A2(n3020), .ZN(n3024) );
  MUX2ND0BWP12T U3320 ( .I0(n3024), .I1(n3023), .S(n3022), .ZN(n3025) );
  AOI21D0BWP12T U3321 ( .A1(b[22]), .A2(n3026), .B(n3025), .ZN(n3027) );
  OAI211D0BWP12T U3322 ( .A1(n3030), .A2(n3029), .B(n3028), .C(n3027), .ZN(
        n3034) );
  NR2D1BWP12T U3323 ( .A1(n3032), .A2(n3031), .ZN(n3033) );
  AOI211XD0BWP12T U3324 ( .A1(n3067), .A2(n3035), .B(n3034), .C(n3033), .ZN(
        n3038) );
  ND2XD0BWP12T U3325 ( .A1(n3036), .A2(n3091), .ZN(n3037) );
  OAI211D1BWP12T U3326 ( .A1(n3040), .A2(n3039), .B(n3038), .C(n3037), .ZN(
        n3041) );
  TPAOI21D0BWP12T U3327 ( .A1(n3042), .A2(n3093), .B(n3041), .ZN(n3045) );
  CKND2D1BWP12T U3328 ( .A1(n3043), .A2(n3082), .ZN(n3044) );
  OAI211D1BWP12T U3329 ( .A1(n3047), .A2(n3046), .B(n3045), .C(n3044), .ZN(
        n3048) );
  AOI21D1BWP12T U3330 ( .A1(n3076), .A2(n3049), .B(n3048), .ZN(n3050) );
  IOA21D1BWP12T U3331 ( .A1(n3051), .A2(n3117), .B(n3050), .ZN(result[22]) );
  AOI22D0BWP12T U3332 ( .A1(n3053), .A2(n3082), .B1(n3091), .B2(n3052), .ZN(
        n3054) );
  IOA21D1BWP12T U3333 ( .A1(n3055), .A2(n382), .B(n3054), .ZN(n3074) );
  AOI22D0BWP12T U3334 ( .A1(n3096), .A2(n3057), .B1(n3056), .B2(n3093), .ZN(
        n3070) );
  MUX2ND0BWP12T U3335 ( .I0(n3102), .I1(n3101), .S(b[13]), .ZN(n3058) );
  CKND2D0BWP12T U3336 ( .A1(n3058), .A2(n3103), .ZN(n3060) );
  MUX2ND0BWP12T U3337 ( .I0(n3060), .I1(n3105), .S(n3059), .ZN(n3063) );
  OAI21D0BWP12T U3338 ( .A1(a[13]), .A2(n3099), .B(n3103), .ZN(n3061) );
  ND2XD0BWP12T U3339 ( .A1(n3061), .A2(b[13]), .ZN(n3062) );
  OAI211D1BWP12T U3340 ( .A1(n3065), .A2(n3064), .B(n3063), .C(n3062), .ZN(
        n3066) );
  AOI21D1BWP12T U3341 ( .A1(n3068), .A2(n3067), .B(n3066), .ZN(n3069) );
  OAI211D1BWP12T U3342 ( .A1(n3072), .A2(n3071), .B(n3070), .C(n3069), .ZN(
        n3073) );
  RCAOI211D0BWP12T U3343 ( .A1(n3076), .A2(n3075), .B(n3074), .C(n3073), .ZN(
        n3077) );
  INVD1BWP12T U3344 ( .I(n3079), .ZN(n3088) );
  AOI22D0BWP12T U3345 ( .A1(n3083), .A2(n3082), .B1(n3081), .B2(n3080), .ZN(
        n3087) );
  ND2XD0BWP12T U3346 ( .A1(n3085), .A2(n3084), .ZN(n3086) );
  OAI211D1BWP12T U3347 ( .A1(n3089), .A2(n3088), .B(n3087), .C(n3086), .ZN(
        n3114) );
  AOI21D0BWP12T U3348 ( .A1(n3092), .A2(n3091), .B(n3090), .ZN(n3111) );
  AOI22D0BWP12T U3349 ( .A1(n3096), .A2(n3095), .B1(n3094), .B2(n3093), .ZN(
        n3110) );
  OAI211D1BWP12T U3350 ( .A1(n3112), .A2(n3111), .B(n3110), .C(n3109), .ZN(
        n3113) );
  RCAOI211D0BWP12T U3351 ( .A1(n382), .A2(n3115), .B(n3114), .C(n3113), .ZN(
        n3116) );
  IOA21D1BWP12T U3352 ( .A1(n3118), .A2(n3117), .B(n3116), .ZN(result[10]) );
  CMPE42D1BWP12T U3353 ( .A(mult_x_18_n601), .B(mult_x_18_n955), .C(
        mult_x_18_n605), .CIX(mult_x_18_n596), .D(mult_x_18_n599), .CO(
        mult_x_18_n592), .COX(mult_x_18_n591), .S(mult_x_18_n593) );
  CMPE42D1BWP12T U3354 ( .A(mult_x_18_n499), .B(mult_x_18_n477), .C(
        mult_x_18_n496), .CIX(mult_x_18_n489), .D(mult_x_18_n493), .CO(
        mult_x_18_n470), .COX(mult_x_18_n469), .S(mult_x_18_n471) );
  CMPE42D1BWP12T U3355 ( .A(mult_x_18_n738), .B(mult_x_18_n809), .C(
        mult_x_18_n625), .CIX(mult_x_18_n613), .D(mult_x_18_n626), .CO(
        mult_x_18_n606), .COX(mult_x_18_n605), .S(mult_x_18_n607) );
  CMPE42D1BWP12T U3356 ( .A(mult_x_18_n857), .B(mult_x_18_n821), .C(
        mult_x_18_n926), .CIX(mult_x_18_n578), .D(mult_x_18_n982), .CO(
        mult_x_18_n567), .COX(mult_x_18_n566), .S(mult_x_18_n568) );
  CMPE42D1BWP12T U3357 ( .A(mult_x_18_n571), .B(mult_x_18_n793), .C(
        mult_x_18_n568), .CIX(mult_x_18_n582), .D(mult_x_18_n565), .CO(
        mult_x_18_n561), .COX(mult_x_18_n560), .S(mult_x_18_n562) );
  CMPE42D1BWP12T U3358 ( .A(mult_x_18_n514), .B(mult_x_18_n500), .C(
        mult_x_18_n517), .CIX(mult_x_18_n507), .D(mult_x_18_n494), .CO(
        mult_x_18_n490), .COX(mult_x_18_n489), .S(mult_x_18_n491) );
  CMPE42D1BWP12T U3359 ( .A(mult_x_18_n862), .B(mult_x_18_n843), .C(
        mult_x_18_n650), .CIX(mult_x_18_n647), .D(mult_x_18_n638), .CO(
        mult_x_18_n632), .COX(mult_x_18_n631), .S(mult_x_18_n633) );
  CMPE42D1BWP12T U3360 ( .A(mult_x_18_n800), .B(mult_x_18_n776), .C(
        mult_x_18_n832), .CIX(mult_x_18_n478), .D(mult_x_18_n851), .CO(
        mult_x_18_n459), .COX(mult_x_18_n458), .S(mult_x_18_n460) );
  CMPE42D1BWP12T U3361 ( .A(mult_x_18_n791), .B(mult_x_18_n876), .C(
        mult_x_18_n951), .CIX(mult_x_18_n552), .D(mult_x_18_n539), .CO(
        mult_x_18_n530), .COX(mult_x_18_n529), .S(mult_x_18_n531) );
  CMPE42D1BWP12T U3362 ( .A(mult_x_18_n898), .B(mult_x_18_n770), .C(
        mult_x_18_n923), .CIX(mult_x_18_n529), .D(mult_x_18_n522), .CO(
        mult_x_18_n517), .COX(mult_x_18_n516), .S(mult_x_18_n518) );
  CMPE42D1BWP12T U3363 ( .A(mult_x_18_n949), .B(mult_x_18_n778), .C(
        mult_x_18_n802), .CIX(mult_x_18_n513), .D(mult_x_18_n834), .CO(
        mult_x_18_n496), .COX(mult_x_18_n495), .S(mult_x_18_n497) );
  CMPE42D1BWP12T U3364 ( .A(mult_x_18_n907), .B(mult_x_18_n884), .C(
        mult_x_18_n932), .CIX(mult_x_18_n655), .D(mult_x_18_n661), .CO(
        mult_x_18_n648), .COX(mult_x_18_n647), .S(mult_x_18_n649) );
  CMPE42D1BWP12T U3365 ( .A(mult_x_18_n921), .B(mult_x_18_n777), .C(
        mult_x_18_n977), .CIX(mult_x_18_n492), .D(mult_x_18_n485), .CO(
        mult_x_18_n482), .COX(mult_x_18_n481), .S(mult_x_18_n483) );
  CMPE42D1BWP12T U3366 ( .A(mult_x_18_n804), .B(mult_x_18_n780), .C(
        mult_x_18_n836), .CIX(mult_x_18_n549), .D(mult_x_18_n855), .CO(
        mult_x_18_n533), .COX(mult_x_18_n532), .S(mult_x_18_n534) );
  CMPE42D1BWP12T U3367 ( .A(mult_x_18_n394), .B(mult_x_18_n397), .C(
        mult_x_18_n391), .CIX(mult_x_18_n406), .D(mult_x_18_n419), .CO(
        mult_x_18_n384), .COX(mult_x_18_n383), .S(mult_x_18_n385) );
  CMPE42D1BWP12T U3368 ( .A(mult_x_18_n437), .B(mult_x_18_n440), .C(
        mult_x_18_n434), .CIX(mult_x_18_n427), .D(mult_x_18_n430), .CO(
        mult_x_18_n407), .COX(mult_x_18_n406), .S(mult_x_18_n408) );
  CMPE42D1BWP12T U3369 ( .A(mult_x_18_n482), .B(mult_x_18_n457), .C(
        mult_x_18_n476), .CIX(mult_x_18_n454), .D(mult_x_18_n479), .CO(
        mult_x_18_n450), .COX(mult_x_18_n449), .S(mult_x_18_n451) );
  CMPE42D1BWP12T U3370 ( .A(mult_x_18_n462), .B(mult_x_18_n435), .C(
        mult_x_18_n459), .CIX(mult_x_18_n453), .D(mult_x_18_n452), .CO(
        mult_x_18_n428), .COX(mult_x_18_n427), .S(mult_x_18_n429) );
  CMPE42D1BWP12T U3371 ( .A(mult_x_18_n533), .B(mult_x_18_n515), .C(
        mult_x_18_n530), .CIX(mult_x_18_n526), .D(mult_x_18_n512), .CO(
        mult_x_18_n508), .COX(mult_x_18_n507), .S(mult_x_18_n509) );
  CMPE42D1BWP12T U3372 ( .A(mult_x_18_n894), .B(mult_x_18_n814), .C(
        mult_x_18_n919), .CIX(mult_x_18_n455), .D(mult_x_18_n445), .CO(
        mult_x_18_n440), .COX(mult_x_18_n439), .S(mult_x_18_n441) );
  CMPE42D1BWP12T U3373 ( .A(mult_x_18_n902), .B(mult_x_18_n794), .C(
        mult_x_18_n927), .CIX(mult_x_18_n594), .D(mult_x_18_n587), .CO(
        mult_x_18_n582), .COX(mult_x_18_n581), .S(mult_x_18_n583) );
  CMPE42D1BWP12T U3374 ( .A(mult_x_18_n757), .B(mult_x_18_n773), .C(
        mult_x_18_n869), .CIX(mult_x_18_n421), .D(mult_x_18_n764), .CO(
        mult_x_18_n390), .COX(mult_x_18_n389), .S(mult_x_18_n391) );
  CMPE42D1BWP12T U3375 ( .A(mult_x_18_n740), .B(mult_x_18_n845), .C(
        mult_x_18_n864), .CIX(mult_x_18_n669), .D(mult_x_18_n908), .CO(
        mult_x_18_n656), .COX(mult_x_18_n655), .S(mult_x_18_n657) );
  CMPE42D1BWP12T U3376 ( .A(mult_x_18_n849), .B(mult_x_18_n753), .C(
        mult_x_18_n893), .CIX(mult_x_18_n433), .D(mult_x_18_n918), .CO(
        mult_x_18_n419), .COX(mult_x_18_n418), .S(mult_x_18_n420) );
  CMPE42D1BWP12T U3377 ( .A(mult_x_18_n929), .B(mult_x_18_n881), .C(
        mult_x_18_n985), .CIX(mult_x_18_n619), .D(mult_x_18_n615), .CO(
        mult_x_18_n612), .COX(mult_x_18_n611), .S(mult_x_18_n613) );
  CMPE42D1BWP12T U3378 ( .A(mult_x_18_n465), .B(mult_x_18_n872), .C(
        mult_x_18_n472), .CIX(mult_x_18_n460), .D(mult_x_18_n463), .CO(
        mult_x_18_n453), .COX(mult_x_18_n452), .S(mult_x_18_n454) );
  CMPE42D1BWP12T U3379 ( .A(mult_x_18_n1009), .B(mult_x_18_n762), .C(
        mult_x_18_n978), .CIX(mult_x_18_n519), .D(mult_x_18_n521), .CO(
        mult_x_18_n502), .COX(mult_x_18_n501), .S(mult_x_18_n503) );
  CMPE42D1BWP12T U3380 ( .A(mult_x_18_n1017), .B(mult_x_18_n810), .C(
        mult_x_18_n986), .CIX(mult_x_18_n637), .D(mult_x_18_n639), .CO(
        mult_x_18_n626), .COX(mult_x_18_n625), .S(mult_x_18_n627) );
  CMPE42D1BWP12T U3381 ( .A(mult_x_18_n585), .B(mult_x_18_n600), .C(
        mult_x_18_n583), .CIX(mult_x_18_n591), .D(mult_x_18_n580), .CO(
        mult_x_18_n576), .COX(mult_x_18_n575), .S(mult_x_18_n577) );
  CMPE42D1BWP12T U3382 ( .A(mult_x_18_n550), .B(mult_x_18_n537), .C(
        mult_x_18_n547), .CIX(mult_x_18_n543), .D(mult_x_18_n531), .CO(
        mult_x_18_n527), .COX(mult_x_18_n526), .S(mult_x_18_n528) );
  CMPE42D1BWP12T U3383 ( .A(mult_x_18_n1025), .B(mult_x_18_n890), .C(
        mult_x_18_n913), .CIX(mult_x_18_n707), .D(mult_x_18_n709), .CO(
        mult_x_18_n702), .COX(mult_x_18_n701), .S(mult_x_18_n703) );
  CMPE42D1BWP12T U3384 ( .A(mult_x_18_n833), .B(mult_x_18_n761), .C(
        mult_x_18_n852), .CIX(mult_x_18_n495), .D(mult_x_18_n896), .CO(
        mult_x_18_n479), .COX(mult_x_18_n478), .S(mult_x_18_n480) );
  CMPE42D1BWP12T U3385 ( .A(mult_x_18_n925), .B(mult_x_18_n736), .C(
        mult_x_18_n981), .CIX(mult_x_18_n563), .D(mult_x_18_n556), .CO(
        mult_x_18_n553), .COX(mult_x_18_n552), .S(mult_x_18_n554) );
  CMPE42D1BWP12T U3386 ( .A(mult_x_18_n937), .B(mult_x_18_n889), .C(
        mult_x_18_n993), .CIX(mult_x_18_n698), .D(mult_x_18_n697), .CO(
        mult_x_18_n694), .COX(mult_x_18_n693), .S(mult_x_18_n695) );
  CMPE42D1BWP12T U3387 ( .A(mult_x_18_n768), .B(mult_x_18_n873), .C(
        mult_x_18_n501), .CIX(mult_x_18_n483), .D(mult_x_18_n502), .CO(
        mult_x_18_n473), .COX(mult_x_18_n472), .S(mult_x_18_n474) );
  CMPE42D1BWP12T U3388 ( .A(mult_x_18_n910), .B(mult_x_18_n866), .C(
        mult_x_18_n935), .CIX(mult_x_18_n685), .D(mult_x_18_n681), .CO(
        mult_x_18_n676), .COX(mult_x_18_n675), .S(mult_x_18_n677) );
  CMPE42D1BWP12T U3389 ( .A(mult_x_18_n870), .B(mult_x_18_n774), .C(
        mult_x_18_n765), .CIX(mult_x_18_n439), .D(mult_x_18_n785), .CO(
        mult_x_18_n413), .COX(mult_x_18_n412), .S(mult_x_18_n414) );
  CMPE42D1BWP12T U3390 ( .A(mult_x_18_n957), .B(mult_x_18_n882), .C(
        mult_x_18_n842), .CIX(mult_x_18_n627), .D(mult_x_18_n631), .CO(
        mult_x_18_n620), .COX(mult_x_18_n619), .S(mult_x_18_n621) );
  CMPE42D1BWP12T U3391 ( .A(mult_x_18_n808), .B(mult_x_18_n880), .C(
        mult_x_18_n840), .CIX(mult_x_18_n611), .D(mult_x_18_n859), .CO(
        mult_x_18_n595), .COX(mult_x_18_n594), .S(mult_x_18_n596) );
  CMPE42D1BWP12T U3392 ( .A(mult_x_18_n792), .B(mult_x_18_n877), .C(
        mult_x_18_n952), .CIX(mult_x_18_n569), .D(mult_x_18_n805), .CO(
        mult_x_18_n547), .COX(mult_x_18_n546), .S(mult_x_18_n548) );
  CMPE42D1BWP12T U3393 ( .A(mult_x_18_n844), .B(mult_x_18_n959), .C(
        mult_x_18_n863), .CIX(mult_x_18_n658), .D(mult_x_18_n651), .CO(
        mult_x_18_n645), .COX(mult_x_18_n644), .S(mult_x_18_n646) );
  CMPE42D1BWP12T U3394 ( .A(mult_x_18_n807), .B(mult_x_18_n954), .C(
        mult_x_18_n839), .CIX(mult_x_18_n597), .D(mult_x_18_n858), .CO(
        mult_x_18_n579), .COX(mult_x_18_n578), .S(mult_x_18_n580) );
  CMPE42D1BWP12T U3395 ( .A(mult_x_18_n400), .B(mult_x_18_n422), .C(
        mult_x_18_n416), .CIX(mult_x_18_n409), .D(mult_x_18_n413), .CO(
        mult_x_18_n387), .COX(mult_x_18_n386), .S(mult_x_18_n388) );
  CMPE42D1BWP12T U3396 ( .A(mult_x_18_n443), .B(mult_x_18_n464), .C(
        mult_x_18_n441), .CIX(mult_x_18_n456), .D(mult_x_18_n438), .CO(
        mult_x_18_n431), .COX(mult_x_18_n430), .S(mult_x_18_n432) );
  CMPE42D1BWP12T U3397 ( .A(mult_x_18_n892), .B(mult_x_18_n749), .C(
        mult_x_18_n973), .CIX(mult_x_18_n412), .D(mult_x_18_n402), .CO(
        mult_x_18_n399), .COX(mult_x_18_n398), .S(mult_x_18_n400) );
  CMPE42D1BWP12T U3398 ( .A(mult_x_18_n1005), .B(mult_x_18_n750), .C(
        mult_x_18_n974), .CIX(mult_x_18_n442), .D(mult_x_18_n444), .CO(
        mult_x_18_n422), .COX(mult_x_18_n421), .S(mult_x_18_n423) );
  CMPE42D1BWP12T U3399 ( .A(mult_x_18_n784), .B(mult_x_18_n812), .C(
        mult_x_18_n944), .CIX(mult_x_18_n418), .D(mult_x_18_n797), .CO(
        mult_x_18_n393), .COX(mult_x_18_n392), .S(mult_x_18_n394) );
  CMPE42D1BWP12T U3400 ( .A(mult_x_18_n423), .B(mult_x_18_n758), .C(
        mult_x_18_n420), .CIX(mult_x_18_n414), .D(mult_x_18_n417), .CO(
        mult_x_18_n410), .COX(mult_x_18_n409), .S(mult_x_18_n411) );
  CMPE42D1BWP12T U3401 ( .A(mult_x_18_n899), .B(mult_x_18_n819), .C(
        mult_x_18_n924), .CIX(mult_x_18_n546), .D(mult_x_18_n555), .CO(
        mult_x_18_n536), .COX(mult_x_18_n535), .S(mult_x_18_n537) );
  CMPE42D1BWP12T U3402 ( .A(mult_x_18_n829), .B(mult_x_18_n752), .C(
        mult_x_18_n848), .CIX(mult_x_18_n415), .D(mult_x_18_n917), .CO(
        mult_x_18_n396), .COX(mult_x_18_n395), .S(mult_x_18_n397) );
  CMPE42D1BWP12T U3403 ( .A(mult_x_18_n841), .B(mult_x_18_n956), .C(
        mult_x_18_n860), .CIX(mult_x_18_n622), .D(mult_x_18_n904), .CO(
        mult_x_18_n609), .COX(mult_x_18_n608), .S(mult_x_18_n610) );
  CMPE42D1BWP12T U3404 ( .A(mult_x_18_n766), .B(mult_x_18_n871), .C(
        mult_x_18_n786), .CIX(mult_x_18_n461), .D(mult_x_18_n946), .CO(
        mult_x_18_n434), .COX(mult_x_18_n433), .S(mult_x_18_n435) );
  CMPE42D1BWP12T U3405 ( .A(mult_x_18_n767), .B(mult_x_18_n760), .C(
        mult_x_18_n787), .CIX(mult_x_18_n481), .D(mult_x_18_n947), .CO(
        mult_x_18_n456), .COX(mult_x_18_n455), .S(mult_x_18_n457) );
  CMPE42D1BWP12T U3406 ( .A(mult_x_18_n803), .B(mult_x_18_n735), .C(
        mult_x_18_n835), .CIX(mult_x_18_n532), .D(mult_x_18_n854), .CO(
        mult_x_18_n514), .COX(mult_x_18_n513), .S(mult_x_18_n515) );
  CMPE42D1BWP12T U3407 ( .A(mult_x_18_n853), .B(mult_x_18_n817), .C(
        mult_x_18_n897), .CIX(mult_x_18_n516), .D(mult_x_18_n922), .CO(
        mult_x_18_n499), .COX(mult_x_18_n498), .S(mult_x_18_n500) );
  CMPE42D1BWP12T U3408 ( .A(mult_x_18_n861), .B(mult_x_18_n825), .C(
        mult_x_18_n905), .CIX(mult_x_18_n634), .D(mult_x_18_n930), .CO(
        mult_x_18_n623), .COX(mult_x_18_n622), .S(mult_x_18_n624) );
  CMPE42D1BWP12T U3409 ( .A(mult_x_18_n788), .B(mult_x_18_n734), .C(
        mult_x_18_n948), .CIX(mult_x_18_n498), .D(mult_x_18_n801), .CO(
        mult_x_18_n476), .COX(mult_x_18_n475), .S(mult_x_18_n477) );
  CMPE42D1BWP12T U3410 ( .A(mult_x_18_n388), .B(mult_x_18_n410), .C(
        mult_x_18_n385), .CIX(mult_x_18_n403), .D(mult_x_18_n407), .CO(
        mult_x_18_n381), .COX(mult_x_18_n380), .S(mult_x_18_n382) );
  CMPE42D1BWP12T U3411 ( .A(mult_x_18_n431), .B(mult_x_18_n411), .C(
        mult_x_18_n408), .CIX(mult_x_18_n424), .D(mult_x_18_n428), .CO(
        mult_x_18_n404), .COX(mult_x_18_n403), .S(mult_x_18_n405) );
  CMPE42D1BWP12T U3412 ( .A(mult_x_18_n903), .B(mult_x_18_n823), .C(
        mult_x_18_n928), .CIX(mult_x_18_n608), .D(mult_x_18_n614), .CO(
        mult_x_18_n598), .COX(mult_x_18_n597), .S(mult_x_18_n599) );
  CMPE42D1BWP12T U3413 ( .A(mult_x_18_n769), .B(mult_x_18_n874), .C(
        mult_x_18_n789), .CIX(mult_x_18_n503), .D(mult_x_18_n510), .CO(
        mult_x_18_n493), .COX(mult_x_18_n492), .S(mult_x_18_n494) );
  CMPE42D1BWP12T U3414 ( .A(mult_x_18_n953), .B(mult_x_18_n878), .C(
        mult_x_18_n806), .CIX(mult_x_18_n581), .D(mult_x_18_n838), .CO(
        mult_x_18_n564), .COX(mult_x_18_n563), .S(mult_x_18_n565) );
  CMPE42D1BWP12T U3415 ( .A(mult_x_18_n945), .B(mult_x_18_n813), .C(
        mult_x_18_n798), .CIX(mult_x_18_n436), .D(mult_x_18_n830), .CO(
        mult_x_18_n416), .COX(mult_x_18_n415), .S(mult_x_18_n417) );
  CMPE42D1BWP12T U3416 ( .A(mult_x_18_n799), .B(mult_x_18_n759), .C(
        mult_x_18_n831), .CIX(mult_x_18_n458), .D(mult_x_18_n850), .CO(
        mult_x_18_n437), .COX(mult_x_18_n436), .S(mult_x_18_n438) );
  CMPE42D1BWP12T U3417 ( .A(mult_x_18_n895), .B(mult_x_18_n815), .C(
        mult_x_18_n920), .CIX(mult_x_18_n475), .D(mult_x_18_n484), .CO(
        mult_x_18_n462), .COX(mult_x_18_n461), .S(mult_x_18_n463) );
  CMPE42D1BWP12T U3418 ( .A(mult_x_18_n950), .B(mult_x_18_n790), .C(
        mult_x_18_n538), .CIX(mult_x_18_n535), .D(mult_x_18_n520), .CO(
        mult_x_18_n511), .COX(mult_x_18_n510), .S(mult_x_18_n512) );
  CMPE42D1BWP12T U3419 ( .A(mult_x_18_n595), .B(mult_x_18_n598), .C(
        mult_x_18_n592), .CIX(mult_x_18_n577), .D(mult_x_18_n588), .CO(
        mult_x_18_n573), .COX(mult_x_18_n572), .S(mult_x_18_n574) );
  CMPE42D1BWP12T U3420 ( .A(mult_x_18_n511), .B(mult_x_18_n497), .C(
        mult_x_18_n491), .CIX(mult_x_18_n504), .D(mult_x_18_n508), .CO(
        mult_x_18_n487), .COX(mult_x_18_n486), .S(mult_x_18_n488) );
  CMPE42D1BWP12T U3421 ( .A(mult_x_18_n744), .B(mult_x_18_n941), .C(
        mult_x_18_n997), .CIX(mult_x_18_n721), .D(mult_x_18_n720), .CO(
        mult_x_18_n717), .COX(mult_x_18_n716), .S(mult_x_18_n718) );
  CMPE42D1BWP12T U3422 ( .A(mult_x_18_n912), .B(mult_x_18_n964), .C(
        mult_x_18_n701), .CIX(mult_x_18_n695), .D(mult_x_18_n702), .CO(
        mult_x_18_n691), .COX(mult_x_18_n690), .S(mult_x_18_n692) );
  CMPE42D1BWP12T U3423 ( .A(mult_x_18_n623), .B(mult_x_18_n610), .C(
        mult_x_18_n620), .CIX(mult_x_18_n616), .D(mult_x_18_n607), .CO(
        mult_x_18_n603), .COX(mult_x_18_n602), .S(mult_x_18_n604) );
  CMPE42D1BWP12T U3424 ( .A(mult_x_18_n609), .B(mult_x_18_n612), .C(
        mult_x_18_n606), .CIX(mult_x_18_n593), .D(mult_x_18_n602), .CO(
        mult_x_18_n589), .COX(mult_x_18_n588), .S(mult_x_18_n590) );
  CMPE42D1BWP12T U3425 ( .A(mult_x_18_n536), .B(mult_x_18_n518), .C(
        mult_x_18_n509), .CIX(mult_x_18_n523), .D(mult_x_18_n527), .CO(
        mult_x_18_n505), .COX(mult_x_18_n504), .S(mult_x_18_n506) );
  CMPE42D1BWP12T U3426 ( .A(mult_x_18_n432), .B(mult_x_18_n449), .C(
        mult_x_18_n429), .CIX(mult_x_18_n446), .D(mult_x_18_n450), .CO(
        mult_x_18_n425), .COX(mult_x_18_n424), .S(mult_x_18_n426) );
  CMPE42D1BWP12T U3427 ( .A(mult_x_18_n553), .B(mult_x_18_n534), .C(
        mult_x_18_n544), .CIX(mult_x_18_n540), .D(mult_x_18_n528), .CO(
        mult_x_18_n524), .COX(mult_x_18_n523), .S(mult_x_18_n525) );
  CMPE42D1BWP12T U3428 ( .A(mult_x_18_n469), .B(mult_x_18_n473), .C(
        mult_x_18_n451), .CIX(mult_x_18_n466), .D(mult_x_18_n470), .CO(
        mult_x_18_n447), .COX(mult_x_18_n446), .S(mult_x_18_n448) );
endmodule


module top7 ( clk, reset, MEM_MEMCTRL_from_mem_data, 
        MEMCTRL_MEM_to_mem_read_enable, MEMCTRL_MEM_to_mem_write_enable, 
        MEMCTRL_MEM_to_mem_mem_enable, MEMCTRL_MEM_to_mem_address, 
        MEMCTRL_MEM_to_mem_data );
  input [15:0] MEM_MEMCTRL_from_mem_data;
  output [11:0] MEMCTRL_MEM_to_mem_address;
  output [15:0] MEMCTRL_MEM_to_mem_data;
  input clk, reset;
  output MEMCTRL_MEM_to_mem_read_enable, MEMCTRL_MEM_to_mem_write_enable,
         MEMCTRL_MEM_to_mem_mem_enable;
  wire   DEC_CPSR_update_flag_n, new_n, ALU_OUT_n, RF_OUT_n,
         DEC_CPSR_update_flag_c, new_c, ALU_OUT_c, RF_OUT_c,
         DEC_CPSR_update_flag_z, new_z, ALU_OUT_z, RF_OUT_z,
         DEC_CPSR_update_flag_v, new_v, ALU_OUT_v, RF_OUT_v,
         DEC_RF_alu_write_to_reg_enable, DEC_RF_memory_write_to_reg_enable,
         DEC_MISC_OUT_memory_address_source_is_reg,
         DEC_MEMCTRL_memorycontroller_sign_extend,
         DEC_MEMCTRL_memory_load_request, DEC_MEMCTRL_memory_store_request,
         DEC_IF_stall_to_instructionfetch, ALU_IN_c, irdecode_inst1_N912,
         irdecode_inst1_N911, irdecode_inst1_N910, irdecode_inst1_N907,
         irdecode_inst1_N906, irdecode_inst1_N707, irdecode_inst1_N706,
         irdecode_inst1_N705, irdecode_inst1_N704, irdecode_inst1_N703,
         irdecode_inst1_N702, irdecode_inst1_N701, irdecode_inst1_N546,
         irdecode_inst1_N545, irdecode_inst1_N544, irdecode_inst1_N543,
         irdecode_inst1_N542, irdecode_inst1_N541, irdecode_inst1_N540,
         irdecode_inst1_N539, irdecode_inst1_split_instruction,
         irdecode_inst1_next_step_0_, irdecode_inst1_next_step_1_,
         irdecode_inst1_next_step_2_, irdecode_inst1_next_step_3_,
         irdecode_inst1_next_step_4_, irdecode_inst1_next_step_5_,
         irdecode_inst1_next_step_6_, irdecode_inst1_next_step_7_,
         irdecode_inst1_itstate_0_, irdecode_inst1_itstate_1_,
         irdecode_inst1_itstate_2_, irdecode_inst1_itstate_3_,
         irdecode_inst1_itstate_4_, irdecode_inst1_itstate_5_,
         irdecode_inst1_itstate_6_, irdecode_inst1_itstate_7_,
         irdecode_inst1_next_alu_write_to_reg_enable,
         irdecode_inst1_next_update_flag_v, irdecode_inst1_next_update_flag_c,
         irdecode_inst1_next_update_flag_n,
         memory_interface_inst1_delayed_is_signed, Instruction_Fetch_inst1_N98,
         Instruction_Fetch_inst1_N97, Instruction_Fetch_inst1_N96,
         Instruction_Fetch_inst1_N95, Instruction_Fetch_inst1_N94,
         Instruction_Fetch_inst1_N93, Instruction_Fetch_inst1_N92,
         Instruction_Fetch_inst1_N91, Instruction_Fetch_inst1_N90,
         Instruction_Fetch_inst1_N89, Instruction_Fetch_inst1_N88,
         Instruction_Fetch_inst1_N87, Instruction_Fetch_inst1_N86,
         Instruction_Fetch_inst1_N85, Instruction_Fetch_inst1_N84,
         Instruction_Fetch_inst1_N83, Instruction_Fetch_inst1_N80,
         Instruction_Fetch_inst1_N79,
         Instruction_Fetch_inst1_first_instruction_fetched,
         Instruction_Fetch_inst1_fetched_instruction_reg_0_,
         Instruction_Fetch_inst1_fetched_instruction_reg_1_,
         Instruction_Fetch_inst1_fetched_instruction_reg_2_,
         Instruction_Fetch_inst1_fetched_instruction_reg_3_,
         Instruction_Fetch_inst1_fetched_instruction_reg_4_,
         Instruction_Fetch_inst1_fetched_instruction_reg_5_,
         Instruction_Fetch_inst1_fetched_instruction_reg_6_,
         Instruction_Fetch_inst1_fetched_instruction_reg_7_,
         Instruction_Fetch_inst1_fetched_instruction_reg_8_,
         Instruction_Fetch_inst1_fetched_instruction_reg_9_,
         Instruction_Fetch_inst1_fetched_instruction_reg_10_,
         Instruction_Fetch_inst1_fetched_instruction_reg_11_,
         Instruction_Fetch_inst1_fetched_instruction_reg_12_,
         Instruction_Fetch_inst1_fetched_instruction_reg_13_,
         Instruction_Fetch_inst1_fetched_instruction_reg_14_,
         Instruction_Fetch_inst1_fetched_instruction_reg_15_,
         Instruction_Fetch_inst1_currentState_0_,
         Instruction_Fetch_inst1_currentState_1_,
         memory_interface_inst1_fsm_N35, memory_interface_inst1_fsm_N34,
         memory_interface_inst1_fsm_N33, memory_interface_inst1_fsm_N32,
         memory_interface_inst1_fsm_state_0_,
         memory_interface_inst1_fsm_state_1_,
         memory_interface_inst1_fsm_state_2_,
         memory_interface_inst1_fsm_state_3_, n754, n777, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1684, n1685, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53;
  wire   [7:0] IF_DEC_instruction;
  wire   [4:0] DEC_RF_operand_a;
  wire   [4:0] DEC_RF_operand_b;
  wire   [31:0] DEC_RF_offset_b;
  wire   [4:0] DEC_ALU_alu_opcode;
  wire   [4:0] DEC_RF_alu_write_to_reg;
  wire   [4:0] DEC_RF_memory_write_to_reg;
  wire   [4:0] DEC_RF_memory_store_data_reg;
  wire   [4:0] DEC_RF_memory_store_address_reg;
  wire   [1:0] DEC_MEMCTRL_load_store_width;
  wire   [31:0] ALU_MISC_OUT_result;
  wire   [31:0] MEMCTRL_RF_IF_data_in;
  wire   [31:0] IF_RF_incremented_pc_out;
  wire   [31:0] RF_ALU_operand_a;
  wire   [31:0] RF_ALU_operand_b;
  wire   [31:0] RF_MEMCTRL_data_reg;
  wire   [12:2] RF_MEMCTRL_address_reg;
  wire   [31:0] RF_pc_out;
  wire   [11:0] MEMCTRL_IN_address;
  wire   [7:0] irdecode_inst1_step;
  wire   [15:0] memory_interface_inst1_delay_first_two_bytes_out;
  wire   [31:0] memory_interface_inst1_delay_data_in32;
  wire   [11:0] memory_interface_inst1_delay_addr_for_adder;

  register_file register_file_inst1 ( .readA_sel(DEC_RF_operand_a), 
        .readB_sel(DEC_RF_operand_b), .readC_sel(DEC_RF_memory_store_data_reg), 
        .readD_sel(DEC_RF_memory_store_address_reg), .write1_sel(
        DEC_RF_alu_write_to_reg), .write2_sel(DEC_RF_memory_write_to_reg), 
        .write1_en(DEC_RF_alu_write_to_reg_enable), .write2_en(
        DEC_RF_memory_write_to_reg_enable), .write1_in(ALU_MISC_OUT_result), 
        .write2_in(MEMCTRL_RF_IF_data_in), .immediate1_in({n864, n864, n864, 
        n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, 
        n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, 
        n864, n864, n864, n864, n864}), .immediate2_in(DEC_RF_offset_b), 
        .next_pc_in({IF_RF_incremented_pc_out[31:2], MEMCTRL_IN_address[0], 
        IF_RF_incremented_pc_out[0]}), .next_cpsr_in({new_n, new_c, new_z, 
        new_v}), .next_sp_in({n864, n864, n864, n864, n864, n864, n864, n864, 
        n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, 
        n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864}), .clk(clk), .reset(reset), .regA_out(RF_ALU_operand_a), .regB_out(
        RF_ALU_operand_b), .regC_out(RF_MEMCTRL_data_reg), .regD_out({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        RF_MEMCTRL_address_reg, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21}), .pc_out(RF_pc_out), .cpsr_out({RF_OUT_n, 
        RF_OUT_c, RF_OUT_z, RF_OUT_v}), .sp_out({SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53}), .next_pc_en_BAR(n754) );
  ALU_VARIABLE ALU_VARIABLE_inst1 ( .a({RF_ALU_operand_a[31:14], n1685, 
        RF_ALU_operand_a[12:0]}), .b(RF_ALU_operand_b), .op(
        DEC_ALU_alu_opcode[3:0]), .c_in(ALU_IN_c), .result(ALU_MISC_OUT_result), .c_out(ALU_OUT_c), .z(ALU_OUT_z), .n(ALU_OUT_n), .v(ALU_OUT_v) );
  CKAN2D2BWP12T irdecode_inst1_C5193 ( .A1(irdecode_inst1_next_step_7_), .A2(
        IF_DEC_instruction[7]), .Z(irdecode_inst1_N539) );
  CKAN2D2BWP12T irdecode_inst1_C5194 ( .A1(irdecode_inst1_next_step_6_), .A2(
        IF_DEC_instruction[6]), .Z(irdecode_inst1_N540) );
  CKAN2D2BWP12T irdecode_inst1_C5195 ( .A1(irdecode_inst1_next_step_5_), .A2(
        IF_DEC_instruction[5]), .Z(irdecode_inst1_N541) );
  CKAN2D2BWP12T irdecode_inst1_C5196 ( .A1(irdecode_inst1_next_step_4_), .A2(
        IF_DEC_instruction[4]), .Z(irdecode_inst1_N542) );
  CKAN2D2BWP12T irdecode_inst1_C5197 ( .A1(irdecode_inst1_next_step_3_), .A2(
        IF_DEC_instruction[3]), .Z(irdecode_inst1_N543) );
  CKAN2D2BWP12T irdecode_inst1_C5198 ( .A1(irdecode_inst1_next_step_2_), .A2(
        IF_DEC_instruction[2]), .Z(irdecode_inst1_N544) );
  CKAN2D2BWP12T irdecode_inst1_C5199 ( .A1(irdecode_inst1_next_step_1_), .A2(
        IF_DEC_instruction[1]), .Z(irdecode_inst1_N545) );
  CKAN2D2BWP12T irdecode_inst1_C5200 ( .A1(irdecode_inst1_next_step_0_), .A2(
        IF_DEC_instruction[0]), .Z(irdecode_inst1_N546) );
  CKAN2D2BWP12T irdecode_inst1_C5280 ( .A1(irdecode_inst1_next_step_6_), .A2(
        IF_DEC_instruction[6]), .Z(irdecode_inst1_N701) );
  CKAN2D2BWP12T irdecode_inst1_C5281 ( .A1(irdecode_inst1_next_step_5_), .A2(
        IF_DEC_instruction[5]), .Z(irdecode_inst1_N702) );
  CKAN2D2BWP12T irdecode_inst1_C5282 ( .A1(irdecode_inst1_next_step_4_), .A2(
        IF_DEC_instruction[4]), .Z(irdecode_inst1_N703) );
  CKAN2D2BWP12T irdecode_inst1_C5283 ( .A1(irdecode_inst1_next_step_3_), .A2(
        IF_DEC_instruction[3]), .Z(irdecode_inst1_N704) );
  CKAN2D2BWP12T irdecode_inst1_C5284 ( .A1(irdecode_inst1_next_step_2_), .A2(
        IF_DEC_instruction[2]), .Z(irdecode_inst1_N705) );
  CKAN2D2BWP12T irdecode_inst1_C5285 ( .A1(irdecode_inst1_next_step_1_), .A2(
        IF_DEC_instruction[1]), .Z(irdecode_inst1_N706) );
  CKAN2D2BWP12T irdecode_inst1_C5286 ( .A1(irdecode_inst1_next_step_0_), .A2(
        IF_DEC_instruction[0]), .Z(irdecode_inst1_N707) );
  CKAN2D2BWP12T irdecode_inst1_C2476 ( .A1(irdecode_inst1_next_step_1_), .A2(
        irdecode_inst1_next_step_0_), .Z(irdecode_inst1_N906) );
  CKAN2D2BWP12T irdecode_inst1_C2482 ( .A1(irdecode_inst1_N907), .A2(
        irdecode_inst1_N910), .Z(irdecode_inst1_N911) );
  OR2XD4BWP12T irdecode_inst1_C2484 ( .A1(irdecode_inst1_next_step_1_), .A2(
        irdecode_inst1_N910), .Z(irdecode_inst1_N912) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_0_ ( .D(
        MEM_MEMCTRL_from_mem_data[8]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[0]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_1_ ( .D(
        MEM_MEMCTRL_from_mem_data[9]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[1]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_2_ ( .D(
        MEM_MEMCTRL_from_mem_data[10]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_3_ ( .D(
        MEM_MEMCTRL_from_mem_data[11]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_4_ ( .D(
        MEM_MEMCTRL_from_mem_data[12]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[4]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_5_ ( .D(
        MEM_MEMCTRL_from_mem_data[13]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[5]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_6_ ( .D(
        MEM_MEMCTRL_from_mem_data[14]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_7_ ( .D(
        MEM_MEMCTRL_from_mem_data[15]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_8_ ( .D(
        MEM_MEMCTRL_from_mem_data[0]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_9_ ( .D(
        MEM_MEMCTRL_from_mem_data[1]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_10_ ( .D(
        MEM_MEMCTRL_from_mem_data[2]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_11_ ( .D(
        MEM_MEMCTRL_from_mem_data[3]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[11]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_12_ ( .D(
        MEM_MEMCTRL_from_mem_data[4]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[12]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_13_ ( .D(
        MEM_MEMCTRL_from_mem_data[5]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[13]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_14_ ( .D(
        MEM_MEMCTRL_from_mem_data[6]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[14]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_15_ ( .D(
        MEM_MEMCTRL_from_mem_data[7]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[15]) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_3_ ( .D(
        memory_interface_inst1_fsm_N35), .CP(clk), .Q(
        memory_interface_inst1_fsm_state_3_) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_31_ ( .D(n777), .CP(clk), .Q(
        DEC_RF_offset_b[31]) );
  DFQD1BWP12T irdecode_inst1_load_store_width_reg_0_ ( .D(n838), .CP(clk), .Q(
        DEC_MEMCTRL_load_store_width[0]) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_1_ ( .D(
        memory_interface_inst1_fsm_N33), .CP(clk), .Q(
        memory_interface_inst1_fsm_state_1_) );
  DFQD1BWP12T Instruction_Fetch_inst1_first_instruction_fetched_reg ( .D(n862), 
        .CP(clk), .Q(Instruction_Fetch_inst1_first_instruction_fetched) );
  DFQD1BWP12T irdecode_inst1_load_store_width_reg_1_ ( .D(n837), .CP(clk), .Q(
        DEC_MEMCTRL_load_store_width[1]) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_0_ ( .D(
        memory_interface_inst1_fsm_N32), .CP(clk), .Q(
        memory_interface_inst1_fsm_state_0_) );
  DFQD1BWP12T irdecode_inst1_memory_load_request_reg ( .D(n861), .CP(clk), .Q(
        DEC_MEMCTRL_memory_load_request) );
  DFQD1BWP12T irdecode_inst1_stall_to_instructionfetch_reg ( .D(n845), .CP(clk), .Q(DEC_IF_stall_to_instructionfetch) );
  DFQD1BWP12T Instruction_Fetch_inst1_currentState_reg_1_ ( .D(
        Instruction_Fetch_inst1_N80), .CP(clk), .Q(
        Instruction_Fetch_inst1_currentState_1_) );
  DFQD1BWP12T Instruction_Fetch_inst1_currentState_reg_0_ ( .D(
        Instruction_Fetch_inst1_N79), .CP(clk), .Q(
        Instruction_Fetch_inst1_currentState_0_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_0_ ( .D(
        MEMCTRL_IN_address[0]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[0]) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_0_ ( .D(
        Instruction_Fetch_inst1_N83), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_0_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_1_ ( .D(
        Instruction_Fetch_inst1_N84), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_1_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_2_ ( .D(
        Instruction_Fetch_inst1_N85), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_2_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_3_ ( .D(
        Instruction_Fetch_inst1_N86), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_3_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_4_ ( .D(
        Instruction_Fetch_inst1_N87), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_4_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_5_ ( .D(
        Instruction_Fetch_inst1_N88), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_5_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_6_ ( .D(
        Instruction_Fetch_inst1_N89), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_6_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_7_ ( .D(
        Instruction_Fetch_inst1_N90), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_7_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_15_ ( .D(
        Instruction_Fetch_inst1_N98), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_15_) );
  DFQD1BWP12T irdecode_inst1_memorycontroller_sign_extend_reg ( .D(n839), .CP(
        clk), .Q(DEC_MEMCTRL_memorycontroller_sign_extend) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_8_ ( .D(
        Instruction_Fetch_inst1_N91), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_8_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_9_ ( .D(
        Instruction_Fetch_inst1_N92), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_9_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_11_ ( .D(
        Instruction_Fetch_inst1_N94), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_11_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_10_ ( .D(
        Instruction_Fetch_inst1_N93), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_10_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_13_ ( .D(
        Instruction_Fetch_inst1_N96), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_13_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_14_ ( .D(
        Instruction_Fetch_inst1_N97), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_14_) );
  DFQD1BWP12T irdecode_inst1_step_reg_1_ ( .D(irdecode_inst1_next_step_1_), 
        .CP(clk), .Q(irdecode_inst1_step[1]) );
  DFQD1BWP12T irdecode_inst1_split_instruction_reg ( .D(n847), .CP(clk), .Q(
        irdecode_inst1_split_instruction) );
  DFQD1BWP12T irdecode_inst1_step_reg_6_ ( .D(irdecode_inst1_next_step_6_), 
        .CP(clk), .Q(irdecode_inst1_step[6]) );
  DFQD1BWP12T irdecode_inst1_step_reg_5_ ( .D(irdecode_inst1_next_step_5_), 
        .CP(clk), .Q(irdecode_inst1_step[5]) );
  DFQD1BWP12T irdecode_inst1_step_reg_0_ ( .D(irdecode_inst1_next_step_0_), 
        .CP(clk), .Q(irdecode_inst1_step[0]) );
  DFQD1BWP12T irdecode_inst1_step_reg_2_ ( .D(irdecode_inst1_next_step_2_), 
        .CP(clk), .Q(irdecode_inst1_step[2]) );
  DFQD1BWP12T irdecode_inst1_step_reg_3_ ( .D(irdecode_inst1_next_step_3_), 
        .CP(clk), .Q(irdecode_inst1_step[3]) );
  DFQD1BWP12T irdecode_inst1_step_reg_4_ ( .D(irdecode_inst1_next_step_4_), 
        .CP(clk), .Q(irdecode_inst1_step[4]) );
  DFQD1BWP12T irdecode_inst1_step_reg_7_ ( .D(irdecode_inst1_next_step_7_), 
        .CP(clk), .Q(irdecode_inst1_step[7]) );
  DFQD1BWP12T irdecode_inst1_memory_store_request_reg ( .D(n852), .CP(clk), 
        .Q(DEC_MEMCTRL_memory_store_request) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_0_ ( .D(n860), .CP(clk), .Q(
        irdecode_inst1_itstate_0_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_1_ ( .D(n859), .CP(clk), .Q(
        irdecode_inst1_itstate_1_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_2_ ( .D(n858), .CP(clk), .Q(
        irdecode_inst1_itstate_2_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_3_ ( .D(n857), .CP(clk), .Q(
        irdecode_inst1_itstate_3_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_4_ ( .D(n856), .CP(clk), .Q(
        irdecode_inst1_itstate_4_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_5_ ( .D(n855), .CP(clk), .Q(
        irdecode_inst1_itstate_5_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_7_ ( .D(n853), .CP(clk), .Q(
        irdecode_inst1_itstate_7_) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_0_ ( .D(n835), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[0]) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_2_ ( .D(n833), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[2]) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_3_ ( .D(n832), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[3]) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_4_ ( .D(n831), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[4]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_0_ ( .D(n830), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[0]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_2_ ( .D(n828), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[2]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_3_ ( .D(n827), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[3]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_4_ ( .D(n826), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[4]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_0_ ( .D(n824), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[0]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_2_ ( .D(n822), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[2]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_4_ ( .D(n848), .CP(clk), .Q(
        DEC_ALU_alu_opcode[4]) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_12_ ( .D(
        Instruction_Fetch_inst1_N95), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_12_) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_3_ ( .D(n821), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[3]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_4_ ( .D(n820), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[4]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_1_ ( .D(n850), .CP(clk), .Q(
        DEC_ALU_alu_opcode[1]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_2_ ( .D(n846), .CP(clk), .Q(
        DEC_ALU_alu_opcode[2]) );
  DFQD1BWP12T irdecode_inst1_update_flag_v_reg ( .D(
        irdecode_inst1_next_update_flag_v), .CP(clk), .Q(
        DEC_CPSR_update_flag_v) );
  DFQD1BWP12T irdecode_inst1_update_flag_c_reg ( .D(
        irdecode_inst1_next_update_flag_c), .CP(clk), .Q(
        DEC_CPSR_update_flag_c) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_0_ ( .D(n851), .CP(clk), .Q(
        DEC_ALU_alu_opcode[0]) );
  DFQD1BWP12T irdecode_inst1_update_flag_n_reg ( .D(
        irdecode_inst1_next_update_flag_n), .CP(clk), .Q(
        DEC_CPSR_update_flag_n) );
  DFQD1BWP12T irdecode_inst1_update_flag_z_reg ( .D(
        irdecode_inst1_next_update_flag_n), .CP(clk), .Q(
        DEC_CPSR_update_flag_z) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_3_ ( .D(n849), .CP(clk), .Q(
        DEC_ALU_alu_opcode[3]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_2_ ( .D(n818), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[2]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_3_ ( .D(n817), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[3]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_4_ ( .D(n815), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[4]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_0_ ( .D(n816), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[0]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_enable_reg ( .D(
        irdecode_inst1_next_alu_write_to_reg_enable), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg_enable) );
  DFQD1BWP12T irdecode_inst1_memory_address_source_is_reg_reg ( .D(n836), .CP(
        clk), .Q(DEC_MISC_OUT_memory_address_source_is_reg) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_1_ ( .D(n834), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[1]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_1_ ( .D(n829), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[1]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_enable_reg ( .D(n825), .CP(
        clk), .Q(DEC_RF_memory_write_to_reg_enable) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_1_ ( .D(n823), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[1]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_1_ ( .D(n819), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[1]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_0_ ( .D(n809), .CP(clk), .Q(
        DEC_RF_offset_b[0]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_1_ ( .D(n808), .CP(clk), .Q(
        DEC_RF_offset_b[1]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_2_ ( .D(n807), .CP(clk), .Q(
        DEC_RF_offset_b[2]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_3_ ( .D(n806), .CP(clk), .Q(
        DEC_RF_offset_b[3]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_4_ ( .D(n805), .CP(clk), .Q(
        DEC_RF_offset_b[4]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_5_ ( .D(n804), .CP(clk), .Q(
        DEC_RF_offset_b[5]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_6_ ( .D(n803), .CP(clk), .Q(
        DEC_RF_offset_b[6]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_7_ ( .D(n802), .CP(clk), .Q(
        DEC_RF_offset_b[7]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_8_ ( .D(n801), .CP(clk), .Q(
        DEC_RF_offset_b[8]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_9_ ( .D(n800), .CP(clk), .Q(
        DEC_RF_offset_b[9]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_10_ ( .D(n799), .CP(clk), .Q(
        DEC_RF_offset_b[10]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_11_ ( .D(n798), .CP(clk), .Q(
        DEC_RF_offset_b[11]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_12_ ( .D(n797), .CP(clk), .Q(
        DEC_RF_offset_b[12]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_13_ ( .D(n796), .CP(clk), .Q(
        DEC_RF_offset_b[13]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_14_ ( .D(n795), .CP(clk), .Q(
        DEC_RF_offset_b[14]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_15_ ( .D(n794), .CP(clk), .Q(
        DEC_RF_offset_b[15]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_16_ ( .D(n793), .CP(clk), .Q(
        DEC_RF_offset_b[16]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_17_ ( .D(n792), .CP(clk), .Q(
        DEC_RF_offset_b[17]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_18_ ( .D(n791), .CP(clk), .Q(
        DEC_RF_offset_b[18]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_19_ ( .D(n790), .CP(clk), .Q(
        DEC_RF_offset_b[19]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_20_ ( .D(n789), .CP(clk), .Q(
        DEC_RF_offset_b[20]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_21_ ( .D(n788), .CP(clk), .Q(
        DEC_RF_offset_b[21]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_22_ ( .D(n787), .CP(clk), .Q(
        DEC_RF_offset_b[22]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_23_ ( .D(n786), .CP(clk), .Q(
        DEC_RF_offset_b[23]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_24_ ( .D(n785), .CP(clk), .Q(
        DEC_RF_offset_b[24]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_25_ ( .D(n784), .CP(clk), .Q(
        DEC_RF_offset_b[25]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_26_ ( .D(n783), .CP(clk), .Q(
        DEC_RF_offset_b[26]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_27_ ( .D(n782), .CP(clk), .Q(
        DEC_RF_offset_b[27]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_28_ ( .D(n781), .CP(clk), .Q(
        DEC_RF_offset_b[28]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_29_ ( .D(n780), .CP(clk), .Q(
        DEC_RF_offset_b[29]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_30_ ( .D(n779), .CP(clk), .Q(
        DEC_RF_offset_b[30]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_0_ ( .D(
        RF_MEMCTRL_data_reg[0]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[0]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_1_ ( .D(
        RF_MEMCTRL_data_reg[1]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[1]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_2_ ( .D(
        RF_MEMCTRL_data_reg[2]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_3_ ( .D(
        RF_MEMCTRL_data_reg[3]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_4_ ( .D(
        RF_MEMCTRL_data_reg[4]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[4]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_5_ ( .D(
        RF_MEMCTRL_data_reg[5]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[5]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_6_ ( .D(
        RF_MEMCTRL_data_reg[6]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_7_ ( .D(
        RF_MEMCTRL_data_reg[7]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_8_ ( .D(
        RF_MEMCTRL_data_reg[8]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_9_ ( .D(
        RF_MEMCTRL_data_reg[9]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_10_ ( .D(
        RF_MEMCTRL_data_reg[10]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_11_ ( .D(
        RF_MEMCTRL_data_reg[11]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[11]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_12_ ( .D(
        RF_MEMCTRL_data_reg[12]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[12]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_13_ ( .D(
        RF_MEMCTRL_data_reg[13]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[13]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_14_ ( .D(
        RF_MEMCTRL_data_reg[14]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[14]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_15_ ( .D(
        RF_MEMCTRL_data_reg[15]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[15]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_16_ ( .D(
        RF_MEMCTRL_data_reg[16]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[16]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_17_ ( .D(
        RF_MEMCTRL_data_reg[17]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[17]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_18_ ( .D(
        RF_MEMCTRL_data_reg[18]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[18]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_19_ ( .D(
        RF_MEMCTRL_data_reg[19]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[19]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_20_ ( .D(
        RF_MEMCTRL_data_reg[20]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[20]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_21_ ( .D(
        RF_MEMCTRL_data_reg[21]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[21]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_22_ ( .D(
        RF_MEMCTRL_data_reg[22]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[22]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_23_ ( .D(
        RF_MEMCTRL_data_reg[23]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[23]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_24_ ( .D(
        RF_MEMCTRL_data_reg[24]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[24]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_25_ ( .D(
        RF_MEMCTRL_data_reg[25]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[25]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_26_ ( .D(
        RF_MEMCTRL_data_reg[26]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[26]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_27_ ( .D(
        RF_MEMCTRL_data_reg[27]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[27]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_28_ ( .D(
        RF_MEMCTRL_data_reg[28]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[28]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_29_ ( .D(
        RF_MEMCTRL_data_reg[29]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[29]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_30_ ( .D(
        RF_MEMCTRL_data_reg[30]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[30]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_31_ ( .D(
        RF_MEMCTRL_data_reg[31]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[31]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_1_ ( .D(
        MEMCTRL_IN_address[1]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[1]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_2_ ( .D(
        MEMCTRL_IN_address[2]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_3_ ( .D(
        MEMCTRL_IN_address[3]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_4_ ( .D(
        MEMCTRL_IN_address[4]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[4]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_5_ ( .D(
        MEMCTRL_IN_address[5]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[5]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_6_ ( .D(
        MEMCTRL_IN_address[6]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_7_ ( .D(
        MEMCTRL_IN_address[7]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_8_ ( .D(
        MEMCTRL_IN_address[8]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_9_ ( .D(
        MEMCTRL_IN_address[9]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_10_ ( .D(
        MEMCTRL_IN_address[10]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_11_ ( .D(
        MEMCTRL_IN_address[11]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[11]) );
  DFQD4BWP12T irdecode_inst1_operand_a_reg_4_ ( .D(n810), .CP(clk), .Q(
        DEC_RF_operand_a[4]) );
  DFQD4BWP12T irdecode_inst1_operand_a_reg_3_ ( .D(n812), .CP(clk), .Q(
        DEC_RF_operand_a[3]) );
  DFQD4BWP12T irdecode_inst1_operand_a_reg_0_ ( .D(n811), .CP(clk), .Q(
        DEC_RF_operand_a[0]) );
  DFQD4BWP12T irdecode_inst1_operand_b_reg_0_ ( .D(n844), .CP(clk), .Q(
        DEC_RF_operand_b[0]) );
  DFQD4BWP12T irdecode_inst1_operand_b_reg_3_ ( .D(n841), .CP(clk), .Q(
        DEC_RF_operand_b[3]) );
  DFQD4BWP12T irdecode_inst1_operand_a_reg_2_ ( .D(n813), .CP(clk), .Q(
        DEC_RF_operand_a[2]) );
  DFQD4BWP12T irdecode_inst1_operand_a_reg_1_ ( .D(n814), .CP(clk), .Q(
        DEC_RF_operand_a[1]) );
  DFQD4BWP12T irdecode_inst1_operand_b_reg_2_ ( .D(n842), .CP(clk), .Q(
        DEC_RF_operand_b[2]) );
  DFQD4BWP12T irdecode_inst1_operand_b_reg_1_ ( .D(n843), .CP(clk), .Q(
        DEC_RF_operand_b[1]) );
  DFQD4BWP12T irdecode_inst1_operand_b_reg_4_ ( .D(n840), .CP(clk), .Q(
        DEC_RF_operand_b[4]) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_6_ ( .D(n854), .CP(clk), .Q(
        irdecode_inst1_itstate_6_) );
  DFXD1BWP12T memory_interface_inst1_delayed_is_signed_reg ( .D(
        DEC_MEMCTRL_memorycontroller_sign_extend), .CP(clk), .Q(
        memory_interface_inst1_delayed_is_signed), .QN(n1684) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_2_ ( .D(
        memory_interface_inst1_fsm_N34), .CP(clk), .Q(
        memory_interface_inst1_fsm_state_2_) );
  TIELBWP12T U1022 ( .ZN(n864) );
  INVD1BWP12T U1023 ( .I(n864), .ZN(MEMCTRL_MEM_to_mem_mem_enable) );
  MUX2ND0BWP12T U1024 ( .I0(n1377), .I1(MEM_MEMCTRL_from_mem_data[15]), .S(
        n1376), .ZN(n1547) );
  HA1D0BWP12T U1025 ( .A(n1198), .B(RF_pc_out[28]), .CO(n1169), .S(n1199) );
  ND2D1BWP12T U1026 ( .A1(n938), .A2(Instruction_Fetch_inst1_currentState_1_), 
        .ZN(n1369) );
  ND2D1BWP12T U1027 ( .A1(n1612), .A2(n994), .ZN(n1057) );
  ND3D0BWP12T U1028 ( .A1(memory_interface_inst1_fsm_state_3_), .A2(n940), 
        .A3(memory_interface_inst1_fsm_state_2_), .ZN(n1386) );
  OR2D0BWP12T U1029 ( .A1(n964), .A2(n1122), .Z(n1619) );
  INR3D0BWP12T U1030 ( .A1(n1000), .B1(n1628), .B2(n1664), .ZN(n1661) );
  INR2D0BWP12T U1031 ( .A1(n1399), .B1(n1557), .ZN(n1448) );
  IOA21D1BWP12T U1032 ( .A1(n1116), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_8_), .B(n1119), .ZN(
        n865) );
  AOI21D1BWP12T U1033 ( .A1(n1422), .A2(MEMCTRL_RF_IF_data_in[8]), .B(n865), 
        .ZN(n1583) );
  IND2D0BWP12T U1034 ( .A1(n1448), .B1(n1472), .ZN(n1465) );
  AOI31D0BWP12T U1035 ( .A1(n1359), .A2(irdecode_inst1_split_instruction), 
        .A3(DEC_IF_stall_to_instructionfetch), .B(n1559), .ZN(n866) );
  INR2D0BWP12T U1036 ( .A1(n995), .B1(n866), .ZN(n1328) );
  IND2D0BWP12T U1037 ( .A1(n1116), .B1(n754), .ZN(n1119) );
  INR2D0BWP12T U1038 ( .A1(n1557), .B1(n1399), .ZN(n1466) );
  AOI21D0BWP12T U1039 ( .A1(n1141), .A2(irdecode_inst1_N706), .B(n1069), .ZN(
        n867) );
  ND3D0BWP12T U1040 ( .A1(n1142), .A2(n867), .A3(n1068), .ZN(n868) );
  OAI31D0BWP12T U1041 ( .A1(n1597), .A2(n1201), .A3(n868), .B(n1595), .ZN(n869) );
  OAI211D0BWP12T U1042 ( .A1(n1647), .A2(n1164), .B(n1273), .C(n869), .ZN(
        n1184) );
  IOA21D0BWP12T U1043 ( .A1(
        Instruction_Fetch_inst1_fetched_instruction_reg_10_), .A2(n1116), .B(
        n1119), .ZN(n870) );
  AO21D0BWP12T U1044 ( .A1(n1422), .A2(MEMCTRL_RF_IF_data_in[10]), .B(n870), 
        .Z(n1656) );
  CKND0BWP12T U1045 ( .I(n1017), .ZN(n871) );
  OAI31D1BWP12T U1046 ( .A1(n1016), .A2(irdecode_inst1_N546), .A3(n871), .B(
        n1064), .ZN(n1024) );
  NR2D1BWP12T U1047 ( .A1(irdecode_inst1_N704), .A2(n1140), .ZN(n872) );
  ND4D1BWP12T U1048 ( .A1(n1004), .A2(n1006), .A3(n1002), .A4(n872), .ZN(n1146) );
  AN3D0BWP12T U1049 ( .A1(n1385), .A2(n1383), .A3(n1384), .Z(n1557) );
  OA211D0BWP12T U1050 ( .A1(n1641), .A2(n1640), .B(n1639), .C(n1638), .Z(n873)
         );
  CKND0BWP12T U1051 ( .I(n1637), .ZN(n874) );
  AOI22D0BWP12T U1052 ( .A1(n1672), .A2(n1636), .B1(n1664), .B2(n874), .ZN(
        n875) );
  OAI211D0BWP12T U1053 ( .A1(n1643), .A2(n1642), .B(n873), .C(n875), .ZN(n876)
         );
  NR3D0BWP12T U1054 ( .A1(n1644), .A2(n1674), .A3(n876), .ZN(n877) );
  MOAI22D0BWP12T U1055 ( .A1(n877), .A2(n1679), .B1(DEC_RF_operand_a[1]), .B2(
        n1682), .ZN(n814) );
  IND4D0BWP12T U1056 ( .A1(n1021), .B1(n1019), .B2(n1020), .B3(n1660), .ZN(
        n878) );
  NR2D0BWP12T U1057 ( .A1(n1025), .A2(n878), .ZN(n1055) );
  INR3D0BWP12T U1058 ( .A1(irdecode_inst1_N705), .B1(irdecode_inst1_N707), 
        .B2(n1007), .ZN(n1144) );
  IAO21D0BWP12T U1059 ( .A1(n1551), .A2(
        memory_interface_inst1_delay_addr_for_adder[0]), .B(n1434), .ZN(n1460)
         );
  CKND0BWP12T U1060 ( .I(n1556), .ZN(n879) );
  CKND0BWP12T U1061 ( .I(n1557), .ZN(n880) );
  AOI32D0BWP12T U1062 ( .A1(n1555), .A2(n1557), .A3(n879), .B1(n1558), .B2(
        n880), .ZN(MEMCTRL_MEM_to_mem_read_enable) );
  AN2D0BWP12T U1063 ( .A1(n1422), .A2(n1343), .Z(IF_RF_incremented_pc_out[13])
         );
  CKND0BWP12T U1064 ( .I(n1582), .ZN(n881) );
  AOI32D0BWP12T U1065 ( .A1(IF_DEC_instruction[7]), .A2(n1600), .A3(n1617), 
        .B1(n1582), .B2(n1600), .ZN(n882) );
  OAI22D0BWP12T U1066 ( .A1(n1088), .A2(n881), .B1(n1290), .B2(n882), .ZN(n883) );
  OAI31D0BWP12T U1067 ( .A1(n1090), .A2(n1586), .A3(n883), .B(n1584), .ZN(n884) );
  IND2D0BWP12T U1068 ( .A1(n1589), .B1(n884), .ZN(
        irdecode_inst1_next_update_flag_v) );
  IIND4D1BWP12T U1069 ( .A1(irdecode_inst1_N540), .A2(irdecode_inst1_N541), 
        .B1(irdecode_inst1_N539), .B2(n1013), .ZN(n1061) );
  CKND0BWP12T U1070 ( .I(n1549), .ZN(n885) );
  AOI21D0BWP12T U1071 ( .A1(
        memory_interface_inst1_delay_first_two_bytes_out[9]), .A2(n885), .B(
        n956), .ZN(n886) );
  OAI21D0BWP12T U1072 ( .A1(n957), .A2(n1443), .B(n886), .ZN(
        MEMCTRL_RF_IF_data_in[9]) );
  CKND0BWP12T U1073 ( .I(n1467), .ZN(n887) );
  AOI222D0BWP12T U1074 ( .A1(n887), .A2(RF_MEMCTRL_data_reg[0]), .B1(n1465), 
        .B2(memory_interface_inst1_delay_data_in32[0]), .C1(n1474), .C2(
        memory_interface_inst1_delay_data_in32[16]), .ZN(n888) );
  IOA21D0BWP12T U1075 ( .A1(n1466), .A2(RF_MEMCTRL_data_reg[16]), .B(n888), 
        .ZN(MEMCTRL_MEM_to_mem_data[8]) );
  AN2D0BWP12T U1076 ( .A1(n1422), .A2(n1341), .Z(IF_RF_incremented_pc_out[14])
         );
  MOAI22D1BWP12T U1077 ( .A1(n754), .A2(n1568), .B1(n1116), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_0_), .ZN(
        IF_DEC_instruction[0]) );
  NR2D0BWP12T U1078 ( .A1(n1375), .A2(memory_interface_inst1_delayed_is_signed), .ZN(n889) );
  NR3D0BWP12T U1079 ( .A1(n889), .A2(n943), .A3(MEM_MEMCTRL_from_mem_data[15]), 
        .ZN(n956) );
  CKND0BWP12T U1080 ( .I(n1467), .ZN(n890) );
  AOI222D0BWP12T U1081 ( .A1(n890), .A2(RF_MEMCTRL_data_reg[1]), .B1(n1465), 
        .B2(memory_interface_inst1_delay_data_in32[1]), .C1(n1474), .C2(
        memory_interface_inst1_delay_data_in32[17]), .ZN(n891) );
  IOA21D0BWP12T U1082 ( .A1(RF_MEMCTRL_data_reg[17]), .A2(n1466), .B(n891), 
        .ZN(MEMCTRL_MEM_to_mem_data[9]) );
  AN2D0BWP12T U1083 ( .A1(n1422), .A2(n1339), .Z(IF_RF_incremented_pc_out[15])
         );
  MOAI22D0BWP12T U1084 ( .A1(n754), .A2(n1565), .B1(n1116), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_1_), .ZN(
        IF_DEC_instruction[1]) );
  IND3D1BWP12T U1085 ( .A1(irdecode_inst1_N541), .B1(irdecode_inst1_N540), 
        .B2(n1013), .ZN(n1510) );
  CKND0BWP12T U1086 ( .I(n1467), .ZN(n892) );
  AOI222D0BWP12T U1087 ( .A1(n892), .A2(RF_MEMCTRL_data_reg[3]), .B1(n1465), 
        .B2(memory_interface_inst1_delay_data_in32[3]), .C1(n1474), .C2(
        memory_interface_inst1_delay_data_in32[19]), .ZN(n893) );
  IOA21D0BWP12T U1088 ( .A1(RF_MEMCTRL_data_reg[19]), .A2(n1466), .B(n893), 
        .ZN(MEMCTRL_MEM_to_mem_data[11]) );
  AN2D0BWP12T U1089 ( .A1(n1422), .A2(n1312), .Z(IF_RF_incremented_pc_out[18])
         );
  MOAI22D0BWP12T U1090 ( .A1(n754), .A2(n1566), .B1(n1116), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_2_), .ZN(
        IF_DEC_instruction[2]) );
  MAOI22D0BWP12T U1091 ( .A1(n990), .A2(n1573), .B1(n1306), .B2(n1290), .ZN(
        n1227) );
  CKND0BWP12T U1092 ( .I(n1467), .ZN(n894) );
  AOI222D0BWP12T U1093 ( .A1(n894), .A2(RF_MEMCTRL_data_reg[2]), .B1(n1465), 
        .B2(memory_interface_inst1_delay_data_in32[2]), .C1(n1474), .C2(
        memory_interface_inst1_delay_data_in32[18]), .ZN(n895) );
  IOA21D0BWP12T U1094 ( .A1(RF_MEMCTRL_data_reg[18]), .A2(n1466), .B(n895), 
        .ZN(MEMCTRL_MEM_to_mem_data[10]) );
  AN2D0BWP12T U1095 ( .A1(n1422), .A2(n1285), .Z(IF_RF_incremented_pc_out[19])
         );
  AOI22D0BWP12T U1096 ( .A1(irdecode_inst1_N707), .A2(n1595), .B1(
        irdecode_inst1_step[1]), .B2(n1682), .ZN(n896) );
  AOI21D0BWP12T U1097 ( .A1(irdecode_inst1_N546), .A2(n1501), .B(n1028), .ZN(
        n897) );
  OAI211D1BWP12T U1098 ( .A1(n1331), .A2(n1057), .B(n896), .C(n897), .ZN(
        irdecode_inst1_next_step_1_) );
  MOAI22D0BWP12T U1099 ( .A1(n754), .A2(n1561), .B1(n1116), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_3_), .ZN(
        IF_DEC_instruction[3]) );
  NR2D0BWP12T U1100 ( .A1(n1144), .A2(n1174), .ZN(n898) );
  ND4D0BWP12T U1101 ( .A1(n1143), .A2(n1173), .A3(n898), .A4(n1142), .ZN(n1659) );
  MOAI22D0BWP12T U1102 ( .A1(n1379), .A2(n1545), .B1(n1379), .B2(
        memory_interface_inst1_delay_first_two_bytes_out[1]), .ZN(
        MEMCTRL_RF_IF_data_in[1]) );
  MOAI22D0BWP12T U1103 ( .A1(n1379), .A2(n1544), .B1(n1379), .B2(
        memory_interface_inst1_delay_first_two_bytes_out[2]), .ZN(
        MEMCTRL_RF_IF_data_in[2]) );
  MOAI22D0BWP12T U1104 ( .A1(n1379), .A2(n1542), .B1(n1379), .B2(
        memory_interface_inst1_delay_first_two_bytes_out[5]), .ZN(
        MEMCTRL_RF_IF_data_in[5]) );
  MOAI22D0BWP12T U1105 ( .A1(n1379), .A2(n1546), .B1(n1379), .B2(
        memory_interface_inst1_delay_first_two_bytes_out[0]), .ZN(
        MEMCTRL_RF_IF_data_in[0]) );
  CKND0BWP12T U1106 ( .I(n1549), .ZN(n899) );
  AOI21D0BWP12T U1107 ( .A1(
        memory_interface_inst1_delay_first_two_bytes_out[8]), .A2(n899), .B(
        n956), .ZN(n900) );
  OAI21D0BWP12T U1108 ( .A1(n957), .A2(n1539), .B(n900), .ZN(
        MEMCTRL_RF_IF_data_in[8]) );
  CKND0BWP12T U1109 ( .I(n1467), .ZN(n901) );
  AOI222D0BWP12T U1110 ( .A1(n901), .A2(RF_MEMCTRL_data_reg[6]), .B1(n1465), 
        .B2(memory_interface_inst1_delay_data_in32[6]), .C1(n1474), .C2(
        memory_interface_inst1_delay_data_in32[22]), .ZN(n902) );
  IOA21D0BWP12T U1111 ( .A1(RF_MEMCTRL_data_reg[22]), .A2(n1466), .B(n902), 
        .ZN(MEMCTRL_MEM_to_mem_data[14]) );
  AN2D0BWP12T U1112 ( .A1(n1422), .A2(n1283), .Z(IF_RF_incremented_pc_out[20])
         );
  MOAI22D0BWP12T U1113 ( .A1(n754), .A2(n1564), .B1(n1116), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_4_), .ZN(
        IF_DEC_instruction[4]) );
  CKND0BWP12T U1114 ( .I(DEC_ALU_alu_opcode[1]), .ZN(n903) );
  OR4D0BWP12T U1115 ( .A1(DEC_ALU_alu_opcode[3]), .A2(n1550), .A3(
        DEC_ALU_alu_opcode[0]), .A4(n903), .Z(n904) );
  MAOI22D0BWP12T U1116 ( .A1(DEC_ALU_alu_opcode[4]), .A2(n904), .B1(
        DEC_ALU_alu_opcode[4]), .B2(RF_OUT_c), .ZN(ALU_IN_c) );
  MOAI22D0BWP12T U1117 ( .A1(n1379), .A2(n1543), .B1(n1379), .B2(
        memory_interface_inst1_delay_first_two_bytes_out[3]), .ZN(
        MEMCTRL_RF_IF_data_in[3]) );
  MOAI22D0BWP12T U1118 ( .A1(n1379), .A2(n1548), .B1(n1379), .B2(
        memory_interface_inst1_delay_first_two_bytes_out[4]), .ZN(
        MEMCTRL_RF_IF_data_in[4]) );
  MOAI22D0BWP12T U1119 ( .A1(n1379), .A2(n1541), .B1(n1379), .B2(
        memory_interface_inst1_delay_first_two_bytes_out[6]), .ZN(
        MEMCTRL_RF_IF_data_in[6]) );
  MOAI22D0BWP12T U1120 ( .A1(n1379), .A2(n1540), .B1(n1379), .B2(
        memory_interface_inst1_delay_first_two_bytes_out[7]), .ZN(
        MEMCTRL_RF_IF_data_in[7]) );
  CKND0BWP12T U1121 ( .I(n1549), .ZN(n905) );
  AOI21D0BWP12T U1122 ( .A1(
        memory_interface_inst1_delay_first_two_bytes_out[10]), .A2(n905), .B(
        n956), .ZN(n906) );
  OAI21D0BWP12T U1123 ( .A1(n957), .A2(n1538), .B(n906), .ZN(
        MEMCTRL_RF_IF_data_in[10]) );
  AOI211D1BWP12T U1124 ( .A1(irdecode_inst1_N911), .A2(n1612), .B(n1212), .C(
        n1037), .ZN(n907) );
  AOI22D0BWP12T U1125 ( .A1(n1210), .A2(n1501), .B1(n1214), .B2(n1595), .ZN(
        n908) );
  OAI211D1BWP12T U1126 ( .A1(n1331), .A2(n907), .B(n1273), .C(n908), .ZN(n1028) );
  CKND0BWP12T U1127 ( .I(n1467), .ZN(n909) );
  AOI222D0BWP12T U1128 ( .A1(n909), .A2(RF_MEMCTRL_data_reg[7]), .B1(n1465), 
        .B2(memory_interface_inst1_delay_data_in32[7]), .C1(n1474), .C2(
        memory_interface_inst1_delay_data_in32[23]), .ZN(n910) );
  IOA21D0BWP12T U1129 ( .A1(RF_MEMCTRL_data_reg[23]), .A2(n1466), .B(n910), 
        .ZN(MEMCTRL_MEM_to_mem_data[15]) );
  AN2D0BWP12T U1130 ( .A1(n1422), .A2(n1366), .Z(IF_RF_incremented_pc_out[2])
         );
  AN2D0BWP12T U1131 ( .A1(n1422), .A2(n1087), .Z(IF_RF_incremented_pc_out[21])
         );
  CKND0BWP12T U1132 ( .I(n1575), .ZN(n911) );
  OAI21D0BWP12T U1133 ( .A1(n1576), .A2(n911), .B(n1584), .ZN(n912) );
  IOA21D0BWP12T U1134 ( .A1(n1578), .A2(n1577), .B(n912), .ZN(
        irdecode_inst1_next_update_flag_n) );
  MOAI22D0BWP12T U1135 ( .A1(n754), .A2(n1560), .B1(n1116), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_5_), .ZN(
        IF_DEC_instruction[5]) );
  INR2D0BWP12T U1136 ( .A1(n1082), .B1(n1275), .ZN(n1070) );
  IND2D0BWP12T U1137 ( .A1(memory_interface_inst1_fsm_state_1_), .B1(n1378), 
        .ZN(n1371) );
  OAI21D0BWP12T U1138 ( .A1(n1131), .A2(RF_pc_out[31]), .B(n1422), .ZN(n913)
         );
  AOI21D0BWP12T U1139 ( .A1(n1131), .A2(RF_pc_out[31]), .B(n913), .ZN(
        IF_RF_incremented_pc_out[31]) );
  CKND0BWP12T U1140 ( .I(n1549), .ZN(n914) );
  AOI21D0BWP12T U1141 ( .A1(
        memory_interface_inst1_delay_first_two_bytes_out[14]), .A2(n914), .B(
        n956), .ZN(n915) );
  OAI21D0BWP12T U1142 ( .A1(n957), .A2(n1426), .B(n915), .ZN(
        MEMCTRL_RF_IF_data_in[14]) );
  CKND0BWP12T U1143 ( .I(n1467), .ZN(n916) );
  AOI222D0BWP12T U1144 ( .A1(n916), .A2(RF_MEMCTRL_data_reg[4]), .B1(n1465), 
        .B2(memory_interface_inst1_delay_data_in32[4]), .C1(n1474), .C2(
        memory_interface_inst1_delay_data_in32[20]), .ZN(n917) );
  IOA21D0BWP12T U1145 ( .A1(RF_MEMCTRL_data_reg[20]), .A2(n1466), .B(n917), 
        .ZN(MEMCTRL_MEM_to_mem_data[12]) );
  AO222D0BWP12T U1146 ( .A1(memory_interface_inst1_delay_addr_for_adder[9]), 
        .A2(n1554), .B1(MEMCTRL_IN_address[9]), .B2(n1551), .C1(n1552), .C2(
        n1553), .Z(MEMCTRL_MEM_to_mem_address[9]) );
  AN2D0BWP12T U1147 ( .A1(n1422), .A2(n1368), .Z(IF_RF_incremented_pc_out[3])
         );
  CKND0BWP12T U1148 ( .I(RF_OUT_c), .ZN(n918) );
  MOAI22D0BWP12T U1149 ( .A1(DEC_CPSR_update_flag_c), .A2(n918), .B1(
        DEC_CPSR_update_flag_c), .B2(ALU_OUT_c), .ZN(new_c) );
  AN2D0BWP12T U1150 ( .A1(n1422), .A2(n1363), .Z(IF_RF_incremented_pc_out[5])
         );
  AN2D0BWP12T U1151 ( .A1(n1422), .A2(n1355), .Z(IF_RF_incremented_pc_out[7])
         );
  AN2D0BWP12T U1152 ( .A1(n1422), .A2(n1351), .Z(IF_RF_incremented_pc_out[9])
         );
  AN2D0BWP12T U1153 ( .A1(n1422), .A2(n1347), .Z(IF_RF_incremented_pc_out[11])
         );
  AN2D0BWP12T U1154 ( .A1(n1422), .A2(n1085), .Z(IF_RF_incremented_pc_out[22])
         );
  AOI21D0BWP12T U1155 ( .A1(n1590), .A2(n1306), .B(n1583), .ZN(n919) );
  ND3D0BWP12T U1156 ( .A1(n1263), .A2(n1625), .A3(n1264), .ZN(n920) );
  AOI211D0BWP12T U1157 ( .A1(n1593), .A2(IF_DEC_instruction[0]), .B(n919), .C(
        n920), .ZN(n921) );
  CKND2D0BWP12T U1158 ( .A1(DEC_RF_alu_write_to_reg[0]), .A2(n1682), .ZN(n922)
         );
  OAI211D0BWP12T U1159 ( .A1(n1331), .A2(n921), .B(n1038), .C(n922), .ZN(n816)
         );
  MOAI22D0BWP12T U1160 ( .A1(n754), .A2(n1563), .B1(n1116), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_6_), .ZN(
        IF_DEC_instruction[6]) );
  IND3D0BWP12T U1161 ( .A1(n1470), .B1(n1383), .B2(n1385), .ZN(n1551) );
  MUX2ND0BWP12T U1162 ( .I0(RF_OUT_n), .I1(n974), .S(RF_OUT_v), .ZN(n1293) );
  CKND0BWP12T U1163 ( .I(n1467), .ZN(n923) );
  AOI222D0BWP12T U1164 ( .A1(n923), .A2(RF_MEMCTRL_data_reg[5]), .B1(n1465), 
        .B2(memory_interface_inst1_delay_data_in32[5]), .C1(n1474), .C2(
        memory_interface_inst1_delay_data_in32[21]), .ZN(n924) );
  IOA21D0BWP12T U1165 ( .A1(RF_MEMCTRL_data_reg[21]), .A2(n1466), .B(n924), 
        .ZN(MEMCTRL_MEM_to_mem_data[13]) );
  AN2D0BWP12T U1166 ( .A1(n1422), .A2(RF_pc_out[0]), .Z(
        IF_RF_incremented_pc_out[0]) );
  AN2D0BWP12T U1167 ( .A1(n1422), .A2(n1365), .Z(IF_RF_incremented_pc_out[4])
         );
  AN2D0BWP12T U1168 ( .A1(n1422), .A2(n1361), .Z(IF_RF_incremented_pc_out[6])
         );
  AN2D0BWP12T U1169 ( .A1(n1422), .A2(n1353), .Z(IF_RF_incremented_pc_out[8])
         );
  AN2D0BWP12T U1170 ( .A1(n1422), .A2(n1349), .Z(IF_RF_incremented_pc_out[10])
         );
  AN2D0BWP12T U1171 ( .A1(n1422), .A2(n1345), .Z(IF_RF_incremented_pc_out[12])
         );
  AN2D0BWP12T U1172 ( .A1(n1422), .A2(n1244), .Z(IF_RF_incremented_pc_out[23])
         );
  CKND0BWP12T U1173 ( .I(n1676), .ZN(n925) );
  AOI222D0BWP12T U1174 ( .A1(n925), .A2(n1674), .B1(IF_DEC_instruction[1]), 
        .B2(n1675), .C1(n1677), .C2(n1678), .ZN(n926) );
  MOAI22D0BWP12T U1175 ( .A1(n1679), .A2(n926), .B1(
        DEC_RF_memory_write_to_reg[1]), .B2(n1682), .ZN(n823) );
  MUX2ND0BWP12T U1176 ( .I0(MEMCTRL_RF_IF_data_in[8]), .I1(
        Instruction_Fetch_inst1_fetched_instruction_reg_8_), .S(n754), .ZN(
        n927) );
  CKND2D0BWP12T U1177 ( .A1(n1359), .A2(n927), .ZN(Instruction_Fetch_inst1_N91) );
  MOAI22D0BWP12T U1178 ( .A1(n754), .A2(n1562), .B1(n1116), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_7_), .ZN(
        IF_DEC_instruction[7]) );
  BUFFD6BWP12T U1179 ( .I(RF_ALU_operand_a[13]), .Z(n1685) );
  OA32D1BWP12T U1180 ( .A1(n1230), .A2(n1203), .A3(n1202), .B1(n1328), .B2(
        n1230), .Z(n928) );
  INVD1BWP12T U1181 ( .I(reset), .ZN(n1359) );
  INVD1BWP12T U1182 ( .I(Instruction_Fetch_inst1_currentState_0_), .ZN(n938)
         );
  INVD4BWP12T U1183 ( .I(n1369), .ZN(n1422) );
  IND2D1BWP12T U1184 ( .A1(memory_interface_inst1_fsm_state_2_), .B1(
        memory_interface_inst1_fsm_state_1_), .ZN(n941) );
  INVD1BWP12T U1185 ( .I(n941), .ZN(n929) );
  NR2D1BWP12T U1186 ( .A1(memory_interface_inst1_fsm_state_0_), .A2(
        memory_interface_inst1_fsm_state_3_), .ZN(n931) );
  ND2D1BWP12T U1187 ( .A1(n929), .A2(n931), .ZN(n1375) );
  INR2D1BWP12T U1188 ( .A1(memory_interface_inst1_fsm_state_2_), .B1(
        memory_interface_inst1_fsm_state_1_), .ZN(n936) );
  INVD1BWP12T U1189 ( .I(n936), .ZN(n930) );
  INR2D2BWP12T U1190 ( .A1(n931), .B1(n930), .ZN(n1379) );
  INVD1BWP12T U1191 ( .I(n1379), .ZN(n933) );
  INR2D1BWP12T U1192 ( .A1(memory_interface_inst1_fsm_state_0_), .B1(
        memory_interface_inst1_fsm_state_1_), .ZN(n940) );
  NR2D1BWP12T U1193 ( .A1(memory_interface_inst1_fsm_state_2_), .A2(
        memory_interface_inst1_fsm_state_3_), .ZN(n1378) );
  CKND2D1BWP12T U1194 ( .A1(n940), .A2(n1378), .ZN(n932) );
  ND2D1BWP12T U1195 ( .A1(n933), .A2(n932), .ZN(n942) );
  INR2D1BWP12T U1196 ( .A1(n1375), .B1(n942), .ZN(n1385) );
  INVD1BWP12T U1197 ( .I(n1385), .ZN(n1480) );
  ND2D1BWP12T U1198 ( .A1(n1422), .A2(n1480), .ZN(n754) );
  NR2D1BWP12T U1199 ( .A1(n754), .A2(reset), .ZN(n1559) );
  CKND1BWP12T U1200 ( .I(memory_interface_inst1_fsm_state_0_), .ZN(n939) );
  TPND2D0BWP12T U1201 ( .A1(n941), .A2(n939), .ZN(n937) );
  OAI21D0BWP12T U1202 ( .A1(n939), .A2(memory_interface_inst1_fsm_state_2_), 
        .B(memory_interface_inst1_fsm_state_3_), .ZN(n934) );
  NR2D1BWP12T U1203 ( .A1(n934), .A2(n940), .ZN(n935) );
  OAI21D1BWP12T U1204 ( .A1(n937), .A2(n936), .B(n935), .ZN(n1383) );
  AOI22D1BWP12T U1205 ( .A1(n1385), .A2(DEC_MEMCTRL_memory_load_request), .B1(
        n1383), .B2(DEC_MEMCTRL_memory_store_request), .ZN(n995) );
  INVD1BWP12T U1206 ( .I(n1328), .ZN(n1331) );
  NR2D1BWP12T U1207 ( .A1(Instruction_Fetch_inst1_currentState_1_), .A2(n938), 
        .ZN(n1116) );
  INR2D1BWP12T U1208 ( .A1(n939), .B1(n1371), .ZN(n1470) );
  INR2D1BWP12T U1209 ( .A1(n1383), .B1(n1470), .ZN(n1373) );
  INR2D1BWP12T U1210 ( .A1(memory_interface_inst1_fsm_state_0_), .B1(n941), 
        .ZN(n1476) );
  INR2D1BWP12T U1211 ( .A1(n1386), .B1(n1476), .ZN(n1384) );
  IND3D1BWP12T U1212 ( .A1(n942), .B1(n1373), .B2(n1384), .ZN(n943) );
  INVD1BWP12T U1213 ( .I(n1379), .ZN(n1549) );
  ND2D1BWP12T U1214 ( .A1(n943), .A2(n1549), .ZN(n957) );
  INVD1BWP12T U1215 ( .I(n956), .ZN(n954) );
  ND2D1BWP12T U1216 ( .A1(n1379), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[12]), .ZN(n944) );
  OAI211D1BWP12T U1217 ( .A1(n957), .A2(n1391), .B(n954), .C(n944), .ZN(
        MEMCTRL_RF_IF_data_in[12]) );
  AN2D0BWP12T U1218 ( .A1(MEMCTRL_RF_IF_data_in[12]), .A2(n1422), .Z(n945) );
  INVD1BWP12T U1219 ( .I(n1119), .ZN(n949) );
  AOI211D1BWP12T U1220 ( .A1(n1116), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_12_), .B(n945), .C(
        n949), .ZN(n1276) );
  ND2D1BWP12T U1221 ( .A1(n1379), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[11]), .ZN(n946) );
  OAI211D1BWP12T U1222 ( .A1(n957), .A2(n1403), .B(n954), .C(n946), .ZN(
        MEMCTRL_RF_IF_data_in[11]) );
  AN2D0BWP12T U1223 ( .A1(MEMCTRL_RF_IF_data_in[11]), .A2(n1422), .Z(n947) );
  AOI211D1BWP12T U1224 ( .A1(n1116), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_11_), .B(n947), .C(
        n949), .ZN(n1672) );
  CKND2D1BWP12T U1225 ( .A1(n1276), .A2(n1672), .ZN(n1032) );
  ND2D1BWP12T U1226 ( .A1(n1379), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[13]), .ZN(n948) );
  OAI211D1BWP12T U1227 ( .A1(n957), .A2(n1387), .B(n954), .C(n948), .ZN(
        MEMCTRL_RF_IF_data_in[13]) );
  AN2D0BWP12T U1228 ( .A1(MEMCTRL_RF_IF_data_in[13]), .A2(n1422), .Z(n950) );
  AOI211D1BWP12T U1229 ( .A1(n1116), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_13_), .B(n950), .C(
        n949), .ZN(n1122) );
  INVD1BWP12T U1230 ( .I(n1122), .ZN(n961) );
  INVD1BWP12T U1231 ( .I(n754), .ZN(n1479) );
  AN2D0BWP12T U1232 ( .A1(n1116), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_14_), .Z(n951) );
  AOI21D1BWP12T U1233 ( .A1(MEMCTRL_RF_IF_data_in[14]), .A2(n1479), .B(n951), 
        .ZN(n992) );
  INVD1BWP12T U1234 ( .I(n992), .ZN(n988) );
  INVD1BWP12T U1235 ( .I(MEM_MEMCTRL_from_mem_data[7]), .ZN(n1372) );
  ND2D1BWP12T U1236 ( .A1(n1379), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[15]), .ZN(n952) );
  OA21D1BWP12T U1237 ( .A1(n957), .A2(n1372), .B(n952), .Z(n953) );
  ND2D1BWP12T U1238 ( .A1(n954), .A2(n953), .ZN(MEMCTRL_RF_IF_data_in[15]) );
  IOA21D1BWP12T U1239 ( .A1(n1116), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_15_), .B(n1119), .ZN(
        n955) );
  AOI21D1BWP12T U1240 ( .A1(n1422), .A2(MEMCTRL_RF_IF_data_in[15]), .B(n955), 
        .ZN(n963) );
  CKND2D1BWP12T U1241 ( .A1(n988), .A2(n963), .ZN(n964) );
  NR2D1BWP12T U1242 ( .A1(n961), .A2(n964), .ZN(n966) );
  INVD1BWP12T U1243 ( .I(n966), .ZN(n989) );
  NR2D1BWP12T U1244 ( .A1(n1032), .A2(n989), .ZN(n1255) );
  ND2D1BWP12T U1245 ( .A1(n1255), .A2(n1656), .ZN(n1306) );
  INVD1BWP12T U1246 ( .I(n1583), .ZN(n1631) );
  TPND2D0BWP12T U1247 ( .A1(n1116), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_9_), .ZN(n958) );
  ND2D1BWP12T U1248 ( .A1(n1119), .A2(n958), .ZN(n959) );
  AOI21D1BWP12T U1249 ( .A1(MEMCTRL_RF_IF_data_in[9]), .A2(n1422), .B(n959), 
        .ZN(n1676) );
  INVD1BWP12T U1250 ( .I(MEM_MEMCTRL_from_mem_data[14]), .ZN(n1541) );
  INVD0BWP12T U1251 ( .I(MEMCTRL_RF_IF_data_in[6]), .ZN(n1563) );
  INVD1BWP12T U1252 ( .I(IF_DEC_instruction[6]), .ZN(n1617) );
  INVD1BWP12T U1253 ( .I(MEM_MEMCTRL_from_mem_data[15]), .ZN(n1540) );
  INVD1BWP12T U1254 ( .I(MEMCTRL_RF_IF_data_in[7]), .ZN(n1562) );
  NR2XD0BWP12T U1255 ( .A1(n1617), .A2(IF_DEC_instruction[7]), .ZN(n1582) );
  INVD1BWP12T U1256 ( .I(n1276), .ZN(n1056) );
  INVD1BWP12T U1257 ( .I(n1656), .ZN(n1628) );
  CKND2D1BWP12T U1258 ( .A1(n1628), .A2(n1672), .ZN(n1300) );
  NR3XD0BWP12T U1259 ( .A1(n1056), .A2(n989), .A3(n1300), .ZN(n1600) );
  OA31XD0BWP12T U1260 ( .A1(n1676), .A2(n1582), .A3(n1631), .B(n1600), .Z(n960) );
  INVD1BWP12T U1261 ( .I(n963), .ZN(n987) );
  NR2D1BWP12T U1262 ( .A1(n988), .A2(n987), .ZN(n996) );
  TPND2D0BWP12T U1263 ( .A1(n1122), .A2(n996), .ZN(n1608) );
  INVD1BWP12T U1264 ( .I(n1608), .ZN(n1604) );
  NR2D1BWP12T U1265 ( .A1(n960), .A2(n1604), .ZN(n1575) );
  OAI21D0BWP12T U1266 ( .A1(n1306), .A2(n1631), .B(n1575), .ZN(n1593) );
  INVD1BWP12T U1267 ( .I(MEM_MEMCTRL_from_mem_data[8]), .ZN(n1546) );
  INVD1BWP12T U1268 ( .I(MEMCTRL_RF_IF_data_in[0]), .ZN(n1568) );
  NR2D1BWP12T U1269 ( .A1(n1672), .A2(n1056), .ZN(n990) );
  INVD1BWP12T U1270 ( .I(n996), .ZN(n1121) );
  NR2D1BWP12T U1271 ( .A1(n1121), .A2(n1122), .ZN(n1573) );
  INVD1BWP12T U1272 ( .I(n1573), .ZN(n1624) );
  TPNR2D0BWP12T U1273 ( .A1(n990), .A2(n1624), .ZN(n1576) );
  NR2XD0BWP12T U1274 ( .A1(n961), .A2(n1056), .ZN(n962) );
  CKND2D1BWP12T U1275 ( .A1(n962), .A2(n987), .ZN(n965) );
  NR2XD0BWP12T U1276 ( .A1(n965), .A2(n992), .ZN(n1653) );
  INVD1BWP12T U1277 ( .I(n1653), .ZN(n1670) );
  NR2D1BWP12T U1278 ( .A1(n963), .A2(n1122), .ZN(n967) );
  CKND2D1BWP12T U1279 ( .A1(n992), .A2(n967), .ZN(n1327) );
  NR2D1BWP12T U1280 ( .A1(n1056), .A2(n1327), .ZN(n1636) );
  INVD1BWP12T U1281 ( .I(n1636), .ZN(n998) );
  CKND2D0BWP12T U1282 ( .A1(n1670), .A2(n998), .ZN(n1044) );
  NR2D1BWP12T U1283 ( .A1(n1576), .A2(n1044), .ZN(n1590) );
  INVD1BWP12T U1284 ( .I(n1619), .ZN(n1632) );
  NR2D1BWP12T U1285 ( .A1(n965), .A2(n988), .ZN(n1657) );
  NR2D1BWP12T U1286 ( .A1(n1632), .A2(n1657), .ZN(n1082) );
  CKND2D1BWP12T U1287 ( .A1(n966), .A2(n1056), .ZN(n1071) );
  CKND2D1BWP12T U1288 ( .A1(n1082), .A2(n1071), .ZN(n1045) );
  NR2D1BWP12T U1289 ( .A1(n1276), .A2(n1327), .ZN(n1000) );
  AOI32D1BWP12T U1290 ( .A1(n1672), .A2(n1676), .A3(n1583), .B1(n1656), .B2(
        n1676), .ZN(n968) );
  ND2D1BWP12T U1291 ( .A1(n967), .A2(n988), .ZN(n993) );
  CKND0BWP12T U1292 ( .I(n993), .ZN(n1043) );
  AOI22D1BWP12T U1293 ( .A1(n1000), .A2(n968), .B1(n1043), .B2(n990), .ZN(
        n1226) );
  NR2D1BWP12T U1294 ( .A1(irdecode_inst1_itstate_6_), .A2(
        irdecode_inst1_itstate_7_), .ZN(n985) );
  AOI22D0BWP12T U1295 ( .A1(irdecode_inst1_itstate_6_), .A2(RF_OUT_v), .B1(
        RF_OUT_c), .B2(n985), .ZN(n970) );
  INVD1BWP12T U1296 ( .I(RF_OUT_n), .ZN(n974) );
  TPOAI21D0BWP12T U1297 ( .A1(irdecode_inst1_itstate_6_), .A2(n1293), .B(
        irdecode_inst1_itstate_7_), .ZN(n969) );
  INVD1BWP12T U1298 ( .I(irdecode_inst1_itstate_5_), .ZN(n1485) );
  AOI21D1BWP12T U1299 ( .A1(n970), .A2(n969), .B(n1485), .ZN(n983) );
  INVD1BWP12T U1300 ( .I(irdecode_inst1_itstate_6_), .ZN(n1486) );
  AOI22D0BWP12T U1301 ( .A1(irdecode_inst1_itstate_6_), .A2(RF_OUT_n), .B1(
        RF_OUT_z), .B2(n1486), .ZN(n973) );
  INR2XD0BWP12T U1302 ( .A1(RF_OUT_c), .B1(RF_OUT_z), .ZN(n1292) );
  INVD1BWP12T U1303 ( .I(RF_OUT_z), .ZN(n979) );
  ND2D1BWP12T U1304 ( .A1(n1293), .A2(n979), .ZN(n1289) );
  NR2D1BWP12T U1305 ( .A1(n1289), .A2(n1486), .ZN(n971) );
  TPAOI31D0BWP12T U1306 ( .A1(n1485), .A2(n1292), .A3(n1486), .B(n971), .ZN(
        n972) );
  INVD1BWP12T U1307 ( .I(irdecode_inst1_itstate_7_), .ZN(n1484) );
  OAI32D0BWP12T U1308 ( .A1(irdecode_inst1_itstate_7_), .A2(
        irdecode_inst1_itstate_5_), .A3(n973), .B1(n972), .B2(n1484), .ZN(n982) );
  TPND2D0BWP12T U1309 ( .A1(irdecode_inst1_itstate_6_), .A2(n1289), .ZN(n977)
         );
  OR2XD0BWP12T U1310 ( .A1(n1292), .A2(irdecode_inst1_itstate_6_), .Z(n976) );
  TPND2D0BWP12T U1311 ( .A1(irdecode_inst1_itstate_6_), .A2(n974), .ZN(n975)
         );
  AOI32D1BWP12T U1312 ( .A1(n977), .A2(irdecode_inst1_itstate_7_), .A3(n976), 
        .B1(n975), .B2(n1484), .ZN(n978) );
  RCAOI211D0BWP12T U1313 ( .A1(n985), .A2(n979), .B(irdecode_inst1_itstate_5_), 
        .C(n978), .ZN(n980) );
  OAI21D1BWP12T U1314 ( .A1(n983), .A2(n980), .B(irdecode_inst1_itstate_4_), 
        .ZN(n981) );
  OAI31D1BWP12T U1315 ( .A1(n983), .A2(irdecode_inst1_itstate_4_), .A3(n982), 
        .B(n981), .ZN(n986) );
  NR2D1BWP12T U1316 ( .A1(irdecode_inst1_itstate_1_), .A2(
        irdecode_inst1_itstate_0_), .ZN(n1333) );
  NR4D0BWP12T U1317 ( .A1(irdecode_inst1_itstate_5_), .A2(
        irdecode_inst1_itstate_4_), .A3(irdecode_inst1_itstate_2_), .A4(
        irdecode_inst1_itstate_3_), .ZN(n984) );
  ND3D1BWP12T U1318 ( .A1(n985), .A2(n1333), .A3(n984), .ZN(n1089) );
  ND2D1BWP12T U1319 ( .A1(n986), .A2(n1089), .ZN(n1072) );
  CKND2D1BWP12T U1320 ( .A1(n1226), .A2(n1072), .ZN(n1233) );
  NR2D1BWP12T U1321 ( .A1(n1045), .A2(n1233), .ZN(n997) );
  ND3D1BWP12T U1322 ( .A1(n1122), .A2(n987), .A3(n1056), .ZN(n991) );
  NR2D1BWP12T U1323 ( .A1(n988), .A2(n991), .ZN(n1665) );
  INVD1BWP12T U1324 ( .I(n990), .ZN(n1607) );
  NR2D1BWP12T U1325 ( .A1(n1607), .A2(n989), .ZN(n1674) );
  NR2D1BWP12T U1326 ( .A1(n1665), .A2(n1674), .ZN(n999) );
  INVD1BWP12T U1327 ( .I(n999), .ZN(n1166) );
  INVD1BWP12T U1328 ( .I(n1676), .ZN(n1664) );
  ND3XD0BWP12T U1329 ( .A1(n1583), .A2(n1600), .A3(n1664), .ZN(n1088) );
  INR2XD0BWP12T U1330 ( .A1(n1676), .B1(n1583), .ZN(n1581) );
  INVD1BWP12T U1331 ( .I(n1581), .ZN(n1290) );
  OAI21D1BWP12T U1332 ( .A1(n1582), .A2(n1088), .B(n1227), .ZN(n1577) );
  INR3XD0BWP12T U1333 ( .A1(n997), .B1(n1166), .B2(n1577), .ZN(n1264) );
  NR2D1BWP12T U1334 ( .A1(n992), .A2(n991), .ZN(n1303) );
  NR2D1BWP12T U1335 ( .A1(n993), .A2(n1032), .ZN(n1301) );
  NR2D1BWP12T U1336 ( .A1(n1303), .A2(n1301), .ZN(n1639) );
  INVD1BWP12T U1337 ( .I(n1639), .ZN(n1261) );
  NR2D1BWP12T U1338 ( .A1(n1276), .A2(n993), .ZN(n1612) );
  INR2D1BWP12T U1339 ( .A1(irdecode_inst1_N912), .B1(irdecode_inst1_N906), 
        .ZN(n1120) );
  INVD1BWP12T U1340 ( .I(n1120), .ZN(n994) );
  INR2D2BWP12T U1341 ( .A1(n1359), .B1(n995), .ZN(n1682) );
  NR2D1BWP12T U1342 ( .A1(n1331), .A2(n1670), .ZN(n1595) );
  ND2D1BWP12T U1343 ( .A1(n1661), .A2(n1328), .ZN(n1509) );
  INVD1BWP12T U1344 ( .I(n1509), .ZN(n1501) );
  NR2D1BWP12T U1345 ( .A1(n996), .A2(n1255), .ZN(n1278) );
  ND3D1BWP12T U1346 ( .A1(n1639), .A2(n997), .A3(n1278), .ZN(n1212) );
  ND2D1BWP12T U1347 ( .A1(n999), .A2(n998), .ZN(n1513) );
  CKND2D1BWP12T U1348 ( .A1(n1583), .A2(n1676), .ZN(n1579) );
  INR3D0BWP12T U1349 ( .A1(n1000), .B1(n1300), .B2(n1579), .ZN(n1601) );
  INVD1BWP12T U1350 ( .I(n1601), .ZN(n1263) );
  IND2D1BWP12T U1351 ( .A1(n1513), .B1(n1263), .ZN(n1634) );
  INVD1BWP12T U1352 ( .I(n1634), .ZN(n1535) );
  CKND2D0BWP12T U1353 ( .A1(n1672), .A2(n1612), .ZN(n1001) );
  ND2D1BWP12T U1354 ( .A1(n1535), .A2(n1001), .ZN(n1037) );
  INVD1BWP12T U1355 ( .I(IF_DEC_instruction[7]), .ZN(n1602) );
  NR4D0BWP12T U1356 ( .A1(irdecode_inst1_N702), .A2(irdecode_inst1_N703), .A3(
        irdecode_inst1_N701), .A4(irdecode_inst1_N706), .ZN(n1003) );
  INVD1BWP12T U1357 ( .I(irdecode_inst1_N704), .ZN(n1067) );
  ND3D1BWP12T U1358 ( .A1(n1602), .A2(n1003), .A3(n1067), .ZN(n1007) );
  NR2D1BWP12T U1359 ( .A1(irdecode_inst1_N707), .A2(irdecode_inst1_N705), .ZN(
        n1004) );
  INVD1BWP12T U1360 ( .I(irdecode_inst1_N706), .ZN(n1140) );
  ND2D1BWP12T U1361 ( .A1(n1004), .A2(n1140), .ZN(n1066) );
  NR2D1BWP12T U1362 ( .A1(irdecode_inst1_N704), .A2(n1066), .ZN(n1005) );
  CKND2D1BWP12T U1363 ( .A1(irdecode_inst1_N703), .A2(n1005), .ZN(n1135) );
  NR4D0BWP12T U1364 ( .A1(irdecode_inst1_N702), .A2(irdecode_inst1_N701), .A3(
        IF_DEC_instruction[7]), .A4(n1135), .ZN(n1136) );
  INVD1BWP12T U1365 ( .I(irdecode_inst1_N707), .ZN(n1139) );
  NR3D1BWP12T U1366 ( .A1(irdecode_inst1_N705), .A2(n1139), .A3(n1007), .ZN(
        n1145) );
  NR2D0BWP12T U1367 ( .A1(irdecode_inst1_N701), .A2(IF_DEC_instruction[7]), 
        .ZN(n1002) );
  IND3D1BWP12T U1368 ( .A1(irdecode_inst1_N703), .B1(irdecode_inst1_N702), 
        .B2(n1005), .ZN(n1065) );
  INR2D1BWP12T U1369 ( .A1(n1002), .B1(n1065), .ZN(n1137) );
  NR2D1BWP12T U1370 ( .A1(irdecode_inst1_N702), .A2(irdecode_inst1_N703), .ZN(
        n1006) );
  AN2XD1BWP12T U1371 ( .A1(n1004), .A2(n1003), .Z(n1008) );
  ND3D1BWP12T U1372 ( .A1(n1602), .A2(irdecode_inst1_N704), .A3(n1008), .ZN(
        n1143) );
  IND3D1BWP12T U1373 ( .A1(n1137), .B1(n1146), .B2(n1143), .ZN(n1069) );
  NR4D0BWP12T U1374 ( .A1(n1144), .A2(n1136), .A3(n1145), .A4(n1069), .ZN(
        n1171) );
  AN3XD1BWP12T U1375 ( .A1(n1006), .A2(irdecode_inst1_N701), .A3(n1005), .Z(
        n1153) );
  ND2D1BWP12T U1376 ( .A1(n1602), .A2(n1153), .ZN(n1009) );
  CKND2D1BWP12T U1377 ( .A1(n1009), .A2(n1171), .ZN(n1138) );
  NR2D1BWP12T U1378 ( .A1(n1138), .A2(irdecode_inst1_N707), .ZN(n1141) );
  INVD1BWP12T U1379 ( .I(n1141), .ZN(n1134) );
  NR2D1BWP12T U1380 ( .A1(n1007), .A2(n1134), .ZN(n1201) );
  ND3D0BWP12T U1381 ( .A1(n1008), .A2(IF_DEC_instruction[7]), .A3(n1067), .ZN(
        n1068) );
  ND2D1BWP12T U1382 ( .A1(n1009), .A2(n1068), .ZN(n1174) );
  NR2D1BWP12T U1383 ( .A1(n1201), .A2(n1174), .ZN(n1156) );
  ND2D1BWP12T U1384 ( .A1(n1171), .A2(n1156), .ZN(n1214) );
  NR3D1BWP12T U1385 ( .A1(irdecode_inst1_N541), .A2(irdecode_inst1_N540), .A3(
        irdecode_inst1_N539), .ZN(n1012) );
  CKND2D1BWP12T U1386 ( .A1(n1583), .A2(n1012), .ZN(n1011) );
  NR2D1BWP12T U1387 ( .A1(irdecode_inst1_N542), .A2(n1011), .ZN(n1015) );
  INVD1BWP12T U1388 ( .I(irdecode_inst1_N543), .ZN(n1026) );
  CKND2D1BWP12T U1389 ( .A1(n1015), .A2(n1026), .ZN(n1014) );
  INVD1BWP12T U1390 ( .I(irdecode_inst1_N544), .ZN(n1016) );
  INVD1BWP12T U1391 ( .I(irdecode_inst1_N546), .ZN(n1062) );
  IND4D1BWP12T U1392 ( .A1(n1014), .B1(n1016), .B2(n1062), .B3(
        irdecode_inst1_N545), .ZN(n1019) );
  NR2D1BWP12T U1393 ( .A1(irdecode_inst1_N545), .A2(irdecode_inst1_N546), .ZN(
        n1050) );
  ND2D1BWP12T U1394 ( .A1(n1016), .A2(n1050), .ZN(n1027) );
  NR2D1BWP12T U1395 ( .A1(n1027), .A2(irdecode_inst1_N543), .ZN(n1010) );
  INR2D1BWP12T U1396 ( .A1(n1010), .B1(irdecode_inst1_N542), .ZN(n1013) );
  ND2D1BWP12T U1397 ( .A1(n1013), .A2(irdecode_inst1_N541), .ZN(n1060) );
  NR4D0BWP12T U1398 ( .A1(irdecode_inst1_N540), .A2(irdecode_inst1_N539), .A3(
        n1060), .A4(n1631), .ZN(n1025) );
  ND2D1BWP12T U1399 ( .A1(irdecode_inst1_N542), .A2(n1010), .ZN(n1499) );
  NR2D1BWP12T U1400 ( .A1(n1499), .A2(n1011), .ZN(n1021) );
  NR3D1BWP12T U1401 ( .A1(irdecode_inst1_N539), .A2(n1510), .A3(n1631), .ZN(
        n1018) );
  ND3D1BWP12T U1402 ( .A1(n1013), .A2(n1012), .A3(n1631), .ZN(n1158) );
  OAI21D1BWP12T U1403 ( .A1(n1631), .A2(n1061), .B(n1158), .ZN(n1023) );
  NR2D1BWP12T U1404 ( .A1(n1014), .A2(irdecode_inst1_N545), .ZN(n1017) );
  NR2D1BWP12T U1405 ( .A1(n1027), .A2(n1026), .ZN(n1049) );
  ND2D1BWP12T U1406 ( .A1(n1049), .A2(n1015), .ZN(n1064) );
  NR3XD0BWP12T U1407 ( .A1(n1018), .A2(n1023), .A3(n1024), .ZN(n1660) );
  ND3D1BWP12T U1408 ( .A1(irdecode_inst1_N546), .A2(n1017), .A3(n1016), .ZN(
        n1020) );
  NR2D1BWP12T U1409 ( .A1(irdecode_inst1_N540), .A2(irdecode_inst1_N539), .ZN(
        n1052) );
  ND2D1BWP12T U1410 ( .A1(n1499), .A2(n1060), .ZN(n1047) );
  INVD1BWP12T U1411 ( .I(n1018), .ZN(n1157) );
  IND4D1BWP12T U1412 ( .A1(n1021), .B1(n1020), .B2(n1157), .B3(n1019), .ZN(
        n1022) );
  NR4D0BWP12T U1413 ( .A1(n1025), .A2(n1024), .A3(n1023), .A4(n1022), .ZN(
        n1054) );
  IND3D1BWP12T U1414 ( .A1(n1027), .B1(n1054), .B2(n1026), .ZN(n1048) );
  NR2D1BWP12T U1415 ( .A1(n1047), .A2(n1048), .ZN(n1161) );
  ND2D1BWP12T U1416 ( .A1(n1052), .A2(n1161), .ZN(n1200) );
  ND2D1BWP12T U1417 ( .A1(n1055), .A2(n1200), .ZN(n1210) );
  INVD1BWP12T U1418 ( .I(n1682), .ZN(n1527) );
  INR2D1BWP12T U1419 ( .A1(n1527), .B1(n1328), .ZN(n1280) );
  INVD1BWP12T U1420 ( .I(n1280), .ZN(n1273) );
  INVD1BWP12T U1421 ( .I(irdecode_inst1_next_step_1_), .ZN(irdecode_inst1_N907) );
  INVD1BWP12T U1422 ( .I(n1612), .ZN(n1638) );
  AOI21D2BWP12T U1423 ( .A1(n1682), .A2(irdecode_inst1_step[0]), .B(n1028), 
        .ZN(irdecode_inst1_N910) );
  INVD2BWP12T U1424 ( .I(irdecode_inst1_N910), .ZN(irdecode_inst1_next_step_0_) );
  NR3D1BWP12T U1425 ( .A1(irdecode_inst1_N907), .A2(n1638), .A3(
        irdecode_inst1_next_step_0_), .ZN(n1041) );
  NR2D2BWP12T U1426 ( .A1(n1261), .A2(n1041), .ZN(n1625) );
  NR2D0BWP12T U1427 ( .A1(n1501), .A2(n1280), .ZN(n1038) );
  INR2D1BWP12T U1428 ( .A1(n1072), .B1(n1331), .ZN(n1578) );
  INVD1BWP12T U1429 ( .I(n1578), .ZN(n1679) );
  ND2D1BWP12T U1430 ( .A1(n1578), .A2(IF_DEC_instruction[7]), .ZN(n1529) );
  INVD1BWP12T U1431 ( .I(n1529), .ZN(n1536) );
  INVD0BWP12T U1432 ( .I(n1625), .ZN(n1029) );
  AOI22D0BWP12T U1433 ( .A1(n1536), .A2(n1029), .B1(n1682), .B2(
        DEC_RF_offset_b[8]), .ZN(n1030) );
  OAI31D0BWP12T U1434 ( .A1(n1617), .A2(n1679), .A3(n1535), .B(n1030), .ZN(
        n801) );
  INVD1BWP12T U1435 ( .I(MEM_MEMCTRL_from_mem_data[10]), .ZN(n1544) );
  INVD1BWP12T U1436 ( .I(MEMCTRL_RF_IF_data_in[2]), .ZN(n1566) );
  INVD1BWP12T U1437 ( .I(MEM_MEMCTRL_from_mem_data[13]), .ZN(n1542) );
  INVD0BWP12T U1438 ( .I(MEMCTRL_RF_IF_data_in[5]), .ZN(n1560) );
  INVD1BWP12T U1439 ( .I(IF_DEC_instruction[5]), .ZN(n1618) );
  OAI22D1BWP12T U1440 ( .A1(n1535), .A2(n1618), .B1(n1617), .B2(n1625), .ZN(
        n1031) );
  AO222D0BWP12T U1441 ( .A1(n1031), .A2(n1578), .B1(n1573), .B2(n1536), .C1(
        n1682), .C2(DEC_RF_offset_b[7]), .Z(n802) );
  INVD1BWP12T U1442 ( .I(DEC_RF_operand_a[0]), .ZN(n1040) );
  INVD1BWP12T U1443 ( .I(MEM_MEMCTRL_from_mem_data[11]), .ZN(n1543) );
  INVD1BWP12T U1444 ( .I(MEMCTRL_RF_IF_data_in[3]), .ZN(n1561) );
  CKND0BWP12T U1445 ( .I(IF_DEC_instruction[3]), .ZN(n1626) );
  ND2XD0BWP12T U1446 ( .A1(n1071), .A2(n1608), .ZN(n1239) );
  INVD1BWP12T U1447 ( .I(n1239), .ZN(n1077) );
  ND2XD0BWP12T U1448 ( .A1(n1077), .A2(n1082), .ZN(n1258) );
  INVD1BWP12T U1449 ( .I(n1258), .ZN(n1643) );
  TPNR2D0BWP12T U1450 ( .A1(n1653), .A2(n1573), .ZN(n1637) );
  OAI21D0BWP12T U1451 ( .A1(n1583), .A2(n1637), .B(n1057), .ZN(n1034) );
  OAI22D0BWP12T U1452 ( .A1(n1306), .A2(n1676), .B1(n1624), .B2(n1032), .ZN(
        n1644) );
  INR2D1BWP12T U1453 ( .A1(n1072), .B1(n1644), .ZN(n1225) );
  CKND2D0BWP12T U1454 ( .A1(n1639), .A2(n1225), .ZN(n1033) );
  RCAOI211D0BWP12T U1455 ( .A1(n1255), .A2(IF_DEC_instruction[0]), .B(n1034), 
        .C(n1033), .ZN(n1035) );
  OAI211D1BWP12T U1456 ( .A1(n1626), .A2(n1643), .B(n1035), .C(n1226), .ZN(
        n1036) );
  OAI21D0BWP12T U1457 ( .A1(n1037), .A2(n1036), .B(n1328), .ZN(n1039) );
  OAI211D0BWP12T U1458 ( .A1(n1527), .A2(n1040), .B(n1039), .C(n1038), .ZN(
        n811) );
  TPOAI21D0BWP12T U1459 ( .A1(n1301), .A2(n1041), .B(n1578), .ZN(n1517) );
  AN2XD1BWP12T U1460 ( .A1(n1303), .A2(n1536), .Z(n1514) );
  INVD1BWP12T U1461 ( .I(n1514), .ZN(n1512) );
  TPND2D0BWP12T U1462 ( .A1(n1682), .A2(DEC_RF_offset_b[10]), .ZN(n1042) );
  OAI211D0BWP12T U1463 ( .A1(n1676), .A2(n1517), .B(n1512), .C(n1042), .ZN(
        n799) );
  OAI211D0BWP12T U1464 ( .A1(n1043), .A2(n1573), .B(n1672), .C(n1056), .ZN(
        n1046) );
  NR4D0BWP12T U1465 ( .A1(n1261), .A2(n1045), .A3(n1166), .A4(n1044), .ZN(
        n1091) );
  OAI211D1BWP12T U1466 ( .A1(n1579), .A2(n1306), .B(n1046), .C(n1091), .ZN(
        n1609) );
  INVD0BWP12T U1467 ( .I(n1050), .ZN(n1211) );
  CKND1BWP12T U1468 ( .I(n1047), .ZN(n1507) );
  NR2D0BWP12T U1469 ( .A1(n1507), .A2(n1048), .ZN(n1053) );
  CKND0BWP12T U1470 ( .I(n1161), .ZN(n1051) );
  CKND2D1BWP12T U1471 ( .A1(n1049), .A2(n1054), .ZN(n1493) );
  TPND3D0BWP12T U1472 ( .A1(n1050), .A2(irdecode_inst1_N544), .A3(n1054), .ZN(
        n1489) );
  OAI211D1BWP12T U1473 ( .A1(n1052), .A2(n1051), .B(n1493), .C(n1489), .ZN(
        n1662) );
  RCAOI211D0BWP12T U1474 ( .A1(n1054), .A2(n1211), .B(n1053), .C(n1662), .ZN(
        n1649) );
  INVD1BWP12T U1475 ( .I(n1661), .ZN(n1648) );
  AOI21D1BWP12T U1476 ( .A1(n1055), .A2(n1649), .B(n1648), .ZN(n1603) );
  INVD1BWP12T U1477 ( .I(n1603), .ZN(n1125) );
  INVD1BWP12T U1478 ( .I(n1672), .ZN(n1677) );
  ND2D1BWP12T U1479 ( .A1(n1056), .A2(n1677), .ZN(n1530) );
  NR2D0BWP12T U1480 ( .A1(n1121), .A2(n1530), .ZN(n1090) );
  TPNR2D0BWP12T U1481 ( .A1(n1601), .A2(n1090), .ZN(n1058) );
  IND4D1BWP12T U1482 ( .A1(n1609), .B1(n1125), .B2(n1058), .B3(n1057), .ZN(
        n1059) );
  AO22XD0BWP12T U1483 ( .A1(n1059), .A2(n1578), .B1(n1682), .B2(
        DEC_ALU_alu_opcode[4]), .Z(n848) );
  AN3D0BWP12T U1484 ( .A1(n1061), .A2(n1060), .A3(n1200), .Z(n1159) );
  CKND2D0BWP12T U1485 ( .A1(irdecode_inst1_N545), .A2(n1062), .ZN(n1063) );
  ND4D1BWP12T U1486 ( .A1(n1159), .A2(n1064), .A3(n1063), .A4(n1493), .ZN(
        n1185) );
  CKND0BWP12T U1487 ( .I(IF_DEC_instruction[0]), .ZN(n1647) );
  NR2D0BWP12T U1488 ( .A1(n1664), .A2(n1071), .ZN(n1275) );
  INVD1BWP12T U1489 ( .I(n1070), .ZN(n1666) );
  CKND2D0BWP12T U1490 ( .A1(n1666), .A2(n1328), .ZN(n1164) );
  NR2D1BWP12T U1491 ( .A1(n1065), .A2(n1134), .ZN(n1597) );
  NR3D1BWP12T U1492 ( .A1(n1067), .A2(n1066), .A3(n1134), .ZN(n1494) );
  CKND0BWP12T U1493 ( .I(n1494), .ZN(n1142) );
  INVD0BWP12T U1494 ( .I(n1665), .ZN(n1194) );
  CKND2D1BWP12T U1495 ( .A1(n1070), .A2(n1194), .ZN(n1148) );
  NR2XD0BWP12T U1496 ( .A1(n1071), .A2(n1676), .ZN(n1655) );
  INVD1BWP12T U1497 ( .I(n1655), .ZN(n1094) );
  NR2D1BWP12T U1498 ( .A1(n1300), .A2(n1094), .ZN(n1671) );
  AOI21D0BWP12T U1499 ( .A1(n1672), .A2(n1148), .B(n1671), .ZN(n1176) );
  ND4D0BWP12T U1500 ( .A1(n1639), .A2(n1226), .A3(n1072), .A4(n1638), .ZN(
        n1079) );
  INR4D0BWP12T U1501 ( .A1(n1278), .B1(n1636), .B2(n1601), .B3(n1079), .ZN(
        n1181) );
  AN2XD1BWP12T U1502 ( .A1(n1176), .A2(n1181), .Z(n1205) );
  NR2XD0BWP12T U1503 ( .A1(n1158), .A2(n1509), .ZN(n1681) );
  INVD1BWP12T U1504 ( .I(n1595), .ZN(n1503) );
  AOI21D0BWP12T U1505 ( .A1(n1509), .A2(n1503), .B(n1677), .ZN(n1165) );
  AOI211D0BWP12T U1506 ( .A1(n1682), .A2(DEC_RF_memory_write_to_reg[0]), .B(
        n1681), .C(n1165), .ZN(n1074) );
  CKND0BWP12T U1507 ( .I(n1300), .ZN(n1195) );
  NR2D1BWP12T U1508 ( .A1(n1195), .A2(n1094), .ZN(n1675) );
  AOI22D0BWP12T U1509 ( .A1(n1675), .A2(IF_DEC_instruction[0]), .B1(n1631), 
        .B2(n1166), .ZN(n1073) );
  AOI32D0BWP12T U1510 ( .A1(n1205), .A2(n1074), .A3(n1073), .B1(n1331), .B2(
        n1074), .ZN(n1075) );
  AO211D0BWP12T U1511 ( .A1(n1501), .A2(n1185), .B(n1184), .C(n1075), .Z(n824)
         );
  INVD1BWP12T U1512 ( .I(MEM_MEMCTRL_from_mem_data[9]), .ZN(n1545) );
  INVD0BWP12T U1513 ( .I(MEMCTRL_RF_IF_data_in[1]), .ZN(n1565) );
  INVD1BWP12T U1514 ( .I(DEC_RF_operand_b[1]), .ZN(n1078) );
  INVD1BWP12T U1515 ( .I(MEM_MEMCTRL_from_mem_data[12]), .ZN(n1548) );
  INVD1BWP12T U1516 ( .I(MEMCTRL_RF_IF_data_in[4]), .ZN(n1564) );
  OAI21D1BWP12T U1517 ( .A1(n1530), .A2(n1656), .B(n1604), .ZN(n1570) );
  NR4D0BWP12T U1518 ( .A1(n1661), .A2(n1612), .A3(n1261), .A4(n1634), .ZN(
        n1246) );
  ND4D1BWP12T U1519 ( .A1(n1082), .A2(n1570), .A3(n1637), .A4(n1246), .ZN(
        n1234) );
  AOI21D0BWP12T U1520 ( .A1(n1255), .A2(IF_DEC_instruction[4]), .B(n1234), 
        .ZN(n1076) );
  OAI222D0BWP12T U1521 ( .A1(n1078), .A2(n1527), .B1(n1529), .B2(n1077), .C1(
        n1679), .C2(n1076), .ZN(n843) );
  CKND0BWP12T U1522 ( .I(DEC_ALU_alu_opcode[2]), .ZN(n1550) );
  TPND2D0BWP12T U1523 ( .A1(n1670), .A2(n1648), .ZN(n1521) );
  NR3D0BWP12T U1524 ( .A1(n1521), .A2(n1634), .A3(n1079), .ZN(n1279) );
  NR2D0BWP12T U1525 ( .A1(n1581), .A2(n1306), .ZN(n1080) );
  AOI211D0BWP12T U1526 ( .A1(n1600), .A2(n1631), .B(n1080), .C(n1576), .ZN(
        n1081) );
  ND4D0BWP12T U1527 ( .A1(n1276), .A2(n1082), .A3(n1279), .A4(n1081), .ZN(
        n1083) );
  CKND2D0BWP12T U1528 ( .A1(n1083), .A2(n1328), .ZN(n1084) );
  OAI211D0BWP12T U1529 ( .A1(n1527), .A2(n1550), .B(n1084), .C(n1273), .ZN(
        n846) );
  HA1D0BWP12T U1530 ( .A(n1086), .B(RF_pc_out[21]), .CO(n1130), .S(n1087) );
  OAI22D0BWP12T U1531 ( .A1(n1227), .A2(n1679), .B1(n1088), .B2(n1529), .ZN(
        n1589) );
  NR2D0BWP12T U1532 ( .A1(n1276), .A2(n1624), .ZN(n1586) );
  TPNR2D0BWP12T U1533 ( .A1(n1331), .A2(n1089), .ZN(n1584) );
  CKND2D1BWP12T U1534 ( .A1(n1612), .A2(n1677), .ZN(n1224) );
  AN4D0BWP12T U1535 ( .A1(n1091), .A2(n1648), .A3(n1224), .A4(n1306), .Z(n1092) );
  CKND0BWP12T U1536 ( .I(DEC_IF_stall_to_instructionfetch), .ZN(n1115) );
  OAI22D0BWP12T U1537 ( .A1(n1092), .A2(n1679), .B1(n1115), .B2(n1527), .ZN(
        n845) );
  TPND2D0BWP12T U1538 ( .A1(n1682), .A2(
        DEC_MEMCTRL_memorycontroller_sign_extend), .ZN(n1093) );
  OAI31D0BWP12T U1539 ( .A1(n1672), .A2(n1679), .A3(n1094), .B(n1093), .ZN(
        n839) );
  INVD1BWP12T U1540 ( .I(RF_pc_out[1]), .ZN(n1370) );
  MAOI22D0BWP12T U1541 ( .A1(RF_pc_out[2]), .A2(n1370), .B1(RF_pc_out[2]), 
        .B2(n1370), .ZN(n1421) );
  OR4D0BWP12T U1542 ( .A1(RF_pc_out[15]), .A2(RF_pc_out[18]), .A3(
        RF_pc_out[20]), .A4(RF_pc_out[19]), .Z(n1095) );
  NR4D0BWP12T U1543 ( .A1(n1421), .A2(RF_pc_out[17]), .A3(RF_pc_out[16]), .A4(
        n1095), .ZN(n1113) );
  NR4D0BWP12T U1544 ( .A1(RF_pc_out[14]), .A2(RF_pc_out[13]), .A3(
        RF_pc_out[27]), .A4(RF_pc_out[26]), .ZN(n1112) );
  NR4D0BWP12T U1545 ( .A1(RF_pc_out[25]), .A2(RF_pc_out[24]), .A3(
        RF_pc_out[23]), .A4(RF_pc_out[22]), .ZN(n1111) );
  NR4D0BWP12T U1546 ( .A1(RF_pc_out[4]), .A2(RF_pc_out[3]), .A3(RF_pc_out[2]), 
        .A4(RF_pc_out[1]), .ZN(n1100) );
  IND2D1BWP12T U1547 ( .A1(RF_pc_out[5]), .B1(n1100), .ZN(n1104) );
  NR2D1BWP12T U1548 ( .A1(RF_pc_out[6]), .A2(n1104), .ZN(n1102) );
  IND2D1BWP12T U1549 ( .A1(RF_pc_out[7]), .B1(n1102), .ZN(n1105) );
  NR2D1BWP12T U1550 ( .A1(RF_pc_out[8]), .A2(n1105), .ZN(n1103) );
  IND2D1BWP12T U1551 ( .A1(RF_pc_out[9]), .B1(n1103), .ZN(n1098) );
  NR2XD0BWP12T U1552 ( .A1(RF_pc_out[10]), .A2(n1098), .ZN(n1097) );
  IND2XD0BWP12T U1553 ( .A1(RF_pc_out[11]), .B1(n1097), .ZN(n1096) );
  MOAI22D0BWP12T U1554 ( .A1(RF_pc_out[12]), .A2(n1096), .B1(RF_pc_out[12]), 
        .B2(n1096), .ZN(n1151) );
  MAOI22D0BWP12T U1555 ( .A1(RF_pc_out[11]), .A2(n1097), .B1(RF_pc_out[11]), 
        .B2(n1097), .ZN(n1189) );
  MOAI22D0BWP12T U1556 ( .A1(RF_pc_out[10]), .A2(n1098), .B1(RF_pc_out[10]), 
        .B2(n1098), .ZN(n1191) );
  NR4D0BWP12T U1557 ( .A1(n1151), .A2(n1189), .A3(n1191), .A4(RF_pc_out[28]), 
        .ZN(n1109) );
  NR4D0BWP12T U1558 ( .A1(RF_pc_out[31]), .A2(RF_pc_out[30]), .A3(
        RF_pc_out[21]), .A4(RF_pc_out[29]), .ZN(n1108) );
  NR2D0BWP12T U1559 ( .A1(RF_pc_out[2]), .A2(RF_pc_out[1]), .ZN(n1099) );
  MAOI22D0BWP12T U1560 ( .A1(RF_pc_out[3]), .A2(n1099), .B1(RF_pc_out[3]), 
        .B2(n1099), .ZN(n1218) );
  MAOI22D0BWP12T U1561 ( .A1(RF_pc_out[5]), .A2(n1100), .B1(RF_pc_out[5]), 
        .B2(n1100), .ZN(n1190) );
  NR3D0BWP12T U1562 ( .A1(RF_pc_out[3]), .A2(RF_pc_out[2]), .A3(RF_pc_out[1]), 
        .ZN(n1101) );
  MAOI22D0BWP12T U1563 ( .A1(RF_pc_out[4]), .A2(n1101), .B1(RF_pc_out[4]), 
        .B2(n1101), .ZN(n1412) );
  NR4D0BWP12T U1564 ( .A1(n1218), .A2(n1190), .A3(n1412), .A4(n1370), .ZN(
        n1107) );
  MAOI22D0BWP12T U1565 ( .A1(RF_pc_out[7]), .A2(n1102), .B1(RF_pc_out[7]), 
        .B2(n1102), .ZN(n1180) );
  MAOI22D0BWP12T U1566 ( .A1(RF_pc_out[9]), .A2(n1103), .B1(RF_pc_out[9]), 
        .B2(n1103), .ZN(n1216) );
  MOAI22D0BWP12T U1567 ( .A1(RF_pc_out[6]), .A2(n1104), .B1(RF_pc_out[6]), 
        .B2(n1104), .ZN(n1219) );
  MOAI22D0BWP12T U1568 ( .A1(RF_pc_out[8]), .A2(n1105), .B1(RF_pc_out[8]), 
        .B2(n1105), .ZN(n1217) );
  NR4D0BWP12T U1569 ( .A1(n1180), .A2(n1216), .A3(n1219), .A4(n1217), .ZN(
        n1106) );
  AN4XD1BWP12T U1570 ( .A1(n1109), .A2(n1108), .A3(n1107), .A4(n1106), .Z(
        n1110) );
  AN4XD1BWP12T U1571 ( .A1(n1113), .A2(n1112), .A3(n1111), .A4(n1110), .Z(
        n1481) );
  TPND3D0BWP12T U1572 ( .A1(n1422), .A2(
        Instruction_Fetch_inst1_first_instruction_fetched), .A3(n1481), .ZN(
        n1118) );
  OAI21D0BWP12T U1573 ( .A1(Instruction_Fetch_inst1_currentState_1_), .A2(
        DEC_IF_stall_to_instructionfetch), .B(
        Instruction_Fetch_inst1_currentState_0_), .ZN(n1114) );
  AOI31D0BWP12T U1574 ( .A1(n1118), .A2(n754), .A3(n1114), .B(reset), .ZN(
        Instruction_Fetch_inst1_N79) );
  CKND2D0BWP12T U1575 ( .A1(n1116), .A2(n1115), .ZN(n1117) );
  AOI31D0BWP12T U1576 ( .A1(n1119), .A2(n1118), .A3(n1117), .B(reset), .ZN(
        Instruction_Fetch_inst1_N80) );
  NR2D1BWP12T U1577 ( .A1(n1479), .A2(reset), .ZN(n1567) );
  AO22XD0BWP12T U1578 ( .A1(MEMCTRL_RF_IF_data_in[14]), .A2(n1559), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_14_), .B2(n1567), .Z(
        Instruction_Fetch_inst1_N97) );
  AO221D0BWP12T U1579 ( .A1(n754), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_12_), .B1(n1479), .B2(
        MEMCTRL_RF_IF_data_in[12]), .C(reset), .Z(Instruction_Fetch_inst1_N95)
         );
  MUX2D1BWP12T U1580 ( .I0(RF_OUT_v), .I1(ALU_OUT_v), .S(
        DEC_CPSR_update_flag_v), .Z(new_v) );
  NR2D1BWP12T U1581 ( .A1(n1120), .A2(n1224), .ZN(n1651) );
  AOI211D0BWP12T U1582 ( .A1(n1122), .A2(n1676), .B(n1121), .C(n1530), .ZN(
        n1123) );
  AOI211D0BWP12T U1583 ( .A1(n1276), .A2(n1604), .B(n1651), .C(n1123), .ZN(
        n1124) );
  TPND2D0BWP12T U1584 ( .A1(n1124), .A2(n1227), .ZN(n1128) );
  NR3XD0BWP12T U1585 ( .A1(n1125), .A2(n1679), .A3(n1677), .ZN(n1179) );
  NR2D0BWP12T U1586 ( .A1(n1600), .A2(n1601), .ZN(n1126) );
  MOAI22D0BWP12T U1587 ( .A1(n1126), .A2(n1529), .B1(n1682), .B2(
        DEC_ALU_alu_opcode[1]), .ZN(n1127) );
  AO211D0BWP12T U1588 ( .A1(n1578), .A2(n1128), .B(n1179), .C(n1127), .Z(n850)
         );
  INVD1BWP12T U1589 ( .I(n1651), .ZN(n1518) );
  AOI21D0BWP12T U1590 ( .A1(n1518), .A2(n1264), .B(n1331), .ZN(n1129) );
  AO211D0BWP12T U1591 ( .A1(n1682), .A2(DEC_RF_alu_write_to_reg[4]), .B(n1129), 
        .C(n1280), .Z(n815) );
  HA1D0BWP12T U1592 ( .A(n1130), .B(RF_pc_out[22]), .CO(n1243), .S(n1085) );
  HA1D0BWP12T U1593 ( .A(n1132), .B(RF_pc_out[30]), .CO(n1131), .S(n1133) );
  CKAN2D0BWP12T U1594 ( .A1(n1133), .A2(n1422), .Z(
        IF_RF_incremented_pc_out[30]) );
  NR2D1BWP12T U1595 ( .A1(n1674), .A2(n1675), .ZN(n1182) );
  NR2D0BWP12T U1596 ( .A1(n1135), .A2(n1134), .ZN(n1172) );
  NR4D0BWP12T U1597 ( .A1(n1137), .A2(n1136), .A3(n1172), .A4(n1597), .ZN(
        n1155) );
  AO21D1BWP12T U1598 ( .A1(n1139), .A2(n1140), .B(n1138), .Z(n1213) );
  AOI32D0BWP12T U1599 ( .A1(n1141), .A2(n1140), .A3(irdecode_inst1_N705), .B1(
        n1153), .B2(n1141), .ZN(n1173) );
  INR3XD0BWP12T U1600 ( .A1(n1146), .B1(n1145), .B2(n1659), .ZN(n1147) );
  AOI31D0BWP12T U1601 ( .A1(n1155), .A2(n1213), .A3(n1147), .B(n1670), .ZN(
        n1149) );
  TPOAI31D0BWP12T U1602 ( .A1(n1149), .A2(n1603), .A3(n1148), .B(n1677), .ZN(
        n1150) );
  AOI21D1BWP12T U1603 ( .A1(n1182), .A2(n1150), .B(n1679), .ZN(n1152) );
  AO21D0BWP12T U1604 ( .A1(n1682), .A2(DEC_MEMCTRL_memory_load_request), .B(
        n1152), .Z(n861) );
  NR2D0BWP12T U1605 ( .A1(n1679), .A2(n1670), .ZN(n1308) );
  AO211D0BWP12T U1606 ( .A1(n1682), .A2(
        DEC_MISC_OUT_memory_address_source_is_reg), .B(n1308), .C(n1179), .Z(
        n836) );
  NR2D1BWP12T U1607 ( .A1(Instruction_Fetch_inst1_currentState_1_), .A2(
        DEC_MISC_OUT_memory_address_source_is_reg), .ZN(n1419) );
  INR2XD0BWP12T U1608 ( .A1(DEC_MISC_OUT_memory_address_source_is_reg), .B1(
        Instruction_Fetch_inst1_currentState_1_), .ZN(n1420) );
  AO222D0BWP12T U1609 ( .A1(n1422), .A2(n1151), .B1(ALU_MISC_OUT_result[12]), 
        .B2(n1419), .C1(n1420), .C2(RF_MEMCTRL_address_reg[12]), .Z(
        MEMCTRL_IN_address[11]) );
  AO21D0BWP12T U1610 ( .A1(n1682), .A2(DEC_RF_memory_write_to_reg_enable), .B(
        n1152), .Z(n825) );
  CKND1BWP12T U1611 ( .I(IF_DEC_instruction[2]), .ZN(n1531) );
  CKND0BWP12T U1612 ( .I(n1153), .ZN(n1154) );
  TPAOI31D0BWP12T U1613 ( .A1(n1156), .A2(n1155), .A3(n1154), .B(n1503), .ZN(
        n1162) );
  ND4D0BWP12T U1614 ( .A1(n1159), .A2(n1499), .A3(n1158), .A4(n1157), .ZN(
        n1160) );
  OAI32D0BWP12T U1615 ( .A1(n1162), .A2(n1161), .A3(n1160), .B1(n1501), .B2(
        n1162), .ZN(n1163) );
  OAI211D0BWP12T U1616 ( .A1(n1531), .A2(n1164), .B(n1273), .C(n1163), .ZN(
        n1196) );
  AOI211D0BWP12T U1617 ( .A1(n1682), .A2(DEC_RF_memory_write_to_reg[2]), .B(
        n1165), .C(n1196), .ZN(n1168) );
  AOI22D0BWP12T U1618 ( .A1(n1166), .A2(n1656), .B1(n1675), .B2(
        IF_DEC_instruction[2]), .ZN(n1167) );
  AOI32D0BWP12T U1619 ( .A1(n1205), .A2(n1168), .A3(n1167), .B1(n1331), .B2(
        n1168), .ZN(n822) );
  HA1D0BWP12T U1620 ( .A(n1169), .B(RF_pc_out[29]), .CO(n1132), .S(n1170) );
  AN2D0BWP12T U1621 ( .A1(n1170), .A2(n1422), .Z(IF_RF_incremented_pc_out[29])
         );
  CKND0BWP12T U1622 ( .I(n1171), .ZN(n1175) );
  NR2D1BWP12T U1623 ( .A1(n1172), .A2(n1494), .ZN(n1497) );
  IND4D1BWP12T U1624 ( .A1(n1597), .B1(n1173), .B2(n1213), .B3(n1497), .ZN(
        n1652) );
  AOI211D0BWP12T U1625 ( .A1(n1672), .A2(n1175), .B(n1174), .C(n1652), .ZN(
        n1177) );
  OAI32D0BWP12T U1626 ( .A1(n1679), .A2(n1177), .A3(n1670), .B1(n1176), .B2(
        n1679), .ZN(n1178) );
  AO211D0BWP12T U1627 ( .A1(n1682), .A2(DEC_MEMCTRL_memory_store_request), .B(
        n1179), .C(n1178), .Z(n852) );
  AO222D0BWP12T U1628 ( .A1(n1422), .A2(n1180), .B1(n1420), .B2(
        RF_MEMCTRL_address_reg[7]), .C1(ALU_MISC_OUT_result[7]), .C2(n1419), 
        .Z(MEMCTRL_IN_address[6]) );
  NR2D0BWP12T U1629 ( .A1(n1583), .A2(n1194), .ZN(n1183) );
  TPND2D0BWP12T U1630 ( .A1(n1182), .A2(n1181), .ZN(n1192) );
  OR2XD1BWP12T U1631 ( .A1(n1192), .A2(n1677), .Z(n1202) );
  AOI211D0BWP12T U1632 ( .A1(n1671), .A2(IF_DEC_instruction[0]), .B(n1183), 
        .C(n1202), .ZN(n1188) );
  CKND2D0BWP12T U1633 ( .A1(n1682), .A2(DEC_RF_memory_store_data_reg[0]), .ZN(
        n1187) );
  AOI21D0BWP12T U1634 ( .A1(n1501), .A2(n1185), .B(n1184), .ZN(n1186) );
  OAI211D0BWP12T U1635 ( .A1(n1188), .A2(n1331), .B(n1187), .C(n1186), .ZN(
        n830) );
  AO222D0BWP12T U1636 ( .A1(n1422), .A2(n1189), .B1(n1420), .B2(
        RF_MEMCTRL_address_reg[11]), .C1(ALU_MISC_OUT_result[11]), .C2(n1419), 
        .Z(MEMCTRL_IN_address[10]) );
  AO222D0BWP12T U1637 ( .A1(n1422), .A2(n1190), .B1(n1420), .B2(
        RF_MEMCTRL_address_reg[5]), .C1(ALU_MISC_OUT_result[5]), .C2(n1419), 
        .Z(MEMCTRL_IN_address[4]) );
  AO222D0BWP12T U1638 ( .A1(n1422), .A2(n1191), .B1(n1420), .B2(
        RF_MEMCTRL_address_reg[10]), .C1(ALU_MISC_OUT_result[10]), .C2(n1419), 
        .Z(MEMCTRL_IN_address[9]) );
  AOI211D0BWP12T U1639 ( .A1(n1671), .A2(IF_DEC_instruction[2]), .B(n1192), 
        .C(n1677), .ZN(n1193) );
  OAI32D0BWP12T U1640 ( .A1(n1331), .A2(n1195), .A3(n1194), .B1(n1193), .B2(
        n1331), .ZN(n1197) );
  AO211D0BWP12T U1641 ( .A1(n1682), .A2(DEC_RF_memory_store_data_reg[2]), .B(
        n1197), .C(n1196), .Z(n828) );
  AN2D0BWP12T U1642 ( .A1(n1199), .A2(n1422), .Z(IF_RF_incremented_pc_out[28])
         );
  OAI21D1BWP12T U1643 ( .A1(n1200), .A2(n1509), .B(n1273), .ZN(n1230) );
  CKND0BWP12T U1644 ( .I(n1201), .ZN(n1204) );
  NR2D0BWP12T U1645 ( .A1(n1204), .A2(n1670), .ZN(n1203) );
  AO21D0BWP12T U1646 ( .A1(n1682), .A2(DEC_RF_memory_store_data_reg[4]), .B(
        n928), .Z(n826) );
  AO211D0BWP12T U1647 ( .A1(n1682), .A2(DEC_RF_memory_store_data_reg[3]), .B(
        n1681), .C(n928), .Z(n827) );
  AOI32D0BWP12T U1648 ( .A1(n1677), .A2(n1205), .A3(n1204), .B1(n1670), .B2(
        n1205), .ZN(n1206) );
  AOI21D0BWP12T U1649 ( .A1(n1328), .A2(n1206), .B(n1230), .ZN(n1207) );
  OAI21D0BWP12T U1650 ( .A1(n1677), .A2(n1509), .B(n1207), .ZN(n1680) );
  AO21D0BWP12T U1651 ( .A1(n1682), .A2(DEC_RF_memory_write_to_reg[4]), .B(
        n1680), .Z(n820) );
  HA1D1BWP12T U1652 ( .A(n1208), .B(RF_pc_out[27]), .CO(n1198), .S(n1209) );
  AN2D0BWP12T U1653 ( .A1(n1209), .A2(n1422), .Z(IF_RF_incremented_pc_out[27])
         );
  NR2XD0BWP12T U1654 ( .A1(n1211), .A2(n1210), .ZN(n1490) );
  OR3D1BWP12T U1655 ( .A1(n1212), .A2(n1612), .A3(n1634), .Z(n1251) );
  RCAOI21D0BWP12T U1656 ( .A1(n1328), .A2(n1251), .B(n1280), .ZN(n1506) );
  IND2XD1BWP12T U1657 ( .A1(n1214), .B1(n1213), .ZN(n1488) );
  AOI22D0BWP12T U1658 ( .A1(n1682), .A2(irdecode_inst1_step[2]), .B1(n1595), 
        .B2(n1488), .ZN(n1215) );
  OAI211D0BWP12T U1659 ( .A1(n1490), .A2(n1509), .B(n1506), .C(n1215), .ZN(
        irdecode_inst1_next_step_2_) );
  AO222D0BWP12T U1660 ( .A1(n1422), .A2(n1216), .B1(n1420), .B2(
        RF_MEMCTRL_address_reg[9]), .C1(ALU_MISC_OUT_result[9]), .C2(n1419), 
        .Z(MEMCTRL_IN_address[8]) );
  AO222D0BWP12T U1661 ( .A1(n1422), .A2(n1217), .B1(n1420), .B2(
        RF_MEMCTRL_address_reg[8]), .C1(ALU_MISC_OUT_result[8]), .C2(n1419), 
        .Z(MEMCTRL_IN_address[7]) );
  AO222D0BWP12T U1662 ( .A1(n1422), .A2(n1218), .B1(n1420), .B2(
        RF_MEMCTRL_address_reg[3]), .C1(ALU_MISC_OUT_result[3]), .C2(n1419), 
        .Z(MEMCTRL_IN_address[2]) );
  AO222D0BWP12T U1663 ( .A1(n1422), .A2(n1219), .B1(n1420), .B2(
        RF_MEMCTRL_address_reg[6]), .C1(ALU_MISC_OUT_result[6]), .C2(n1419), 
        .Z(MEMCTRL_IN_address[5]) );
  HA1D1BWP12T U1664 ( .A(n1220), .B(RF_pc_out[26]), .CO(n1208), .S(n1221) );
  AN2D0BWP12T U1665 ( .A1(n1221), .A2(n1422), .Z(IF_RF_incremented_pc_out[26])
         );
  HA1D0BWP12T U1666 ( .A(n1222), .B(RF_pc_out[25]), .CO(n1220), .S(n1223) );
  CKAN2D1BWP12T U1667 ( .A1(n1223), .A2(n1422), .Z(
        IF_RF_incremented_pc_out[25]) );
  CKND2D0BWP12T U1668 ( .A1(n1600), .A2(n1664), .ZN(n1228) );
  INR2XD0BWP12T U1669 ( .A1(irdecode_inst1_N911), .B1(n1224), .ZN(n1571) );
  TPND2D0BWP12T U1670 ( .A1(n1226), .A2(n1225), .ZN(n1247) );
  NR2D1BWP12T U1671 ( .A1(n1571), .A2(n1247), .ZN(n1274) );
  AOI31D0BWP12T U1672 ( .A1(n1228), .A2(n1274), .A3(n1227), .B(n1331), .ZN(
        n1229) );
  AO211D0BWP12T U1673 ( .A1(n1682), .A2(DEC_ALU_alu_opcode[3]), .B(n1230), .C(
        n1229), .Z(n849) );
  HA1D0BWP12T U1674 ( .A(n1231), .B(RF_pc_out[24]), .CO(n1222), .S(n1232) );
  CKAN2D1BWP12T U1675 ( .A1(n1232), .A2(n1422), .Z(
        IF_RF_incremented_pc_out[24]) );
  AOI22D0BWP12T U1676 ( .A1(n1255), .A2(IF_DEC_instruction[3]), .B1(
        IF_DEC_instruction[6]), .B2(n1239), .ZN(n1237) );
  OAI21D0BWP12T U1677 ( .A1(n1234), .A2(n1233), .B(n1328), .ZN(n1235) );
  CKND2D1BWP12T U1678 ( .A1(n1235), .A2(n1273), .ZN(n1245) );
  INVD1BWP12T U1679 ( .I(n1245), .ZN(n1241) );
  ND2D1BWP12T U1680 ( .A1(n1682), .A2(DEC_RF_operand_b[0]), .ZN(n1236) );
  OAI211D0BWP12T U1681 ( .A1(n1237), .A2(n1331), .B(n1241), .C(n1236), .ZN(
        n844) );
  NR2D0BWP12T U1682 ( .A1(n1306), .A2(n1331), .ZN(n1248) );
  AOI22D0BWP12T U1683 ( .A1(n1248), .A2(IF_DEC_instruction[6]), .B1(n1682), 
        .B2(DEC_RF_operand_b[3]), .ZN(n1238) );
  CKND2D1BWP12T U1684 ( .A1(n1241), .A2(n1238), .ZN(n841) );
  AOI22D0BWP12T U1685 ( .A1(n1255), .A2(IF_DEC_instruction[5]), .B1(n1631), 
        .B2(n1239), .ZN(n1242) );
  ND2D1BWP12T U1686 ( .A1(n1682), .A2(DEC_RF_operand_b[2]), .ZN(n1240) );
  OAI211D0BWP12T U1687 ( .A1(n1242), .A2(n1331), .B(n1241), .C(n1240), .ZN(
        n842) );
  HA1D0BWP12T U1688 ( .A(n1243), .B(RF_pc_out[23]), .CO(n1231), .S(n1244) );
  AO21D0BWP12T U1689 ( .A1(n1682), .A2(DEC_RF_operand_b[4]), .B(n1245), .Z(
        n840) );
  IND2XD1BWP12T U1690 ( .A1(n1247), .B1(n1246), .ZN(n1257) );
  INVD1BWP12T U1691 ( .I(n1257), .ZN(n1250) );
  AOI21D0BWP12T U1692 ( .A1(IF_DEC_instruction[7]), .A2(n1248), .B(n1280), 
        .ZN(n1266) );
  ND2D1BWP12T U1693 ( .A1(n1682), .A2(DEC_RF_operand_a[3]), .ZN(n1249) );
  OAI211D0BWP12T U1694 ( .A1(n1331), .A2(n1250), .B(n1266), .C(n1249), .ZN(
        n812) );
  OAI32D0BWP12T U1695 ( .A1(n1280), .A2(n1661), .A3(n1251), .B1(n1328), .B2(
        n1280), .ZN(n1254) );
  AOI22D0BWP12T U1696 ( .A1(n1682), .A2(DEC_RF_memory_store_address_reg[0]), 
        .B1(n1595), .B2(n1631), .ZN(n1252) );
  TPND2D0BWP12T U1697 ( .A1(n1254), .A2(n1252), .ZN(n835) );
  AOI22D0BWP12T U1698 ( .A1(DEC_RF_memory_store_address_reg[2]), .A2(n1682), 
        .B1(n1595), .B2(n1656), .ZN(n1253) );
  TPND2D0BWP12T U1699 ( .A1(n1254), .A2(n1253), .ZN(n833) );
  IOA21D0BWP12T U1700 ( .A1(n1682), .A2(DEC_RF_memory_store_address_reg[3]), 
        .B(n1254), .ZN(n832) );
  IOA21D0BWP12T U1701 ( .A1(n1682), .A2(DEC_RF_memory_store_address_reg[4]), 
        .B(n1506), .ZN(n831) );
  CKND0BWP12T U1702 ( .I(n1255), .ZN(n1640) );
  OAI22D0BWP12T U1703 ( .A1(n1640), .A2(n1531), .B1(n1628), .B2(n1637), .ZN(
        n1256) );
  AOI211XD0BWP12T U1704 ( .A1(IF_DEC_instruction[5]), .A2(n1258), .B(n1257), 
        .C(n1256), .ZN(n1260) );
  ND2D1BWP12T U1705 ( .A1(n1682), .A2(DEC_RF_operand_a[2]), .ZN(n1259) );
  OAI211D0BWP12T U1706 ( .A1(n1331), .A2(n1260), .B(n1273), .C(n1259), .ZN(
        n813) );
  NR2D0BWP12T U1707 ( .A1(n1612), .A2(n1261), .ZN(n1262) );
  OAI31D0BWP12T U1708 ( .A1(n1583), .A2(n1676), .A3(n1306), .B(n1262), .ZN(
        n1591) );
  IND4D0BWP12T U1709 ( .A1(n1591), .B1(n1264), .B2(n1263), .B3(n1648), .ZN(
        n1268) );
  CKND0BWP12T U1710 ( .I(n1268), .ZN(n1267) );
  CKND2D0BWP12T U1711 ( .A1(n1682), .A2(DEC_RF_alu_write_to_reg[3]), .ZN(n1265) );
  OAI211D0BWP12T U1712 ( .A1(n1331), .A2(n1267), .B(n1266), .C(n1265), .ZN(
        n817) );
  NR2D0BWP12T U1713 ( .A1(n1590), .A2(n1628), .ZN(n1269) );
  AOI211D0BWP12T U1714 ( .A1(n1593), .A2(IF_DEC_instruction[2]), .B(n1269), 
        .C(n1268), .ZN(n1271) );
  CKND2D0BWP12T U1715 ( .A1(n1682), .A2(DEC_RF_alu_write_to_reg[2]), .ZN(n1270) );
  OAI211D0BWP12T U1716 ( .A1(n1331), .A2(n1271), .B(n1273), .C(n1270), .ZN(
        n818) );
  ND2D1BWP12T U1717 ( .A1(n1682), .A2(DEC_RF_operand_a[4]), .ZN(n1272) );
  OAI211D0BWP12T U1718 ( .A1(n1274), .A2(n1331), .B(n1273), .C(n1272), .ZN(
        n810) );
  AOI22D0BWP12T U1719 ( .A1(n1276), .A2(n1632), .B1(n1628), .B2(n1275), .ZN(
        n1277) );
  AOI31D0BWP12T U1720 ( .A1(n1279), .A2(n1278), .A3(n1277), .B(n1331), .ZN(
        n1281) );
  AO211D0BWP12T U1721 ( .A1(n1682), .A2(DEC_MEMCTRL_load_store_width[1]), .B(
        n1281), .C(n1280), .Z(n837) );
  HA1D0BWP12T U1722 ( .A(n1282), .B(RF_pc_out[20]), .CO(n1086), .S(n1283) );
  HA1D2BWP12T U1723 ( .A(n1284), .B(RF_pc_out[19]), .CO(n1282), .S(n1285) );
  AOI22D0BWP12T U1724 ( .A1(n1676), .A2(RF_OUT_z), .B1(RF_OUT_c), .B2(n1664), 
        .ZN(n1286) );
  MAOI22D0BWP12T U1725 ( .A1(n1286), .A2(n1631), .B1(n1286), .B2(n1631), .ZN(
        n1299) );
  AOI22D0BWP12T U1726 ( .A1(n1676), .A2(RF_OUT_n), .B1(RF_OUT_v), .B2(n1664), 
        .ZN(n1288) );
  AOI211D0BWP12T U1727 ( .A1(n1288), .A2(n1583), .B(n1628), .C(n1677), .ZN(
        n1287) );
  OAI21D0BWP12T U1728 ( .A1(n1288), .A2(n1583), .B(n1287), .ZN(n1298) );
  CKND0BWP12T U1729 ( .I(n1289), .ZN(n1291) );
  AOI22D0BWP12T U1730 ( .A1(n1291), .A2(n1579), .B1(n1290), .B2(n1289), .ZN(
        n1296) );
  MUX2ND0BWP12T U1731 ( .I0(n1293), .I1(n1292), .S(n1676), .ZN(n1294) );
  MAOI22D0BWP12T U1732 ( .A1(n1583), .A2(n1294), .B1(n1583), .B2(n1294), .ZN(
        n1295) );
  OAI221D0BWP12T U1733 ( .A1(n1628), .A2(n1296), .B1(n1656), .B2(n1295), .C(
        n1677), .ZN(n1297) );
  OAI211D0BWP12T U1734 ( .A1(n1300), .A2(n1299), .B(n1298), .C(n1297), .ZN(
        n1302) );
  AOI211D0BWP12T U1735 ( .A1(n1303), .A2(n1302), .B(n1601), .C(n1301), .ZN(
        n1305) );
  NR2D0BWP12T U1736 ( .A1(n1661), .A2(n1612), .ZN(n1304) );
  OA211D0BWP12T U1737 ( .A1(n1581), .A2(n1306), .B(n1305), .C(n1304), .Z(n1307) );
  AOI31D0BWP12T U1738 ( .A1(n1575), .A2(n1590), .A3(n1307), .B(n1679), .ZN(
        irdecode_inst1_next_alu_write_to_reg_enable) );
  AO22XD0BWP12T U1739 ( .A1(DEC_RF_memory_store_address_reg[1]), .A2(n1682), 
        .B1(n1308), .B2(n1664), .Z(n834) );
  CKND2D0BWP12T U1740 ( .A1(n1578), .A2(n1672), .ZN(n1309) );
  NR2D1BWP12T U1741 ( .A1(n1638), .A2(n1309), .ZN(n1322) );
  AOI22D0BWP12T U1742 ( .A1(n1322), .A2(IF_DEC_instruction[0]), .B1(n1682), 
        .B2(DEC_RF_offset_b[12]), .ZN(n1310) );
  TPND2D0BWP12T U1743 ( .A1(n1512), .A2(n1310), .ZN(n797) );
  HA1D2BWP12T U1744 ( .A(n1311), .B(RF_pc_out[18]), .CO(n1284), .S(n1312) );
  AOI22D0BWP12T U1745 ( .A1(n1322), .A2(IF_DEC_instruction[1]), .B1(n1682), 
        .B2(DEC_RF_offset_b[13]), .ZN(n1313) );
  TPND2D0BWP12T U1746 ( .A1(n1512), .A2(n1313), .ZN(n796) );
  AOI22D0BWP12T U1747 ( .A1(n1322), .A2(IF_DEC_instruction[2]), .B1(n1682), 
        .B2(DEC_RF_offset_b[14]), .ZN(n1314) );
  TPND2D0BWP12T U1748 ( .A1(n1512), .A2(n1314), .ZN(n795) );
  AOI22D0BWP12T U1749 ( .A1(n1322), .A2(IF_DEC_instruction[3]), .B1(n1682), 
        .B2(DEC_RF_offset_b[15]), .ZN(n1315) );
  TPND2D0BWP12T U1750 ( .A1(n1512), .A2(n1315), .ZN(n794) );
  AOI22D0BWP12T U1751 ( .A1(n1322), .A2(IF_DEC_instruction[4]), .B1(n1682), 
        .B2(DEC_RF_offset_b[16]), .ZN(n1316) );
  TPND2D0BWP12T U1752 ( .A1(n1512), .A2(n1316), .ZN(n793) );
  AOI22D0BWP12T U1753 ( .A1(n1322), .A2(IF_DEC_instruction[5]), .B1(n1682), 
        .B2(DEC_RF_offset_b[17]), .ZN(n1317) );
  TPND2D0BWP12T U1754 ( .A1(n1512), .A2(n1317), .ZN(n792) );
  AOI22D0BWP12T U1755 ( .A1(n1322), .A2(IF_DEC_instruction[6]), .B1(n1682), 
        .B2(DEC_RF_offset_b[18]), .ZN(n1318) );
  TPND2D0BWP12T U1756 ( .A1(n1512), .A2(n1318), .ZN(n791) );
  AOI22D0BWP12T U1757 ( .A1(n1322), .A2(IF_DEC_instruction[7]), .B1(n1682), 
        .B2(DEC_RF_offset_b[19]), .ZN(n1319) );
  TPND2D0BWP12T U1758 ( .A1(n1512), .A2(n1319), .ZN(n790) );
  AOI22D0BWP12T U1759 ( .A1(n1322), .A2(n1631), .B1(n1682), .B2(
        DEC_RF_offset_b[20]), .ZN(n1320) );
  TPND2D0BWP12T U1760 ( .A1(n1512), .A2(n1320), .ZN(n789) );
  AOI22D0BWP12T U1761 ( .A1(n1322), .A2(n1664), .B1(n1682), .B2(
        DEC_RF_offset_b[21]), .ZN(n1321) );
  TPND2D0BWP12T U1762 ( .A1(n1512), .A2(n1321), .ZN(n788) );
  AOI22D0BWP12T U1763 ( .A1(n1322), .A2(n1656), .B1(n1682), .B2(
        DEC_RF_offset_b[22]), .ZN(n1323) );
  TPND2D0BWP12T U1764 ( .A1(n1512), .A2(n1323), .ZN(n787) );
  AO21D0BWP12T U1765 ( .A1(n1682), .A2(DEC_RF_offset_b[30]), .B(n1514), .Z(
        n779) );
  AO21D0BWP12T U1766 ( .A1(n1682), .A2(DEC_RF_offset_b[29]), .B(n1514), .Z(
        n780) );
  AO21D0BWP12T U1767 ( .A1(n1682), .A2(DEC_RF_offset_b[28]), .B(n1514), .Z(
        n781) );
  AO21D0BWP12T U1768 ( .A1(n1682), .A2(DEC_RF_offset_b[27]), .B(n1514), .Z(
        n782) );
  AO21D0BWP12T U1769 ( .A1(n1682), .A2(DEC_RF_offset_b[26]), .B(n1514), .Z(
        n783) );
  AO21D0BWP12T U1770 ( .A1(n1682), .A2(DEC_RF_offset_b[25]), .B(n1514), .Z(
        n784) );
  AO21D0BWP12T U1771 ( .A1(n1682), .A2(DEC_RF_offset_b[24]), .B(n1514), .Z(
        n785) );
  AO21D0BWP12T U1772 ( .A1(n1682), .A2(DEC_RF_offset_b[23]), .B(n1514), .Z(
        n786) );
  HA1D0BWP12T U1773 ( .A(n1324), .B(RF_pc_out[17]), .CO(n1311), .S(n1325) );
  AN2XD0BWP12T U1774 ( .A1(n1325), .A2(n1422), .Z(IF_RF_incremented_pc_out[17]) );
  AO21D0BWP12T U1775 ( .A1(n1682), .A2(DEC_RF_offset_b[31]), .B(n1514), .Z(
        n777) );
  NR4D0BWP12T U1776 ( .A1(IF_DEC_instruction[1]), .A2(IF_DEC_instruction[2]), 
        .A3(IF_DEC_instruction[0]), .A4(IF_DEC_instruction[3]), .ZN(n1329) );
  TPND2D0BWP12T U1777 ( .A1(n1664), .A2(n1631), .ZN(n1326) );
  NR4D0BWP12T U1778 ( .A1(n1628), .A2(n1327), .A3(n1530), .A4(n1326), .ZN(
        n1332) );
  IND3D1BWP12T U1779 ( .A1(n1329), .B1(n1328), .B2(n1332), .ZN(n1646) );
  INVD1BWP12T U1780 ( .I(n1646), .ZN(n1335) );
  AOI21D0BWP12T U1781 ( .A1(n1329), .A2(n1332), .B(n1331), .ZN(n1330) );
  NR2D1BWP12T U1782 ( .A1(n1330), .A2(reset), .ZN(n1645) );
  INR2D0BWP12T U1783 ( .A1(irdecode_inst1_itstate_3_), .B1(
        irdecode_inst1_itstate_2_), .ZN(n1334) );
  AOI211XD0BWP12T U1784 ( .A1(n1334), .A2(n1333), .B(n1332), .C(n1331), .ZN(
        n1483) );
  AO222D0BWP12T U1785 ( .A1(IF_DEC_instruction[1]), .A2(n1335), .B1(n1645), 
        .B2(irdecode_inst1_itstate_1_), .C1(n1483), .C2(
        irdecode_inst1_itstate_0_), .Z(n859) );
  AO222D0BWP12T U1786 ( .A1(IF_DEC_instruction[2]), .A2(n1335), .B1(n1645), 
        .B2(irdecode_inst1_itstate_2_), .C1(n1483), .C2(
        irdecode_inst1_itstate_1_), .Z(n858) );
  AO222D0BWP12T U1787 ( .A1(IF_DEC_instruction[3]), .A2(n1335), .B1(n1645), 
        .B2(irdecode_inst1_itstate_3_), .C1(irdecode_inst1_itstate_2_), .C2(
        n1483), .Z(n857) );
  AO222D0BWP12T U1788 ( .A1(IF_DEC_instruction[4]), .A2(n1335), .B1(n1645), 
        .B2(irdecode_inst1_itstate_4_), .C1(irdecode_inst1_itstate_3_), .C2(
        n1483), .Z(n856) );
  HA1D0BWP12T U1789 ( .A(n1336), .B(RF_pc_out[16]), .CO(n1324), .S(n1337) );
  AN2XD0BWP12T U1790 ( .A1(n1337), .A2(n1422), .Z(IF_RF_incremented_pc_out[16]) );
  HA1D2BWP12T U1791 ( .A(n1338), .B(RF_pc_out[15]), .CO(n1336), .S(n1339) );
  HA1D1BWP12T U1792 ( .A(n1340), .B(RF_pc_out[14]), .CO(n1338), .S(n1341) );
  HA1D0BWP12T U1793 ( .A(n1342), .B(RF_pc_out[13]), .CO(n1340), .S(n1343) );
  HA1D0BWP12T U1794 ( .A(n1344), .B(RF_pc_out[12]), .CO(n1342), .S(n1345) );
  HA1D0BWP12T U1795 ( .A(n1346), .B(RF_pc_out[11]), .CO(n1344), .S(n1347) );
  HA1D0BWP12T U1796 ( .A(n1348), .B(RF_pc_out[10]), .CO(n1346), .S(n1349) );
  HA1D0BWP12T U1797 ( .A(n1350), .B(RF_pc_out[9]), .CO(n1348), .S(n1351) );
  HA1D0BWP12T U1798 ( .A(n1352), .B(RF_pc_out[8]), .CO(n1350), .S(n1353) );
  HA1D0BWP12T U1799 ( .A(n1354), .B(RF_pc_out[7]), .CO(n1352), .S(n1355) );
  NR2D1BWP12T U1800 ( .A1(DEC_MEMCTRL_load_store_width[1]), .A2(
        DEC_MEMCTRL_load_store_width[0]), .ZN(n1556) );
  NR2D0BWP12T U1801 ( .A1(Instruction_Fetch_inst1_currentState_1_), .A2(
        DEC_MEMCTRL_memory_load_request), .ZN(n1555) );
  CKND0BWP12T U1802 ( .I(n1470), .ZN(n1356) );
  AOI211XD0BWP12T U1803 ( .A1(DEC_MEMCTRL_load_store_width[0]), .A2(
        DEC_MEMCTRL_load_store_width[1]), .B(n1356), .C(reset), .ZN(n1357) );
  CKND0BWP12T U1804 ( .I(n1357), .ZN(n1358) );
  ND3XD0BWP12T U1805 ( .A1(n1357), .A2(DEC_MEMCTRL_memory_store_request), .A3(
        n1555), .ZN(n1478) );
  OAI31D0BWP12T U1806 ( .A1(n1556), .A2(n1555), .A3(n1358), .B(n1478), .ZN(
        memory_interface_inst1_fsm_N32) );
  ND2D1BWP12T U1807 ( .A1(n1476), .A2(memory_interface_inst1_fsm_state_3_), 
        .ZN(n1472) );
  CKND2D0BWP12T U1808 ( .A1(n1472), .A2(n1386), .ZN(n1416) );
  IOA21D0BWP12T U1809 ( .A1(n1359), .A2(n1416), .B(n1478), .ZN(
        memory_interface_inst1_fsm_N35) );
  HA1D1BWP12T U1810 ( .A(n1360), .B(RF_pc_out[6]), .CO(n1354), .S(n1361) );
  HA1D2BWP12T U1811 ( .A(n1362), .B(RF_pc_out[5]), .CO(n1360), .S(n1363) );
  HA1D0BWP12T U1812 ( .A(n1364), .B(RF_pc_out[4]), .CO(n1362), .S(n1365) );
  HA1D0BWP12T U1813 ( .A(RF_pc_out[1]), .B(RF_pc_out[2]), .CO(n1367), .S(n1366) );
  HA1D0BWP12T U1814 ( .A(n1367), .B(RF_pc_out[3]), .CO(n1364), .S(n1368) );
  INR2D0BWP12T U1815 ( .A1(n1370), .B1(n1369), .ZN(MEMCTRL_IN_address[0]) );
  INR3XD0BWP12T U1816 ( .A1(memory_interface_inst1_delayed_is_signed), .B1(
        n1372), .B2(n1371), .ZN(n1377) );
  AN2XD1BWP12T U1817 ( .A1(n1384), .A2(n1373), .Z(n1374) );
  OAI21D1BWP12T U1818 ( .A1(n1375), .A2(n1684), .B(n1374), .ZN(n1376) );
  OAI21D1BWP12T U1819 ( .A1(n1372), .A2(n1549), .B(n1547), .ZN(
        MEMCTRL_RF_IF_data_in[31]) );
  INVD1BWP12T U1820 ( .I(MEM_MEMCTRL_from_mem_data[6]), .ZN(n1426) );
  OAI21D1BWP12T U1821 ( .A1(n1426), .A2(n1549), .B(n1547), .ZN(
        MEMCTRL_RF_IF_data_in[30]) );
  INVD1BWP12T U1822 ( .I(MEM_MEMCTRL_from_mem_data[5]), .ZN(n1387) );
  OAI21D1BWP12T U1823 ( .A1(n1387), .A2(n1549), .B(n1547), .ZN(
        MEMCTRL_RF_IF_data_in[29]) );
  INVD1BWP12T U1824 ( .I(MEM_MEMCTRL_from_mem_data[4]), .ZN(n1391) );
  OAI21D1BWP12T U1825 ( .A1(n1391), .A2(n1549), .B(n1547), .ZN(
        MEMCTRL_RF_IF_data_in[28]) );
  INVD1BWP12T U1826 ( .I(MEM_MEMCTRL_from_mem_data[3]), .ZN(n1403) );
  OAI21D1BWP12T U1827 ( .A1(n1403), .A2(n1549), .B(n1547), .ZN(
        MEMCTRL_RF_IF_data_in[27]) );
  INVD1BWP12T U1828 ( .I(MEM_MEMCTRL_from_mem_data[1]), .ZN(n1443) );
  OAI21D1BWP12T U1829 ( .A1(n1443), .A2(n1549), .B(n1547), .ZN(
        MEMCTRL_RF_IF_data_in[25]) );
  INVD1BWP12T U1830 ( .I(memory_interface_inst1_delay_addr_for_adder[10]), 
        .ZN(n1397) );
  NR2D1BWP12T U1831 ( .A1(n1379), .A2(n1378), .ZN(n1558) );
  CKND2D0BWP12T U1832 ( .A1(n1383), .A2(n1558), .ZN(n1399) );
  INR2D1BWP12T U1833 ( .A1(n1386), .B1(n1399), .ZN(n1434) );
  NR2D1BWP12T U1834 ( .A1(n1434), .A2(n1551), .ZN(n1418) );
  ND3D1BWP12T U1835 ( .A1(memory_interface_inst1_delay_addr_for_adder[0]), 
        .A2(memory_interface_inst1_delay_addr_for_adder[1]), .A3(
        memory_interface_inst1_delay_addr_for_adder[2]), .ZN(n1415) );
  INVD1BWP12T U1836 ( .I(n1415), .ZN(n1411) );
  ND2D1BWP12T U1837 ( .A1(n1411), .A2(
        memory_interface_inst1_delay_addr_for_adder[3]), .ZN(n1459) );
  IND2D1BWP12T U1838 ( .A1(n1459), .B1(
        memory_interface_inst1_delay_addr_for_adder[4]), .ZN(n1438) );
  INVD1BWP12T U1839 ( .I(n1438), .ZN(n1435) );
  ND2D1BWP12T U1840 ( .A1(n1435), .A2(
        memory_interface_inst1_delay_addr_for_adder[5]), .ZN(n1442) );
  IND2D1BWP12T U1841 ( .A1(n1442), .B1(
        memory_interface_inst1_delay_addr_for_adder[6]), .ZN(n1410) );
  INVD1BWP12T U1842 ( .I(n1410), .ZN(n1407) );
  ND2D1BWP12T U1843 ( .A1(n1407), .A2(
        memory_interface_inst1_delay_addr_for_adder[7]), .ZN(n1455) );
  INR2D1BWP12T U1844 ( .A1(memory_interface_inst1_delay_addr_for_adder[8]), 
        .B1(n1455), .ZN(n1380) );
  AN2D1BWP12T U1845 ( .A1(n1418), .A2(n1380), .Z(n1552) );
  ND2D1BWP12T U1846 ( .A1(memory_interface_inst1_delay_addr_for_adder[9]), 
        .A2(n1552), .ZN(n1398) );
  INVD1BWP12T U1847 ( .I(n1418), .ZN(n1464) );
  INVD1BWP12T U1848 ( .I(memory_interface_inst1_delay_addr_for_adder[9]), .ZN(
        n1553) );
  INVD1BWP12T U1849 ( .I(n1434), .ZN(n1447) );
  OAI21D1BWP12T U1850 ( .A1(n1380), .A2(n1464), .B(n1447), .ZN(n1554) );
  AOI21D1BWP12T U1851 ( .A1(n1418), .A2(n1553), .B(n1554), .ZN(n1396) );
  OAI21D1BWP12T U1852 ( .A1(memory_interface_inst1_delay_addr_for_adder[10]), 
        .A2(n1464), .B(n1396), .ZN(n1381) );
  AOI22D1BWP12T U1853 ( .A1(memory_interface_inst1_delay_addr_for_adder[11]), 
        .A2(n1381), .B1(MEMCTRL_IN_address[11]), .B2(n1551), .ZN(n1382) );
  OAI31D1BWP12T U1854 ( .A1(memory_interface_inst1_delay_addr_for_adder[11]), 
        .A2(n1397), .A3(n1398), .B(n1382), .ZN(MEMCTRL_MEM_to_mem_address[11])
         );
  INVD1BWP12T U1855 ( .I(RF_MEMCTRL_data_reg[13]), .ZN(n1390) );
  ND2D1BWP12T U1856 ( .A1(n1557), .A2(n1399), .ZN(n1467) );
  CKND1BWP12T U1857 ( .I(n1386), .ZN(n1474) );
  MAOI22D0BWP12T U1858 ( .A1(n1474), .A2(
        memory_interface_inst1_delay_data_in32[29]), .B1(n1387), .B2(n1447), 
        .ZN(n1389) );
  ND2D1BWP12T U1859 ( .A1(n1448), .A2(
        memory_interface_inst1_delay_data_in32[13]), .ZN(n1388) );
  OAI211D1BWP12T U1860 ( .A1(n1390), .A2(n1467), .B(n1389), .C(n1388), .ZN(
        MEMCTRL_MEM_to_mem_data[5]) );
  INVD1BWP12T U1861 ( .I(RF_MEMCTRL_data_reg[12]), .ZN(n1394) );
  MAOI22D0BWP12T U1862 ( .A1(n1474), .A2(
        memory_interface_inst1_delay_data_in32[28]), .B1(n1391), .B2(n1447), 
        .ZN(n1393) );
  ND2D1BWP12T U1863 ( .A1(n1448), .A2(
        memory_interface_inst1_delay_data_in32[12]), .ZN(n1392) );
  OAI211D1BWP12T U1864 ( .A1(n1394), .A2(n1467), .B(n1393), .C(n1392), .ZN(
        MEMCTRL_MEM_to_mem_data[4]) );
  ND2D1BWP12T U1865 ( .A1(MEMCTRL_IN_address[10]), .A2(n1551), .ZN(n1395) );
  OAI221D1BWP12T U1866 ( .A1(memory_interface_inst1_delay_addr_for_adder[10]), 
        .A2(n1398), .B1(n1397), .B2(n1396), .C(n1395), .ZN(
        MEMCTRL_MEM_to_mem_address[10]) );
  INVD1BWP12T U1867 ( .I(RF_MEMCTRL_data_reg[15]), .ZN(n1402) );
  MAOI22D0BWP12T U1868 ( .A1(n1474), .A2(
        memory_interface_inst1_delay_data_in32[31]), .B1(n1372), .B2(n1447), 
        .ZN(n1401) );
  ND2D1BWP12T U1869 ( .A1(n1448), .A2(
        memory_interface_inst1_delay_data_in32[15]), .ZN(n1400) );
  OAI211D1BWP12T U1870 ( .A1(n1402), .A2(n1467), .B(n1401), .C(n1400), .ZN(
        MEMCTRL_MEM_to_mem_data[7]) );
  INVD1BWP12T U1871 ( .I(RF_MEMCTRL_data_reg[11]), .ZN(n1406) );
  MAOI22D0BWP12T U1872 ( .A1(n1474), .A2(
        memory_interface_inst1_delay_data_in32[27]), .B1(n1403), .B2(n1447), 
        .ZN(n1405) );
  ND2D1BWP12T U1873 ( .A1(n1448), .A2(
        memory_interface_inst1_delay_data_in32[11]), .ZN(n1404) );
  OAI211D1BWP12T U1874 ( .A1(n1406), .A2(n1467), .B(n1405), .C(n1404), .ZN(
        MEMCTRL_MEM_to_mem_data[3]) );
  RCIAO21D0BWP12T U1875 ( .A1(n1407), .A2(n1551), .B(n1434), .ZN(n1452) );
  INVD1BWP12T U1876 ( .I(n1452), .ZN(n1408) );
  AOI22D1BWP12T U1877 ( .A1(memory_interface_inst1_delay_addr_for_adder[7]), 
        .A2(n1408), .B1(MEMCTRL_IN_address[7]), .B2(n1551), .ZN(n1409) );
  OAI31D1BWP12T U1878 ( .A1(memory_interface_inst1_delay_addr_for_adder[7]), 
        .A2(n1464), .A3(n1410), .B(n1409), .ZN(MEMCTRL_MEM_to_mem_address[7])
         );
  RCIAO21D0BWP12T U1879 ( .A1(n1411), .A2(n1551), .B(n1434), .ZN(n1456) );
  INVD1BWP12T U1880 ( .I(n1456), .ZN(n1413) );
  AO222D1BWP12T U1881 ( .A1(n1422), .A2(n1412), .B1(n1420), .B2(
        RF_MEMCTRL_address_reg[4]), .C1(ALU_MISC_OUT_result[4]), .C2(n1419), 
        .Z(MEMCTRL_IN_address[3]) );
  AOI22D1BWP12T U1882 ( .A1(memory_interface_inst1_delay_addr_for_adder[3]), 
        .A2(n1413), .B1(MEMCTRL_IN_address[3]), .B2(n1551), .ZN(n1414) );
  OAI31D1BWP12T U1883 ( .A1(memory_interface_inst1_delay_addr_for_adder[3]), 
        .A2(n1464), .A3(n1415), .B(n1414), .ZN(MEMCTRL_MEM_to_mem_address[3])
         );
  INVD1BWP12T U1884 ( .I(n1556), .ZN(n1417) );
  AO31D1BWP12T U1885 ( .A1(n1557), .A2(DEC_MEMCTRL_memory_store_request), .A3(
        n1417), .B(n1416), .Z(MEMCTRL_MEM_to_mem_write_enable) );
  INVD1BWP12T U1886 ( .I(memory_interface_inst1_delay_addr_for_adder[1]), .ZN(
        n1425) );
  ND3D1BWP12T U1887 ( .A1(n1418), .A2(
        memory_interface_inst1_delay_addr_for_adder[0]), .A3(n1425), .ZN(n1424) );
  AO222D1BWP12T U1888 ( .A1(n1422), .A2(n1421), .B1(n1420), .B2(
        RF_MEMCTRL_address_reg[2]), .C1(ALU_MISC_OUT_result[2]), .C2(n1419), 
        .Z(MEMCTRL_IN_address[1]) );
  ND2D1BWP12T U1889 ( .A1(MEMCTRL_IN_address[1]), .A2(n1551), .ZN(n1423) );
  OAI211D1BWP12T U1890 ( .A1(n1460), .A2(n1425), .B(n1424), .C(n1423), .ZN(
        MEMCTRL_MEM_to_mem_address[1]) );
  INVD1BWP12T U1891 ( .I(RF_MEMCTRL_data_reg[14]), .ZN(n1429) );
  MAOI22D0BWP12T U1892 ( .A1(n1474), .A2(
        memory_interface_inst1_delay_data_in32[30]), .B1(n1426), .B2(n1447), 
        .ZN(n1428) );
  ND2D1BWP12T U1893 ( .A1(n1448), .A2(
        memory_interface_inst1_delay_data_in32[14]), .ZN(n1427) );
  OAI211D1BWP12T U1894 ( .A1(n1429), .A2(n1467), .B(n1428), .C(n1427), .ZN(
        MEMCTRL_MEM_to_mem_data[6]) );
  AOI22D1BWP12T U1895 ( .A1(n1434), .A2(
        memory_interface_inst1_delay_addr_for_adder[0]), .B1(
        MEMCTRL_IN_address[0]), .B2(n1551), .ZN(n1430) );
  OAI21D1BWP12T U1896 ( .A1(memory_interface_inst1_delay_addr_for_adder[0]), 
        .A2(n1464), .B(n1430), .ZN(MEMCTRL_MEM_to_mem_address[0]) );
  INVD1BWP12T U1897 ( .I(RF_MEMCTRL_data_reg[10]), .ZN(n1433) );
  INVD1BWP12T U1898 ( .I(MEM_MEMCTRL_from_mem_data[2]), .ZN(n1538) );
  MAOI22D0BWP12T U1899 ( .A1(n1474), .A2(
        memory_interface_inst1_delay_data_in32[26]), .B1(n1538), .B2(n1447), 
        .ZN(n1432) );
  ND2D1BWP12T U1900 ( .A1(n1448), .A2(
        memory_interface_inst1_delay_data_in32[10]), .ZN(n1431) );
  OAI211D1BWP12T U1901 ( .A1(n1433), .A2(n1467), .B(n1432), .C(n1431), .ZN(
        MEMCTRL_MEM_to_mem_data[2]) );
  RCIAO21D0BWP12T U1902 ( .A1(n1435), .A2(n1551), .B(n1434), .ZN(n1439) );
  INVD1BWP12T U1903 ( .I(n1439), .ZN(n1436) );
  AOI22D1BWP12T U1904 ( .A1(memory_interface_inst1_delay_addr_for_adder[5]), 
        .A2(n1436), .B1(MEMCTRL_IN_address[5]), .B2(n1551), .ZN(n1437) );
  OAI31D1BWP12T U1905 ( .A1(memory_interface_inst1_delay_addr_for_adder[5]), 
        .A2(n1464), .A3(n1438), .B(n1437), .ZN(MEMCTRL_MEM_to_mem_address[5])
         );
  OAI21D1BWP12T U1906 ( .A1(memory_interface_inst1_delay_addr_for_adder[5]), 
        .A2(n1551), .B(n1439), .ZN(n1440) );
  AOI22D1BWP12T U1907 ( .A1(memory_interface_inst1_delay_addr_for_adder[6]), 
        .A2(n1440), .B1(MEMCTRL_IN_address[6]), .B2(n1551), .ZN(n1441) );
  OAI31D1BWP12T U1908 ( .A1(memory_interface_inst1_delay_addr_for_adder[6]), 
        .A2(n1464), .A3(n1442), .B(n1441), .ZN(MEMCTRL_MEM_to_mem_address[6])
         );
  INVD1BWP12T U1909 ( .I(RF_MEMCTRL_data_reg[9]), .ZN(n1446) );
  MAOI22D0BWP12T U1910 ( .A1(n1474), .A2(
        memory_interface_inst1_delay_data_in32[25]), .B1(n1443), .B2(n1447), 
        .ZN(n1445) );
  ND2D1BWP12T U1911 ( .A1(n1448), .A2(
        memory_interface_inst1_delay_data_in32[9]), .ZN(n1444) );
  OAI211D1BWP12T U1912 ( .A1(n1446), .A2(n1467), .B(n1445), .C(n1444), .ZN(
        MEMCTRL_MEM_to_mem_data[1]) );
  INVD1BWP12T U1913 ( .I(RF_MEMCTRL_data_reg[8]), .ZN(n1451) );
  INVD1BWP12T U1914 ( .I(MEM_MEMCTRL_from_mem_data[0]), .ZN(n1539) );
  MAOI22D0BWP12T U1915 ( .A1(n1474), .A2(
        memory_interface_inst1_delay_data_in32[24]), .B1(n1539), .B2(n1447), 
        .ZN(n1450) );
  ND2D1BWP12T U1916 ( .A1(n1448), .A2(
        memory_interface_inst1_delay_data_in32[8]), .ZN(n1449) );
  OAI211D1BWP12T U1917 ( .A1(n1451), .A2(n1467), .B(n1450), .C(n1449), .ZN(
        MEMCTRL_MEM_to_mem_data[0]) );
  OAI21D1BWP12T U1918 ( .A1(memory_interface_inst1_delay_addr_for_adder[7]), 
        .A2(n1551), .B(n1452), .ZN(n1453) );
  AOI22D1BWP12T U1919 ( .A1(memory_interface_inst1_delay_addr_for_adder[8]), 
        .A2(n1453), .B1(MEMCTRL_IN_address[8]), .B2(n1551), .ZN(n1454) );
  OAI31D1BWP12T U1920 ( .A1(memory_interface_inst1_delay_addr_for_adder[8]), 
        .A2(n1464), .A3(n1455), .B(n1454), .ZN(MEMCTRL_MEM_to_mem_address[8])
         );
  OAI21D1BWP12T U1921 ( .A1(memory_interface_inst1_delay_addr_for_adder[3]), 
        .A2(n1551), .B(n1456), .ZN(n1457) );
  AOI22D1BWP12T U1922 ( .A1(memory_interface_inst1_delay_addr_for_adder[4]), 
        .A2(n1457), .B1(MEMCTRL_IN_address[4]), .B2(n1551), .ZN(n1458) );
  OAI31D1BWP12T U1923 ( .A1(memory_interface_inst1_delay_addr_for_adder[4]), 
        .A2(n1464), .A3(n1459), .B(n1458), .ZN(MEMCTRL_MEM_to_mem_address[4])
         );
  ND2D1BWP12T U1924 ( .A1(memory_interface_inst1_delay_addr_for_adder[0]), 
        .A2(memory_interface_inst1_delay_addr_for_adder[1]), .ZN(n1463) );
  OAI21D1BWP12T U1925 ( .A1(memory_interface_inst1_delay_addr_for_adder[1]), 
        .A2(n1551), .B(n1460), .ZN(n1461) );
  AOI22D1BWP12T U1926 ( .A1(memory_interface_inst1_delay_addr_for_adder[2]), 
        .A2(n1461), .B1(MEMCTRL_IN_address[2]), .B2(n1551), .ZN(n1462) );
  OAI31D1BWP12T U1927 ( .A1(memory_interface_inst1_delay_addr_for_adder[2]), 
        .A2(n1464), .A3(n1463), .B(n1462), .ZN(MEMCTRL_MEM_to_mem_address[2])
         );
  CKND0BWP12T U1928 ( .I(DEC_MEMCTRL_load_store_width[0]), .ZN(n1471) );
  CKND0BWP12T U1929 ( .I(DEC_MEMCTRL_memory_store_request), .ZN(n1468) );
  OAI21D0BWP12T U1930 ( .A1(DEC_MEMCTRL_load_store_width[1]), .A2(n1468), .B(
        n1555), .ZN(n1469) );
  OAI211D0BWP12T U1931 ( .A1(n1555), .A2(n1471), .B(n1470), .C(n1469), .ZN(
        n1473) );
  AOI21D1BWP12T U1932 ( .A1(n1473), .A2(n1472), .B(reset), .ZN(
        memory_interface_inst1_fsm_N33) );
  INVD1BWP12T U1933 ( .I(memory_interface_inst1_fsm_state_3_), .ZN(n1475) );
  AOI21D0BWP12T U1934 ( .A1(n1476), .A2(n1475), .B(n1474), .ZN(n1477) );
  OAI22D1BWP12T U1935 ( .A1(n1478), .A2(n1556), .B1(reset), .B2(n1477), .ZN(
        memory_interface_inst1_fsm_N34) );
  AO221D1BWP12T U1936 ( .A1(n1479), .A2(MEMCTRL_RF_IF_data_in[10]), .B1(n754), 
        .B2(Instruction_Fetch_inst1_fetched_instruction_reg_10_), .C(reset), 
        .Z(Instruction_Fetch_inst1_N93) );
  AO221D1BWP12T U1937 ( .A1(n754), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_13_), .B1(n1479), .B2(
        MEMCTRL_RF_IF_data_in[13]), .C(reset), .Z(Instruction_Fetch_inst1_N96)
         );
  AO221D1BWP12T U1938 ( .A1(n754), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_11_), .B1(n1479), .B2(
        MEMCTRL_RF_IF_data_in[11]), .C(reset), .Z(Instruction_Fetch_inst1_N94)
         );
  AO221D1BWP12T U1939 ( .A1(n754), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_9_), .B1(n1479), .B2(
        MEMCTRL_RF_IF_data_in[9]), .C(reset), .Z(Instruction_Fetch_inst1_N92)
         );
  AO221D1BWP12T U1940 ( .A1(n754), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_15_), .B1(n1479), .B2(
        MEMCTRL_RF_IF_data_in[15]), .C(reset), .Z(Instruction_Fetch_inst1_N98)
         );
  AOI21D0BWP12T U1941 ( .A1(n1481), .A2(n1480), .B(
        Instruction_Fetch_inst1_first_instruction_fetched), .ZN(n1482) );
  NR2D1BWP12T U1942 ( .A1(reset), .A2(n1482), .ZN(n862) );
  NR2D1BWP12T U1943 ( .A1(n1645), .A2(n1483), .ZN(n1487) );
  OAI22D1BWP12T U1944 ( .A1(n1602), .A2(n1646), .B1(n1487), .B2(n1484), .ZN(
        n853) );
  OAI22D1BWP12T U1945 ( .A1(n1618), .A2(n1646), .B1(n1487), .B2(n1485), .ZN(
        n855) );
  OAI22D1BWP12T U1946 ( .A1(n1617), .A2(n1646), .B1(n1487), .B2(n1486), .ZN(
        n854) );
  NR2D1BWP12T U1947 ( .A1(irdecode_inst1_N705), .A2(n1488), .ZN(n1498) );
  OA21XD1BWP12T U1948 ( .A1(n1498), .A2(n1503), .B(n1506), .Z(n1496) );
  CKND2D1BWP12T U1949 ( .A1(n1490), .A2(n1489), .ZN(n1492) );
  AOI22D0BWP12T U1950 ( .A1(n1682), .A2(irdecode_inst1_step[3]), .B1(n1501), 
        .B2(n1492), .ZN(n1491) );
  ND2D1BWP12T U1951 ( .A1(n1496), .A2(n1491), .ZN(irdecode_inst1_next_step_3_)
         );
  INR2D1BWP12T U1952 ( .A1(n1493), .B1(n1492), .ZN(n1505) );
  AOI22D0BWP12T U1953 ( .A1(n1682), .A2(irdecode_inst1_step[4]), .B1(n1595), 
        .B2(n1494), .ZN(n1495) );
  OAI211D1BWP12T U1954 ( .A1(n1505), .A2(n1509), .B(n1496), .C(n1495), .ZN(
        irdecode_inst1_next_step_4_) );
  ND2D1BWP12T U1955 ( .A1(n1498), .A2(n1497), .ZN(n1596) );
  INVD1BWP12T U1956 ( .I(n1596), .ZN(n1504) );
  ND2XD0BWP12T U1957 ( .A1(n1505), .A2(n1499), .ZN(n1500) );
  AOI22D0BWP12T U1958 ( .A1(n1682), .A2(irdecode_inst1_step[5]), .B1(n1501), 
        .B2(n1500), .ZN(n1502) );
  OAI211D1BWP12T U1959 ( .A1(n1504), .A2(n1503), .B(n1506), .C(n1502), .ZN(
        irdecode_inst1_next_step_5_) );
  AOI32D0BWP12T U1960 ( .A1(n1507), .A2(n1506), .A3(n1505), .B1(n1509), .B2(
        n1506), .ZN(n1598) );
  AOI211D0BWP12T U1961 ( .A1(n1682), .A2(irdecode_inst1_step[7]), .B(n1595), 
        .C(n1598), .ZN(n1508) );
  OAI21D1BWP12T U1962 ( .A1(n1510), .A2(n1509), .B(n1508), .ZN(
        irdecode_inst1_next_step_7_) );
  TPND2D0BWP12T U1963 ( .A1(n1682), .A2(DEC_RF_offset_b[11]), .ZN(n1511) );
  OAI211D1BWP12T U1964 ( .A1(n1628), .A2(n1517), .B(n1512), .C(n1511), .ZN(
        n798) );
  CKND2D0BWP12T U1965 ( .A1(n1513), .A2(n1536), .ZN(n1516) );
  AOI21D0BWP12T U1966 ( .A1(n1682), .A2(DEC_RF_offset_b[9]), .B(n1514), .ZN(
        n1515) );
  OAI211D1BWP12T U1967 ( .A1(n1583), .A2(n1517), .B(n1516), .C(n1515), .ZN(
        n800) );
  MUX2D1BWP12T U1968 ( .I0(RF_OUT_n), .I1(ALU_OUT_n), .S(
        DEC_CPSR_update_flag_n), .Z(new_n) );
  CKND2D0BWP12T U1969 ( .A1(n1573), .A2(IF_DEC_instruction[1]), .ZN(n1519) );
  OAI211D1BWP12T U1970 ( .A1(n1647), .A2(n1625), .B(n1519), .C(n1518), .ZN(
        n1520) );
  AOI211D1BWP12T U1971 ( .A1(n1657), .A2(IF_DEC_instruction[6]), .B(n1521), 
        .C(n1520), .ZN(n1523) );
  CKND0BWP12T U1972 ( .I(DEC_RF_offset_b[1]), .ZN(n1522) );
  OAI222D1BWP12T U1973 ( .A1(n1570), .A2(n1529), .B1(n1679), .B2(n1523), .C1(
        n1527), .C2(n1522), .ZN(n808) );
  INVD1BWP12T U1974 ( .I(n1657), .ZN(n1623) );
  INVD0BWP12T U1975 ( .I(IF_DEC_instruction[1]), .ZN(n1641) );
  OAI22D1BWP12T U1976 ( .A1(n1619), .A2(n1617), .B1(n1641), .B2(n1625), .ZN(
        n1525) );
  OAI22D0BWP12T U1977 ( .A1(n1624), .A2(n1531), .B1(n1583), .B2(n1570), .ZN(
        n1524) );
  AOI211D1BWP12T U1978 ( .A1(n1634), .A2(IF_DEC_instruction[0]), .B(n1525), 
        .C(n1524), .ZN(n1528) );
  CKND0BWP12T U1979 ( .I(DEC_RF_offset_b[2]), .ZN(n1526) );
  OAI222D1BWP12T U1980 ( .A1(n1623), .A2(n1529), .B1(n1679), .B2(n1528), .C1(
        n1527), .C2(n1526), .ZN(n807) );
  MUX2D1BWP12T U1981 ( .I0(RF_OUT_z), .I1(ALU_OUT_z), .S(
        DEC_CPSR_update_flag_z), .Z(new_z) );
  NR2XD0BWP12T U1982 ( .A1(n1623), .A2(n1583), .ZN(n1533) );
  CKND2D1BWP12T U1983 ( .A1(n1604), .A2(n1530), .ZN(n1627) );
  OAI22D1BWP12T U1984 ( .A1(n1676), .A2(n1627), .B1(n1531), .B2(n1625), .ZN(
        n1532) );
  AOI211D1BWP12T U1985 ( .A1(n1573), .A2(IF_DEC_instruction[3]), .B(n1533), 
        .C(n1532), .ZN(n1534) );
  OAI21D1BWP12T U1986 ( .A1(n1535), .A2(n1641), .B(n1534), .ZN(n1537) );
  AO222D1BWP12T U1987 ( .A1(n1537), .A2(n1578), .B1(n1536), .B2(n1632), .C1(
        n1682), .C2(DEC_RF_offset_b[3]), .Z(n806) );
  OAI21D1BWP12T U1988 ( .A1(n1538), .A2(n1549), .B(n1547), .ZN(
        MEMCTRL_RF_IF_data_in[26]) );
  OAI21D1BWP12T U1989 ( .A1(n1539), .A2(n1549), .B(n1547), .ZN(
        MEMCTRL_RF_IF_data_in[24]) );
  OAI21D1BWP12T U1990 ( .A1(n1549), .A2(n1540), .B(n1547), .ZN(
        MEMCTRL_RF_IF_data_in[23]) );
  OAI21D1BWP12T U1991 ( .A1(n1541), .A2(n1549), .B(n1547), .ZN(
        MEMCTRL_RF_IF_data_in[22]) );
  OAI21D1BWP12T U1992 ( .A1(n1542), .A2(n1549), .B(n1547), .ZN(
        MEMCTRL_RF_IF_data_in[21]) );
  OAI21D1BWP12T U1993 ( .A1(n1549), .A2(n1543), .B(n1547), .ZN(
        MEMCTRL_RF_IF_data_in[19]) );
  OAI21D1BWP12T U1994 ( .A1(n1549), .A2(n1544), .B(n1547), .ZN(
        MEMCTRL_RF_IF_data_in[18]) );
  OAI21D1BWP12T U1995 ( .A1(n1549), .A2(n1545), .B(n1547), .ZN(
        MEMCTRL_RF_IF_data_in[17]) );
  OAI21D1BWP12T U1996 ( .A1(n1549), .A2(n1546), .B(n1547), .ZN(
        MEMCTRL_RF_IF_data_in[16]) );
  OAI21D1BWP12T U1997 ( .A1(n1549), .A2(n1548), .B(n1547), .ZN(
        MEMCTRL_RF_IF_data_in[20]) );
  CKND0BWP12T U1998 ( .I(n1559), .ZN(n1569) );
  MOAI22D0BWP12T U1999 ( .A1(n1569), .A2(n1560), .B1(n1567), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_5_), .ZN(
        Instruction_Fetch_inst1_N88) );
  MOAI22D0BWP12T U2000 ( .A1(n1569), .A2(n1561), .B1(n1567), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_3_), .ZN(
        Instruction_Fetch_inst1_N86) );
  MOAI22D0BWP12T U2001 ( .A1(n1569), .A2(n1562), .B1(n1567), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_7_), .ZN(
        Instruction_Fetch_inst1_N90) );
  MOAI22D0BWP12T U2002 ( .A1(n1569), .A2(n1563), .B1(n1567), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_6_), .ZN(
        Instruction_Fetch_inst1_N89) );
  MOAI22D0BWP12T U2003 ( .A1(n1569), .A2(n1564), .B1(n1567), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_4_), .ZN(
        Instruction_Fetch_inst1_N87) );
  MOAI22D0BWP12T U2004 ( .A1(n1569), .A2(n1565), .B1(n1567), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_1_), .ZN(
        Instruction_Fetch_inst1_N84) );
  MOAI22D0BWP12T U2005 ( .A1(n1569), .A2(n1566), .B1(n1567), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_2_), .ZN(
        Instruction_Fetch_inst1_N85) );
  MOAI22D0BWP12T U2006 ( .A1(n1569), .A2(n1568), .B1(n1567), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_0_), .ZN(
        Instruction_Fetch_inst1_N83) );
  NR2D0BWP12T U2007 ( .A1(n1570), .A2(n1617), .ZN(n1572) );
  AOI211D0BWP12T U2008 ( .A1(n1573), .A2(IF_DEC_instruction[0]), .B(n1572), 
        .C(n1571), .ZN(n1574) );
  MOAI22D0BWP12T U2009 ( .A1(n1574), .A2(n1679), .B1(n1682), .B2(
        DEC_RF_offset_b[0]), .ZN(n809) );
  CKND0BWP12T U2010 ( .I(n1579), .ZN(n1580) );
  ND4D0BWP12T U2011 ( .A1(n1600), .A2(n1580), .A3(n1584), .A4(
        IF_DEC_instruction[7]), .ZN(n1588) );
  AO32D0BWP12T U2012 ( .A1(n1600), .A2(n1583), .A3(n1582), .B1(n1581), .B2(
        n1600), .Z(n1585) );
  OAI31D0BWP12T U2013 ( .A1(n1604), .A2(n1586), .A3(n1585), .B(n1584), .ZN(
        n1587) );
  IND3D1BWP12T U2014 ( .A1(n1589), .B1(n1588), .B2(n1587), .ZN(
        irdecode_inst1_next_update_flag_c) );
  NR2D0BWP12T U2015 ( .A1(n1590), .A2(n1676), .ZN(n1592) );
  AOI211D0BWP12T U2016 ( .A1(n1593), .A2(IF_DEC_instruction[1]), .B(n1592), 
        .C(n1591), .ZN(n1594) );
  MOAI22D0BWP12T U2017 ( .A1(n1594), .A2(n1679), .B1(n1682), .B2(
        DEC_RF_alu_write_to_reg[1]), .ZN(n819) );
  OAI32D0BWP12T U2018 ( .A1(n1598), .A2(n1597), .A3(n1596), .B1(n1595), .B2(
        n1598), .ZN(n1599) );
  IOA21D1BWP12T U2019 ( .A1(n1682), .A2(irdecode_inst1_step[6]), .B(n1599), 
        .ZN(irdecode_inst1_next_step_6_) );
  NR2D0BWP12T U2020 ( .A1(irdecode_inst1_N907), .A2(
        irdecode_inst1_next_step_0_), .ZN(n1611) );
  AOI22D0BWP12T U2021 ( .A1(n1602), .A2(n1601), .B1(n1600), .B2(
        IF_DEC_instruction[6]), .ZN(n1606) );
  AOI32D0BWP12T U2022 ( .A1(n1676), .A2(n1677), .A3(n1604), .B1(n1603), .B2(
        n1677), .ZN(n1605) );
  OAI211D0BWP12T U2023 ( .A1(n1608), .A2(n1607), .B(n1606), .C(n1605), .ZN(
        n1610) );
  AOI211XD0BWP12T U2024 ( .A1(n1612), .A2(n1611), .B(n1610), .C(n1609), .ZN(
        n1613) );
  MOAI22D0BWP12T U2025 ( .A1(n1613), .A2(n1679), .B1(DEC_ALU_alu_opcode[0]), 
        .B2(n1682), .ZN(n851) );
  INVD0BWP12T U2026 ( .I(IF_DEC_instruction[4]), .ZN(n1642) );
  OAI22D1BWP12T U2027 ( .A1(n1619), .A2(n1676), .B1(n1642), .B2(n1625), .ZN(
        n1615) );
  OAI22D0BWP12T U2028 ( .A1(n1624), .A2(n1618), .B1(n1623), .B2(n1628), .ZN(
        n1614) );
  AOI211D1BWP12T U2029 ( .A1(n1634), .A2(IF_DEC_instruction[3]), .B(n1615), 
        .C(n1614), .ZN(n1616) );
  MOAI22D0BWP12T U2030 ( .A1(n1616), .A2(n1679), .B1(n1682), .B2(
        DEC_RF_offset_b[5]), .ZN(n804) );
  NR2XD0BWP12T U2031 ( .A1(n1624), .A2(n1617), .ZN(n1621) );
  OAI22D1BWP12T U2032 ( .A1(n1619), .A2(n1628), .B1(n1618), .B2(n1625), .ZN(
        n1620) );
  AOI211D1BWP12T U2033 ( .A1(n1634), .A2(IF_DEC_instruction[4]), .B(n1621), 
        .C(n1620), .ZN(n1622) );
  MOAI22D0BWP12T U2034 ( .A1(n1622), .A2(n1679), .B1(n1682), .B2(
        DEC_RF_offset_b[6]), .ZN(n803) );
  OAI22D0BWP12T U2035 ( .A1(n1624), .A2(n1642), .B1(n1623), .B2(n1676), .ZN(
        n1630) );
  OAI22D1BWP12T U2036 ( .A1(n1628), .A2(n1627), .B1(n1626), .B2(n1625), .ZN(
        n1629) );
  AO211D1BWP12T U2037 ( .A1(n1632), .A2(n1631), .B(n1630), .C(n1629), .Z(n1633) );
  RCAOI21D0BWP12T U2038 ( .A1(IF_DEC_instruction[2]), .A2(n1634), .B(n1633), 
        .ZN(n1635) );
  MOAI22D0BWP12T U2039 ( .A1(n1635), .A2(n1679), .B1(n1682), .B2(
        DEC_RF_offset_b[4]), .ZN(n805) );
  MOAI22D0BWP12T U2040 ( .A1(n1647), .A2(n1646), .B1(irdecode_inst1_itstate_0_), .B2(n1645), .ZN(n860) );
  NR2D0BWP12T U2041 ( .A1(n1649), .A2(n1648), .ZN(n1650) );
  AOI211D0BWP12T U2042 ( .A1(n1653), .A2(n1652), .B(n1651), .C(n1650), .ZN(
        n1654) );
  MOAI22D0BWP12T U2043 ( .A1(n1654), .A2(n1679), .B1(
        irdecode_inst1_split_instruction), .B2(n1682), .ZN(n847) );
  OAI32D0BWP12T U2044 ( .A1(n1657), .A2(n1672), .A3(n1656), .B1(n1655), .B2(
        n1657), .ZN(n1658) );
  MOAI22D0BWP12T U2045 ( .A1(n1658), .A2(n1679), .B1(n1682), .B2(
        DEC_MEMCTRL_load_store_width[0]), .ZN(n838) );
  INVD1BWP12T U2046 ( .I(n1659), .ZN(n1669) );
  CKND0BWP12T U2047 ( .I(n1660), .ZN(n1663) );
  OAI21D0BWP12T U2048 ( .A1(n1663), .A2(n1662), .B(n1661), .ZN(n1668) );
  AOI22D0BWP12T U2049 ( .A1(n1666), .A2(IF_DEC_instruction[1]), .B1(n1665), 
        .B2(n1664), .ZN(n1667) );
  OAI211D1BWP12T U2050 ( .A1(n1670), .A2(n1669), .B(n1668), .C(n1667), .ZN(
        n1678) );
  AOI22D0BWP12T U2051 ( .A1(n1678), .A2(n1672), .B1(n1671), .B2(
        IF_DEC_instruction[1]), .ZN(n1673) );
  MOAI22D0BWP12T U2052 ( .A1(n1673), .A2(n1679), .B1(n1682), .B2(
        DEC_RF_memory_store_data_reg[1]), .ZN(n829) );
  AO211D0BWP12T U2053 ( .A1(n1682), .A2(DEC_RF_memory_write_to_reg[3]), .B(
        n1681), .C(n1680), .Z(n821) );
endmodule

