// AUTHORS: Group 06 / Julian Käuser
// Wed 08/09/2017


module memory_interface (


  );

  endmodule
