
module register_file ( readA_sel, readB_sel, readC_sel, readD_sel, write1_sel, 
        write2_sel, write1_en, write2_en, write1_in, write2_in, immediate1_in, 
        immediate2_in, next_pc_in, next_cpsr_in, next_sp_in, clk, reset, 
        regA_out, regB_out, regC_out, regD_out, pc_out, cpsr_out, sp_out, 
        next_pc_en_BAR );
  input [4:0] readA_sel;
  input [4:0] readB_sel;
  input [4:0] readC_sel;
  input [4:0] readD_sel;
  input [4:0] write1_sel;
  input [4:0] write2_sel;
  input [31:0] write1_in;
  input [31:0] write2_in;
  input [31:0] immediate1_in;
  input [31:0] immediate2_in;
  input [31:0] next_pc_in;
  input [3:0] next_cpsr_in;
  input [31:0] next_sp_in;
  output [31:0] regA_out;
  output [31:0] regB_out;
  output [31:0] regC_out;
  output [31:0] regD_out;
  output [31:0] pc_out;
  output [3:0] cpsr_out;
  output [31:0] sp_out;
  input write1_en, write2_en, clk, reset, next_pc_en_BAR;
  wire   n3668, n2136, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2137, n2167, n2294, n2326,
         n2327, n2455, n2487, n2519, n2550, n2551, n2583, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667;
  wire   [3669:3700] n;
  wire   [31:0] r0;
  wire   [31:0] r1;
  wire   [31:0] r2;
  wire   [31:0] r3;
  wire   [31:0] r4;
  wire   [31:0] r5;
  wire   [31:0] r6;
  wire   [31:0] r7;
  wire   [31:0] r8;
  wire   [31:0] r9;
  wire   [31:0] r10;
  wire   [31:0] r11;
  wire   [31:0] r12;
  wire   [31:0] lr;
  wire   [31:0] tmp1;
  wire   [31:0] spin;
  wire   [3:2] cpsrin;

  DFQD1BWP12T r0_reg_31_ ( .D(n2648), .CP(clk), .Q(r0[31]) );
  DFQD1BWP12T r0_reg_28_ ( .D(n2645), .CP(clk), .Q(r0[28]) );
  DFQD1BWP12T r0_reg_27_ ( .D(n2644), .CP(clk), .Q(r0[27]) );
  DFQD1BWP12T r0_reg_26_ ( .D(n2643), .CP(clk), .Q(r0[26]) );
  DFQD1BWP12T r0_reg_25_ ( .D(n2642), .CP(clk), .Q(r0[25]) );
  DFQD1BWP12T r0_reg_24_ ( .D(n2641), .CP(clk), .Q(r0[24]) );
  DFQD1BWP12T r0_reg_23_ ( .D(n2640), .CP(clk), .Q(r0[23]) );
  DFQD1BWP12T r0_reg_22_ ( .D(n2639), .CP(clk), .Q(r0[22]) );
  DFQD1BWP12T r0_reg_21_ ( .D(n2638), .CP(clk), .Q(r0[21]) );
  DFQD1BWP12T r0_reg_20_ ( .D(n2637), .CP(clk), .Q(r0[20]) );
  DFQD1BWP12T r0_reg_19_ ( .D(n2636), .CP(clk), .Q(r0[19]) );
  DFQD1BWP12T r0_reg_18_ ( .D(n2635), .CP(clk), .Q(r0[18]) );
  DFQD1BWP12T r0_reg_17_ ( .D(n2634), .CP(clk), .Q(r0[17]) );
  DFQD1BWP12T r0_reg_16_ ( .D(n2633), .CP(clk), .Q(r0[16]) );
  DFQD1BWP12T r0_reg_15_ ( .D(n2632), .CP(clk), .Q(r0[15]) );
  DFQD1BWP12T r0_reg_14_ ( .D(n2631), .CP(clk), .Q(r0[14]) );
  DFQD1BWP12T r0_reg_13_ ( .D(n2630), .CP(clk), .Q(r0[13]) );
  DFQD1BWP12T r0_reg_12_ ( .D(n2629), .CP(clk), .Q(r0[12]) );
  DFQD1BWP12T r0_reg_11_ ( .D(n2628), .CP(clk), .Q(r0[11]) );
  DFQD1BWP12T r0_reg_10_ ( .D(n2627), .CP(clk), .Q(r0[10]) );
  DFQD1BWP12T r0_reg_9_ ( .D(n2626), .CP(clk), .Q(r0[9]) );
  DFQD1BWP12T r0_reg_8_ ( .D(n2625), .CP(clk), .Q(r0[8]) );
  DFQD1BWP12T r0_reg_7_ ( .D(n2624), .CP(clk), .Q(r0[7]) );
  DFQD1BWP12T r0_reg_6_ ( .D(n2623), .CP(clk), .Q(r0[6]) );
  DFQD1BWP12T r0_reg_5_ ( .D(n2622), .CP(clk), .Q(r0[5]) );
  DFQD1BWP12T r0_reg_4_ ( .D(n2621), .CP(clk), .Q(r0[4]) );
  DFQD1BWP12T r0_reg_3_ ( .D(n2620), .CP(clk), .Q(r0[3]) );
  DFQD1BWP12T r0_reg_2_ ( .D(n2619), .CP(clk), .Q(r0[2]) );
  DFQD1BWP12T r0_reg_1_ ( .D(n2618), .CP(clk), .Q(r0[1]) );
  DFQD1BWP12T r0_reg_0_ ( .D(n2617), .CP(clk), .Q(r0[0]) );
  DFQD1BWP12T r1_reg_31_ ( .D(n2616), .CP(clk), .Q(r1[31]) );
  DFQD1BWP12T r1_reg_28_ ( .D(n2613), .CP(clk), .Q(r1[28]) );
  DFQD1BWP12T r1_reg_27_ ( .D(n2612), .CP(clk), .Q(r1[27]) );
  DFQD1BWP12T r1_reg_26_ ( .D(n2611), .CP(clk), .Q(r1[26]) );
  DFQD1BWP12T r1_reg_24_ ( .D(n2609), .CP(clk), .Q(r1[24]) );
  DFQD1BWP12T r1_reg_23_ ( .D(n2608), .CP(clk), .Q(r1[23]) );
  DFQD1BWP12T r1_reg_22_ ( .D(n2607), .CP(clk), .Q(r1[22]) );
  DFQD1BWP12T r1_reg_21_ ( .D(n2606), .CP(clk), .Q(r1[21]) );
  DFQD1BWP12T r1_reg_20_ ( .D(n2605), .CP(clk), .Q(r1[20]) );
  DFQD1BWP12T r1_reg_19_ ( .D(n2604), .CP(clk), .Q(r1[19]) );
  DFQD1BWP12T r1_reg_18_ ( .D(n2603), .CP(clk), .Q(r1[18]) );
  DFQD1BWP12T r1_reg_17_ ( .D(n2602), .CP(clk), .Q(r1[17]) );
  DFQD1BWP12T r1_reg_16_ ( .D(n2601), .CP(clk), .Q(r1[16]) );
  DFQD1BWP12T r1_reg_15_ ( .D(n2600), .CP(clk), .Q(r1[15]) );
  DFQD1BWP12T r1_reg_14_ ( .D(n2599), .CP(clk), .Q(r1[14]) );
  DFQD1BWP12T r1_reg_13_ ( .D(n2598), .CP(clk), .Q(r1[13]) );
  DFQD1BWP12T r1_reg_11_ ( .D(n2596), .CP(clk), .Q(r1[11]) );
  DFQD1BWP12T r1_reg_10_ ( .D(n2595), .CP(clk), .Q(r1[10]) );
  DFQD1BWP12T r1_reg_9_ ( .D(n2594), .CP(clk), .Q(r1[9]) );
  DFQD1BWP12T r1_reg_8_ ( .D(n2593), .CP(clk), .Q(r1[8]) );
  DFQD1BWP12T r1_reg_7_ ( .D(n2592), .CP(clk), .Q(r1[7]) );
  DFQD1BWP12T r1_reg_6_ ( .D(n2591), .CP(clk), .Q(r1[6]) );
  DFQD1BWP12T r1_reg_5_ ( .D(n2590), .CP(clk), .Q(r1[5]) );
  DFQD1BWP12T r1_reg_4_ ( .D(n2589), .CP(clk), .Q(r1[4]) );
  DFQD1BWP12T r1_reg_2_ ( .D(n2587), .CP(clk), .Q(r1[2]) );
  DFQD1BWP12T r1_reg_1_ ( .D(n2586), .CP(clk), .Q(r1[1]) );
  DFQD1BWP12T r1_reg_0_ ( .D(n2585), .CP(clk), .Q(r1[0]) );
  DFQD1BWP12T r2_reg_31_ ( .D(n2584), .CP(clk), .Q(r2[31]) );
  DFQD1BWP12T r2_reg_29_ ( .D(n2582), .CP(clk), .Q(r2[29]) );
  DFQD1BWP12T r2_reg_28_ ( .D(n2581), .CP(clk), .Q(r2[28]) );
  DFQD1BWP12T r2_reg_27_ ( .D(n2580), .CP(clk), .Q(r2[27]) );
  DFQD1BWP12T r2_reg_26_ ( .D(n2579), .CP(clk), .Q(r2[26]) );
  DFQD1BWP12T r2_reg_25_ ( .D(n2578), .CP(clk), .Q(r2[25]) );
  DFQD1BWP12T r2_reg_24_ ( .D(n2577), .CP(clk), .Q(r2[24]) );
  DFQD1BWP12T r2_reg_23_ ( .D(n2576), .CP(clk), .Q(r2[23]) );
  DFQD1BWP12T r2_reg_22_ ( .D(n2575), .CP(clk), .Q(r2[22]) );
  DFQD1BWP12T r2_reg_21_ ( .D(n2574), .CP(clk), .Q(r2[21]) );
  DFQD1BWP12T r2_reg_20_ ( .D(n2573), .CP(clk), .Q(r2[20]) );
  DFQD1BWP12T r2_reg_19_ ( .D(n2572), .CP(clk), .Q(r2[19]) );
  DFQD1BWP12T r2_reg_18_ ( .D(n2571), .CP(clk), .Q(r2[18]) );
  DFQD1BWP12T r2_reg_17_ ( .D(n2570), .CP(clk), .Q(r2[17]) );
  DFQD1BWP12T r2_reg_16_ ( .D(n2569), .CP(clk), .Q(r2[16]) );
  DFQD1BWP12T r2_reg_15_ ( .D(n2568), .CP(clk), .Q(r2[15]) );
  DFQD1BWP12T r2_reg_14_ ( .D(n2567), .CP(clk), .Q(r2[14]) );
  DFQD1BWP12T r2_reg_13_ ( .D(n2566), .CP(clk), .Q(r2[13]) );
  DFQD1BWP12T r2_reg_11_ ( .D(n2564), .CP(clk), .Q(r2[11]) );
  DFQD1BWP12T r2_reg_10_ ( .D(n2563), .CP(clk), .Q(r2[10]) );
  DFQD1BWP12T r2_reg_9_ ( .D(n2562), .CP(clk), .Q(r2[9]) );
  DFQD1BWP12T r2_reg_8_ ( .D(n2561), .CP(clk), .Q(r2[8]) );
  DFQD1BWP12T r2_reg_7_ ( .D(n2560), .CP(clk), .Q(r2[7]) );
  DFQD1BWP12T r2_reg_6_ ( .D(n2559), .CP(clk), .Q(r2[6]) );
  DFQD1BWP12T r2_reg_5_ ( .D(n2558), .CP(clk), .Q(r2[5]) );
  DFQD1BWP12T r2_reg_4_ ( .D(n2557), .CP(clk), .Q(r2[4]) );
  DFQD1BWP12T r2_reg_3_ ( .D(n2556), .CP(clk), .Q(r2[3]) );
  DFQD1BWP12T r2_reg_2_ ( .D(n2555), .CP(clk), .Q(r2[2]) );
  DFQD1BWP12T r2_reg_1_ ( .D(n2554), .CP(clk), .Q(r2[1]) );
  DFQD1BWP12T r2_reg_0_ ( .D(n2553), .CP(clk), .Q(r2[0]) );
  DFQD1BWP12T r3_reg_31_ ( .D(n2552), .CP(clk), .Q(r3[31]) );
  DFQD1BWP12T r3_reg_28_ ( .D(n2549), .CP(clk), .Q(r3[28]) );
  DFQD1BWP12T r3_reg_27_ ( .D(n2548), .CP(clk), .Q(r3[27]) );
  DFQD1BWP12T r3_reg_26_ ( .D(n2547), .CP(clk), .Q(r3[26]) );
  DFQD1BWP12T r3_reg_25_ ( .D(n2546), .CP(clk), .Q(r3[25]) );
  DFQD1BWP12T r3_reg_24_ ( .D(n2545), .CP(clk), .Q(r3[24]) );
  DFQD1BWP12T r3_reg_23_ ( .D(n2544), .CP(clk), .Q(r3[23]) );
  DFQD1BWP12T r3_reg_22_ ( .D(n2543), .CP(clk), .Q(r3[22]) );
  DFQD1BWP12T r3_reg_21_ ( .D(n2542), .CP(clk), .Q(r3[21]) );
  DFQD1BWP12T r3_reg_20_ ( .D(n2541), .CP(clk), .Q(r3[20]) );
  DFQD1BWP12T r3_reg_19_ ( .D(n2540), .CP(clk), .Q(r3[19]) );
  DFQD1BWP12T r3_reg_18_ ( .D(n2539), .CP(clk), .Q(r3[18]) );
  DFQD1BWP12T r3_reg_17_ ( .D(n2538), .CP(clk), .Q(r3[17]) );
  DFQD1BWP12T r3_reg_16_ ( .D(n2537), .CP(clk), .Q(r3[16]) );
  DFQD1BWP12T r3_reg_15_ ( .D(n2536), .CP(clk), .Q(r3[15]) );
  DFQD1BWP12T r3_reg_14_ ( .D(n2535), .CP(clk), .Q(r3[14]) );
  DFQD1BWP12T r3_reg_13_ ( .D(n2534), .CP(clk), .Q(r3[13]) );
  DFQD1BWP12T r3_reg_12_ ( .D(n2533), .CP(clk), .Q(r3[12]) );
  DFQD1BWP12T r3_reg_11_ ( .D(n2532), .CP(clk), .Q(r3[11]) );
  DFQD1BWP12T r3_reg_10_ ( .D(n2531), .CP(clk), .Q(r3[10]) );
  DFQD1BWP12T r3_reg_9_ ( .D(n2530), .CP(clk), .Q(r3[9]) );
  DFQD1BWP12T r3_reg_8_ ( .D(n2529), .CP(clk), .Q(r3[8]) );
  DFQD1BWP12T r3_reg_7_ ( .D(n2528), .CP(clk), .Q(r3[7]) );
  DFQD1BWP12T r3_reg_6_ ( .D(n2527), .CP(clk), .Q(r3[6]) );
  DFQD1BWP12T r3_reg_5_ ( .D(n2526), .CP(clk), .Q(r3[5]) );
  DFQD1BWP12T r3_reg_4_ ( .D(n2525), .CP(clk), .Q(r3[4]) );
  DFQD1BWP12T r3_reg_3_ ( .D(n2524), .CP(clk), .Q(r3[3]) );
  DFQD1BWP12T r3_reg_1_ ( .D(n2522), .CP(clk), .Q(r3[1]) );
  DFQD1BWP12T r3_reg_0_ ( .D(n2521), .CP(clk), .Q(r3[0]) );
  DFQD1BWP12T r4_reg_31_ ( .D(n2520), .CP(clk), .Q(r4[31]) );
  DFQD1BWP12T r4_reg_28_ ( .D(n2517), .CP(clk), .Q(r4[28]) );
  DFQD1BWP12T r4_reg_26_ ( .D(n2515), .CP(clk), .Q(r4[26]) );
  DFQD1BWP12T r4_reg_25_ ( .D(n2514), .CP(clk), .Q(r4[25]) );
  DFQD1BWP12T r4_reg_24_ ( .D(n2513), .CP(clk), .Q(r4[24]) );
  DFQD1BWP12T r4_reg_23_ ( .D(n2512), .CP(clk), .Q(r4[23]) );
  DFQD1BWP12T r4_reg_22_ ( .D(n2511), .CP(clk), .Q(r4[22]) );
  DFQD1BWP12T r4_reg_21_ ( .D(n2510), .CP(clk), .Q(r4[21]) );
  DFQD1BWP12T r4_reg_20_ ( .D(n2509), .CP(clk), .Q(r4[20]) );
  DFQD1BWP12T r4_reg_19_ ( .D(n2508), .CP(clk), .Q(r4[19]) );
  DFQD1BWP12T r4_reg_18_ ( .D(n2507), .CP(clk), .Q(r4[18]) );
  DFQD1BWP12T r4_reg_16_ ( .D(n2505), .CP(clk), .Q(r4[16]) );
  DFQD1BWP12T r4_reg_15_ ( .D(n2504), .CP(clk), .Q(r4[15]) );
  DFQD1BWP12T r4_reg_14_ ( .D(n2503), .CP(clk), .Q(r4[14]) );
  DFQD1BWP12T r4_reg_13_ ( .D(n2502), .CP(clk), .Q(r4[13]) );
  DFQD1BWP12T r4_reg_12_ ( .D(n2501), .CP(clk), .Q(r4[12]) );
  DFQD1BWP12T r4_reg_11_ ( .D(n2500), .CP(clk), .Q(r4[11]) );
  DFQD1BWP12T r4_reg_10_ ( .D(n2499), .CP(clk), .Q(r4[10]) );
  DFQD1BWP12T r4_reg_8_ ( .D(n2497), .CP(clk), .Q(r4[8]) );
  DFQD1BWP12T r4_reg_7_ ( .D(n2496), .CP(clk), .Q(r4[7]) );
  DFQD1BWP12T r4_reg_6_ ( .D(n2495), .CP(clk), .Q(r4[6]) );
  DFQD1BWP12T r4_reg_5_ ( .D(n2494), .CP(clk), .Q(r4[5]) );
  DFQD1BWP12T r4_reg_4_ ( .D(n2493), .CP(clk), .Q(r4[4]) );
  DFQD1BWP12T r4_reg_3_ ( .D(n2492), .CP(clk), .Q(r4[3]) );
  DFQD1BWP12T r4_reg_2_ ( .D(n2491), .CP(clk), .Q(r4[2]) );
  DFQD1BWP12T r4_reg_1_ ( .D(n2490), .CP(clk), .Q(r4[1]) );
  DFQD1BWP12T r4_reg_0_ ( .D(n2489), .CP(clk), .Q(r4[0]) );
  DFQD1BWP12T r5_reg_31_ ( .D(n2488), .CP(clk), .Q(r5[31]) );
  DFQD1BWP12T r5_reg_29_ ( .D(n2486), .CP(clk), .Q(r5[29]) );
  DFQD1BWP12T r5_reg_28_ ( .D(n2485), .CP(clk), .Q(r5[28]) );
  DFQD1BWP12T r5_reg_27_ ( .D(n2484), .CP(clk), .Q(r5[27]) );
  DFQD1BWP12T r5_reg_26_ ( .D(n2483), .CP(clk), .Q(r5[26]) );
  DFQD1BWP12T r5_reg_25_ ( .D(n2482), .CP(clk), .Q(r5[25]) );
  DFQD1BWP12T r5_reg_24_ ( .D(n2481), .CP(clk), .Q(r5[24]) );
  DFQD1BWP12T r5_reg_23_ ( .D(n2480), .CP(clk), .Q(r5[23]) );
  DFQD1BWP12T r5_reg_22_ ( .D(n2479), .CP(clk), .Q(r5[22]) );
  DFQD1BWP12T r5_reg_21_ ( .D(n2478), .CP(clk), .Q(r5[21]) );
  DFQD1BWP12T r5_reg_20_ ( .D(n2477), .CP(clk), .Q(r5[20]) );
  DFQD1BWP12T r5_reg_19_ ( .D(n2476), .CP(clk), .Q(r5[19]) );
  DFQD1BWP12T r5_reg_18_ ( .D(n2475), .CP(clk), .Q(r5[18]) );
  DFQD1BWP12T r5_reg_17_ ( .D(n2474), .CP(clk), .Q(r5[17]) );
  DFQD1BWP12T r5_reg_16_ ( .D(n2473), .CP(clk), .Q(r5[16]) );
  DFQD1BWP12T r5_reg_15_ ( .D(n2472), .CP(clk), .Q(r5[15]) );
  DFQD1BWP12T r5_reg_14_ ( .D(n2471), .CP(clk), .Q(r5[14]) );
  DFQD1BWP12T r5_reg_13_ ( .D(n2470), .CP(clk), .Q(r5[13]) );
  DFQD1BWP12T r5_reg_12_ ( .D(n2469), .CP(clk), .Q(r5[12]) );
  DFQD1BWP12T r5_reg_11_ ( .D(n2468), .CP(clk), .Q(r5[11]) );
  DFQD1BWP12T r5_reg_10_ ( .D(n2467), .CP(clk), .Q(r5[10]) );
  DFQD1BWP12T r5_reg_9_ ( .D(n2466), .CP(clk), .Q(r5[9]) );
  DFQD1BWP12T r5_reg_8_ ( .D(n2465), .CP(clk), .Q(r5[8]) );
  DFQD1BWP12T r5_reg_7_ ( .D(n2464), .CP(clk), .Q(r5[7]) );
  DFQD1BWP12T r5_reg_6_ ( .D(n2463), .CP(clk), .Q(r5[6]) );
  DFQD1BWP12T r5_reg_5_ ( .D(n2462), .CP(clk), .Q(r5[5]) );
  DFQD1BWP12T r5_reg_4_ ( .D(n2461), .CP(clk), .Q(r5[4]) );
  DFQD1BWP12T r5_reg_3_ ( .D(n2460), .CP(clk), .Q(r5[3]) );
  DFQD1BWP12T r5_reg_2_ ( .D(n2459), .CP(clk), .Q(r5[2]) );
  DFQD1BWP12T r5_reg_1_ ( .D(n2458), .CP(clk), .Q(r5[1]) );
  DFQD1BWP12T r5_reg_0_ ( .D(n2457), .CP(clk), .Q(r5[0]) );
  DFQD1BWP12T r6_reg_31_ ( .D(n2456), .CP(clk), .Q(r6[31]) );
  DFQD1BWP12T r6_reg_29_ ( .D(n2454), .CP(clk), .Q(r6[29]) );
  DFQD1BWP12T r6_reg_28_ ( .D(n2453), .CP(clk), .Q(r6[28]) );
  DFQD1BWP12T r6_reg_27_ ( .D(n2452), .CP(clk), .Q(r6[27]) );
  DFQD1BWP12T r6_reg_25_ ( .D(n2450), .CP(clk), .Q(r6[25]) );
  DFQD1BWP12T r6_reg_24_ ( .D(n2449), .CP(clk), .Q(r6[24]) );
  DFQD1BWP12T r6_reg_23_ ( .D(n2448), .CP(clk), .Q(r6[23]) );
  DFQD1BWP12T r6_reg_22_ ( .D(n2447), .CP(clk), .Q(r6[22]) );
  DFQD1BWP12T r6_reg_21_ ( .D(n2446), .CP(clk), .Q(r6[21]) );
  DFQD1BWP12T r6_reg_20_ ( .D(n2445), .CP(clk), .Q(r6[20]) );
  DFQD1BWP12T r6_reg_19_ ( .D(n2444), .CP(clk), .Q(r6[19]) );
  DFQD1BWP12T r6_reg_18_ ( .D(n2443), .CP(clk), .Q(r6[18]) );
  DFQD1BWP12T r6_reg_17_ ( .D(n2442), .CP(clk), .Q(r6[17]) );
  DFQD1BWP12T r6_reg_16_ ( .D(n2441), .CP(clk), .Q(r6[16]) );
  DFQD1BWP12T r6_reg_15_ ( .D(n2440), .CP(clk), .Q(r6[15]) );
  DFQD1BWP12T r6_reg_14_ ( .D(n2439), .CP(clk), .Q(r6[14]) );
  DFQD1BWP12T r6_reg_13_ ( .D(n2438), .CP(clk), .Q(r6[13]) );
  DFQD1BWP12T r6_reg_12_ ( .D(n2437), .CP(clk), .Q(r6[12]) );
  DFQD1BWP12T r6_reg_11_ ( .D(n2436), .CP(clk), .Q(r6[11]) );
  DFQD1BWP12T r6_reg_10_ ( .D(n2435), .CP(clk), .Q(r6[10]) );
  DFQD1BWP12T r6_reg_9_ ( .D(n2434), .CP(clk), .Q(r6[9]) );
  DFQD1BWP12T r6_reg_8_ ( .D(n2433), .CP(clk), .Q(r6[8]) );
  DFQD1BWP12T r6_reg_7_ ( .D(n2432), .CP(clk), .Q(r6[7]) );
  DFQD1BWP12T r6_reg_6_ ( .D(n2431), .CP(clk), .Q(r6[6]) );
  DFQD1BWP12T r6_reg_5_ ( .D(n2430), .CP(clk), .Q(r6[5]) );
  DFQD1BWP12T r6_reg_4_ ( .D(n2429), .CP(clk), .Q(r6[4]) );
  DFQD1BWP12T r6_reg_3_ ( .D(n2428), .CP(clk), .Q(r6[3]) );
  DFQD1BWP12T r6_reg_2_ ( .D(n2427), .CP(clk), .Q(r6[2]) );
  DFQD1BWP12T r6_reg_1_ ( .D(n2426), .CP(clk), .Q(r6[1]) );
  DFQD1BWP12T r6_reg_0_ ( .D(n2425), .CP(clk), .Q(r6[0]) );
  DFQD1BWP12T r7_reg_31_ ( .D(n2424), .CP(clk), .Q(r7[31]) );
  DFQD1BWP12T r7_reg_29_ ( .D(n2422), .CP(clk), .Q(r7[29]) );
  DFQD1BWP12T r7_reg_28_ ( .D(n2421), .CP(clk), .Q(r7[28]) );
  DFQD1BWP12T r7_reg_27_ ( .D(n2420), .CP(clk), .Q(r7[27]) );
  DFQD1BWP12T r7_reg_26_ ( .D(n2419), .CP(clk), .Q(r7[26]) );
  DFQD1BWP12T r7_reg_25_ ( .D(n2418), .CP(clk), .Q(r7[25]) );
  DFQD1BWP12T r7_reg_24_ ( .D(n2417), .CP(clk), .Q(r7[24]) );
  DFQD1BWP12T r7_reg_23_ ( .D(n2416), .CP(clk), .Q(r7[23]) );
  DFQD1BWP12T r7_reg_22_ ( .D(n2415), .CP(clk), .Q(r7[22]) );
  DFQD1BWP12T r7_reg_21_ ( .D(n2414), .CP(clk), .Q(r7[21]) );
  DFQD1BWP12T r7_reg_20_ ( .D(n2413), .CP(clk), .Q(r7[20]) );
  DFQD1BWP12T r7_reg_19_ ( .D(n2412), .CP(clk), .Q(r7[19]) );
  DFQD1BWP12T r7_reg_18_ ( .D(n2411), .CP(clk), .Q(r7[18]) );
  DFQD1BWP12T r7_reg_17_ ( .D(n2410), .CP(clk), .Q(r7[17]) );
  DFQD1BWP12T r7_reg_16_ ( .D(n2409), .CP(clk), .Q(r7[16]) );
  DFQD1BWP12T r7_reg_14_ ( .D(n2407), .CP(clk), .Q(r7[14]) );
  DFQD1BWP12T r7_reg_13_ ( .D(n2406), .CP(clk), .Q(r7[13]) );
  DFQD1BWP12T r7_reg_12_ ( .D(n2405), .CP(clk), .Q(r7[12]) );
  DFQD1BWP12T r7_reg_11_ ( .D(n2404), .CP(clk), .Q(r7[11]) );
  DFQD1BWP12T r7_reg_10_ ( .D(n2403), .CP(clk), .Q(r7[10]) );
  DFQD1BWP12T r7_reg_8_ ( .D(n2401), .CP(clk), .Q(r7[8]) );
  DFQD1BWP12T r7_reg_7_ ( .D(n2400), .CP(clk), .Q(r7[7]) );
  DFQD1BWP12T r7_reg_6_ ( .D(n2399), .CP(clk), .Q(r7[6]) );
  DFQD1BWP12T r7_reg_5_ ( .D(n2398), .CP(clk), .Q(r7[5]) );
  DFQD1BWP12T r7_reg_4_ ( .D(n2397), .CP(clk), .Q(r7[4]) );
  DFQD1BWP12T r7_reg_3_ ( .D(n2396), .CP(clk), .Q(r7[3]) );
  DFQD1BWP12T r7_reg_2_ ( .D(n2395), .CP(clk), .Q(r7[2]) );
  DFQD1BWP12T r7_reg_1_ ( .D(n2394), .CP(clk), .Q(r7[1]) );
  DFQD1BWP12T r7_reg_0_ ( .D(n2393), .CP(clk), .Q(r7[0]) );
  DFQD1BWP12T r8_reg_31_ ( .D(n2392), .CP(clk), .Q(r8[31]) );
  DFQD1BWP12T r8_reg_28_ ( .D(n2389), .CP(clk), .Q(r8[28]) );
  DFQD1BWP12T r8_reg_26_ ( .D(n2387), .CP(clk), .Q(r8[26]) );
  DFQD1BWP12T r8_reg_24_ ( .D(n2385), .CP(clk), .Q(r8[24]) );
  DFQD1BWP12T r8_reg_23_ ( .D(n2384), .CP(clk), .Q(r8[23]) );
  DFQD1BWP12T r8_reg_22_ ( .D(n2383), .CP(clk), .Q(r8[22]) );
  DFQD1BWP12T r8_reg_21_ ( .D(n2382), .CP(clk), .Q(r8[21]) );
  DFQD1BWP12T r8_reg_20_ ( .D(n2381), .CP(clk), .Q(r8[20]) );
  DFQD1BWP12T r8_reg_19_ ( .D(n2380), .CP(clk), .Q(r8[19]) );
  DFQD1BWP12T r8_reg_18_ ( .D(n2379), .CP(clk), .Q(r8[18]) );
  DFQD1BWP12T r8_reg_17_ ( .D(n2378), .CP(clk), .Q(r8[17]) );
  DFQD1BWP12T r8_reg_16_ ( .D(n2377), .CP(clk), .Q(r8[16]) );
  DFQD1BWP12T r8_reg_15_ ( .D(n2376), .CP(clk), .Q(r8[15]) );
  DFQD1BWP12T r8_reg_14_ ( .D(n2375), .CP(clk), .Q(r8[14]) );
  DFQD1BWP12T r8_reg_13_ ( .D(n2374), .CP(clk), .Q(r8[13]) );
  DFQD1BWP12T r8_reg_12_ ( .D(n2373), .CP(clk), .Q(r8[12]) );
  DFQD1BWP12T r8_reg_10_ ( .D(n2371), .CP(clk), .Q(r8[10]) );
  DFQD1BWP12T r8_reg_9_ ( .D(n2370), .CP(clk), .Q(r8[9]) );
  DFQD1BWP12T r8_reg_8_ ( .D(n2369), .CP(clk), .Q(r8[8]) );
  DFQD1BWP12T r8_reg_7_ ( .D(n2368), .CP(clk), .Q(r8[7]) );
  DFQD1BWP12T r8_reg_6_ ( .D(n2367), .CP(clk), .Q(r8[6]) );
  DFQD1BWP12T r8_reg_5_ ( .D(n2366), .CP(clk), .Q(r8[5]) );
  DFQD1BWP12T r8_reg_4_ ( .D(n2365), .CP(clk), .Q(r8[4]) );
  DFQD1BWP12T r8_reg_3_ ( .D(n2364), .CP(clk), .Q(r8[3]) );
  DFQD1BWP12T r8_reg_2_ ( .D(n2363), .CP(clk), .Q(r8[2]) );
  DFQD1BWP12T r8_reg_1_ ( .D(n2362), .CP(clk), .Q(r8[1]) );
  DFQD1BWP12T r8_reg_0_ ( .D(n2361), .CP(clk), .Q(r8[0]) );
  DFQD1BWP12T r9_reg_31_ ( .D(n2360), .CP(clk), .Q(r9[31]) );
  DFQD1BWP12T r9_reg_29_ ( .D(n2358), .CP(clk), .Q(r9[29]) );
  DFQD1BWP12T r9_reg_28_ ( .D(n2357), .CP(clk), .Q(r9[28]) );
  DFQD1BWP12T r9_reg_27_ ( .D(n2356), .CP(clk), .Q(r9[27]) );
  DFQD1BWP12T r9_reg_26_ ( .D(n2355), .CP(clk), .Q(r9[26]) );
  DFQD1BWP12T r9_reg_25_ ( .D(n2354), .CP(clk), .Q(r9[25]) );
  DFQD1BWP12T r9_reg_24_ ( .D(n2353), .CP(clk), .Q(r9[24]) );
  DFQD1BWP12T r9_reg_23_ ( .D(n2352), .CP(clk), .Q(r9[23]) );
  DFQD1BWP12T r9_reg_22_ ( .D(n2351), .CP(clk), .Q(r9[22]) );
  DFQD1BWP12T r9_reg_21_ ( .D(n2350), .CP(clk), .Q(r9[21]) );
  DFQD1BWP12T r9_reg_20_ ( .D(n2349), .CP(clk), .Q(r9[20]) );
  DFQD1BWP12T r9_reg_19_ ( .D(n2348), .CP(clk), .Q(r9[19]) );
  DFQD1BWP12T r9_reg_18_ ( .D(n2347), .CP(clk), .Q(r9[18]) );
  DFQD1BWP12T r9_reg_17_ ( .D(n2346), .CP(clk), .Q(r9[17]) );
  DFQD1BWP12T r9_reg_16_ ( .D(n2345), .CP(clk), .Q(r9[16]) );
  DFQD1BWP12T r9_reg_14_ ( .D(n2343), .CP(clk), .Q(r9[14]) );
  DFQD1BWP12T r9_reg_13_ ( .D(n2342), .CP(clk), .Q(r9[13]) );
  DFQD1BWP12T r9_reg_12_ ( .D(n2341), .CP(clk), .Q(r9[12]) );
  DFQD1BWP12T r9_reg_11_ ( .D(n2340), .CP(clk), .Q(r9[11]) );
  DFQD1BWP12T r9_reg_10_ ( .D(n2339), .CP(clk), .Q(r9[10]) );
  DFQD1BWP12T r9_reg_8_ ( .D(n2337), .CP(clk), .Q(r9[8]) );
  DFQD1BWP12T r9_reg_7_ ( .D(n2336), .CP(clk), .Q(r9[7]) );
  DFQD1BWP12T r9_reg_6_ ( .D(n2335), .CP(clk), .Q(r9[6]) );
  DFQD1BWP12T r9_reg_5_ ( .D(n2334), .CP(clk), .Q(r9[5]) );
  DFQD1BWP12T r9_reg_4_ ( .D(n2333), .CP(clk), .Q(r9[4]) );
  DFQD1BWP12T r9_reg_3_ ( .D(n2332), .CP(clk), .Q(r9[3]) );
  DFQD1BWP12T r9_reg_2_ ( .D(n2331), .CP(clk), .Q(r9[2]) );
  DFQD1BWP12T r9_reg_1_ ( .D(n2330), .CP(clk), .Q(r9[1]) );
  DFQD1BWP12T r9_reg_0_ ( .D(n2329), .CP(clk), .Q(r9[0]) );
  DFQD1BWP12T r10_reg_31_ ( .D(n2328), .CP(clk), .Q(r10[31]) );
  DFQD1BWP12T r10_reg_28_ ( .D(n2325), .CP(clk), .Q(r10[28]) );
  DFQD1BWP12T r10_reg_27_ ( .D(n2324), .CP(clk), .Q(r10[27]) );
  DFQD1BWP12T r10_reg_26_ ( .D(n2323), .CP(clk), .Q(r10[26]) );
  DFQD1BWP12T r10_reg_25_ ( .D(n2322), .CP(clk), .Q(r10[25]) );
  DFQD1BWP12T r10_reg_24_ ( .D(n2321), .CP(clk), .Q(r10[24]) );
  DFQD1BWP12T r10_reg_23_ ( .D(n2320), .CP(clk), .Q(r10[23]) );
  DFQD1BWP12T r10_reg_22_ ( .D(n2319), .CP(clk), .Q(r10[22]) );
  DFQD1BWP12T r10_reg_21_ ( .D(n2318), .CP(clk), .Q(r10[21]) );
  DFQD1BWP12T r10_reg_20_ ( .D(n2317), .CP(clk), .Q(r10[20]) );
  DFQD1BWP12T r10_reg_19_ ( .D(n2316), .CP(clk), .Q(r10[19]) );
  DFQD1BWP12T r10_reg_18_ ( .D(n2315), .CP(clk), .Q(r10[18]) );
  DFQD1BWP12T r10_reg_17_ ( .D(n2314), .CP(clk), .Q(r10[17]) );
  DFQD1BWP12T r10_reg_16_ ( .D(n2313), .CP(clk), .Q(r10[16]) );
  DFQD1BWP12T r10_reg_15_ ( .D(n2312), .CP(clk), .Q(r10[15]) );
  DFQD1BWP12T r10_reg_14_ ( .D(n2311), .CP(clk), .Q(r10[14]) );
  DFQD1BWP12T r10_reg_13_ ( .D(n2310), .CP(clk), .Q(r10[13]) );
  DFQD1BWP12T r10_reg_12_ ( .D(n2309), .CP(clk), .Q(r10[12]) );
  DFQD1BWP12T r10_reg_11_ ( .D(n2308), .CP(clk), .Q(r10[11]) );
  DFQD1BWP12T r10_reg_10_ ( .D(n2307), .CP(clk), .Q(r10[10]) );
  DFQD1BWP12T r10_reg_9_ ( .D(n2306), .CP(clk), .Q(r10[9]) );
  DFQD1BWP12T r10_reg_8_ ( .D(n2305), .CP(clk), .Q(r10[8]) );
  DFQD1BWP12T r10_reg_7_ ( .D(n2304), .CP(clk), .Q(r10[7]) );
  DFQD1BWP12T r10_reg_6_ ( .D(n2303), .CP(clk), .Q(r10[6]) );
  DFQD1BWP12T r10_reg_5_ ( .D(n2302), .CP(clk), .Q(r10[5]) );
  DFQD1BWP12T r10_reg_4_ ( .D(n2301), .CP(clk), .Q(r10[4]) );
  DFQD1BWP12T r10_reg_3_ ( .D(n2300), .CP(clk), .Q(r10[3]) );
  DFQD1BWP12T r10_reg_2_ ( .D(n2299), .CP(clk), .Q(r10[2]) );
  DFQD1BWP12T r10_reg_0_ ( .D(n2297), .CP(clk), .Q(r10[0]) );
  DFQD1BWP12T r11_reg_31_ ( .D(n2296), .CP(clk), .Q(r11[31]) );
  DFQD1BWP12T r11_reg_28_ ( .D(n2293), .CP(clk), .Q(r11[28]) );
  DFQD1BWP12T r11_reg_27_ ( .D(n2292), .CP(clk), .Q(r11[27]) );
  DFQD1BWP12T r11_reg_26_ ( .D(n2291), .CP(clk), .Q(r11[26]) );
  DFQD1BWP12T r11_reg_25_ ( .D(n2290), .CP(clk), .Q(r11[25]) );
  DFQD1BWP12T r11_reg_24_ ( .D(n2289), .CP(clk), .Q(r11[24]) );
  DFQD1BWP12T r11_reg_23_ ( .D(n2288), .CP(clk), .Q(r11[23]) );
  DFQD1BWP12T r11_reg_22_ ( .D(n2287), .CP(clk), .Q(r11[22]) );
  DFQD1BWP12T r11_reg_21_ ( .D(n2286), .CP(clk), .Q(r11[21]) );
  DFQD1BWP12T r11_reg_20_ ( .D(n2285), .CP(clk), .Q(r11[20]) );
  DFQD1BWP12T r11_reg_19_ ( .D(n2284), .CP(clk), .Q(r11[19]) );
  DFQD1BWP12T r11_reg_18_ ( .D(n2283), .CP(clk), .Q(r11[18]) );
  DFQD1BWP12T r11_reg_17_ ( .D(n2282), .CP(clk), .Q(r11[17]) );
  DFQD1BWP12T r11_reg_16_ ( .D(n2281), .CP(clk), .Q(r11[16]) );
  DFQD1BWP12T r11_reg_15_ ( .D(n2280), .CP(clk), .Q(r11[15]) );
  DFQD1BWP12T r11_reg_14_ ( .D(n2279), .CP(clk), .Q(r11[14]) );
  DFQD1BWP12T r11_reg_13_ ( .D(n2278), .CP(clk), .Q(r11[13]) );
  DFQD1BWP12T r11_reg_11_ ( .D(n2276), .CP(clk), .Q(r11[11]) );
  DFQD1BWP12T r11_reg_10_ ( .D(n2275), .CP(clk), .Q(r11[10]) );
  DFQD1BWP12T r11_reg_9_ ( .D(n2274), .CP(clk), .Q(r11[9]) );
  DFQD1BWP12T r11_reg_8_ ( .D(n2273), .CP(clk), .Q(r11[8]) );
  DFQD1BWP12T r11_reg_7_ ( .D(n2272), .CP(clk), .Q(r11[7]) );
  DFQD1BWP12T r11_reg_6_ ( .D(n2271), .CP(clk), .Q(r11[6]) );
  DFQD1BWP12T r11_reg_5_ ( .D(n2270), .CP(clk), .Q(r11[5]) );
  DFQD1BWP12T r11_reg_4_ ( .D(n2269), .CP(clk), .Q(r11[4]) );
  DFQD1BWP12T r11_reg_3_ ( .D(n2268), .CP(clk), .Q(r11[3]) );
  DFQD1BWP12T r11_reg_2_ ( .D(n2267), .CP(clk), .Q(r11[2]) );
  DFQD1BWP12T r11_reg_0_ ( .D(n2265), .CP(clk), .Q(r11[0]) );
  DFQD1BWP12T r12_reg_31_ ( .D(n2264), .CP(clk), .Q(r12[31]) );
  DFQD1BWP12T r12_reg_29_ ( .D(n2262), .CP(clk), .Q(r12[29]) );
  DFQD1BWP12T r12_reg_28_ ( .D(n2261), .CP(clk), .Q(r12[28]) );
  DFQD1BWP12T r12_reg_27_ ( .D(n2260), .CP(clk), .Q(r12[27]) );
  DFQD1BWP12T r12_reg_26_ ( .D(n2259), .CP(clk), .Q(r12[26]) );
  DFQD1BWP12T r12_reg_25_ ( .D(n2258), .CP(clk), .Q(r12[25]) );
  DFQD1BWP12T r12_reg_24_ ( .D(n2257), .CP(clk), .Q(r12[24]) );
  DFQD1BWP12T r12_reg_23_ ( .D(n2256), .CP(clk), .Q(r12[23]) );
  DFQD1BWP12T r12_reg_22_ ( .D(n2255), .CP(clk), .Q(r12[22]) );
  DFQD1BWP12T r12_reg_21_ ( .D(n2254), .CP(clk), .Q(r12[21]) );
  DFQD1BWP12T r12_reg_20_ ( .D(n2253), .CP(clk), .Q(r12[20]) );
  DFQD1BWP12T r12_reg_19_ ( .D(n2252), .CP(clk), .Q(r12[19]) );
  DFQD1BWP12T r12_reg_18_ ( .D(n2251), .CP(clk), .Q(r12[18]) );
  DFQD1BWP12T r12_reg_17_ ( .D(n2250), .CP(clk), .Q(r12[17]) );
  DFQD1BWP12T r12_reg_16_ ( .D(n2249), .CP(clk), .Q(r12[16]) );
  DFQD1BWP12T r12_reg_15_ ( .D(n2248), .CP(clk), .Q(r12[15]) );
  DFQD1BWP12T r12_reg_14_ ( .D(n2247), .CP(clk), .Q(r12[14]) );
  DFQD1BWP12T r12_reg_13_ ( .D(n2246), .CP(clk), .Q(r12[13]) );
  DFQD1BWP12T r12_reg_12_ ( .D(n2245), .CP(clk), .Q(r12[12]) );
  DFQD1BWP12T r12_reg_11_ ( .D(n2244), .CP(clk), .Q(r12[11]) );
  DFQD1BWP12T r12_reg_10_ ( .D(n2243), .CP(clk), .Q(r12[10]) );
  DFQD1BWP12T r12_reg_9_ ( .D(n2242), .CP(clk), .Q(r12[9]) );
  DFQD1BWP12T r12_reg_8_ ( .D(n2241), .CP(clk), .Q(r12[8]) );
  DFQD1BWP12T r12_reg_7_ ( .D(n2240), .CP(clk), .Q(r12[7]) );
  DFQD1BWP12T r12_reg_6_ ( .D(n2239), .CP(clk), .Q(r12[6]) );
  DFQD1BWP12T r12_reg_5_ ( .D(n2238), .CP(clk), .Q(r12[5]) );
  DFQD1BWP12T r12_reg_4_ ( .D(n2237), .CP(clk), .Q(r12[4]) );
  DFQD1BWP12T r12_reg_3_ ( .D(n2236), .CP(clk), .Q(r12[3]) );
  DFQD1BWP12T r12_reg_2_ ( .D(n2235), .CP(clk), .Q(r12[2]) );
  DFQD1BWP12T r12_reg_0_ ( .D(n2233), .CP(clk), .Q(r12[0]) );
  DFQD1BWP12T lr_reg_31_ ( .D(n2232), .CP(clk), .Q(lr[31]) );
  DFQD1BWP12T lr_reg_29_ ( .D(n2230), .CP(clk), .Q(lr[29]) );
  DFQD1BWP12T lr_reg_28_ ( .D(n2229), .CP(clk), .Q(lr[28]) );
  DFQD1BWP12T lr_reg_27_ ( .D(n2228), .CP(clk), .Q(lr[27]) );
  DFQD1BWP12T lr_reg_26_ ( .D(n2227), .CP(clk), .Q(lr[26]) );
  DFQD1BWP12T lr_reg_25_ ( .D(n2226), .CP(clk), .Q(lr[25]) );
  DFQD1BWP12T lr_reg_24_ ( .D(n2225), .CP(clk), .Q(lr[24]) );
  DFQD1BWP12T lr_reg_23_ ( .D(n2224), .CP(clk), .Q(lr[23]) );
  DFQD1BWP12T lr_reg_22_ ( .D(n2223), .CP(clk), .Q(lr[22]) );
  DFQD1BWP12T lr_reg_21_ ( .D(n2222), .CP(clk), .Q(lr[21]) );
  DFQD1BWP12T lr_reg_20_ ( .D(n2221), .CP(clk), .Q(lr[20]) );
  DFQD1BWP12T lr_reg_19_ ( .D(n2220), .CP(clk), .Q(lr[19]) );
  DFQD1BWP12T lr_reg_18_ ( .D(n2219), .CP(clk), .Q(lr[18]) );
  DFQD1BWP12T lr_reg_17_ ( .D(n2218), .CP(clk), .Q(lr[17]) );
  DFQD1BWP12T lr_reg_16_ ( .D(n2217), .CP(clk), .Q(lr[16]) );
  DFQD1BWP12T lr_reg_15_ ( .D(n2216), .CP(clk), .Q(lr[15]) );
  DFQD1BWP12T lr_reg_14_ ( .D(n2215), .CP(clk), .Q(lr[14]) );
  DFQD1BWP12T lr_reg_13_ ( .D(n2214), .CP(clk), .Q(lr[13]) );
  DFQD1BWP12T lr_reg_12_ ( .D(n2213), .CP(clk), .Q(lr[12]) );
  DFQD1BWP12T lr_reg_11_ ( .D(n2212), .CP(clk), .Q(lr[11]) );
  DFQD1BWP12T lr_reg_10_ ( .D(n2211), .CP(clk), .Q(lr[10]) );
  DFQD1BWP12T lr_reg_9_ ( .D(n2210), .CP(clk), .Q(lr[9]) );
  DFQD1BWP12T lr_reg_8_ ( .D(n2209), .CP(clk), .Q(lr[8]) );
  DFQD1BWP12T lr_reg_7_ ( .D(n2208), .CP(clk), .Q(lr[7]) );
  DFQD1BWP12T lr_reg_6_ ( .D(n2207), .CP(clk), .Q(lr[6]) );
  DFQD1BWP12T lr_reg_5_ ( .D(n2206), .CP(clk), .Q(lr[5]) );
  DFQD1BWP12T lr_reg_4_ ( .D(n2205), .CP(clk), .Q(lr[4]) );
  DFQD1BWP12T lr_reg_3_ ( .D(n2204), .CP(clk), .Q(lr[3]) );
  DFQD1BWP12T lr_reg_2_ ( .D(n2203), .CP(clk), .Q(lr[2]) );
  DFQD1BWP12T lr_reg_1_ ( .D(n2202), .CP(clk), .Q(lr[1]) );
  DFQD1BWP12T lr_reg_0_ ( .D(n2201), .CP(clk), .Q(lr[0]) );
  DFQD1BWP12T sp_reg_31_ ( .D(spin[31]), .CP(clk), .Q(n[3669]) );
  DFQD1BWP12T sp_reg_29_ ( .D(spin[29]), .CP(clk), .Q(n[3671]) );
  DFQD1BWP12T sp_reg_28_ ( .D(spin[28]), .CP(clk), .Q(n[3672]) );
  DFQD1BWP12T sp_reg_27_ ( .D(spin[27]), .CP(clk), .Q(n[3673]) );
  DFQD1BWP12T sp_reg_26_ ( .D(spin[26]), .CP(clk), .Q(n[3674]) );
  DFQD1BWP12T sp_reg_25_ ( .D(spin[25]), .CP(clk), .Q(n[3675]) );
  DFQD1BWP12T sp_reg_24_ ( .D(spin[24]), .CP(clk), .Q(n[3676]) );
  DFQD1BWP12T sp_reg_23_ ( .D(spin[23]), .CP(clk), .Q(n[3677]) );
  DFQD1BWP12T sp_reg_22_ ( .D(spin[22]), .CP(clk), .Q(n[3678]) );
  DFQD1BWP12T sp_reg_21_ ( .D(spin[21]), .CP(clk), .Q(n[3679]) );
  DFQD1BWP12T sp_reg_20_ ( .D(spin[20]), .CP(clk), .Q(n[3680]) );
  DFQD1BWP12T sp_reg_19_ ( .D(spin[19]), .CP(clk), .Q(n[3681]) );
  DFQD1BWP12T sp_reg_18_ ( .D(spin[18]), .CP(clk), .Q(n[3682]) );
  DFQD1BWP12T sp_reg_17_ ( .D(spin[17]), .CP(clk), .Q(n[3683]) );
  DFQD1BWP12T sp_reg_16_ ( .D(spin[16]), .CP(clk), .Q(n[3684]) );
  DFQD1BWP12T sp_reg_15_ ( .D(spin[15]), .CP(clk), .Q(n[3685]) );
  DFQD1BWP12T sp_reg_14_ ( .D(spin[14]), .CP(clk), .Q(n[3686]) );
  DFQD1BWP12T sp_reg_13_ ( .D(spin[13]), .CP(clk), .Q(n[3687]) );
  DFQD1BWP12T sp_reg_12_ ( .D(spin[12]), .CP(clk), .Q(n[3688]) );
  DFQD1BWP12T sp_reg_11_ ( .D(spin[11]), .CP(clk), .Q(n[3689]) );
  DFQD1BWP12T sp_reg_10_ ( .D(spin[10]), .CP(clk), .Q(n[3690]) );
  DFQD1BWP12T sp_reg_8_ ( .D(spin[8]), .CP(clk), .Q(n[3692]) );
  DFQD1BWP12T sp_reg_7_ ( .D(spin[7]), .CP(clk), .Q(n[3693]) );
  DFQD1BWP12T sp_reg_6_ ( .D(spin[6]), .CP(clk), .Q(n[3694]) );
  DFQD1BWP12T sp_reg_5_ ( .D(spin[5]), .CP(clk), .Q(n[3695]) );
  DFQD1BWP12T sp_reg_4_ ( .D(spin[4]), .CP(clk), .Q(n[3696]) );
  DFQD1BWP12T sp_reg_3_ ( .D(spin[3]), .CP(clk), .Q(n[3697]) );
  DFQD1BWP12T sp_reg_2_ ( .D(spin[2]), .CP(clk), .Q(n[3698]) );
  DFQD1BWP12T sp_reg_1_ ( .D(spin[1]), .CP(clk), .Q(n[3699]) );
  DFQD1BWP12T sp_reg_0_ ( .D(spin[0]), .CP(clk), .Q(n[3700]) );
  DFQD1BWP12T pc_reg_21_ ( .D(n2190), .CP(clk), .Q(pc_out[21]) );
  DFQD1BWP12T pc_reg_18_ ( .D(n2187), .CP(clk), .Q(pc_out[18]) );
  DFQD1BWP12T pc_reg_17_ ( .D(n2186), .CP(clk), .Q(pc_out[17]) );
  DFQD1BWP12T pc_reg_16_ ( .D(n2185), .CP(clk), .Q(pc_out[16]) );
  DFQD1BWP12T pc_reg_14_ ( .D(n2183), .CP(clk), .Q(pc_out[14]) );
  DFQD1BWP12T pc_reg_13_ ( .D(n2182), .CP(clk), .Q(pc_out[13]) );
  DFQD1BWP12T pc_reg_12_ ( .D(n2181), .CP(clk), .Q(pc_out[12]) );
  DFQD1BWP12T pc_reg_10_ ( .D(n2179), .CP(clk), .Q(pc_out[10]) );
  DFQD1BWP12T pc_reg_8_ ( .D(n2177), .CP(clk), .Q(pc_out[8]) );
  DFQD1BWP12T pc_reg_6_ ( .D(n2175), .CP(clk), .Q(pc_out[6]) );
  DFQD1BWP12T pc_reg_4_ ( .D(n2173), .CP(clk), .Q(pc_out[4]) );
  DFQD1BWP12T pc_reg_3_ ( .D(n2172), .CP(clk), .Q(pc_out[3]) );
  DFQD1BWP12T pc_reg_2_ ( .D(n2171), .CP(clk), .Q(pc_out[2]) );
  DFQD1BWP12T pc_reg_1_ ( .D(n2170), .CP(clk), .Q(pc_out[1]) );
  DFQD1BWP12T pc_reg_0_ ( .D(n2169), .CP(clk), .Q(pc_out[0]) );
  DFQD1BWP12T cpsr_reg_3_ ( .D(cpsrin[3]), .CP(clk), .Q(cpsr_out[3]) );
  DFQD1BWP12T cpsr_reg_2_ ( .D(cpsrin[2]), .CP(clk), .Q(cpsr_out[2]) );
  DFQD1BWP12T tmp1_reg_31_ ( .D(n2168), .CP(clk), .Q(tmp1[31]) );
  DFQD1BWP12T tmp1_reg_29_ ( .D(n2166), .CP(clk), .Q(tmp1[29]) );
  DFQD1BWP12T tmp1_reg_28_ ( .D(n2165), .CP(clk), .Q(tmp1[28]) );
  DFQD1BWP12T tmp1_reg_27_ ( .D(n2164), .CP(clk), .Q(tmp1[27]) );
  DFQD1BWP12T tmp1_reg_26_ ( .D(n2163), .CP(clk), .Q(tmp1[26]) );
  DFQD1BWP12T tmp1_reg_25_ ( .D(n2162), .CP(clk), .Q(tmp1[25]) );
  DFQD1BWP12T tmp1_reg_24_ ( .D(n2161), .CP(clk), .Q(tmp1[24]) );
  DFQD1BWP12T tmp1_reg_23_ ( .D(n2160), .CP(clk), .Q(tmp1[23]) );
  DFQD1BWP12T tmp1_reg_22_ ( .D(n2159), .CP(clk), .Q(tmp1[22]) );
  DFQD1BWP12T tmp1_reg_21_ ( .D(n2158), .CP(clk), .Q(tmp1[21]) );
  DFQD1BWP12T tmp1_reg_20_ ( .D(n2157), .CP(clk), .Q(tmp1[20]) );
  DFQD1BWP12T tmp1_reg_19_ ( .D(n2156), .CP(clk), .Q(tmp1[19]) );
  DFQD1BWP12T tmp1_reg_18_ ( .D(n2155), .CP(clk), .Q(tmp1[18]) );
  DFQD1BWP12T tmp1_reg_17_ ( .D(n2154), .CP(clk), .Q(tmp1[17]) );
  DFQD1BWP12T tmp1_reg_16_ ( .D(n2153), .CP(clk), .Q(tmp1[16]) );
  DFQD1BWP12T tmp1_reg_15_ ( .D(n2152), .CP(clk), .Q(tmp1[15]) );
  DFQD1BWP12T tmp1_reg_14_ ( .D(n2151), .CP(clk), .Q(tmp1[14]) );
  DFQD1BWP12T tmp1_reg_13_ ( .D(n2150), .CP(clk), .Q(tmp1[13]) );
  DFQD1BWP12T tmp1_reg_12_ ( .D(n2149), .CP(clk), .Q(tmp1[12]) );
  DFQD1BWP12T tmp1_reg_11_ ( .D(n2148), .CP(clk), .Q(tmp1[11]) );
  DFQD1BWP12T tmp1_reg_10_ ( .D(n2147), .CP(clk), .Q(tmp1[10]) );
  DFQD1BWP12T tmp1_reg_9_ ( .D(n2146), .CP(clk), .Q(tmp1[9]) );
  DFQD1BWP12T tmp1_reg_8_ ( .D(n2145), .CP(clk), .Q(tmp1[8]) );
  DFQD1BWP12T tmp1_reg_7_ ( .D(n2144), .CP(clk), .Q(tmp1[7]) );
  DFQD1BWP12T tmp1_reg_6_ ( .D(n2143), .CP(clk), .Q(tmp1[6]) );
  DFQD1BWP12T tmp1_reg_5_ ( .D(n2142), .CP(clk), .Q(tmp1[5]) );
  DFQD1BWP12T tmp1_reg_4_ ( .D(n2141), .CP(clk), .Q(tmp1[4]) );
  DFQD1BWP12T tmp1_reg_3_ ( .D(n2140), .CP(clk), .Q(tmp1[3]) );
  DFQD1BWP12T tmp1_reg_2_ ( .D(n2139), .CP(clk), .Q(tmp1[2]) );
  DFQD1BWP12T tmp1_reg_1_ ( .D(n2138), .CP(clk), .Q(tmp1[1]) );
  DFQD1BWP12T tmp1_reg_0_ ( .D(n2136), .CP(clk), .Q(tmp1[0]) );
  DFQD4BWP12T pc_reg_7_ ( .D(n2176), .CP(clk), .Q(pc_out[7]) );
  DFQD4BWP12T pc_reg_9_ ( .D(n2178), .CP(clk), .Q(pc_out[9]) );
  DFQD4BWP12T r11_reg_12_ ( .D(n2277), .CP(clk), .Q(r11[12]) );
  DFQD4BWP12T r9_reg_15_ ( .D(n2344), .CP(clk), .Q(r9[15]) );
  DFQD4BWP12T r8_reg_11_ ( .D(n2372), .CP(clk), .Q(r8[11]) );
  DFQD1BWP12T pc_reg_23_ ( .D(n2192), .CP(clk), .Q(pc_out[23]) );
  DFQD2BWP12T r11_reg_1_ ( .D(n2266), .CP(clk), .Q(r11[1]) );
  DFKCNXD1BWP12T cpsr_reg_0_ ( .CN(n3621), .D(next_cpsr_in[0]), .CP(clk), .Q(
        cpsr_out[0]) );
  DFKCSND1BWP12T r10_reg_30_ ( .D(n3619), .SN(n3627), .CN(n3637), .CP(clk), 
        .Q(n3657), .QN(r10[30]) );
  DFKCSND1BWP12T r3_reg_30_ ( .D(n3619), .SN(n3624), .CN(n3634), .CP(clk), .Q(
        n3661), .QN(r3[30]) );
  DFKCSND1BWP12T r2_reg_30_ ( .D(n3619), .SN(n3625), .CN(n3636), .CP(clk), 
        .QN(r2[30]) );
  DFXD1BWP12T pc_reg_24_ ( .D(n2193), .CP(clk), .Q(pc_out[24]), .QN(n3644) );
  DFXD1BWP12T pc_reg_19_ ( .D(n2188), .CP(clk), .Q(pc_out[19]), .QN(n3641) );
  DFKCNXD1BWP12T cpsr_reg_1_ ( .CN(n3621), .D(next_cpsr_in[1]), .CP(clk), .Q(
        cpsr_out[1]) );
  DFXD1BWP12T pc_reg_31_ ( .D(n2200), .CP(clk), .Q(pc_out[31]), .QN(n3667) );
  DFXD1BWP12T pc_reg_27_ ( .D(n2196), .CP(clk), .Q(pc_out[27]), .QN(n3647) );
  DFXD1BWP12T pc_reg_26_ ( .D(n2195), .CP(clk), .Q(pc_out[26]), .QN(n3646) );
  DFXD1BWP12T pc_reg_30_ ( .D(n2199), .CP(clk), .Q(pc_out[30]), .QN(n3659) );
  DFXD1BWP12T pc_reg_20_ ( .D(n2189), .CP(clk), .Q(pc_out[20]), .QN(n3642) );
  DFXD1BWP12T pc_reg_29_ ( .D(n2198), .CP(clk), .Q(pc_out[29]), .QN(n3650) );
  DFXD1BWP12T pc_reg_22_ ( .D(n2191), .CP(clk), .Q(pc_out[22]), .QN(n3643) );
  DFXD1BWP12T pc_reg_28_ ( .D(n2197), .CP(clk), .Q(pc_out[28]), .QN(n3648) );
  DFKCSND1BWP12T r6_reg_30_ ( .D(n3619), .SN(n3628), .CN(n3632), .CP(clk), .Q(
        n3658), .QN(r6[30]) );
  DFXD1BWP12T pc_reg_25_ ( .D(n2194), .CP(clk), .Q(pc_out[25]), .QN(n3645) );
  DFKCSND1BWP12T r5_reg_30_ ( .D(n3619), .SN(n3622), .CN(n3633), .CP(clk), .Q(
        n3662), .QN(r5[30]) );
  DFKCSND1BWP12T r4_reg_30_ ( .D(n3619), .SN(n3623), .CN(n3635), .CP(clk), .Q(
        n3654), .QN(r4[30]) );
  DFXD1BWP12T r1_reg_30_ ( .D(n2615), .CP(clk), .Q(r1[30]), .QN(n3666) );
  DFXD1BWP12T r0_reg_30_ ( .D(n2647), .CP(clk), .Q(r0[30]), .QN(n3653) );
  DFXD1BWP12T r7_reg_30_ ( .D(n2423), .CP(clk), .Q(r7[30]), .QN(n3660) );
  DFXD1BWP12T sp_reg_30_ ( .D(spin[30]), .CP(clk), .Q(n[3670]), .QN(n3664) );
  DFXD1BWP12T r9_reg_30_ ( .D(n2359), .CP(clk), .Q(r9[30]), .QN(n3640) );
  DFXD1BWP12T r11_reg_30_ ( .D(n2295), .CP(clk), .Q(r11[30]), .QN(n3663) );
  DFXD1BWP12T lr_reg_30_ ( .D(n2231), .CP(clk), .Q(lr[30]), .QN(n3656) );
  DFXD1BWP12T r12_reg_30_ ( .D(n2263), .CP(clk), .Q(r12[30]), .QN(n3665) );
  DFXD1BWP12T r8_reg_30_ ( .D(n2391), .CP(clk), .Q(r8[30]), .QN(n3655) );
  DFKCSND1BWP12T r10_reg_29_ ( .D(n3620), .SN(n3627), .CN(n3631), .CP(clk), 
        .Q(n3649), .QN(r10[29]) );
  DFKCSND1BWP12T r3_reg_29_ ( .D(n3620), .SN(n3624), .CN(n3629), .CP(clk), .Q(
        n3651), .QN(r3[29]) );
  DFQD4BWP12T r10_reg_1_ ( .D(n2298), .CP(clk), .Q(r10[1]) );
  DFKCSND1BWP12T r11_reg_29_ ( .D(n241), .SN(n3626), .CN(n3630), .CP(clk), .Q(
        n3652), .QN(r11[29]) );
  DFKCSND1BWP12T tmp1_reg_30_ ( .D(n3619), .SN(n3638), .CN(n3639), .CP(clk), 
        .QN(tmp1[30]) );
  DFQD4BWP12T r1_reg_12_ ( .D(n2597), .CP(clk), .Q(r1[12]) );
  DFQD4BWP12T r12_reg_1_ ( .D(n2234), .CP(clk), .Q(r12[1]) );
  DFQD4BWP12T r2_reg_12_ ( .D(n2565), .CP(clk), .Q(r2[12]) );
  DFQD4BWP12T r1_reg_3_ ( .D(n2588), .CP(clk), .Q(r1[3]) );
  DFQD4BWP12T r4_reg_17_ ( .D(n2506), .CP(clk), .Q(r4[17]) );
  DFQD4BWP12T r3_reg_2_ ( .D(n2523), .CP(clk), .Q(r3[2]) );
  DFQD4BWP12T r9_reg_9_ ( .D(n2338), .CP(clk), .Q(r9[9]) );
  DFQD4BWP12T pc_reg_11_ ( .D(n2180), .CP(clk), .Q(pc_out[11]) );
  DFQD4BWP12T pc_reg_5_ ( .D(n2174), .CP(clk), .Q(pc_out[5]) );
  DFQD4BWP12T sp_reg_9_ ( .D(spin[9]), .CP(clk), .Q(n[3691]) );
  DFQD4BWP12T r4_reg_9_ ( .D(n2498), .CP(clk), .Q(r4[9]) );
  DFQD4BWP12T r7_reg_9_ ( .D(n2402), .CP(clk), .Q(r7[9]) );
  DFQD4BWP12T r7_reg_15_ ( .D(n2408), .CP(clk), .Q(r7[15]) );
  DFQD4BWP12T r1_reg_25_ ( .D(n2610), .CP(clk), .Q(r1[25]) );
  DFQD4BWP12T r8_reg_27_ ( .D(n2388), .CP(clk), .Q(r8[27]) );
  DFQD4BWP12T r8_reg_25_ ( .D(n2386), .CP(clk), .Q(r8[25]) );
  DFQD4BWP12T r4_reg_27_ ( .D(n2516), .CP(clk), .Q(r4[27]) );
  DFQD1BWP12T r6_reg_26_ ( .D(n2451), .CP(clk), .Q(r6[26]) );
  DFQD2BWP12T pc_reg_15_ ( .D(n2184), .CP(clk), .Q(pc_out[15]) );
  DFQD2BWP12T r0_reg_29_ ( .D(n2646), .CP(clk), .Q(r0[29]) );
  DFQD2BWP12T r1_reg_29_ ( .D(n2614), .CP(clk), .Q(r1[29]) );
  DFQD2BWP12T r4_reg_29_ ( .D(n2518), .CP(clk), .Q(r4[29]) );
  DFQD2BWP12T r8_reg_29_ ( .D(n2390), .CP(clk), .Q(r8[29]) );
  CKND2BWP12T U3 ( .I(lr[5]), .ZN(n2327) );
  CKND2BWP12T U4 ( .I(n[3695]), .ZN(n1418) );
  INVD16BWP12T U5 ( .I(n338), .ZN(n3472) );
  IOA22D4BWP12T U6 ( .B1(n3648), .B2(n3399), .A1(next_pc_in[28]), .A2(n3398), 
        .ZN(n441) );
  TPOAI21D1BWP12T U7 ( .A1(n3488), .A2(n1739), .B(n1262), .ZN(n1266) );
  TPND2D1BWP12T U8 ( .A1(n1950), .A2(r7[12]), .ZN(n1954) );
  TPND2D1BWP12T U9 ( .A1(n1950), .A2(r7[1]), .ZN(n1263) );
  TPND2D1BWP12T U10 ( .A1(n1264), .A2(n1263), .ZN(n1265) );
  OR2D4BWP12T U11 ( .A1(n1666), .A2(n1249), .Z(n1252) );
  INVD2BWP12T U12 ( .I(n236), .ZN(n237) );
  ND2XD4BWP12T U13 ( .A1(n434), .A2(n845), .ZN(n435) );
  BUFFXD8BWP12T U14 ( .I(n349), .Z(n3422) );
  INVD2BWP12T U15 ( .I(n[3678]), .ZN(n2715) );
  TPNR2D2BWP12T U16 ( .A1(n2), .A2(n1), .ZN(n1445) );
  IND2D2BWP12T U17 ( .A1(n1431), .B1(n1433), .ZN(n1) );
  TPND3D2BWP12T U18 ( .A1(n1432), .A2(n3), .A3(n1434), .ZN(n2) );
  CKND3BWP12T U19 ( .I(n1430), .ZN(n3) );
  TPOAI22D2BWP12T U20 ( .A1(n3489), .A2(n1713), .B1(n3488), .B2(n1712), .ZN(
        n1720) );
  TPND2D2BWP12T U21 ( .A1(n1633), .A2(r8[1]), .ZN(n1246) );
  CKND2D2BWP12T U22 ( .A1(n1247), .A2(n1246), .ZN(n236) );
  TPOAI22D2BWP12T U23 ( .A1(n3489), .A2(n1095), .B1(n1806), .B2(n3488), .ZN(
        n1096) );
  INVD9BWP12T U24 ( .I(n1952), .ZN(n3492) );
  INVD8BWP12T U25 ( .I(n1952), .ZN(n3437) );
  TPND2D2BWP12T U26 ( .A1(n1924), .A2(r8[10]), .ZN(n334) );
  ND4D2BWP12T U27 ( .A1(n1607), .A2(n1606), .A3(n5), .A4(n4), .ZN(regB_out[12]) );
  TPNR2D1BWP12T U28 ( .A1(n1597), .A2(n1595), .ZN(n4) );
  TPNR2D2BWP12T U29 ( .A1(n1594), .A2(n1596), .ZN(n5) );
  AOI22D2BWP12T U30 ( .A1(n3592), .A2(r5[0]), .B1(n3580), .B2(immediate2_in[0]), .ZN(n977) );
  BUFFXD8BWP12T U31 ( .I(n1945), .Z(n6) );
  ND3XD3BWP12T U32 ( .A1(n797), .A2(n8), .A3(n7), .ZN(regB_out[15]) );
  TPNR2D1BWP12T U33 ( .A1(n786), .A2(n787), .ZN(n7) );
  TPNR2D1BWP12T U34 ( .A1(n789), .A2(n788), .ZN(n8) );
  ND4D4BWP12T U35 ( .A1(n12), .A2(n11), .A3(n10), .A4(n9), .ZN(regA_out[23])
         );
  NR2XD2BWP12T U36 ( .A1(n1789), .A2(n1802), .ZN(n9) );
  NR2XD2BWP12T U37 ( .A1(n1790), .A2(n1788), .ZN(n10) );
  NR2XD2BWP12T U38 ( .A1(n1799), .A2(n1800), .ZN(n11) );
  NR2XD2BWP12T U39 ( .A1(n1791), .A2(n1801), .ZN(n12) );
  NR2D1BWP12T U40 ( .A1(n1024), .A2(n1023), .ZN(n1027) );
  CKND2D2BWP12T U41 ( .A1(n1924), .A2(r8[2]), .ZN(n1462) );
  INR2D4BWP12T U42 ( .A1(n1462), .B1(n1461), .ZN(n1467) );
  INVD12BWP12T U43 ( .I(n316), .ZN(n328) );
  INVD8BWP12T U44 ( .I(n1272), .ZN(n1942) );
  TPOAI22D2BWP12T U45 ( .A1(n3478), .A2(n2700), .B1(n3477), .B2(n2699), .ZN(
        n1707) );
  CKND2D4BWP12T U46 ( .A1(n329), .A2(n328), .ZN(n1468) );
  NR2D3BWP12T U47 ( .A1(n1257), .A2(n1256), .ZN(n1261) );
  INVD1BWP12T U48 ( .I(n982), .ZN(n13) );
  INVD2BWP12T U49 ( .I(n983), .ZN(n14) );
  CKND2D2BWP12T U50 ( .A1(n14), .A2(n13), .ZN(n990) );
  TPNR2D1BWP12T U51 ( .A1(n1363), .A2(n15), .ZN(n1377) );
  ND3D2BWP12T U52 ( .A1(n1360), .A2(n1361), .A3(n16), .ZN(n15) );
  INVD1BWP12T U53 ( .I(n1362), .ZN(n16) );
  CKND2D2BWP12T U54 ( .A1(n1653), .A2(lr[1]), .ZN(n1247) );
  TPND2D2BWP12T U55 ( .A1(n1942), .A2(r5[1]), .ZN(n1262) );
  TPNR2D2BWP12T U56 ( .A1(n1093), .A2(n1092), .ZN(n1101) );
  ND2D1BWP12T U57 ( .A1(n1946), .A2(n[3690]), .ZN(n341) );
  TPNR3D4BWP12T U58 ( .A1(n360), .A2(n358), .A3(n359), .ZN(n372) );
  OAI22D2BWP12T U59 ( .A1(n3491), .A2(n2784), .B1(n3490), .B2(n1429), .ZN(
        n1210) );
  INVD4BWP12T U60 ( .I(n1286), .ZN(n34) );
  TPND2D2BWP12T U61 ( .A1(n1849), .A2(n1848), .ZN(n1853) );
  AOI22D2BWP12T U62 ( .A1(r9[20]), .A2(n3471), .B1(n3472), .B2(tmp1[20]), .ZN(
        n1486) );
  IOA21D2BWP12T U63 ( .A1(n3474), .A2(r2[20]), .B(n1486), .ZN(n1488) );
  TPOAI21D1BWP12T U64 ( .A1(n234), .A2(n1944), .B(n1943), .ZN(n1957) );
  OR2D2BWP12T U65 ( .A1(n1901), .A2(n1900), .Z(n1902) );
  OAI21D0BWP12T U66 ( .A1(n3586), .A2(n1903), .B(n1902), .ZN(n1904) );
  ND4D2BWP12T U67 ( .A1(n1102), .A2(n1101), .A3(n1100), .A4(n17), .ZN(
        regA_out[28]) );
  TPNR2D2BWP12T U68 ( .A1(n1096), .A2(n1097), .ZN(n17) );
  INVD18BWP12T U69 ( .I(n[3699]), .ZN(n18) );
  TPNR2D1BWP12T U70 ( .A1(n381), .A2(n18), .ZN(n1257) );
  TPND2D1BWP12T U71 ( .A1(n3534), .A2(n3533), .ZN(regB_out[30]) );
  TPND2D1BWP12T U72 ( .A1(n1857), .A2(n3335), .ZN(n1858) );
  ND2D4BWP12T U73 ( .A1(n1946), .A2(n[3683]), .ZN(n1151) );
  TPOAI22D2BWP12T U74 ( .A1(n3487), .A2(n1094), .B1(n3486), .B2(n3648), .ZN(
        n1097) );
  INR2D4BWP12T U75 ( .A1(r11[1]), .B1(n3490), .ZN(n1256) );
  INVD3BWP12T U76 ( .I(n39), .ZN(n1658) );
  AOI22D1BWP12T U77 ( .A1(r12[2]), .A2(n1952), .B1(n1642), .B2(r6[2]), .ZN(
        n1479) );
  TPND2D1BWP12T U78 ( .A1(n3444), .A2(n3443), .ZN(regA_out[27]) );
  OR2D4BWP12T U79 ( .A1(n920), .A2(n919), .Z(n925) );
  NR2D4BWP12T U80 ( .A1(n925), .A2(n924), .ZN(n926) );
  OAI22D1BWP12T U81 ( .A1(n1195), .A2(n3463), .B1(n3492), .B2(n1196), .ZN(n384) );
  OAI22D2BWP12T U82 ( .A1(n3481), .A2(n1507), .B1(n1492), .B2(n3422), .ZN(
        n1493) );
  NR2D2BWP12T U83 ( .A1(n1494), .A2(n1493), .ZN(n1499) );
  ND2D4BWP12T U84 ( .A1(n328), .A2(n34), .ZN(n1337) );
  INR3XD2BWP12T U85 ( .A1(n370), .B1(n369), .B2(n368), .ZN(n371) );
  TPND2D3BWP12T U86 ( .A1(n301), .A2(n280), .ZN(n281) );
  BUFFXD8BWP12T U87 ( .I(n281), .Z(n3582) );
  OAI22D1BWP12T U88 ( .A1(n3656), .A2(n3571), .B1(n3607), .B2(n3661), .ZN(
        n3530) );
  NR3D3BWP12T U89 ( .A1(n1478), .A2(n1474), .A3(n1473), .ZN(n1484) );
  TPND2D8BWP12T U90 ( .A1(n309), .A2(readA_sel[1]), .ZN(n316) );
  TPNR2D1BWP12T U91 ( .A1(n396), .A2(n3381), .ZN(n397) );
  ND3D2BWP12T U92 ( .A1(n237), .A2(n19), .A3(n20), .ZN(n1255) );
  INVD2BWP12T U93 ( .I(n1245), .ZN(n19) );
  TPND2D2BWP12T U94 ( .A1(n1642), .A2(r6[1]), .ZN(n20) );
  TPOAI22D1BWP12T U95 ( .A1(n3586), .A2(n1621), .B1(n1901), .B2(n287), .ZN(
        n288) );
  TPND2D2BWP12T U96 ( .A1(n3472), .A2(tmp1[1]), .ZN(n1250) );
  INVD9BWP12T U97 ( .I(n1633), .ZN(n3477) );
  TPOAI22D1BWP12T U98 ( .A1(n1884), .A2(n2700), .B1(n1913), .B2(n1712), .ZN(
        n787) );
  ND3D1BWP12T U99 ( .A1(n3371), .A2(n3370), .A3(n21), .ZN(n2198) );
  OA21D1BWP12T U100 ( .A1(n3366), .A2(n3367), .B(n167), .Z(n21) );
  NR2XD2BWP12T U101 ( .A1(n1967), .A2(n1966), .ZN(n1895) );
  TPNR2D1BWP12T U102 ( .A1(n22), .A2(n1810), .ZN(n210) );
  OR3D2BWP12T U103 ( .A1(n1808), .A2(n1809), .A3(n23), .Z(n22) );
  TPOAI22D1BWP12T U104 ( .A1(n3571), .A2(n2677), .B1(n3607), .B2(n1806), .ZN(
        n23) );
  ND2XD8BWP12T U105 ( .A1(write1_in[24]), .A2(n47), .ZN(n46) );
  INVD8BWP12T U106 ( .I(readA_sel[0]), .ZN(n335) );
  INVD3BWP12T U107 ( .I(n330), .ZN(n1272) );
  TPOAI22D1BWP12T U108 ( .A1(n3586), .A2(n1526), .B1(n3588), .B2(n1525), .ZN(
        n1527) );
  TPND2D2BWP12T U109 ( .A1(n353), .A2(n24), .ZN(n360) );
  CKAN2D2BWP12T U110 ( .A1(n351), .A2(n352), .Z(n24) );
  TPOAI22D2BWP12T U111 ( .A1(n3584), .A2(n969), .B1(n3582), .B2(n968), .ZN(
        n973) );
  DCCKND4BWP12T U112 ( .I(n3344), .ZN(n3333) );
  OR2D4BWP12T U113 ( .A1(n1960), .A2(n1891), .Z(n1967) );
  CKND4BWP12T U114 ( .I(n[3677]), .ZN(n1796) );
  INVD4BWP12T U115 ( .I(write1_in[27]), .ZN(n43) );
  ND2D2BWP12T U116 ( .A1(n450), .A2(n449), .ZN(n2197) );
  TPNR3D2BWP12T U117 ( .A1(n1626), .A2(n1625), .A3(n1624), .ZN(n1641) );
  TPOAI22D2BWP12T U118 ( .A1(n3489), .A2(n1833), .B1(n1832), .B2(n3488), .ZN(
        n1838) );
  NR4D3BWP12T U119 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .ZN(n348) );
  ND3XD4BWP12T U120 ( .A1(n348), .A2(n347), .A3(n346), .ZN(regA_out[10]) );
  INVD1BWP12T U121 ( .I(n25), .ZN(n399) );
  TPNR2D2BWP12T U122 ( .A1(n3340), .A2(n398), .ZN(n25) );
  TPAOI21D8BWP12T U123 ( .A1(write1_in[26]), .A2(n3381), .B(n397), .ZN(n3340)
         );
  ND3D1BWP12T U124 ( .A1(n29), .A2(n26), .A3(n3332), .ZN(n2194) );
  TPAOI31D1BWP12T U125 ( .A1(n3323), .A2(n45), .A3(n27), .B(n3330), .ZN(n26)
         );
  TPNR2D2BWP12T U126 ( .A1(n28), .A2(n3344), .ZN(n27) );
  INVD1BWP12T U127 ( .I(n3322), .ZN(n28) );
  INVD1BWP12T U128 ( .I(n3331), .ZN(n29) );
  BUFFXD6BWP12T U129 ( .I(write1_in[31]), .Z(n3259) );
  TPNR2D2BWP12T U130 ( .A1(n1241), .A2(n30), .ZN(n1242) );
  ND3D2BWP12T U131 ( .A1(n1238), .A2(n31), .A3(n1237), .ZN(n30) );
  INVD1BWP12T U132 ( .I(n32), .ZN(n31) );
  INR2D2BWP12T U133 ( .A1(n33), .B1(n3437), .ZN(n32) );
  INVD1BWP12T U134 ( .I(n2866), .ZN(n33) );
  ND2XD4BWP12T U135 ( .A1(n3390), .A2(n447), .ZN(n3366) );
  ND2D8BWP12T U136 ( .A1(write1_in[28]), .A2(n3381), .ZN(n3390) );
  INR2D1BWP12T U137 ( .A1(n3381), .B1(write1_in[27]), .ZN(n256) );
  TPND2D3BWP12T U138 ( .A1(n3324), .A2(n1865), .ZN(n3348) );
  TPND2D3BWP12T U139 ( .A1(n3322), .A2(n3320), .ZN(n3324) );
  ND2XD3BWP12T U140 ( .A1(write1_in[25]), .A2(n1856), .ZN(n3322) );
  TPAOI31D1BWP12T U141 ( .A1(write1_in[27]), .A2(write1_in[26]), .A3(n1856), 
        .B(n3356), .ZN(n3358) );
  TPND2D3BWP12T U142 ( .A1(n34), .A2(n1291), .ZN(n1700) );
  CKND2D2BWP12T U143 ( .A1(n1274), .A2(n1273), .ZN(n1284) );
  TPNR3D4BWP12T U144 ( .A1(n1284), .A2(n1283), .A3(n1282), .ZN(n1304) );
  TPOAI22D1BWP12T U145 ( .A1(n3584), .A2(n1699), .B1(n3582), .B2(n1703), .ZN(
        n791) );
  NR2D2BWP12T U146 ( .A1(n791), .A2(n790), .ZN(n796) );
  TPAOI21D2BWP12T U147 ( .A1(n1926), .A2(r6[8]), .B(n1364), .ZN(n1367) );
  TPND3D2BWP12T U148 ( .A1(n1367), .A2(n1366), .A3(n1365), .ZN(n1375) );
  TPND2D1BWP12T U149 ( .A1(n3498), .A2(n3497), .ZN(regA_out[31]) );
  TPND2D1BWP12T U150 ( .A1(n1953), .A2(n1954), .ZN(n1955) );
  TPND2D4BWP12T U151 ( .A1(n1118), .A2(n1117), .ZN(regA_out[13]) );
  AOI22D2BWP12T U152 ( .A1(r9[28]), .A2(n3471), .B1(n3472), .B2(tmp1[28]), 
        .ZN(n1087) );
  IOA21D2BWP12T U153 ( .A1(n3474), .A2(r2[28]), .B(n1087), .ZN(n1088) );
  INR2D4BWP12T U154 ( .A1(r10[11]), .B1(n3422), .ZN(n1662) );
  INVD2BWP12T U155 ( .I(n3347), .ZN(n3342) );
  BUFFXD12BWP12T U156 ( .I(n374), .Z(n3448) );
  CKND3BWP12T U157 ( .I(write1_in[29]), .ZN(n3620) );
  CKND2D4BWP12T U158 ( .A1(n1304), .A2(n1303), .ZN(regA_out[9]) );
  ND2D2BWP12T U159 ( .A1(n35), .A2(n1136), .ZN(n1137) );
  ND2D2BWP12T U160 ( .A1(n1131), .A2(n36), .ZN(n35) );
  INVD2BWP12T U161 ( .I(n37), .ZN(n36) );
  OAI21D1BWP12T U162 ( .A1(write1_in[30]), .A2(n1134), .B(n38), .ZN(n37) );
  AN2XD2BWP12T U163 ( .A1(n1133), .A2(n3363), .Z(n38) );
  ND2D8BWP12T U164 ( .A1(write1_in[29]), .A2(n3381), .ZN(n1131) );
  ND2D3BWP12T U165 ( .A1(write1_in[31]), .A2(n3381), .ZN(n3385) );
  MAOI22D1BWP12T U166 ( .A1(n544), .A2(n64), .B1(n64), .B2(n544), .ZN(n65) );
  TPND2D2BWP12T U167 ( .A1(n665), .A2(n512), .ZN(n1960) );
  TPND2D2BWP12T U168 ( .A1(n3162), .A2(n3161), .ZN(n2226) );
  MOAI22D1BWP12T U169 ( .A1(n1960), .A2(n1961), .B1(n1960), .B2(n1961), .ZN(
        n195) );
  INVD3BWP12T U170 ( .I(n508), .ZN(n509) );
  TPND2D1BWP12T U171 ( .A1(n247), .A2(n3628), .ZN(n496) );
  TPNR2D3BWP12T U172 ( .A1(n728), .A2(n729), .ZN(n731) );
  MUX2ND4BWP12T U173 ( .I0(write1_in[6]), .I1(n2921), .S(n3393), .ZN(n728) );
  TPND2D3BWP12T U174 ( .A1(n733), .A2(n732), .ZN(n729) );
  RCOAI21D1BWP12T U175 ( .A1(n1965), .A2(n3394), .B(n1964), .ZN(n2186) );
  TPOAI21D1BWP12T U176 ( .A1(n65), .A2(n3394), .B(n66), .ZN(n2184) );
  XNR2D1BWP12T U177 ( .A1(n1974), .A2(n1973), .ZN(n1976) );
  TPND2D2BWP12T U178 ( .A1(n479), .A2(n478), .ZN(spin[26]) );
  TPNR2D3BWP12T U179 ( .A1(n2944), .A2(n2943), .ZN(n733) );
  TPND2D2BWP12T U180 ( .A1(n484), .A2(n483), .ZN(n2419) );
  TPND2D2BWP12T U181 ( .A1(n3300), .A2(n3299), .ZN(n2323) );
  TPND2D2BWP12T U182 ( .A1(n3302), .A2(n3301), .ZN(n2579) );
  TPND2D2BWP12T U183 ( .A1(n3305), .A2(n3304), .ZN(n2547) );
  TPND2D2BWP12T U184 ( .A1(n3309), .A2(n3308), .ZN(n2291) );
  TPND2D2BWP12T U185 ( .A1(n507), .A2(n506), .ZN(n2355) );
  TPND2D2BWP12T U186 ( .A1(n3283), .A2(n3282), .ZN(n2515) );
  TPND2D2BWP12T U187 ( .A1(n3275), .A2(n3274), .ZN(n2483) );
  TPND2D2BWP12T U188 ( .A1(n3288), .A2(n3287), .ZN(n2643) );
  TPND2D2BWP12T U189 ( .A1(n489), .A2(n488), .ZN(n2387) );
  TPND2D2BWP12T U190 ( .A1(n455), .A2(n454), .ZN(n2259) );
  TPND2D2BWP12T U191 ( .A1(n474), .A2(n473), .ZN(n2227) );
  TPND2D2BWP12T U192 ( .A1(n3293), .A2(n3292), .ZN(n2611) );
  TPND2D2BWP12T U193 ( .A1(n3279), .A2(n3278), .ZN(n2163) );
  TPNR2D2BWP12T U194 ( .A1(n1970), .A2(n1977), .ZN(n811) );
  TPND3D3BWP12T U195 ( .A1(n1613), .A2(readA_sel[0]), .A3(readA_sel[3]), .ZN(
        n39) );
  TPND3D3BWP12T U196 ( .A1(n1613), .A2(readA_sel[0]), .A3(readA_sel[3]), .ZN(
        n1286) );
  TPND2D2BWP12T U197 ( .A1(n3208), .A2(n3207), .ZN(n2424) );
  OR2D2BWP12T U198 ( .A1(n3396), .A2(n575), .Z(n3208) );
  ND2D4BWP12T U199 ( .A1(n1698), .A2(n1697), .ZN(regB_out[2]) );
  TPND2D1BWP12T U200 ( .A1(n3175), .A2(n3229), .ZN(n3117) );
  CKND2D2BWP12T U201 ( .A1(n3117), .A2(n3116), .ZN(spin[27]) );
  INVD1BWP12T U202 ( .I(n3396), .ZN(n232) );
  TPND2D2BWP12T U203 ( .A1(n3247), .A2(n3246), .ZN(n2456) );
  TPND2D1BWP12T U204 ( .A1(n3175), .A2(n3627), .ZN(n3177) );
  CKND2D2BWP12T U205 ( .A1(n3177), .A2(n3176), .ZN(n2324) );
  TPND2D1BWP12T U206 ( .A1(n3175), .A2(n3625), .ZN(n3172) );
  CKND2D2BWP12T U207 ( .A1(n3172), .A2(n3171), .ZN(n2580) );
  TPND2D1BWP12T U208 ( .A1(n3175), .A2(n3624), .ZN(n3170) );
  CKND2D2BWP12T U209 ( .A1(n3170), .A2(n3169), .ZN(n2548) );
  TPND2D1BWP12T U210 ( .A1(n3175), .A2(n3241), .ZN(n3142) );
  CKND2D2BWP12T U211 ( .A1(n3142), .A2(n3141), .ZN(n2420) );
  TPND2D1BWP12T U212 ( .A1(n3175), .A2(n3626), .ZN(n3168) );
  CKND2D2BWP12T U213 ( .A1(n3168), .A2(n3167), .ZN(n2292) );
  TPND2D1BWP12T U214 ( .A1(n3175), .A2(n3248), .ZN(n3144) );
  CKND2D2BWP12T U215 ( .A1(n3144), .A2(n3143), .ZN(n2356) );
  TPND2D1BWP12T U216 ( .A1(n3175), .A2(n3622), .ZN(n3136) );
  CKND2D2BWP12T U217 ( .A1(n3136), .A2(n3135), .ZN(n2484) );
  TPND2D1BWP12T U218 ( .A1(n3175), .A2(n3628), .ZN(n3166) );
  CKND2D2BWP12T U219 ( .A1(n3166), .A2(n3165), .ZN(n2452) );
  TPND2D1BWP12T U220 ( .A1(n3175), .A2(n3284), .ZN(n3132) );
  CKND2D2BWP12T U221 ( .A1(n3132), .A2(n3131), .ZN(n2644) );
  TPND2D1BWP12T U222 ( .A1(n3175), .A2(n3216), .ZN(n3128) );
  CKND2D2BWP12T U223 ( .A1(n3128), .A2(n3127), .ZN(n2260) );
  TPND2D1BWP12T U224 ( .A1(n3175), .A2(n3234), .ZN(n3140) );
  CKND2D2BWP12T U225 ( .A1(n3140), .A2(n3139), .ZN(n2228) );
  TPND2D1BWP12T U226 ( .A1(n3175), .A2(n3289), .ZN(n3130) );
  CKND2D2BWP12T U227 ( .A1(n3130), .A2(n3129), .ZN(n2612) );
  TPND2D1BWP12T U228 ( .A1(n3175), .A2(n3638), .ZN(n3138) );
  CKND2D2BWP12T U229 ( .A1(n3138), .A2(n3137), .ZN(n2164) );
  TPND2D2BWP12T U230 ( .A1(n3134), .A2(n3133), .ZN(n2516) );
  TPND2D1BWP12T U231 ( .A1(n3175), .A2(n3623), .ZN(n3134) );
  TPND2D1BWP12T U232 ( .A1(n3184), .A2(n3229), .ZN(n3158) );
  TPND2D1BWP12T U233 ( .A1(n3184), .A2(n3638), .ZN(n3160) );
  TPND2D1BWP12T U234 ( .A1(n3184), .A2(n3624), .ZN(n3186) );
  TPND2D1BWP12T U235 ( .A1(n3184), .A2(n3248), .ZN(n3174) );
  TPND2D1BWP12T U236 ( .A1(n3184), .A2(n3622), .ZN(n3156) );
  TPND2D1BWP12T U237 ( .A1(n3184), .A2(n3623), .ZN(n3152) );
  TPND2D1BWP12T U238 ( .A1(n3184), .A2(n3284), .ZN(n3154) );
  TPND2D1BWP12T U239 ( .A1(n3184), .A2(n3216), .ZN(n3148) );
  TPND2D1BWP12T U240 ( .A1(n3184), .A2(n3234), .ZN(n3162) );
  TPND2D2BWP12T U241 ( .A1(n3146), .A2(n3145), .ZN(n2386) );
  TPND2D1BWP12T U242 ( .A1(n3184), .A2(n3211), .ZN(n3146) );
  TPND2D2BWP12T U243 ( .A1(n3123), .A2(n3122), .ZN(n2388) );
  TPND2D1BWP12T U244 ( .A1(n3175), .A2(n3211), .ZN(n3123) );
  TPND2D2BWP12T U245 ( .A1(n496), .A2(n495), .ZN(n2451) );
  RCAOI21D1BWP12T U246 ( .A1(n3325), .A2(n3316), .B(n3315), .ZN(n3317) );
  INR3D2BWP12T U247 ( .A1(n3321), .B1(n238), .B2(n3325), .ZN(n3323) );
  NR2XD3BWP12T U248 ( .A1(n909), .A2(n908), .ZN(n910) );
  OR2D4BWP12T U249 ( .A1(n904), .A2(n903), .Z(n909) );
  TPND2D2BWP12T U250 ( .A1(n1377), .A2(n1376), .ZN(regA_out[8]) );
  ND2XD8BWP12T U251 ( .A1(n1351), .A2(n1350), .ZN(regA_out[14]) );
  NR2D4BWP12T U252 ( .A1(write1_in[19]), .A2(n3393), .ZN(n436) );
  TPND2D2BWP12T U253 ( .A1(n643), .A2(n642), .ZN(spin[30]) );
  TPND2D2BWP12T U254 ( .A1(n639), .A2(n638), .ZN(n2423) );
  TPND2D2BWP12T U255 ( .A1(n832), .A2(n831), .ZN(n2359) );
  TPND2D2BWP12T U256 ( .A1(n637), .A2(n636), .ZN(n2647) );
  TPND2D2BWP12T U257 ( .A1(n826), .A2(n825), .ZN(n2391) );
  TPND2D2BWP12T U258 ( .A1(n641), .A2(n640), .ZN(n2615) );
  TPND2D2BWP12T U259 ( .A1(n828), .A2(n827), .ZN(n2263) );
  NR2XD2BWP12T U260 ( .A1(n2924), .A2(n2925), .ZN(n2930) );
  XNR2XD0BWP12T U261 ( .A1(n2924), .A2(n2925), .ZN(n2927) );
  INVD4BWP12T U262 ( .I(n261), .ZN(n1685) );
  TPND2D1BWP12T U263 ( .A1(n3344), .A2(n3312), .ZN(n3318) );
  ND3XD4BWP12T U264 ( .A1(n811), .A2(n1971), .A3(n812), .ZN(n3344) );
  TPND2D2BWP12T U265 ( .A1(n462), .A2(n461), .ZN(n2518) );
  TPND2D3BWP12T U266 ( .A1(n664), .A2(n544), .ZN(n511) );
  TPND2D2BWP12T U267 ( .A1(n501), .A2(n500), .ZN(n2646) );
  TPND2D2BWP12T U268 ( .A1(n491), .A2(n490), .ZN(n2390) );
  TPNR2D2BWP12T U269 ( .A1(write1_in[17]), .A2(n3362), .ZN(n409) );
  ND2D3BWP12T U270 ( .A1(n299), .A2(n298), .ZN(n792) );
  TPND2D2BWP12T U271 ( .A1(n469), .A2(n468), .ZN(n2614) );
  INVD1BWP12T U272 ( .I(write1_in[2]), .ZN(n40) );
  INVD1BWP12T U273 ( .I(n40), .ZN(n41) );
  DEL025D1BWP12T U274 ( .I(write1_in[13]), .Z(n42) );
  DCCKND4BWP12T U275 ( .I(n3619), .ZN(n249) );
  TPND2D2BWP12T U276 ( .A1(n830), .A2(n829), .ZN(n2231) );
  DCCKND4BWP12T U277 ( .I(n511), .ZN(n512) );
  MAOI22D1BWP12T U278 ( .A1(n700), .A2(n99), .B1(n700), .B2(n99), .ZN(n100) );
  TPND2D3BWP12T U279 ( .A1(n844), .A2(n700), .ZN(n508) );
  TPOAI21D4BWP12T U280 ( .A1(n421), .A2(n3379), .B(n420), .ZN(n700) );
  INVD2BWP12T U281 ( .I(n3329), .ZN(n3328) );
  TPND2D2BWP12T U282 ( .A1(n3256), .A2(n3255), .ZN(n2552) );
  TPND2D2BWP12T U283 ( .A1(n3254), .A2(n3253), .ZN(n2328) );
  TPND2D2BWP12T U284 ( .A1(n3258), .A2(n3257), .ZN(n2584) );
  TPND2D2BWP12T U285 ( .A1(n3261), .A2(n3260), .ZN(n2296) );
  TPOAI21D4BWP12T U286 ( .A1(n430), .A2(n429), .B(n428), .ZN(n2929) );
  INVD2BWP12T U287 ( .I(write1_in[3]), .ZN(n430) );
  AN2XD2BWP12T U288 ( .A1(n1867), .A2(n3352), .Z(n1868) );
  INR3D1BWP12T U289 ( .A1(n3354), .B1(n3353), .B2(n240), .ZN(n3361) );
  ND2D3BWP12T U290 ( .A1(n1942), .A2(r5[8]), .ZN(n1357) );
  INVD2BWP12T U291 ( .I(n1359), .ZN(n1360) );
  TPOAI22D1BWP12T U292 ( .A1(n3584), .A2(n1055), .B1(n3582), .B2(n1240), .ZN(
        n1059) );
  INR3D2BWP12T U293 ( .A1(n1155), .B1(n1154), .B2(n1153), .ZN(n1164) );
  OAI211D1BWP12T U294 ( .A1(n3478), .A2(n2795), .B(n1152), .C(n1151), .ZN(
        n1153) );
  INVD12BWP12T U295 ( .I(n1942), .ZN(n3489) );
  TPND2D2BWP12T U296 ( .A1(n1942), .A2(r5[17]), .ZN(n1146) );
  OAI22D2BWP12T U297 ( .A1(n3448), .A2(n1523), .B1(n3476), .B2(n1525), .ZN(
        n1115) );
  OAI22D1BWP12T U298 ( .A1(n1503), .A2(n3463), .B1(n3492), .B2(n1502), .ZN(
        n1487) );
  TPOAI22D1BWP12T U299 ( .A1(n3588), .A2(n1072), .B1(n3586), .B2(n1073), .ZN(
        n217) );
  NR4D1BWP12T U300 ( .A1(n1084), .A2(n1083), .A3(n1082), .A4(n1081), .ZN(n1085) );
  TPOAI22D1BWP12T U301 ( .A1(n3612), .A2(n1080), .B1(n3611), .B2(n1079), .ZN(
        n1081) );
  TPOAI22D1BWP12T U302 ( .A1(n3478), .A2(n1787), .B1(n3477), .B2(n2689), .ZN(
        n1788) );
  TPNR2D2BWP12T U303 ( .A1(n438), .A2(n1978), .ZN(n44) );
  TPNR2D2BWP12T U304 ( .A1(n438), .A2(n1978), .ZN(n3377) );
  BUFFXD3BWP12T U305 ( .I(write1_in[25]), .Z(n3184) );
  TPND2D2BWP12T U306 ( .A1(n3150), .A2(n3149), .ZN(n2610) );
  TPND2D1BWP12T U307 ( .A1(n3184), .A2(n3289), .ZN(n3150) );
  TPOAI21D1BWP12T U308 ( .A1(n3463), .A2(n1533), .B(n1105), .ZN(n1106) );
  DCCKBD4BWP12T U309 ( .I(n3335), .Z(n45) );
  ND2D8BWP12T U310 ( .A1(n46), .A2(n815), .ZN(n3335) );
  DCCKND4BWP12T U311 ( .I(n3362), .ZN(n47) );
  ND2XD3BWP12T U312 ( .A1(write1_in[15]), .A2(n3381), .ZN(n417) );
  CKND2D2BWP12T U313 ( .A1(n274), .A2(n280), .ZN(n275) );
  TPND2D2BWP12T U314 ( .A1(n3475), .A2(n251), .ZN(n252) );
  TPND2D4BWP12T U315 ( .A1(n317), .A2(n311), .ZN(n374) );
  IOA21D2BWP12T U316 ( .A1(n1950), .A2(r7[15]), .B(n1714), .ZN(n1719) );
  INR2D8BWP12T U317 ( .A1(n297), .B1(n296), .ZN(n3580) );
  TPNR2D4BWP12T U318 ( .A1(n39), .A2(n1287), .ZN(n1945) );
  IAO22D1BWP12T U319 ( .B1(n1950), .B2(r7[9]), .A1(n1271), .A2(n1272), .ZN(
        n1273) );
  TPND2D2BWP12T U320 ( .A1(n1950), .A2(r7[10]), .ZN(n322) );
  BUFFXD4BWP12T U321 ( .I(readB_sel[0]), .Z(n298) );
  INVD2BWP12T U322 ( .I(n3337), .ZN(n3338) );
  TPOAI22D1BWP12T U323 ( .A1(n3491), .A2(n1561), .B1(n3490), .B2(n1560), .ZN(
        n1564) );
  CKND2D2BWP12T U324 ( .A1(n301), .A2(n300), .ZN(n302) );
  TPOAI22D1BWP12T U325 ( .A1(n3586), .A2(n1710), .B1(n3588), .B2(n1702), .ZN(
        n790) );
  TPND2D2BWP12T U326 ( .A1(n252), .A2(n1248), .ZN(n1254) );
  CKND2D2BWP12T U327 ( .A1(n3160), .A2(n3159), .ZN(n2162) );
  TPNR2D3BWP12T U328 ( .A1(n3340), .A2(n3394), .ZN(n3347) );
  TPOAI22D1BWP12T U329 ( .A1(n3509), .A2(n3463), .B1(n3437), .B2(n3510), .ZN(
        n1013) );
  TPNR3D2BWP12T U330 ( .A1(n1267), .A2(n1266), .A3(n1265), .ZN(n1268) );
  ND2D1BWP12T U331 ( .A1(n313), .A2(n312), .ZN(n325) );
  NR2D1BWP12T U332 ( .A1(n3562), .A2(n3561), .ZN(n3565) );
  NR2D2BWP12T U333 ( .A1(n1259), .A2(n1258), .ZN(n1260) );
  IND2D1BWP12T U334 ( .A1(n3344), .B1(n3326), .ZN(n3327) );
  TPND2D1BWP12T U335 ( .A1(n1472), .A2(n1471), .ZN(n1473) );
  CKND2D0BWP12T U336 ( .A1(n235), .A2(r0[2]), .ZN(n1477) );
  OAI22D1BWP12T U337 ( .A1(n3478), .A2(n1552), .B1(n3477), .B2(n1551), .ZN(
        n1553) );
  ND3D1BWP12T U338 ( .A1(n1650), .A2(n1649), .A3(n1648), .ZN(n1657) );
  ND2D1BWP12T U339 ( .A1(n235), .A2(r0[11]), .ZN(n1649) );
  ND2D1BWP12T U340 ( .A1(write2_in[29]), .A2(n3379), .ZN(n3363) );
  NR2D0BWP12T U341 ( .A1(n3325), .A2(n238), .ZN(n3326) );
  ND2D1BWP12T U342 ( .A1(n3335), .A2(n3310), .ZN(n1864) );
  INR2D1BWP12T U343 ( .A1(write1_sel[1]), .B1(write1_sel[2]), .ZN(n538) );
  INVD1BWP12T U344 ( .I(write1_sel[0]), .ZN(n457) );
  INR2D1BWP12T U345 ( .A1(write1_en), .B1(write1_sel[4]), .ZN(n456) );
  NR2D1BWP12T U346 ( .A1(n238), .A2(n3394), .ZN(n1857) );
  INR2D1BWP12T U347 ( .A1(n457), .B1(n463), .ZN(n539) );
  INR2D1BWP12T U348 ( .A1(write1_sel[0]), .B1(n463), .ZN(n583) );
  ND2D1BWP12T U349 ( .A1(n538), .A2(n3621), .ZN(n534) );
  CKND2D0BWP12T U350 ( .A1(next_pc_en_BAR), .A2(n440), .ZN(n3399) );
  IND2D1BWP12T U351 ( .A1(n1961), .B1(n1962), .ZN(n1891) );
  TPOAI21D1BWP12T U352 ( .A1(write1_in[18]), .A2(n3393), .B(n1893), .ZN(n1966)
         );
  INVD1BWP12T U353 ( .I(n3399), .ZN(n2989) );
  AOI22D1BWP12T U354 ( .A1(n3471), .A2(r9[13]), .B1(n3472), .B2(tmp1[13]), 
        .ZN(n1111) );
  ND2D1BWP12T U355 ( .A1(n3474), .A2(r2[13]), .ZN(n1110) );
  TPOAI22D1BWP12T U356 ( .A1(n3478), .A2(n2845), .B1(n3477), .B2(n1535), .ZN(
        n1114) );
  ND2D1BWP12T U357 ( .A1(n3474), .A2(r2[2]), .ZN(n1472) );
  ND2D1BWP12T U358 ( .A1(n3475), .A2(r4[2]), .ZN(n1471) );
  TPOAI22D1BWP12T U359 ( .A1(n3487), .A2(n1104), .B1(n3486), .B2(n1539), .ZN(
        n1107) );
  ND2D1BWP12T U360 ( .A1(n1952), .A2(r12[13]), .ZN(n1105) );
  TPOAI22D1BWP12T U361 ( .A1(n3481), .A2(n3610), .B1(n3479), .B2(n913), .ZN(
        n914) );
  INR2D1BWP12T U362 ( .A1(write2_en), .B1(write2_sel[4]), .ZN(n451) );
  INR2D1BWP12T U363 ( .A1(n451), .B1(write2_sel[0]), .ZN(n458) );
  OAI22D1BWP12T U364 ( .A1(n3481), .A2(n1773), .B1(n3422), .B2(n897), .ZN(n898) );
  TPOAI22D1BWP12T U365 ( .A1(n3481), .A2(n1404), .B1(n3422), .B2(n1403), .ZN(
        n1410) );
  TPOAI22D1BWP12T U366 ( .A1(n3611), .A2(n1392), .B1(n3612), .B2(n2727), .ZN(
        n1397) );
  OAI22D1BWP12T U367 ( .A1(n1389), .A2(n3600), .B1(n3599), .B2(n2074), .ZN(
        n1390) );
  ND4D1BWP12T U368 ( .A1(n1501), .A2(n1500), .A3(n1499), .A4(n1498), .ZN(
        regA_out[20]) );
  CKND2D0BWP12T U369 ( .A1(n1946), .A2(n[3698]), .ZN(n1463) );
  ND3D1BWP12T U370 ( .A1(n1477), .A2(n1476), .A3(n1475), .ZN(n1478) );
  AN2D1BWP12T U371 ( .A1(write2_sel[0]), .A2(n451), .Z(n465) );
  INVD1BWP12T U372 ( .I(n520), .ZN(n485) );
  ND2D1BWP12T U373 ( .A1(n458), .A2(n464), .ZN(n492) );
  ND2D3BWP12T U374 ( .A1(n1018), .A2(n1017), .ZN(regA_out[25]) );
  AN2D1BWP12T U375 ( .A1(n465), .A2(n464), .Z(n585) );
  INVD1BWP12T U376 ( .I(n492), .ZN(n537) );
  NR2D1BWP12T U377 ( .A1(write2_sel[2]), .A2(write2_sel[1]), .ZN(n503) );
  OAI22D1BWP12T U378 ( .A1(n3481), .A2(n1550), .B1(n3422), .B2(n1549), .ZN(
        n1554) );
  AOI22D1BWP12T U379 ( .A1(r9[6]), .A2(n3471), .B1(n3472), .B2(tmp1[6]), .ZN(
        n1213) );
  TPNR2D1BWP12T U380 ( .A1(n1218), .A2(n1217), .ZN(n1219) );
  ND2D1BWP12T U381 ( .A1(n3474), .A2(r2[23]), .ZN(n1781) );
  TPND3D1BWP12T U382 ( .A1(n1384), .A2(n1383), .A3(n1382), .ZN(n1385) );
  AOI22D1BWP12T U383 ( .A1(r10[3]), .A2(n3591), .B1(n3592), .B2(r5[3]), .ZN(
        n1382) );
  AOI22D1BWP12T U384 ( .A1(tmp1[15]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[15]), .ZN(n795) );
  AOI22D1BWP12T U385 ( .A1(n3592), .A2(r5[15]), .B1(n1327), .B2(r7[15]), .ZN(
        n793) );
  ND2D1BWP12T U386 ( .A1(n3475), .A2(r4[11]), .ZN(n1664) );
  OAI21D1BWP12T U387 ( .A1(n3463), .A2(n2969), .B(n1654), .ZN(n1655) );
  ND2D1BWP12T U388 ( .A1(n235), .A2(r0[3]), .ZN(n356) );
  ND2D1BWP12T U389 ( .A1(n3474), .A2(r2[3]), .ZN(n354) );
  AOI22D1BWP12T U390 ( .A1(r10[11]), .A2(n3591), .B1(n3592), .B2(r5[11]), .ZN(
        n934) );
  OAI22D1BWP12T U391 ( .A1(n3605), .A2(n2738), .B1(n3603), .B2(n938), .ZN(n941) );
  OAI22D1BWP12T U392 ( .A1(n3612), .A2(n943), .B1(n3611), .B2(n942), .ZN(n944)
         );
  OAI22D1BWP12T U393 ( .A1(n3489), .A2(n956), .B1(n3488), .B2(n980), .ZN(n961)
         );
  OAI21D1BWP12T U394 ( .A1(n3487), .A2(n958), .B(n957), .ZN(n960) );
  CKND0BWP12T U395 ( .I(r7[0]), .ZN(n958) );
  CKND2D0BWP12T U396 ( .A1(n1945), .A2(pc_out[0]), .ZN(n957) );
  OAI22D1BWP12T U397 ( .A1(n3422), .A2(n2664), .B1(n3481), .B2(n986), .ZN(n953) );
  INR2D1BWP12T U398 ( .A1(write1_sel[2]), .B1(n390), .ZN(n470) );
  ND2D1BWP12T U399 ( .A1(n3363), .A2(n3362), .ZN(n3364) );
  INVD1BWP12T U400 ( .I(n3381), .ZN(n3379) );
  ND2D1BWP12T U401 ( .A1(n2914), .A2(n3621), .ZN(n439) );
  INVD1BWP12T U402 ( .I(n528), .ZN(n531) );
  ND2D1BWP12T U403 ( .A1(n465), .A2(write2_sel[3]), .ZN(n528) );
  NR2D1BWP12T U404 ( .A1(n520), .A2(n527), .ZN(n523) );
  INR3D0BWP12T U405 ( .A1(n3621), .B1(write1_sel[2]), .B2(write1_sel[1]), .ZN(
        n502) );
  NR2D1BWP12T U406 ( .A1(n3628), .A2(reset), .ZN(n493) );
  INVD1BWP12T U407 ( .I(n502), .ZN(n497) );
  OR2XD1BWP12T U408 ( .A1(readC_sel[0]), .A2(readC_sel[1]), .Z(n1986) );
  INVD1BWP12T U409 ( .I(n475), .ZN(n582) );
  ND2D1BWP12T U410 ( .A1(n470), .A2(n3621), .ZN(n550) );
  AN2D1BWP12T U411 ( .A1(write2_in[20]), .A2(n3393), .Z(n412) );
  INVD1BWP12T U412 ( .I(n3333), .ZN(n3334) );
  TPND2D1BWP12T U413 ( .A1(n3397), .A2(n3402), .ZN(n3406) );
  INVD2BWP12T U414 ( .I(n3392), .ZN(n3397) );
  AN2D1BWP12T U415 ( .A1(write2_in[23]), .A2(n3393), .Z(n239) );
  TPND2D1BWP12T U416 ( .A1(n817), .A2(n822), .ZN(n820) );
  INVD1BWP12T U417 ( .I(n816), .ZN(n817) );
  CKND2D2BWP12T U418 ( .A1(n3333), .A2(n1865), .ZN(n822) );
  INVD1BWP12T U419 ( .I(n521), .ZN(n519) );
  NR2D1BWP12T U420 ( .A1(n554), .A2(n553), .ZN(n3277) );
  TPOAI21D1BWP12T U421 ( .A1(write1_in[16]), .A2(n3393), .B(n513), .ZN(n1961)
         );
  INVD1BWP12T U422 ( .I(n3231), .ZN(n2938) );
  NR2D1BWP12T U423 ( .A1(n476), .A2(n477), .ZN(n3231) );
  NR2D1BWP12T U424 ( .A1(n471), .A2(n472), .ZN(n3236) );
  NR2D1BWP12T U425 ( .A1(n452), .A2(n453), .ZN(n3218) );
  NR3D1BWP12T U426 ( .A1(n528), .A2(n530), .A3(n527), .ZN(n3307) );
  AN2D1BWP12T U427 ( .A1(n523), .A2(n522), .Z(n3298) );
  NR2D1BWP12T U428 ( .A1(n504), .A2(n505), .ZN(n3250) );
  NR2D1BWP12T U429 ( .A1(n486), .A2(n487), .ZN(n3213) );
  NR2D1BWP12T U430 ( .A1(n481), .A2(n482), .ZN(n3243) );
  INVD3BWP12T U431 ( .I(write1_in[31]), .ZN(n3396) );
  AN2D1BWP12T U432 ( .A1(n494), .A2(n493), .Z(n3263) );
  NR2D1BWP12T U433 ( .A1(n586), .A2(n587), .ZN(n3273) );
  NR2D1BWP12T U434 ( .A1(n459), .A2(n460), .ZN(n3281) );
  AN3XD1BWP12T U435 ( .A1(n516), .A2(n3621), .A3(n515), .Z(n3303) );
  AN3XD1BWP12T U436 ( .A1(n541), .A2(n3621), .A3(n540), .Z(n3373) );
  NR2D1BWP12T U437 ( .A1(n466), .A2(n467), .ZN(n3291) );
  BUFFXD3BWP12T U438 ( .I(write1_in[0]), .Z(n782) );
  BUFFXD0BWP12T U439 ( .I(write2_in[1]), .Z(n892) );
  BUFFXD0BWP12T U440 ( .I(write2_in[2]), .Z(n2882) );
  BUFFXD0BWP12T U441 ( .I(write2_in[3]), .Z(n2913) );
  BUFFXD0BWP12T U442 ( .I(write2_in[4]), .Z(n2887) );
  BUFFXD0BWP12T U443 ( .I(write2_in[5]), .Z(n2900) );
  BUFFXD0BWP12T U444 ( .I(write2_in[6]), .Z(n2921) );
  BUFFXD0BWP12T U445 ( .I(write2_in[8]), .Z(n866) );
  BUFFXD0BWP12T U446 ( .I(write2_in[9]), .Z(n2937) );
  BUFFXD0BWP12T U447 ( .I(write2_in[10]), .Z(n2951) );
  BUFFXD0BWP12T U448 ( .I(write2_in[11]), .Z(n2971) );
  BUFFXD0BWP12T U449 ( .I(write2_in[12]), .Z(n727) );
  BUFFXD0BWP12T U450 ( .I(write2_in[13]), .Z(n2972) );
  BUFFXD0BWP12T U451 ( .I(write2_in[14]), .Z(n2973) );
  BUFFXD0BWP12T U452 ( .I(write2_in[15]), .Z(n843) );
  NR2D1BWP12T U453 ( .A1(n498), .A2(n499), .ZN(n3286) );
  OR2XD1BWP12T U454 ( .A1(n1988), .A2(n1981), .Z(n2711) );
  OR2XD1BWP12T U455 ( .A1(n1984), .A2(n1981), .Z(n2827) );
  OR2XD1BWP12T U456 ( .A1(n1988), .A2(n1989), .Z(n2822) );
  OR2XD1BWP12T U457 ( .A1(n1990), .A2(n1981), .Z(n2653) );
  NR2D1BWP12T U458 ( .A1(n1990), .A2(n1989), .ZN(n2875) );
  NR2D1BWP12T U459 ( .A1(n1990), .A2(n1987), .ZN(n2857) );
  NR2D1BWP12T U460 ( .A1(n1987), .A2(n1986), .ZN(n2859) );
  NR2D1BWP12T U461 ( .A1(n1984), .A2(n1987), .ZN(n2856) );
  NR2D1BWP12T U462 ( .A1(n1985), .A2(n1984), .ZN(n2855) );
  NR2D1BWP12T U463 ( .A1(n1985), .A2(n1988), .ZN(n2854) );
  NR2D1BWP12T U464 ( .A1(n1985), .A2(n1986), .ZN(n2853) );
  NR2D1BWP12T U465 ( .A1(n1984), .A2(n1989), .ZN(n2869) );
  INVD1BWP12T U466 ( .I(n2653), .ZN(n2871) );
  NR2D1BWP12T U467 ( .A1(n1986), .A2(n1981), .ZN(n2873) );
  INVD1BWP12T U468 ( .I(n2822), .ZN(n2874) );
  INVD1BWP12T U469 ( .I(n2711), .ZN(n2870) );
  INVD1BWP12T U470 ( .I(n2827), .ZN(n2872) );
  NR2D1BWP12T U471 ( .A1(n1986), .A2(n1989), .ZN(n2848) );
  INVD1BWP12T U472 ( .I(readC_sel[4]), .ZN(n2864) );
  INVD1BWP12T U473 ( .I(readD_sel[4]), .ZN(n2970) );
  ND2D1BWP12T U474 ( .A1(n456), .A2(n391), .ZN(n526) );
  INVD16BWP12T U475 ( .I(n1666), .ZN(n3474) );
  BUFFXD4BWP12T U476 ( .I(n1394), .Z(n3571) );
  NR2D1BWP12T U477 ( .A1(n534), .A2(n526), .ZN(n3626) );
  INR2D1BWP12T U478 ( .A1(n539), .B1(n550), .ZN(n3628) );
  OAI21D1BWP12T U479 ( .A1(n1141), .A2(n3403), .B(n1140), .ZN(n1142) );
  AOI21D1BWP12T U480 ( .A1(n1863), .A2(n1867), .B(n1862), .ZN(n1871) );
  NR2D1BWP12T U481 ( .A1(n535), .A2(n534), .ZN(n3625) );
  NR2D1BWP12T U482 ( .A1(n514), .A2(n534), .ZN(n3624) );
  NR2D1BWP12T U483 ( .A1(n534), .A2(n519), .ZN(n3627) );
  RCOAI21D1BWP12T U484 ( .A1(n1969), .A2(n3394), .B(n1968), .ZN(n2187) );
  RCOAI21D1BWP12T U485 ( .A1(n1980), .A2(n3394), .B(n1979), .ZN(n2190) );
  ND2D1BWP12T U486 ( .A1(n3474), .A2(r2[7]), .ZN(n1848) );
  ND2D1BWP12T U487 ( .A1(n3474), .A2(r2[10]), .ZN(n319) );
  INVD1BWP12T U488 ( .I(n3471), .ZN(n233) );
  OAI22D1BWP12T U489 ( .A1(n2817), .A2(n3608), .B1(n1740), .B2(n1629), .ZN(
        n269) );
  AOI22D1BWP12T U490 ( .A1(r5[4]), .A2(n3592), .B1(n3591), .B2(r10[4]), .ZN(
        n306) );
  AOI22D2BWP12T U491 ( .A1(n295), .A2(tmp1[4]), .B1(immediate2_in[4]), .B2(
        n3580), .ZN(n304) );
  CKND2D0BWP12T U492 ( .A1(n1653), .A2(lr[10]), .ZN(n313) );
  ND2D1BWP12T U493 ( .A1(n3475), .A2(r4[10]), .ZN(n312) );
  ND2D1BWP12T U494 ( .A1(n235), .A2(r0[10]), .ZN(n343) );
  AOI22D0BWP12T U495 ( .A1(r9[29]), .A2(n3471), .B1(n3472), .B2(tmp1[29]), 
        .ZN(n993) );
  OAI22D1BWP12T U496 ( .A1(n3481), .A2(n1807), .B1(n1090), .B2(n3422), .ZN(
        n1093) );
  INR2D2BWP12T U497 ( .A1(r12[1]), .B1(n3437), .ZN(n1259) );
  OAI21D1BWP12T U498 ( .A1(n3492), .A2(n1297), .B(n1296), .ZN(n1301) );
  ND2D1BWP12T U499 ( .A1(n1946), .A2(n[3691]), .ZN(n1299) );
  OAI22D1BWP12T U500 ( .A1(n3571), .A2(n1552), .B1(n3607), .B2(n1557), .ZN(
        n1315) );
  AOI22D1BWP12T U501 ( .A1(tmp1[4]), .A2(n3472), .B1(n1617), .B2(n1616), .ZN(
        n1619) );
  CKND2D0BWP12T U502 ( .A1(n1945), .A2(pc_out[15]), .ZN(n1714) );
  AOI22D1BWP12T U503 ( .A1(r10[1]), .A2(n3591), .B1(n3592), .B2(r5[1]), .ZN(
        n1731) );
  OAI22D1BWP12T U504 ( .A1(n2821), .A2(n3600), .B1(n3599), .B2(n1736), .ZN(
        n1745) );
  AOI22D0BWP12T U505 ( .A1(tmp1[30]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[30]), .ZN(n3528) );
  NR4D0BWP12T U506 ( .A1(n1204), .A2(n1203), .A3(n1202), .A4(n1201), .ZN(n1205) );
  TPND3D1BWP12T U507 ( .A1(n1731), .A2(n1732), .A3(n1733), .ZN(n1734) );
  ND3D1BWP12T U508 ( .A1(n343), .A2(n342), .A3(n341), .ZN(n344) );
  NR2D1BWP12T U509 ( .A1(n1729), .A2(n1728), .ZN(n1735) );
  NR2D2BWP12T U510 ( .A1(n973), .A2(n972), .ZN(n974) );
  AN4XD1BWP12T U511 ( .A1(n3566), .A2(n3565), .A3(n3564), .A4(n3563), .Z(n3579) );
  AN2D1BWP12T U512 ( .A1(n1599), .A2(n1598), .Z(n1607) );
  CKND2D2BWP12T U513 ( .A1(n1935), .A2(n1934), .ZN(n1938) );
  AO222D0BWP12T U514 ( .A1(n3241), .A2(n2936), .B1(r7[9]), .B2(n3242), .C1(
        n3243), .C2(n2937), .Z(n2402) );
  MOAI22D0BWP12T U515 ( .A1(n845), .A2(n844), .B1(n845), .B2(n844), .ZN(n48)
         );
  AOI22D0BWP12T U516 ( .A1(pc_out[11]), .A2(n2989), .B1(next_pc_in[11]), .B2(
        n3398), .ZN(n49) );
  OAI21D1BWP12T U517 ( .A1(n3394), .A2(n48), .B(n49), .ZN(n2180) );
  AO222D0BWP12T U518 ( .A1(n3627), .A2(write1_in[1]), .B1(r10[1]), .B2(n3297), 
        .C1(n3298), .C2(n892), .Z(n2298) );
  AO222D0BWP12T U519 ( .A1(n3248), .A2(write1_in[15]), .B1(r9[15]), .B2(n3249), 
        .C1(n3250), .C2(n843), .Z(n2344) );
  AO222D0BWP12T U520 ( .A1(n3626), .A2(write1_in[12]), .B1(r11[12]), .B2(n3306), .C1(n3307), .C2(n727), .Z(n2277) );
  AO222D0BWP12T U521 ( .A1(n3638), .A2(write1_in[3]), .B1(tmp1[3]), .B2(n3276), 
        .C1(n3277), .C2(n2913), .Z(n2140) );
  AO222D0BWP12T U522 ( .A1(n3638), .A2(write1_in[11]), .B1(tmp1[11]), .B2(
        n3276), .C1(n3277), .C2(n2971), .Z(n2148) );
  AO222D0BWP12T U523 ( .A1(n3638), .A2(write1_in[14]), .B1(tmp1[14]), .B2(
        n3276), .C1(n3277), .C2(n2973), .Z(n2151) );
  CKND0BWP12T U524 ( .I(n866), .ZN(n50) );
  AOI21D0BWP12T U525 ( .A1(n[3692]), .A2(n3230), .B(reset), .ZN(n51) );
  CKND2D0BWP12T U526 ( .A1(n3229), .A2(write1_in[8]), .ZN(n52) );
  OAI211D1BWP12T U527 ( .A1(n2938), .A2(n50), .B(n51), .C(n52), .ZN(spin[8])
         );
  AO222D0BWP12T U528 ( .A1(n3234), .A2(write1_in[5]), .B1(lr[5]), .B2(n3235), 
        .C1(n3236), .C2(n2900), .Z(n2206) );
  AO222D0BWP12T U529 ( .A1(n3234), .A2(n2920), .B1(lr[6]), .B2(n3235), .C1(
        n3236), .C2(n2921), .Z(n2207) );
  AO222D0BWP12T U530 ( .A1(n3628), .A2(write1_in[13]), .B1(r6[13]), .B2(n3262), 
        .C1(n3263), .C2(n2972), .Z(n2438) );
  AO222D0BWP12T U531 ( .A1(n3289), .A2(write1_in[16]), .B1(r1[16]), .B2(n3290), 
        .C1(n3291), .C2(write2_in[16]), .Z(n2601) );
  AO222D0BWP12T U532 ( .A1(n3284), .A2(n782), .B1(r0[0]), .B2(n3285), .C1(
        write2_in[0]), .C2(n3286), .Z(n2617) );
  AOI22D0BWP12T U533 ( .A1(r4[2]), .A2(n2953), .B1(r8[2]), .B2(n2954), .ZN(n53) );
  AOI22D0BWP12T U534 ( .A1(n[3698]), .A2(n2956), .B1(r10[2]), .B2(n2955), .ZN(
        n54) );
  AOI22D0BWP12T U535 ( .A1(r2[2]), .A2(n2964), .B1(r3[2]), .B2(n2965), .ZN(n55) );
  AOI22D0BWP12T U536 ( .A1(pc_out[2]), .A2(n2966), .B1(r0[2]), .B2(n2967), 
        .ZN(n56) );
  OAI211D0BWP12T U537 ( .A1(n2088), .A2(n2968), .B(n55), .C(n56), .ZN(n57) );
  AOI22D0BWP12T U538 ( .A1(lr[2]), .A2(n2960), .B1(r9[2]), .B2(n2959), .ZN(n58) );
  AOI22D0BWP12T U539 ( .A1(r7[2]), .A2(n2958), .B1(r5[2]), .B2(n2957), .ZN(n59) );
  AOI22D0BWP12T U540 ( .A1(r11[2]), .A2(n2961), .B1(r6[2]), .B2(n2962), .ZN(
        n60) );
  ND3D0BWP12T U541 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n61) );
  AOI211D0BWP12T U542 ( .A1(r12[2]), .A2(n2963), .B(n57), .C(n61), .ZN(n62) );
  CKND0BWP12T U543 ( .I(n2970), .ZN(n63) );
  AOI31D0BWP12T U544 ( .A1(n53), .A2(n54), .A3(n62), .B(n63), .ZN(regD_out[2])
         );
  AO222D0BWP12T U545 ( .A1(n3623), .A2(n2936), .B1(r4[9]), .B2(n3280), .C1(
        n3281), .C2(n2937), .Z(n2498) );
  ND2D1BWP12T U546 ( .A1(n665), .A2(n664), .ZN(n64) );
  AOI22D0BWP12T U547 ( .A1(next_pc_in[15]), .A2(n3398), .B1(n2989), .B2(
        pc_out[15]), .ZN(n66) );
  AO222D0BWP12T U548 ( .A1(write1_in[15]), .A2(n3638), .B1(tmp1[15]), .B2(
        n3276), .C1(n3277), .C2(n843), .Z(n2152) );
  CKND0BWP12T U549 ( .I(n2924), .ZN(n67) );
  NR2D0BWP12T U550 ( .A1(n2915), .A2(n3399), .ZN(n68) );
  AOI211D0BWP12T U551 ( .A1(next_pc_in[1]), .A2(n3398), .B(n68), .C(reset), 
        .ZN(n69) );
  OAI21D1BWP12T U552 ( .A1(n2914), .A2(n67), .B(n69), .ZN(n2170) );
  CKND0BWP12T U553 ( .I(n2971), .ZN(n70) );
  AOI21D0BWP12T U554 ( .A1(n[3689]), .A2(n3230), .B(reset), .ZN(n71) );
  CKND2D0BWP12T U555 ( .A1(n3229), .A2(write1_in[11]), .ZN(n72) );
  OAI211D1BWP12T U556 ( .A1(n2938), .A2(n70), .B(n71), .C(n72), .ZN(spin[11])
         );
  AO222D0BWP12T U557 ( .A1(n3229), .A2(write1_in[14]), .B1(n[3686]), .B2(n3230), .C1(n3231), .C2(n2973), .Z(spin[14]) );
  AO222D0BWP12T U558 ( .A1(n3234), .A2(write1_in[2]), .B1(lr[2]), .B2(n3235), 
        .C1(n3236), .C2(n2882), .Z(n2203) );
  AO222D0BWP12T U559 ( .A1(n3234), .A2(write1_in[3]), .B1(lr[3]), .B2(n3235), 
        .C1(n3236), .C2(n2913), .Z(n2204) );
  AO222D0BWP12T U560 ( .A1(n3234), .A2(write1_in[8]), .B1(lr[8]), .B2(n3235), 
        .C1(n3236), .C2(n866), .Z(n2209) );
  AO222D0BWP12T U561 ( .A1(n3216), .A2(write1_in[5]), .B1(r12[5]), .B2(n3217), 
        .C1(n3218), .C2(n2900), .Z(n2238) );
  AO222D0BWP12T U562 ( .A1(n3216), .A2(n2920), .B1(r12[6]), .B2(n3217), .C1(
        n3218), .C2(n2921), .Z(n2239) );
  AO222D0BWP12T U563 ( .A1(n3626), .A2(write1_in[10]), .B1(r11[10]), .B2(n3306), .C1(n3307), .C2(n2951), .Z(n2275) );
  AO222D0BWP12T U564 ( .A1(write1_in[4]), .A2(n3622), .B1(r5[4]), .B2(n3272), 
        .C1(n3273), .C2(n2887), .Z(n2461) );
  AO222D0BWP12T U565 ( .A1(n3289), .A2(write1_in[17]), .B1(r1[17]), .B2(n3290), 
        .C1(n3291), .C2(write2_in[17]), .Z(n2602) );
  AOI22D0BWP12T U566 ( .A1(r4[12]), .A2(n2953), .B1(r8[12]), .B2(n2954), .ZN(
        n73) );
  AOI22D0BWP12T U567 ( .A1(r10[12]), .A2(n2955), .B1(n[3688]), .B2(n2956), 
        .ZN(n74) );
  AOI22D0BWP12T U568 ( .A1(r3[12]), .A2(n2965), .B1(r2[12]), .B2(n2964), .ZN(
        n75) );
  AOI22D0BWP12T U569 ( .A1(pc_out[12]), .A2(n2966), .B1(r0[12]), .B2(n2967), 
        .ZN(n76) );
  OAI211D0BWP12T U570 ( .A1(n2952), .A2(n2968), .B(n75), .C(n76), .ZN(n77) );
  AOI22D0BWP12T U571 ( .A1(r9[12]), .A2(n2959), .B1(lr[12]), .B2(n2960), .ZN(
        n78) );
  AOI22D0BWP12T U572 ( .A1(r7[12]), .A2(n2958), .B1(r5[12]), .B2(n2957), .ZN(
        n79) );
  AOI22D0BWP12T U573 ( .A1(r6[12]), .A2(n2962), .B1(r11[12]), .B2(n2961), .ZN(
        n80) );
  ND3D0BWP12T U574 ( .A1(n78), .A2(n79), .A3(n80), .ZN(n81) );
  AOI211D0BWP12T U575 ( .A1(r12[12]), .A2(n2963), .B(n77), .C(n81), .ZN(n82)
         );
  CKND0BWP12T U576 ( .I(n2970), .ZN(n83) );
  AOI31D0BWP12T U577 ( .A1(n73), .A2(n74), .A3(n82), .B(n83), .ZN(regD_out[12]) );
  AO222D0BWP12T U578 ( .A1(n3248), .A2(n2936), .B1(r9[9]), .B2(n3249), .C1(
        n3250), .C2(n2937), .Z(n2338) );
  AO222D0BWP12T U579 ( .A1(n3626), .A2(write1_in[1]), .B1(r11[1]), .B2(n3306), 
        .C1(n3307), .C2(n892), .Z(n2266) );
  AO222D0BWP12T U580 ( .A1(n3638), .A2(write1_in[12]), .B1(tmp1[12]), .B2(
        n3276), .C1(n3277), .C2(n727), .Z(n2149) );
  MOAI22D0BWP12T U581 ( .A1(n729), .A2(n728), .B1(n729), .B2(n728), .ZN(n84)
         );
  AOI22D0BWP12T U582 ( .A1(n3398), .A2(next_pc_in[6]), .B1(pc_out[6]), .B2(
        n2989), .ZN(n85) );
  OAI21D1BWP12T U583 ( .A1(n3394), .A2(n84), .B(n85), .ZN(n2175) );
  AO222D0BWP12T U584 ( .A1(n3229), .A2(write1_in[15]), .B1(n[3685]), .B2(n3230), .C1(n3231), .C2(n843), .Z(spin[15]) );
  AO222D0BWP12T U585 ( .A1(n3234), .A2(write1_in[14]), .B1(lr[14]), .B2(n3235), 
        .C1(n3236), .C2(n2973), .Z(n2215) );
  AO222D0BWP12T U586 ( .A1(n3216), .A2(write1_in[2]), .B1(r12[2]), .B2(n3217), 
        .C1(n3218), .C2(n2882), .Z(n2235) );
  AO222D0BWP12T U587 ( .A1(n3216), .A2(write1_in[3]), .B1(r12[3]), .B2(n3217), 
        .C1(n3218), .C2(n2913), .Z(n2236) );
  AO222D0BWP12T U588 ( .A1(n3216), .A2(write1_in[8]), .B1(r12[8]), .B2(n3217), 
        .C1(n3218), .C2(n866), .Z(n2241) );
  AO222D0BWP12T U589 ( .A1(n3626), .A2(write1_in[5]), .B1(r11[5]), .B2(n3306), 
        .C1(n3307), .C2(n2900), .Z(n2270) );
  AO222D0BWP12T U590 ( .A1(n3627), .A2(write1_in[10]), .B1(r10[10]), .B2(n3297), .C1(n3298), .C2(n2951), .Z(n2307) );
  AO222D0BWP12T U591 ( .A1(n3622), .A2(write1_in[13]), .B1(r5[13]), .B2(n3272), 
        .C1(n3273), .C2(n2972), .Z(n2470) );
  AO222D0BWP12T U592 ( .A1(n3289), .A2(write1_in[18]), .B1(r1[18]), .B2(n3290), 
        .C1(n3291), .C2(write2_in[18]), .Z(n2603) );
  AOI22D0BWP12T U593 ( .A1(r4[11]), .A2(n2953), .B1(r8[11]), .B2(n2954), .ZN(
        n86) );
  AOI22D0BWP12T U594 ( .A1(n[3689]), .A2(n2956), .B1(r10[11]), .B2(n2955), 
        .ZN(n87) );
  AOI22D0BWP12T U595 ( .A1(r3[11]), .A2(n2965), .B1(r2[11]), .B2(n2964), .ZN(
        n88) );
  AOI22D0BWP12T U596 ( .A1(pc_out[11]), .A2(n2966), .B1(r0[11]), .B2(n2967), 
        .ZN(n89) );
  OAI211D0BWP12T U597 ( .A1(n2969), .A2(n2968), .B(n88), .C(n89), .ZN(n90) );
  AOI22D0BWP12T U598 ( .A1(r9[11]), .A2(n2959), .B1(lr[11]), .B2(n2960), .ZN(
        n91) );
  AOI22D0BWP12T U599 ( .A1(r5[11]), .A2(n2957), .B1(r7[11]), .B2(n2958), .ZN(
        n92) );
  AOI22D0BWP12T U600 ( .A1(r11[11]), .A2(n2961), .B1(r6[11]), .B2(n2962), .ZN(
        n93) );
  ND3D0BWP12T U601 ( .A1(n91), .A2(n92), .A3(n93), .ZN(n94) );
  AOI211D0BWP12T U602 ( .A1(r12[11]), .A2(n2963), .B(n90), .C(n94), .ZN(n95)
         );
  CKND0BWP12T U603 ( .I(n2970), .ZN(n96) );
  AOI31D0BWP12T U604 ( .A1(n86), .A2(n87), .A3(n95), .B(n96), .ZN(regD_out[11]) );
  MOAI22D0BWP12T U605 ( .A1(n733), .A2(n732), .B1(n733), .B2(n732), .ZN(n97)
         );
  AOI22D0BWP12T U606 ( .A1(pc_out[5]), .A2(n2989), .B1(next_pc_in[5]), .B2(
        n3398), .ZN(n98) );
  OAI21D1BWP12T U607 ( .A1(n3394), .A2(n97), .B(n98), .ZN(n2174) );
  AO222D0BWP12T U608 ( .A1(n3289), .A2(write1_in[12]), .B1(r1[12]), .B2(n3290), 
        .C1(n3291), .C2(n727), .Z(n2597) );
  AO222D0BWP12T U609 ( .A1(n3638), .A2(n2936), .B1(tmp1[9]), .B2(n3276), .C1(
        n3277), .C2(n2937), .Z(n2146) );
  CKND2D0BWP12T U610 ( .A1(n844), .A2(n845), .ZN(n99) );
  AOI22D0BWP12T U611 ( .A1(pc_out[12]), .A2(n2989), .B1(next_pc_in[12]), .B2(
        n3398), .ZN(n101) );
  OAI21D1BWP12T U612 ( .A1(n3394), .A2(n100), .B(n101), .ZN(n2181) );
  AO222D0BWP12T U613 ( .A1(n3234), .A2(write1_in[1]), .B1(lr[1]), .B2(n3235), 
        .C1(n3236), .C2(n892), .Z(n2202) );
  AO222D0BWP12T U614 ( .A1(n3234), .A2(write1_in[11]), .B1(lr[11]), .B2(n3235), 
        .C1(n3236), .C2(n2971), .Z(n2212) );
  AO222D0BWP12T U615 ( .A1(n3234), .A2(write1_in[15]), .B1(lr[15]), .B2(n3235), 
        .C1(n3236), .C2(n843), .Z(n2216) );
  AO222D0BWP12T U616 ( .A1(n3216), .A2(write1_in[14]), .B1(r12[14]), .B2(n3217), .C1(n3218), .C2(n2973), .Z(n2247) );
  AO222D0BWP12T U617 ( .A1(n3626), .A2(write1_in[2]), .B1(r11[2]), .B2(n3306), 
        .C1(n3307), .C2(n2882), .Z(n2267) );
  AO222D0BWP12T U618 ( .A1(n3626), .A2(write1_in[3]), .B1(r11[3]), .B2(n3306), 
        .C1(n3307), .C2(n2913), .Z(n2268) );
  AO222D0BWP12T U619 ( .A1(n3626), .A2(n2920), .B1(r11[6]), .B2(n3306), .C1(
        n3307), .C2(n2921), .Z(n2271) );
  AO222D0BWP12T U620 ( .A1(n3626), .A2(write1_in[8]), .B1(r11[8]), .B2(n3306), 
        .C1(n3307), .C2(n866), .Z(n2273) );
  AO222D0BWP12T U621 ( .A1(write1_in[4]), .A2(n3623), .B1(r4[4]), .B2(n3280), 
        .C1(n3281), .C2(n2887), .Z(n2493) );
  AO222D0BWP12T U622 ( .A1(n3289), .A2(write1_in[19]), .B1(r1[19]), .B2(n3290), 
        .C1(n3291), .C2(write2_in[19]), .Z(n2604) );
  AOI22D0BWP12T U623 ( .A1(r4[10]), .A2(n2953), .B1(r8[10]), .B2(n2954), .ZN(
        n102) );
  AOI22D0BWP12T U624 ( .A1(n[3690]), .A2(n2956), .B1(r10[10]), .B2(n2955), 
        .ZN(n103) );
  AOI22D0BWP12T U625 ( .A1(r2[10]), .A2(n2964), .B1(r3[10]), .B2(n2965), .ZN(
        n104) );
  AOI22D0BWP12T U626 ( .A1(pc_out[10]), .A2(n2966), .B1(r0[10]), .B2(n2967), 
        .ZN(n105) );
  OAI211D0BWP12T U627 ( .A1(n2931), .A2(n2968), .B(n104), .C(n105), .ZN(n106)
         );
  AOI22D0BWP12T U628 ( .A1(r9[10]), .A2(n2959), .B1(lr[10]), .B2(n2960), .ZN(
        n107) );
  AOI22D0BWP12T U629 ( .A1(r7[10]), .A2(n2958), .B1(r5[10]), .B2(n2957), .ZN(
        n108) );
  AOI22D0BWP12T U630 ( .A1(r11[10]), .A2(n2961), .B1(r6[10]), .B2(n2962), .ZN(
        n109) );
  ND3D0BWP12T U631 ( .A1(n107), .A2(n108), .A3(n109), .ZN(n110) );
  AOI211D0BWP12T U632 ( .A1(r12[10]), .A2(n2963), .B(n106), .C(n110), .ZN(n111) );
  CKND0BWP12T U633 ( .I(n2970), .ZN(n112) );
  AOI31D0BWP12T U634 ( .A1(n102), .A2(n103), .A3(n111), .B(n112), .ZN(
        regD_out[10]) );
  CKND0BWP12T U635 ( .I(n727), .ZN(n113) );
  AOI21D0BWP12T U636 ( .A1(n[3688]), .A2(n3230), .B(reset), .ZN(n114) );
  CKND2D0BWP12T U637 ( .A1(n3229), .A2(write1_in[12]), .ZN(n115) );
  OAI211D1BWP12T U638 ( .A1(n2938), .A2(n113), .B(n114), .C(n115), .ZN(
        spin[12]) );
  AO222D0BWP12T U639 ( .A1(n3216), .A2(write1_in[11]), .B1(r12[11]), .B2(n3217), .C1(n3218), .C2(n2971), .Z(n2244) );
  AO222D0BWP12T U640 ( .A1(n3216), .A2(write1_in[15]), .B1(r12[15]), .B2(n3217), .C1(n3218), .C2(n843), .Z(n2248) );
  AO222D0BWP12T U641 ( .A1(n3626), .A2(write1_in[14]), .B1(r11[14]), .B2(n3306), .C1(n3307), .C2(n2973), .Z(n2279) );
  AO222D0BWP12T U642 ( .A1(n3627), .A2(write1_in[2]), .B1(r10[2]), .B2(n3297), 
        .C1(n3298), .C2(n2882), .Z(n2299) );
  AO222D0BWP12T U643 ( .A1(n3627), .A2(write1_in[3]), .B1(r10[3]), .B2(n3297), 
        .C1(n3298), .C2(n2913), .Z(n2300) );
  AO222D0BWP12T U644 ( .A1(n3627), .A2(write1_in[5]), .B1(r10[5]), .B2(n3297), 
        .C1(n3298), .C2(n2900), .Z(n2302) );
  AO222D0BWP12T U645 ( .A1(n3627), .A2(n2920), .B1(r10[6]), .B2(n3297), .C1(
        n3298), .C2(n2921), .Z(n2303) );
  AO222D0BWP12T U646 ( .A1(n3627), .A2(write1_in[8]), .B1(r10[8]), .B2(n3297), 
        .C1(n3298), .C2(n866), .Z(n2305) );
  AO222D0BWP12T U647 ( .A1(n3248), .A2(write1_in[1]), .B1(r9[1]), .B2(n3249), 
        .C1(n3250), .C2(n892), .Z(n2330) );
  AO222D0BWP12T U648 ( .A1(n3248), .A2(write1_in[10]), .B1(r9[10]), .B2(n3249), 
        .C1(n3250), .C2(n2951), .Z(n2339) );
  AO222D0BWP12T U649 ( .A1(n3289), .A2(n3051), .B1(r1[20]), .B2(n3290), .C1(
        n3291), .C2(write2_in[20]), .Z(n2605) );
  AOI22D0BWP12T U650 ( .A1(r8[9]), .A2(n2954), .B1(r4[9]), .B2(n2953), .ZN(
        n116) );
  AOI22D0BWP12T U651 ( .A1(r10[9]), .A2(n2955), .B1(n[3691]), .B2(n2956), .ZN(
        n117) );
  AOI22D0BWP12T U652 ( .A1(r3[9]), .A2(n2965), .B1(r2[9]), .B2(n2964), .ZN(
        n118) );
  AOI22D0BWP12T U653 ( .A1(pc_out[9]), .A2(n2966), .B1(r0[9]), .B2(n2967), 
        .ZN(n119) );
  OAI211D0BWP12T U654 ( .A1(n2923), .A2(n2968), .B(n118), .C(n119), .ZN(n120)
         );
  AOI22D0BWP12T U655 ( .A1(lr[9]), .A2(n2960), .B1(r9[9]), .B2(n2959), .ZN(
        n121) );
  AOI22D0BWP12T U656 ( .A1(r5[9]), .A2(n2957), .B1(r7[9]), .B2(n2958), .ZN(
        n122) );
  AOI22D0BWP12T U657 ( .A1(r11[9]), .A2(n2961), .B1(r6[9]), .B2(n2962), .ZN(
        n123) );
  ND3D0BWP12T U658 ( .A1(n121), .A2(n122), .A3(n123), .ZN(n124) );
  AOI211D0BWP12T U659 ( .A1(r12[9]), .A2(n2963), .B(n120), .C(n124), .ZN(n125)
         );
  CKND0BWP12T U660 ( .I(n2970), .ZN(n126) );
  AOI31D0BWP12T U661 ( .A1(n116), .A2(n117), .A3(n125), .B(n126), .ZN(
        regD_out[9]) );
  MOAI22D0BWP12T U662 ( .A1(n2930), .A2(n2929), .B1(n2930), .B2(n2929), .ZN(
        n127) );
  AOI22D0BWP12T U663 ( .A1(pc_out[3]), .A2(n2989), .B1(next_pc_in[3]), .B2(
        n3398), .ZN(n128) );
  OAI21D1BWP12T U664 ( .A1(n3394), .A2(n127), .B(n128), .ZN(n2172) );
  MOAI22D0BWP12T U665 ( .A1(n665), .A2(n664), .B1(n665), .B2(n664), .ZN(n129)
         );
  AOI22D0BWP12T U666 ( .A1(n3398), .A2(next_pc_in[14]), .B1(pc_out[14]), .B2(
        n2989), .ZN(n130) );
  OAI21D1BWP12T U667 ( .A1(n129), .A2(n3394), .B(n130), .ZN(n2183) );
  AO222D0BWP12T U668 ( .A1(n3234), .A2(n2936), .B1(lr[9]), .B2(n3235), .C1(
        n3236), .C2(n2937), .Z(n2210) );
  AO222D0BWP12T U669 ( .A1(n3234), .A2(write1_in[12]), .B1(lr[12]), .B2(n3235), 
        .C1(n3236), .C2(n727), .Z(n2213) );
  AO222D0BWP12T U670 ( .A1(n3626), .A2(write1_in[11]), .B1(r11[11]), .B2(n3306), .C1(n3307), .C2(n2971), .Z(n2276) );
  AO222D0BWP12T U671 ( .A1(n3626), .A2(write1_in[15]), .B1(r11[15]), .B2(n3306), .C1(n3307), .C2(n843), .Z(n2280) );
  AO222D0BWP12T U672 ( .A1(n3627), .A2(write1_in[14]), .B1(r10[14]), .B2(n3297), .C1(n3298), .C2(n2973), .Z(n2311) );
  AO222D0BWP12T U673 ( .A1(n3248), .A2(write1_in[2]), .B1(r9[2]), .B2(n3249), 
        .C1(n3250), .C2(n2882), .Z(n2331) );
  AO222D0BWP12T U674 ( .A1(n3248), .A2(write1_in[5]), .B1(r9[5]), .B2(n3249), 
        .C1(n3250), .C2(n2900), .Z(n2334) );
  AO222D0BWP12T U675 ( .A1(n3248), .A2(n2920), .B1(r9[6]), .B2(n3249), .C1(
        n3250), .C2(n2921), .Z(n2335) );
  AO222D0BWP12T U676 ( .A1(n3211), .A2(write1_in[1]), .B1(r8[1]), .B2(n3212), 
        .C1(n3213), .C2(n892), .Z(n2362) );
  AO222D0BWP12T U677 ( .A1(n3211), .A2(write1_in[10]), .B1(r8[10]), .B2(n3212), 
        .C1(n3213), .C2(n2951), .Z(n2371) );
  AO222D0BWP12T U678 ( .A1(n3623), .A2(write1_in[13]), .B1(r4[13]), .B2(n3280), 
        .C1(n3281), .C2(n2972), .Z(n2502) );
  AO222D0BWP12T U679 ( .A1(n3289), .A2(write1_in[21]), .B1(r1[21]), .B2(n3290), 
        .C1(n3291), .C2(write2_in[21]), .Z(n2606) );
  AOI22D0BWP12T U680 ( .A1(r4[8]), .A2(n2953), .B1(r8[8]), .B2(n2954), .ZN(
        n131) );
  AOI22D0BWP12T U681 ( .A1(r10[8]), .A2(n2955), .B1(n[3692]), .B2(n2956), .ZN(
        n132) );
  AOI22D0BWP12T U682 ( .A1(r3[8]), .A2(n2965), .B1(r2[8]), .B2(n2964), .ZN(
        n133) );
  AOI22D0BWP12T U683 ( .A1(pc_out[8]), .A2(n2966), .B1(r0[8]), .B2(n2967), 
        .ZN(n134) );
  OAI211D0BWP12T U684 ( .A1(n2928), .A2(n2968), .B(n133), .C(n134), .ZN(n135)
         );
  AOI22D0BWP12T U685 ( .A1(r9[8]), .A2(n2959), .B1(lr[8]), .B2(n2960), .ZN(
        n136) );
  AOI22D0BWP12T U686 ( .A1(r5[8]), .A2(n2957), .B1(r7[8]), .B2(n2958), .ZN(
        n137) );
  AOI22D0BWP12T U687 ( .A1(r11[8]), .A2(n2961), .B1(r6[8]), .B2(n2962), .ZN(
        n138) );
  ND3D0BWP12T U688 ( .A1(n136), .A2(n137), .A3(n138), .ZN(n139) );
  AOI211D0BWP12T U689 ( .A1(r12[8]), .A2(n2963), .B(n135), .C(n139), .ZN(n140)
         );
  CKND0BWP12T U690 ( .I(n2970), .ZN(n141) );
  AOI31D0BWP12T U691 ( .A1(n131), .A2(n132), .A3(n140), .B(n141), .ZN(
        regD_out[8]) );
  CKND0BWP12T U692 ( .I(r7[21]), .ZN(n142) );
  TPOAI22D1BWP12T U693 ( .A1(n3487), .A2(n142), .B1(n3486), .B2(n1559), .ZN(
        n1565) );
  MAOI22D0BWP12T U694 ( .A1(next_pc_in[26]), .A2(n3398), .B1(n3646), .B2(n3399), .ZN(n3341) );
  AO222D0BWP12T U695 ( .A1(n3216), .A2(n2936), .B1(r12[9]), .B2(n3217), .C1(
        n3218), .C2(n2937), .Z(n2242) );
  AO222D0BWP12T U696 ( .A1(n3216), .A2(write1_in[12]), .B1(r12[12]), .B2(n3217), .C1(n3218), .C2(n727), .Z(n2245) );
  AO222D0BWP12T U697 ( .A1(n3627), .A2(write1_in[11]), .B1(r10[11]), .B2(n3297), .C1(n3298), .C2(n2971), .Z(n2308) );
  AO222D0BWP12T U698 ( .A1(n3627), .A2(write1_in[15]), .B1(r10[15]), .B2(n3297), .C1(n3298), .C2(n843), .Z(n2312) );
  AO222D0BWP12T U699 ( .A1(n3248), .A2(write1_in[3]), .B1(r9[3]), .B2(n3249), 
        .C1(n3250), .C2(n2913), .Z(n2332) );
  AO222D0BWP12T U700 ( .A1(n3248), .A2(write1_in[8]), .B1(r9[8]), .B2(n3249), 
        .C1(n3250), .C2(n866), .Z(n2337) );
  AO222D0BWP12T U701 ( .A1(n3248), .A2(write1_in[14]), .B1(r9[14]), .B2(n3249), 
        .C1(n3250), .C2(n2973), .Z(n2343) );
  AO222D0BWP12T U702 ( .A1(n3211), .A2(write1_in[5]), .B1(r8[5]), .B2(n3212), 
        .C1(n3213), .C2(n2900), .Z(n2366) );
  AO222D0BWP12T U703 ( .A1(n3211), .A2(n2920), .B1(r8[6]), .B2(n3212), .C1(
        n3213), .C2(n2921), .Z(n2367) );
  AO222D0BWP12T U704 ( .A1(n3241), .A2(write1_in[1]), .B1(r7[1]), .B2(n3242), 
        .C1(n3243), .C2(n892), .Z(n2394) );
  AO222D0BWP12T U705 ( .A1(n3289), .A2(write1_in[22]), .B1(r1[22]), .B2(n3290), 
        .C1(n3291), .C2(write2_in[22]), .Z(n2607) );
  MOAI22D0BWP12T U706 ( .A1(n3645), .A2(n3399), .B1(next_pc_in[25]), .B2(n3398), .ZN(n3330) );
  AO222D0BWP12T U707 ( .A1(n3626), .A2(n2936), .B1(r11[9]), .B2(n3306), .C1(
        n3307), .C2(n2937), .Z(n2274) );
  AO222D0BWP12T U708 ( .A1(n3627), .A2(write1_in[12]), .B1(r10[12]), .B2(n3297), .C1(n3298), .C2(n727), .Z(n2309) );
  AO222D0BWP12T U709 ( .A1(n3248), .A2(write1_in[11]), .B1(r9[11]), .B2(n3249), 
        .C1(n3250), .C2(n2971), .Z(n2340) );
  AO222D0BWP12T U710 ( .A1(n3211), .A2(write1_in[3]), .B1(r8[3]), .B2(n3212), 
        .C1(n3213), .C2(n2913), .Z(n2364) );
  AO222D0BWP12T U711 ( .A1(n3211), .A2(write1_in[8]), .B1(r8[8]), .B2(n3212), 
        .C1(n3213), .C2(n866), .Z(n2369) );
  AO222D0BWP12T U712 ( .A1(n3211), .A2(write1_in[14]), .B1(r8[14]), .B2(n3212), 
        .C1(n3213), .C2(n2973), .Z(n2375) );
  AO222D0BWP12T U713 ( .A1(n3211), .A2(write1_in[15]), .B1(r8[15]), .B2(n3212), 
        .C1(n3213), .C2(n843), .Z(n2376) );
  AO222D0BWP12T U714 ( .A1(n3241), .A2(write1_in[5]), .B1(r7[5]), .B2(n3242), 
        .C1(n3243), .C2(n2900), .Z(n2398) );
  AO222D0BWP12T U715 ( .A1(n3241), .A2(n2920), .B1(r7[6]), .B2(n3242), .C1(
        n3243), .C2(n2921), .Z(n2399) );
  AO222D0BWP12T U716 ( .A1(n3628), .A2(write1_in[1]), .B1(r6[1]), .B2(n3262), 
        .C1(n3263), .C2(n892), .Z(n2426) );
  AO222D0BWP12T U717 ( .A1(n3624), .A2(write1_in[4]), .B1(n3028), .B2(n2887), 
        .C1(r3[4]), .C2(n3303), .Z(n2525) );
  AO222D0BWP12T U718 ( .A1(n3289), .A2(write1_in[24]), .B1(r1[24]), .B2(n3290), 
        .C1(n3291), .C2(write2_in[24]), .Z(n2609) );
  AOI22D0BWP12T U719 ( .A1(r4[7]), .A2(n2953), .B1(r8[7]), .B2(n2954), .ZN(
        n143) );
  AOI22D0BWP12T U720 ( .A1(r10[7]), .A2(n2955), .B1(n[3693]), .B2(n2956), .ZN(
        n144) );
  AOI22D0BWP12T U721 ( .A1(r3[7]), .A2(n2965), .B1(r2[7]), .B2(n2964), .ZN(
        n145) );
  AOI22D0BWP12T U722 ( .A1(pc_out[7]), .A2(n2966), .B1(r0[7]), .B2(n2967), 
        .ZN(n146) );
  OAI211D0BWP12T U723 ( .A1(n2922), .A2(n2968), .B(n145), .C(n146), .ZN(n147)
         );
  AOI22D0BWP12T U724 ( .A1(r9[7]), .A2(n2959), .B1(lr[7]), .B2(n2960), .ZN(
        n148) );
  AOI22D0BWP12T U725 ( .A1(r5[7]), .A2(n2957), .B1(r7[7]), .B2(n2958), .ZN(
        n149) );
  AOI22D0BWP12T U726 ( .A1(r6[7]), .A2(n2962), .B1(r11[7]), .B2(n2961), .ZN(
        n150) );
  ND3D0BWP12T U727 ( .A1(n148), .A2(n149), .A3(n150), .ZN(n151) );
  AOI211D0BWP12T U728 ( .A1(r12[7]), .A2(n2963), .B(n147), .C(n151), .ZN(n152)
         );
  CKND0BWP12T U729 ( .I(n2970), .ZN(n153) );
  AOI31D0BWP12T U730 ( .A1(n143), .A2(n144), .A3(n152), .B(n153), .ZN(
        regD_out[7]) );
  AOI21D0BWP12T U731 ( .A1(n[3699]), .A2(n3230), .B(reset), .ZN(n154) );
  CKND2D0BWP12T U732 ( .A1(n3229), .A2(write1_in[1]), .ZN(n155) );
  OAI211D0BWP12T U733 ( .A1(n891), .A2(n2938), .B(n154), .C(n155), .ZN(spin[1]) );
  AO222D0BWP12T U734 ( .A1(n3627), .A2(n2936), .B1(r10[9]), .B2(n3297), .C1(
        n3298), .C2(n2937), .Z(n2306) );
  AO222D0BWP12T U735 ( .A1(n3248), .A2(write1_in[12]), .B1(r9[12]), .B2(n3249), 
        .C1(n3250), .C2(n727), .Z(n2341) );
  AO222D0BWP12T U736 ( .A1(n3211), .A2(write1_in[2]), .B1(r8[2]), .B2(n3212), 
        .C1(n3213), .C2(n2882), .Z(n2363) );
  AO222D0BWP12T U737 ( .A1(n3241), .A2(write1_in[3]), .B1(r7[3]), .B2(n3242), 
        .C1(n3243), .C2(n2913), .Z(n2396) );
  AO222D0BWP12T U738 ( .A1(n3241), .A2(write1_in[8]), .B1(r7[8]), .B2(n3242), 
        .C1(n3243), .C2(n866), .Z(n2401) );
  AO222D0BWP12T U739 ( .A1(n3241), .A2(write1_in[10]), .B1(r7[10]), .B2(n3242), 
        .C1(n3243), .C2(n2951), .Z(n2403) );
  AO222D0BWP12T U740 ( .A1(n3241), .A2(write1_in[11]), .B1(r7[11]), .B2(n3242), 
        .C1(n3243), .C2(n2971), .Z(n2404) );
  AO222D0BWP12T U741 ( .A1(n3241), .A2(write1_in[14]), .B1(r7[14]), .B2(n3242), 
        .C1(n3243), .C2(n2973), .Z(n2407) );
  AO222D0BWP12T U742 ( .A1(n3241), .A2(write1_in[15]), .B1(r7[15]), .B2(n3242), 
        .C1(n3243), .C2(n843), .Z(n2408) );
  AO222D0BWP12T U743 ( .A1(n3628), .A2(write1_in[5]), .B1(r6[5]), .B2(n3262), 
        .C1(n3263), .C2(n2900), .Z(n2430) );
  AO222D0BWP12T U744 ( .A1(n3628), .A2(n2920), .B1(r6[6]), .B2(n3262), .C1(
        n3263), .C2(n2921), .Z(n2431) );
  AO222D0BWP12T U745 ( .A1(n3284), .A2(write1_in[16]), .B1(r0[16]), .B2(n3285), 
        .C1(n3286), .C2(write2_in[16]), .Z(n2633) );
  AOI22D0BWP12T U746 ( .A1(r4[4]), .A2(n2953), .B1(r8[4]), .B2(n2954), .ZN(
        n156) );
  AOI22D0BWP12T U747 ( .A1(n[3696]), .A2(n2956), .B1(r10[4]), .B2(n2955), .ZN(
        n157) );
  AOI22D0BWP12T U748 ( .A1(r2[4]), .A2(n2964), .B1(r3[4]), .B2(n2965), .ZN(
        n158) );
  AOI22D0BWP12T U749 ( .A1(pc_out[4]), .A2(n2966), .B1(r0[4]), .B2(n2967), 
        .ZN(n159) );
  OAI211D0BWP12T U750 ( .A1(n2778), .A2(n2968), .B(n158), .C(n159), .ZN(n160)
         );
  AOI22D0BWP12T U751 ( .A1(r9[4]), .A2(n2959), .B1(lr[4]), .B2(n2960), .ZN(
        n161) );
  AOI22D0BWP12T U752 ( .A1(r7[4]), .A2(n2958), .B1(r5[4]), .B2(n2957), .ZN(
        n162) );
  AOI22D0BWP12T U753 ( .A1(r11[4]), .A2(n2961), .B1(r6[4]), .B2(n2962), .ZN(
        n163) );
  ND3D0BWP12T U754 ( .A1(n161), .A2(n162), .A3(n163), .ZN(n164) );
  AOI211D0BWP12T U755 ( .A1(r12[4]), .A2(n2963), .B(n160), .C(n164), .ZN(n165)
         );
  CKND0BWP12T U756 ( .I(n2970), .ZN(n166) );
  AOI31D0BWP12T U757 ( .A1(n156), .A2(n157), .A3(n165), .B(n166), .ZN(
        regD_out[4]) );
  MAOI22D0BWP12T U758 ( .A1(next_pc_in[29]), .A2(n3398), .B1(n3650), .B2(n3399), .ZN(n167) );
  MOAI22D0BWP12T U759 ( .A1(n2943), .A2(n2944), .B1(n2944), .B2(n2943), .ZN(
        n168) );
  AOI22D0BWP12T U760 ( .A1(n2989), .A2(pc_out[4]), .B1(next_pc_in[4]), .B2(
        n3398), .ZN(n169) );
  OAI21D1BWP12T U761 ( .A1(n3394), .A2(n168), .B(n169), .ZN(n2173) );
  AO222D0BWP12T U762 ( .A1(n3211), .A2(n2936), .B1(r8[9]), .B2(n3212), .C1(
        n3213), .C2(n2937), .Z(n2370) );
  AO222D0BWP12T U763 ( .A1(n3211), .A2(write1_in[12]), .B1(r8[12]), .B2(n3212), 
        .C1(n3213), .C2(n727), .Z(n2373) );
  AO222D0BWP12T U764 ( .A1(n3241), .A2(write1_in[2]), .B1(r7[2]), .B2(n3242), 
        .C1(n3243), .C2(n2882), .Z(n2395) );
  AO222D0BWP12T U765 ( .A1(n3628), .A2(write1_in[3]), .B1(r6[3]), .B2(n3262), 
        .C1(n3263), .C2(n2913), .Z(n2428) );
  AO222D0BWP12T U766 ( .A1(n3628), .A2(write1_in[8]), .B1(r6[8]), .B2(n3262), 
        .C1(n3263), .C2(n866), .Z(n2433) );
  AO222D0BWP12T U767 ( .A1(n3628), .A2(write1_in[10]), .B1(r6[10]), .B2(n3262), 
        .C1(n3263), .C2(n2951), .Z(n2435) );
  AO222D0BWP12T U768 ( .A1(n3628), .A2(write1_in[11]), .B1(r6[11]), .B2(n3262), 
        .C1(n3263), .C2(n2971), .Z(n2436) );
  AO222D0BWP12T U769 ( .A1(n3628), .A2(write1_in[14]), .B1(r6[14]), .B2(n3262), 
        .C1(n3263), .C2(n2973), .Z(n2439) );
  AO222D0BWP12T U770 ( .A1(write1_in[15]), .A2(n3628), .B1(r6[15]), .B2(n3262), 
        .C1(n3263), .C2(n843), .Z(n2440) );
  AO222D0BWP12T U771 ( .A1(n3622), .A2(write1_in[1]), .B1(r5[1]), .B2(n3272), 
        .C1(n3273), .C2(n892), .Z(n2458) );
  AO222D0BWP12T U772 ( .A1(n3622), .A2(n2920), .B1(r5[6]), .B2(n3272), .C1(
        n3273), .C2(n2921), .Z(n2463) );
  AO222D0BWP12T U773 ( .A1(n3624), .A2(write1_in[13]), .B1(r3[13]), .B2(n3303), 
        .C1(n3028), .C2(n2972), .Z(n2534) );
  AO222D0BWP12T U774 ( .A1(n3284), .A2(write1_in[17]), .B1(r0[17]), .B2(n3285), 
        .C1(n3286), .C2(write2_in[17]), .Z(n2634) );
  CKND0BWP12T U775 ( .I(pc_out[16]), .ZN(n170) );
  CKND0BWP12T U776 ( .I(r6[16]), .ZN(n171) );
  OAI22D1BWP12T U777 ( .A1(n3612), .A2(n170), .B1(n3611), .B2(n171), .ZN(n1065) );
  MOAI22D0BWP12T U778 ( .A1(n3647), .A2(n3399), .B1(next_pc_in[27]), .B2(n3398), .ZN(n1862) );
  AO222D0BWP12T U779 ( .A1(n3241), .A2(write1_in[12]), .B1(r7[12]), .B2(n3242), 
        .C1(n3243), .C2(n727), .Z(n2405) );
  AO222D0BWP12T U780 ( .A1(n3628), .A2(write1_in[2]), .B1(r6[2]), .B2(n3262), 
        .C1(n3263), .C2(n2882), .Z(n2427) );
  AO222D0BWP12T U781 ( .A1(n3628), .A2(n2936), .B1(r6[9]), .B2(n3262), .C1(
        n3263), .C2(n2937), .Z(n2434) );
  AO222D0BWP12T U782 ( .A1(n3622), .A2(write1_in[3]), .B1(r5[3]), .B2(n3272), 
        .C1(n3273), .C2(n2913), .Z(n2460) );
  AO222D0BWP12T U783 ( .A1(n3622), .A2(write1_in[5]), .B1(r5[5]), .B2(n3272), 
        .C1(n3273), .C2(n2900), .Z(n2462) );
  AO222D0BWP12T U784 ( .A1(n3622), .A2(write1_in[8]), .B1(r5[8]), .B2(n3272), 
        .C1(n3273), .C2(n866), .Z(n2465) );
  AO222D0BWP12T U785 ( .A1(n3622), .A2(write1_in[10]), .B1(r5[10]), .B2(n3272), 
        .C1(n3273), .C2(n2951), .Z(n2467) );
  AO222D0BWP12T U786 ( .A1(n3622), .A2(write1_in[11]), .B1(r5[11]), .B2(n3272), 
        .C1(n3273), .C2(n2971), .Z(n2468) );
  AO222D0BWP12T U787 ( .A1(n3622), .A2(write1_in[14]), .B1(r5[14]), .B2(n3272), 
        .C1(n3273), .C2(n2973), .Z(n2471) );
  AO222D0BWP12T U788 ( .A1(n3622), .A2(write1_in[15]), .B1(r5[15]), .B2(n3272), 
        .C1(n3273), .C2(n843), .Z(n2472) );
  AO222D0BWP12T U789 ( .A1(n3623), .A2(write1_in[1]), .B1(r4[1]), .B2(n3280), 
        .C1(n3281), .C2(n892), .Z(n2490) );
  AO222D0BWP12T U790 ( .A1(n3623), .A2(n2920), .B1(r4[6]), .B2(n3280), .C1(
        n3281), .C2(n2921), .Z(n2495) );
  AO222D0BWP12T U791 ( .A1(n3625), .A2(write1_in[4]), .B1(n2887), .B2(n3374), 
        .C1(r2[4]), .C2(n3373), .Z(n2557) );
  AO222D0BWP12T U792 ( .A1(n3284), .A2(write1_in[7]), .B1(r0[7]), .B2(n3285), 
        .C1(n3286), .C2(write2_in[7]), .Z(n2624) );
  AO222D0BWP12T U793 ( .A1(n3284), .A2(write1_in[18]), .B1(r0[18]), .B2(n3285), 
        .C1(n3286), .C2(write2_in[18]), .Z(n2635) );
  NR2D0BWP12T U794 ( .A1(write2_sel[2]), .A2(n529), .ZN(n172) );
  AOI211D1BWP12T U795 ( .A1(n531), .A2(n172), .B(n530), .C(reset), .ZN(n3306)
         );
  MOAI22D0BWP12T U796 ( .A1(n731), .A2(n730), .B1(n731), .B2(n730), .ZN(n173)
         );
  AOI22D0BWP12T U797 ( .A1(n2989), .A2(pc_out[7]), .B1(next_pc_in[7]), .B2(
        n3398), .ZN(n174) );
  OAI21D1BWP12T U798 ( .A1(n3394), .A2(n173), .B(n174), .ZN(n2176) );
  AO222D0BWP12T U799 ( .A1(n3628), .A2(write1_in[12]), .B1(r6[12]), .B2(n3262), 
        .C1(n3263), .C2(n727), .Z(n2437) );
  AO222D0BWP12T U800 ( .A1(n3622), .A2(write1_in[2]), .B1(r5[2]), .B2(n3272), 
        .C1(n3273), .C2(n2882), .Z(n2459) );
  AO222D0BWP12T U801 ( .A1(n3622), .A2(n2936), .B1(r5[9]), .B2(n3272), .C1(
        n3273), .C2(n2937), .Z(n2466) );
  AO222D0BWP12T U802 ( .A1(n3623), .A2(write1_in[3]), .B1(r4[3]), .B2(n3280), 
        .C1(n3281), .C2(n2913), .Z(n2492) );
  AO222D0BWP12T U803 ( .A1(n3623), .A2(write1_in[5]), .B1(r4[5]), .B2(n3280), 
        .C1(n3281), .C2(n2900), .Z(n2494) );
  AO222D0BWP12T U804 ( .A1(n3623), .A2(write1_in[8]), .B1(r4[8]), .B2(n3280), 
        .C1(n3281), .C2(n866), .Z(n2497) );
  AO222D0BWP12T U805 ( .A1(n3623), .A2(write1_in[10]), .B1(r4[10]), .B2(n3280), 
        .C1(n3281), .C2(n2951), .Z(n2499) );
  AO222D0BWP12T U806 ( .A1(n3623), .A2(write1_in[11]), .B1(r4[11]), .B2(n3280), 
        .C1(n3281), .C2(n2971), .Z(n2500) );
  AO222D0BWP12T U807 ( .A1(n3623), .A2(write1_in[14]), .B1(r4[14]), .B2(n3280), 
        .C1(n3281), .C2(n2973), .Z(n2503) );
  AO222D0BWP12T U808 ( .A1(n3623), .A2(write1_in[15]), .B1(r4[15]), .B2(n3280), 
        .C1(n3281), .C2(n843), .Z(n2504) );
  AO222D0BWP12T U809 ( .A1(n3624), .A2(write1_in[1]), .B1(n3028), .B2(n892), 
        .C1(r3[1]), .C2(n3303), .Z(n2522) );
  AO222D0BWP12T U810 ( .A1(n3624), .A2(n2920), .B1(n3028), .B2(n2921), .C1(
        r3[6]), .C2(n3303), .Z(n2527) );
  AO222D0BWP12T U811 ( .A1(n3625), .A2(write1_in[13]), .B1(r2[13]), .B2(n3373), 
        .C1(n3374), .C2(n2972), .Z(n2566) );
  AO222D0BWP12T U812 ( .A1(n3284), .A2(write1_in[19]), .B1(r0[19]), .B2(n3285), 
        .C1(n3286), .C2(write2_in[19]), .Z(n2636) );
  OAI22D0BWP12T U813 ( .A1(n3603), .A2(n3425), .B1(n1738), .B2(n3435), .ZN(
        n175) );
  OAI22D1BWP12T U814 ( .A1(n3611), .A2(n3424), .B1(n3612), .B2(n3647), .ZN(
        n176) );
  NR4D0BWP12T U815 ( .A1(n806), .A2(n805), .A3(n175), .A4(n176), .ZN(n807) );
  CKND0BWP12T U816 ( .I(r7[25]), .ZN(n177) );
  OAI22D1BWP12T U817 ( .A1(n3487), .A2(n177), .B1(n3486), .B2(n3645), .ZN(
        n1016) );
  MOAI22D0BWP12T U818 ( .A1(n3667), .A2(n3399), .B1(next_pc_in[31]), .B2(n3398), .ZN(n3400) );
  INR2D0BWP12T U819 ( .A1(n504), .B1(n505), .ZN(n3249) );
  INR2D0BWP12T U820 ( .A1(n586), .B1(n587), .ZN(n3272) );
  MOAI22D0BWP12T U821 ( .A1(n568), .A2(n567), .B1(n568), .B2(n567), .ZN(n178)
         );
  AOI22D0BWP12T U822 ( .A1(pc_out[13]), .A2(n2989), .B1(n3398), .B2(
        next_pc_in[13]), .ZN(n179) );
  OAI21D1BWP12T U823 ( .A1(n3394), .A2(n178), .B(n179), .ZN(n2182) );
  AO222D0BWP12T U824 ( .A1(n3622), .A2(write1_in[12]), .B1(r5[12]), .B2(n3272), 
        .C1(n3273), .C2(n727), .Z(n2469) );
  AO222D0BWP12T U825 ( .A1(n3623), .A2(write1_in[2]), .B1(r4[2]), .B2(n3280), 
        .C1(n3281), .C2(n2882), .Z(n2491) );
  AO222D0BWP12T U826 ( .A1(n3624), .A2(write1_in[3]), .B1(n3028), .B2(n2913), 
        .C1(r3[3]), .C2(n3303), .Z(n2524) );
  AO222D0BWP12T U827 ( .A1(n3624), .A2(write1_in[5]), .B1(n3028), .B2(n2900), 
        .C1(r3[5]), .C2(n3303), .Z(n2526) );
  AO222D0BWP12T U828 ( .A1(n3624), .A2(write1_in[8]), .B1(r3[8]), .B2(n3303), 
        .C1(n3028), .C2(n866), .Z(n2529) );
  AO222D0BWP12T U829 ( .A1(n3624), .A2(n2936), .B1(r3[9]), .B2(n3303), .C1(
        n3028), .C2(n2937), .Z(n2530) );
  AO222D0BWP12T U830 ( .A1(n3624), .A2(write1_in[10]), .B1(r3[10]), .B2(n3303), 
        .C1(n3028), .C2(n2951), .Z(n2531) );
  AO222D0BWP12T U831 ( .A1(n3624), .A2(write1_in[11]), .B1(r3[11]), .B2(n3303), 
        .C1(n3028), .C2(n2971), .Z(n2532) );
  AO222D0BWP12T U832 ( .A1(n3624), .A2(write1_in[14]), .B1(r3[14]), .B2(n3303), 
        .C1(n3028), .C2(n2973), .Z(n2535) );
  AO222D0BWP12T U833 ( .A1(n3624), .A2(write1_in[15]), .B1(r3[15]), .B2(n3303), 
        .C1(n3028), .C2(n843), .Z(n2536) );
  AO222D0BWP12T U834 ( .A1(n3625), .A2(write1_in[1]), .B1(n892), .B2(n3374), 
        .C1(r2[1]), .C2(n3373), .Z(n2554) );
  AO222D0BWP12T U835 ( .A1(n3289), .A2(write1_in[4]), .B1(r1[4]), .B2(n3290), 
        .C1(n3291), .C2(n2887), .Z(n2589) );
  AO222D0BWP12T U836 ( .A1(n3284), .A2(n3051), .B1(r0[20]), .B2(n3285), .C1(
        n3286), .C2(write2_in[20]), .Z(n2637) );
  AOI22D0BWP12T U837 ( .A1(r9[26]), .A2(n2871), .B1(r8[26]), .B2(n2873), .ZN(
        n180) );
  AOI22D0BWP12T U838 ( .A1(lr[26]), .A2(n2869), .B1(r12[26]), .B2(n2848), .ZN(
        n181) );
  AOI22D0BWP12T U839 ( .A1(r11[26]), .A2(n2870), .B1(r10[26]), .B2(n2872), 
        .ZN(n182) );
  AOI22D0BWP12T U840 ( .A1(r4[26]), .A2(n2853), .B1(r7[26]), .B2(n2854), .ZN(
        n183) );
  AOI22D0BWP12T U841 ( .A1(r6[26]), .A2(n2855), .B1(r2[26]), .B2(n2856), .ZN(
        n184) );
  AOI22D0BWP12T U842 ( .A1(r1[26]), .A2(n2857), .B1(r5[26]), .B2(n2757), .ZN(
        n185) );
  AOI22D0BWP12T U843 ( .A1(r0[26]), .A2(n2859), .B1(r3[26]), .B2(n2858), .ZN(
        n186) );
  ND4D0BWP12T U844 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(n187) );
  OAI22D0BWP12T U845 ( .A1(n2822), .A2(n3646), .B1(n1991), .B2(n2832), .ZN(
        n188) );
  AOI21D0BWP12T U846 ( .A1(n2864), .A2(n187), .B(n188), .ZN(n189) );
  ND4D0BWP12T U847 ( .A1(n180), .A2(n181), .A3(n182), .A4(n189), .ZN(
        regC_out[26]) );
  CKND0BWP12T U848 ( .I(pc_out[17]), .ZN(n190) );
  CKND0BWP12T U849 ( .I(r6[17]), .ZN(n191) );
  OAI22D1BWP12T U850 ( .A1(n3612), .A2(n190), .B1(n3611), .B2(n191), .ZN(n1885) );
  CKND0BWP12T U851 ( .I(r7[31]), .ZN(n192) );
  OAI22D0BWP12T U852 ( .A1(n3487), .A2(n192), .B1(n3486), .B2(n3667), .ZN(
        n3496) );
  NR4D0BWP12T U853 ( .A1(n1457), .A2(n1456), .A3(n1455), .A4(n1454), .ZN(n193)
         );
  TPND2D2BWP12T U854 ( .A1(n1458), .A2(n193), .ZN(regB_out[23]) );
  MOAI22D1BWP12T U855 ( .A1(n3488), .A2(n1393), .B1(r5[3]), .B2(n1942), .ZN(
        n369) );
  IND2D0BWP12T U856 ( .A1(write1_sel[3]), .B1(n456), .ZN(n463) );
  NR2D0BWP12T U857 ( .A1(write2_sel[0]), .A2(n552), .ZN(n194) );
  ND4D0BWP12T U858 ( .A1(write2_en), .A2(write2_sel[4]), .A3(write2_sel[3]), 
        .A4(n194), .ZN(n553) );
  MOAI22D0BWP12T U859 ( .A1(n3644), .A2(n3399), .B1(next_pc_in[24]), .B2(n3398), .ZN(n818) );
  INR3D0BWP12T U860 ( .A1(n522), .B1(n523), .B2(reset), .ZN(n3297) );
  INR2D0BWP12T U861 ( .A1(n486), .B1(n487), .ZN(n3212) );
  INR2D0BWP12T U862 ( .A1(n481), .B1(n482), .ZN(n3242) );
  INR2D0BWP12T U863 ( .A1(n459), .B1(n460), .ZN(n3280) );
  AO222D0BWP12T U864 ( .A1(n3638), .A2(write1_in[1]), .B1(tmp1[1]), .B2(n3276), 
        .C1(n3277), .C2(n892), .Z(n2138) );
  AOI22D0BWP12T U865 ( .A1(n3398), .A2(next_pc_in[16]), .B1(pc_out[16]), .B2(
        n2989), .ZN(n196) );
  OAI21D1BWP12T U866 ( .A1(n3394), .A2(n195), .B(n196), .ZN(n2185) );
  AO222D0BWP12T U867 ( .A1(n3623), .A2(write1_in[12]), .B1(r4[12]), .B2(n3280), 
        .C1(n3281), .C2(n727), .Z(n2501) );
  AO222D0BWP12T U868 ( .A1(n3625), .A2(write1_in[2]), .B1(n2882), .B2(n3374), 
        .C1(r2[2]), .C2(n3373), .Z(n2555) );
  AO222D0BWP12T U869 ( .A1(n3625), .A2(write1_in[5]), .B1(n2900), .B2(n3374), 
        .C1(r2[5]), .C2(n3373), .Z(n2558) );
  AO222D0BWP12T U870 ( .A1(n3625), .A2(n2920), .B1(n2921), .B2(n3374), .C1(
        r2[6]), .C2(n3373), .Z(n2559) );
  AO222D0BWP12T U871 ( .A1(n3625), .A2(write1_in[8]), .B1(r2[8]), .B2(n3373), 
        .C1(n3374), .C2(n866), .Z(n2561) );
  AO222D0BWP12T U872 ( .A1(n3625), .A2(n2936), .B1(r2[9]), .B2(n3373), .C1(
        n3374), .C2(n2937), .Z(n2562) );
  AO222D0BWP12T U873 ( .A1(n3625), .A2(write1_in[10]), .B1(r2[10]), .B2(n3373), 
        .C1(n3374), .C2(n2951), .Z(n2563) );
  AO222D0BWP12T U874 ( .A1(n3625), .A2(write1_in[11]), .B1(r2[11]), .B2(n3373), 
        .C1(n3374), .C2(n2971), .Z(n2564) );
  AO222D0BWP12T U875 ( .A1(n3625), .A2(write1_in[14]), .B1(r2[14]), .B2(n3373), 
        .C1(n3374), .C2(n2973), .Z(n2567) );
  AO222D0BWP12T U876 ( .A1(n3625), .A2(write1_in[15]), .B1(r2[15]), .B2(n3373), 
        .C1(n3374), .C2(n843), .Z(n2568) );
  AO222D0BWP12T U877 ( .A1(n3289), .A2(write1_in[13]), .B1(r1[13]), .B2(n3290), 
        .C1(n3291), .C2(n2972), .Z(n2598) );
  AO222D0BWP12T U878 ( .A1(n3284), .A2(write1_in[21]), .B1(r0[21]), .B2(n3285), 
        .C1(n3286), .C2(write2_in[21]), .Z(n2638) );
  AOI22D0BWP12T U879 ( .A1(r4[1]), .A2(n2853), .B1(r7[1]), .B2(n2854), .ZN(
        n197) );
  AOI22D0BWP12T U880 ( .A1(r6[1]), .A2(n2855), .B1(r2[1]), .B2(n2856), .ZN(
        n198) );
  AOI22D0BWP12T U881 ( .A1(r1[1]), .A2(n2857), .B1(r5[1]), .B2(n2757), .ZN(
        n199) );
  AOI22D0BWP12T U882 ( .A1(r0[1]), .A2(n2859), .B1(r3[1]), .B2(n2858), .ZN(
        n200) );
  ND4D0BWP12T U883 ( .A1(n197), .A2(n198), .A3(n199), .A4(n200), .ZN(n201) );
  OAI22D0BWP12T U884 ( .A1(n2819), .A2(n2830), .B1(n2820), .B2(n2846), .ZN(
        n202) );
  OAI22D0BWP12T U885 ( .A1(n2867), .A2(n2821), .B1(n2822), .B2(n2915), .ZN(
        n203) );
  AOI211D0BWP12T U886 ( .A1(n2864), .A2(n201), .B(n202), .C(n203), .ZN(n204)
         );
  AOI22D0BWP12T U887 ( .A1(n[3699]), .A2(n2875), .B1(r10[1]), .B2(n2872), .ZN(
        n205) );
  AOI22D0BWP12T U888 ( .A1(r11[1]), .A2(n2870), .B1(r9[1]), .B2(n2871), .ZN(
        n206) );
  ND3D0BWP12T U889 ( .A1(n204), .A2(n205), .A3(n206), .ZN(regC_out[1]) );
  CKND0BWP12T U890 ( .I(n[3684]), .ZN(n207) );
  CKND0BWP12T U891 ( .I(r8[16]), .ZN(n208) );
  TPOAI22D1BWP12T U892 ( .A1(n3605), .A2(n207), .B1(n3603), .B2(n208), .ZN(
        n1067) );
  AN4XD1BWP12T U893 ( .A1(n1817), .A2(n1818), .A3(n1819), .A4(n1820), .Z(n209)
         );
  TPND2D2BWP12T U894 ( .A1(n209), .A2(n210), .ZN(regB_out[28]) );
  OAI22D0BWP12T U895 ( .A1(n3588), .A2(n3446), .B1(n3586), .B2(n3460), .ZN(
        n211) );
  OAI22D1BWP12T U896 ( .A1(n3584), .A2(n1748), .B1(n3582), .B2(n3447), .ZN(
        n212) );
  TPNR2D1BWP12T U897 ( .A1(n211), .A2(n212), .ZN(n1751) );
  CKND0BWP12T U898 ( .I(r8[17]), .ZN(n213) );
  TPOAI22D1BWP12T U899 ( .A1(n3605), .A2(n2796), .B1(n3603), .B2(n213), .ZN(
        n1887) );
  CKND0BWP12T U900 ( .I(r5[31]), .ZN(n214) );
  OAI22D0BWP12T U901 ( .A1(n3489), .A2(n214), .B1(n3549), .B2(n3488), .ZN(
        n3495) );
  OAI22D1BWP12T U902 ( .A1(n3588), .A2(n1380), .B1(n3586), .B2(n1381), .ZN(
        n215) );
  TPOAI22D1BWP12T U903 ( .A1(n3584), .A2(n1379), .B1(n3582), .B2(n1378), .ZN(
        n216) );
  NR2D1BWP12T U904 ( .A1(n215), .A2(n216), .ZN(n1386) );
  OAI22D1BWP12T U905 ( .A1(n3584), .A2(n2038), .B1(n3582), .B2(n1071), .ZN(
        n218) );
  TPNR2D1BWP12T U906 ( .A1(n217), .A2(n218), .ZN(n1076) );
  IND2D0BWP12T U907 ( .A1(n3638), .B1(n3621), .ZN(n554) );
  INR3D0BWP12T U908 ( .A1(write1_sel[2]), .B1(write1_sel[1]), .B2(reset), .ZN(
        n475) );
  IND2D0BWP12T U909 ( .A1(n3216), .B1(n3621), .ZN(n453) );
  IND2D0BWP12T U910 ( .A1(n3284), .B1(n3621), .ZN(n499) );
  IAO21D0BWP12T U911 ( .A1(n528), .A2(n552), .B(n3381), .ZN(n2914) );
  INR2D1BWP12T U912 ( .A1(n476), .B1(n477), .ZN(n3230) );
  INR2D0BWP12T U913 ( .A1(n471), .B1(n472), .ZN(n3235) );
  INR2D0BWP12T U914 ( .A1(n540), .B1(n541), .ZN(n3374) );
  INR2D0BWP12T U915 ( .A1(n466), .B1(n467), .ZN(n3290) );
  AO222D0BWP12T U916 ( .A1(n3624), .A2(write1_in[12]), .B1(r3[12]), .B2(n3303), 
        .C1(n3028), .C2(n727), .Z(n2533) );
  AO222D0BWP12T U917 ( .A1(n3625), .A2(write1_in[3]), .B1(n2913), .B2(n3374), 
        .C1(r2[3]), .C2(n3373), .Z(n2556) );
  AO222D0BWP12T U918 ( .A1(n3289), .A2(write1_in[1]), .B1(r1[1]), .B2(n3290), 
        .C1(n3291), .C2(n892), .Z(n2586) );
  AO222D0BWP12T U919 ( .A1(n3289), .A2(write1_in[2]), .B1(r1[2]), .B2(n3290), 
        .C1(n3291), .C2(n2882), .Z(n2587) );
  AO222D0BWP12T U920 ( .A1(n3289), .A2(write1_in[5]), .B1(r1[5]), .B2(n3290), 
        .C1(n3291), .C2(n2900), .Z(n2590) );
  AO222D0BWP12T U921 ( .A1(n3289), .A2(n2920), .B1(r1[6]), .B2(n3290), .C1(
        n3291), .C2(n2921), .Z(n2591) );
  AO222D0BWP12T U922 ( .A1(n3289), .A2(write1_in[8]), .B1(r1[8]), .B2(n3290), 
        .C1(n3291), .C2(n866), .Z(n2593) );
  AO222D0BWP12T U923 ( .A1(n3289), .A2(n2936), .B1(r1[9]), .B2(n3290), .C1(
        n3291), .C2(n2937), .Z(n2594) );
  AO222D0BWP12T U924 ( .A1(n3289), .A2(write1_in[10]), .B1(r1[10]), .B2(n3290), 
        .C1(n3291), .C2(n2951), .Z(n2595) );
  AO222D0BWP12T U925 ( .A1(n3289), .A2(write1_in[11]), .B1(r1[11]), .B2(n3290), 
        .C1(n3291), .C2(n2971), .Z(n2596) );
  AO222D0BWP12T U926 ( .A1(n3289), .A2(write1_in[14]), .B1(r1[14]), .B2(n3290), 
        .C1(n3291), .C2(n2973), .Z(n2599) );
  AO222D0BWP12T U927 ( .A1(n3289), .A2(write1_in[15]), .B1(r1[15]), .B2(n3290), 
        .C1(n3291), .C2(n843), .Z(n2600) );
  AO222D0BWP12T U928 ( .A1(n3284), .A2(write1_in[4]), .B1(r0[4]), .B2(n3285), 
        .C1(n3286), .C2(n2887), .Z(n2621) );
  AO222D0BWP12T U929 ( .A1(n3284), .A2(write1_in[22]), .B1(r0[22]), .B2(n3285), 
        .C1(n3286), .C2(write2_in[22]), .Z(n2639) );
  CKND0BWP12T U930 ( .I(r1[16]), .ZN(n219) );
  OAI22D0BWP12T U931 ( .A1(n2866), .A2(n3600), .B1(n3599), .B2(n219), .ZN(
        n1068) );
  CKND0BWP12T U932 ( .I(r1[17]), .ZN(n220) );
  CKND0BWP12T U933 ( .I(r12[17]), .ZN(n221) );
  OAI22D0BWP12T U934 ( .A1(n3599), .A2(n220), .B1(n3600), .B2(n221), .ZN(n1888) );
  ND3D0BWP12T U935 ( .A1(n1659), .A2(n1658), .A3(n[3689]), .ZN(n1661) );
  AN2D0BWP12T U936 ( .A1(n1950), .A2(r7[2]), .Z(n1480) );
  MOAI22D0BWP12T U937 ( .A1(n3476), .A2(n3537), .B1(r4[31]), .B2(n3475), .ZN(
        n3484) );
  IND2D0BWP12T U938 ( .A1(n3229), .B1(n3621), .ZN(n477) );
  IND2D0BWP12T U939 ( .A1(n3234), .B1(n3621), .ZN(n472) );
  NR2D0BWP12T U940 ( .A1(write1_sel[4]), .A2(n549), .ZN(n521) );
  IND2D0BWP12T U941 ( .A1(n3248), .B1(n3621), .ZN(n505) );
  IND2D0BWP12T U942 ( .A1(n3211), .B1(n3621), .ZN(n487) );
  IND2D0BWP12T U943 ( .A1(n3622), .B1(n3621), .ZN(n587) );
  IND2D0BWP12T U944 ( .A1(n3623), .B1(n3621), .ZN(n460) );
  IND2D0BWP12T U945 ( .A1(n3289), .B1(n3621), .ZN(n467) );
  MOAI22D0BWP12T U946 ( .A1(n3314), .A2(n3399), .B1(next_pc_in[23]), .B2(n3398), .ZN(n3315) );
  INR2D0BWP12T U947 ( .A1(n553), .B1(n554), .ZN(n3276) );
  INR2D0BWP12T U948 ( .A1(n452), .B1(n453), .ZN(n3217) );
  INR2D0BWP12T U949 ( .A1(n493), .B1(n494), .ZN(n3262) );
  INR2D0BWP12T U950 ( .A1(n515), .B1(n516), .ZN(n3028) );
  INR2D0BWP12T U951 ( .A1(n498), .B1(n499), .ZN(n3285) );
  AO222D0BWP12T U952 ( .A1(n3284), .A2(write1_in[1]), .B1(r0[1]), .B2(n3285), 
        .C1(n3286), .C2(n892), .Z(n2618) );
  AO222D0BWP12T U953 ( .A1(n3284), .A2(write1_in[2]), .B1(r0[2]), .B2(n3285), 
        .C1(n3286), .C2(n2882), .Z(n2619) );
  AO222D0BWP12T U954 ( .A1(n3284), .A2(write1_in[3]), .B1(r0[3]), .B2(n3285), 
        .C1(n3286), .C2(n2913), .Z(n2620) );
  AO222D0BWP12T U955 ( .A1(n3284), .A2(write1_in[5]), .B1(r0[5]), .B2(n3285), 
        .C1(n3286), .C2(n2900), .Z(n2622) );
  AO222D0BWP12T U956 ( .A1(n3284), .A2(n2920), .B1(r0[6]), .B2(n3285), .C1(
        n3286), .C2(n2921), .Z(n2623) );
  AO222D0BWP12T U957 ( .A1(n3284), .A2(write1_in[8]), .B1(r0[8]), .B2(n3285), 
        .C1(n3286), .C2(n866), .Z(n2625) );
  AO222D0BWP12T U958 ( .A1(n3284), .A2(n2936), .B1(r0[9]), .B2(n3285), .C1(
        n3286), .C2(n2937), .Z(n2626) );
  AO222D0BWP12T U959 ( .A1(n3284), .A2(write1_in[10]), .B1(r0[10]), .B2(n3285), 
        .C1(n3286), .C2(n2951), .Z(n2627) );
  AO222D0BWP12T U960 ( .A1(n3284), .A2(write1_in[11]), .B1(r0[11]), .B2(n3285), 
        .C1(n3286), .C2(n2971), .Z(n2628) );
  AO222D0BWP12T U961 ( .A1(n3284), .A2(write1_in[12]), .B1(r0[12]), .B2(n3285), 
        .C1(n3286), .C2(n727), .Z(n2629) );
  AO222D0BWP12T U962 ( .A1(n3284), .A2(write1_in[13]), .B1(r0[13]), .B2(n3285), 
        .C1(n3286), .C2(n2972), .Z(n2630) );
  AO222D0BWP12T U963 ( .A1(n3284), .A2(write1_in[14]), .B1(r0[14]), .B2(n3285), 
        .C1(n3286), .C2(n2973), .Z(n2631) );
  AO222D0BWP12T U964 ( .A1(n3284), .A2(write1_in[15]), .B1(r0[15]), .B2(n3285), 
        .C1(n3286), .C2(n843), .Z(n2632) );
  AO222D0BWP12T U965 ( .A1(n3284), .A2(write1_in[24]), .B1(r0[24]), .B2(n3285), 
        .C1(n3286), .C2(write2_in[24]), .Z(n2641) );
  AOI22D0BWP12T U966 ( .A1(r10[4]), .A2(n2872), .B1(r8[4]), .B2(n2873), .ZN(
        n222) );
  AOI22D0BWP12T U967 ( .A1(r12[4]), .A2(n2848), .B1(n[3696]), .B2(n2875), .ZN(
        n223) );
  AOI22D0BWP12T U968 ( .A1(r11[4]), .A2(n2870), .B1(r9[4]), .B2(n2871), .ZN(
        n224) );
  AOI22D0BWP12T U969 ( .A1(r4[4]), .A2(n2853), .B1(r7[4]), .B2(n2854), .ZN(
        n225) );
  AOI22D0BWP12T U970 ( .A1(r6[4]), .A2(n2855), .B1(r2[4]), .B2(n2856), .ZN(
        n226) );
  AOI22D0BWP12T U971 ( .A1(r1[4]), .A2(n2857), .B1(r5[4]), .B2(n2757), .ZN(
        n227) );
  AOI22D0BWP12T U972 ( .A1(r0[4]), .A2(n2859), .B1(r3[4]), .B2(n2858), .ZN(
        n228) );
  ND4D0BWP12T U973 ( .A1(n225), .A2(n226), .A3(n227), .A4(n228), .ZN(n229) );
  OAI22D0BWP12T U974 ( .A1(n2822), .A2(n2818), .B1(n2846), .B2(n2817), .ZN(
        n230) );
  AOI21D0BWP12T U975 ( .A1(n2864), .A2(n229), .B(n230), .ZN(n231) );
  ND4D0BWP12T U976 ( .A1(n222), .A2(n223), .A3(n224), .A4(n231), .ZN(
        regC_out[4]) );
  MAOI22D1BWP12T U977 ( .A1(n3472), .A2(tmp1[15]), .B1(n1700), .B2(n1699), 
        .ZN(n1701) );
  RCOAI22D0BWP12T U978 ( .A1(n3481), .A2(n1438), .B1(n3479), .B2(n1216), .ZN(
        n1218) );
  TPOAI22D1BWP12T U979 ( .A1(n3489), .A2(n902), .B1(n3488), .B2(n1771), .ZN(
        n903) );
  IOA21D1BWP12T U980 ( .A1(n3474), .A2(r2[22]), .B(n1821), .ZN(n1829) );
  CKND2D2BWP12T U981 ( .A1(n3579), .A2(n3578), .ZN(regB_out[29]) );
  BUFFXD8BWP12T U982 ( .I(n1730), .Z(n3593) );
  BUFFXD8BWP12T U983 ( .I(n349), .Z(n3479) );
  TPND2D2BWP12T U984 ( .A1(n1261), .A2(n1260), .ZN(n1267) );
  INR2D8BWP12T U985 ( .A1(n1291), .B1(n339), .ZN(n235) );
  NR2XD1BWP12T U986 ( .A1(n3334), .A2(n3348), .ZN(n3339) );
  TPNR2D2BWP12T U987 ( .A1(n3383), .A2(n3382), .ZN(n3384) );
  NR4D1BWP12T U988 ( .A1(n380), .A2(n379), .A3(n378), .A4(n377), .ZN(n389) );
  TPND2D1BWP12T U989 ( .A1(n232), .A2(n3628), .ZN(n3247) );
  IOA21D1BWP12T U990 ( .A1(r2[19]), .A2(n3474), .B(n912), .ZN(n917) );
  IOA21D1BWP12T U991 ( .A1(n3474), .A2(r2[27]), .B(n3419), .ZN(n3430) );
  INVD9BWP12T U992 ( .I(n1700), .ZN(n3471) );
  CKND2D2BWP12T U993 ( .A1(write1_in[27]), .A2(n3381), .ZN(n445) );
  MOAI22D1BWP12T U994 ( .A1(n3487), .A2(n905), .B1(n6), .B2(pc_out[18]), .ZN(
        n907) );
  INVD4BWP12T U995 ( .I(n1945), .ZN(n3486) );
  INVD2BWP12T U996 ( .I(pc_out[18]), .ZN(n1774) );
  ND3D2BWP12T U997 ( .A1(n300), .A2(n299), .A3(n298), .ZN(n981) );
  BUFFXD12BWP12T U998 ( .I(write1_in[28]), .Z(n3294) );
  TPND2D2BWP12T U999 ( .A1(n845), .A2(n509), .ZN(n567) );
  DCCKND4BWP12T U1000 ( .I(readB_sel[3]), .ZN(n291) );
  ND2XD0BWP12T U1001 ( .A1(n1633), .A2(r8[3]), .ZN(n351) );
  TPNR2D3BWP12T U1002 ( .A1(readB_sel[0]), .A2(readB_sel[4]), .ZN(n257) );
  TPND2D1BWP12T U1003 ( .A1(n1924), .A2(r8[12]), .ZN(n1929) );
  BUFFXD8BWP12T U1004 ( .I(n1633), .Z(n1924) );
  INVD1BWP12T U1005 ( .I(n1470), .ZN(n234) );
  INR2D4BWP12T U1006 ( .A1(n1291), .B1(n339), .ZN(n375) );
  NR2XD1BWP12T U1007 ( .A1(n1858), .A2(n3340), .ZN(n1859) );
  CKND2D2BWP12T U1008 ( .A1(n1005), .A2(n1004), .ZN(regA_out[29]) );
  ND2XD0BWP12T U1009 ( .A1(n1653), .A2(lr[12]), .ZN(n1930) );
  INR2D2BWP12T U1010 ( .A1(r10[1]), .B1(n3479), .ZN(n1245) );
  TPNR3D2BWP12T U1011 ( .A1(n1302), .A2(n1301), .A3(n1300), .ZN(n1303) );
  TPOAI21D2BWP12T U1012 ( .A1(write1_in[29]), .A2(n3388), .B(n1128), .ZN(n1129) );
  RCAOI21D8BWP12T U1013 ( .A1(write1_in[23]), .A2(n3381), .B(n239), .ZN(n238)
         );
  INVD12BWP12T U1014 ( .I(n238), .ZN(n3310) );
  TPND2D2BWP12T U1015 ( .A1(n3202), .A2(n3201), .ZN(spin[31]) );
  ND2XD3BWP12T U1016 ( .A1(n1131), .A2(n3363), .ZN(n240) );
  AOI22D2BWP12T U1017 ( .A1(r12[10]), .A2(n1952), .B1(n1642), .B2(r6[10]), 
        .ZN(n318) );
  TPOAI22D1BWP12T U1018 ( .A1(n3448), .A2(n1703), .B1(n3476), .B2(n1702), .ZN(
        n1708) );
  INVD9BWP12T U1019 ( .I(n275), .ZN(n3592) );
  NR2XD1BWP12T U1020 ( .A1(n3387), .A2(n3386), .ZN(n3391) );
  NR2D1BWP12T U1021 ( .A1(n3401), .A2(n3394), .ZN(n1140) );
  CKND0BWP12T U1022 ( .I(write1_in[29]), .ZN(n241) );
  TPND2D2BWP12T U1023 ( .A1(n3210), .A2(n3209), .ZN(n2360) );
  TPND2D1BWP12T U1024 ( .A1(n3470), .A2(n3469), .ZN(regA_out[24]) );
  INVD4BWP12T U1025 ( .I(n261), .ZN(n242) );
  BUFFD2BWP12T U1026 ( .I(n1653), .Z(n1923) );
  TPND2D1BWP12T U1027 ( .A1(n243), .A2(n244), .ZN(n245) );
  CKND2D2BWP12T U1028 ( .A1(n245), .A2(n1239), .ZN(n1241) );
  INVD2BWP12T U1029 ( .I(n3448), .ZN(n243) );
  CKND0BWP12T U1030 ( .I(n1240), .ZN(n244) );
  DCCKND4BWP12T U1031 ( .I(readA_sel[3]), .ZN(n246) );
  INVD2BWP12T U1032 ( .I(r4[16]), .ZN(n1240) );
  TPND2D2BWP12T U1033 ( .A1(n235), .A2(r0[16]), .ZN(n1239) );
  TPAOI21D4BWP12T U1034 ( .A1(write1_in[20]), .A2(n1856), .B(n412), .ZN(n1973)
         );
  DCCKND4BWP12T U1035 ( .I(readA_sel[3]), .ZN(n1608) );
  TPOAI21D1BWP12T U1036 ( .A1(write1_in[29]), .A2(n3388), .B(n3365), .ZN(n3367) );
  TPAOI22D2BWP12T U1037 ( .A1(n1906), .A2(r2[15]), .B1(n3591), .B2(r10[15]), 
        .ZN(n794) );
  BUFFXD8BWP12T U1038 ( .I(n1642), .Z(n1926) );
  CKND2D2BWP12T U1039 ( .A1(write1_in[26]), .A2(write1_in[24]), .ZN(n1124) );
  BUFFXD3BWP12T U1040 ( .I(write1_in[26]), .Z(n247) );
  INVD2BWP12T U1041 ( .I(n3390), .ZN(n395) );
  CKND2D2BWP12T U1042 ( .A1(n3238), .A2(n3237), .ZN(n2229) );
  TPND2D2BWP12T U1043 ( .A1(n1040), .A2(n1039), .ZN(regB_out[10]) );
  TPND2D2BWP12T U1044 ( .A1(n1086), .A2(n1085), .ZN(regB_out[9]) );
  IND2D1BWP12T U1045 ( .A1(n1071), .B1(n3475), .ZN(n248) );
  DCCKND4BWP12T U1046 ( .I(r4[9]), .ZN(n1071) );
  DCCKBD4BWP12T U1047 ( .I(n981), .Z(n1913) );
  BUFFD2BWP12T U1048 ( .I(n981), .Z(n1740) );
  TPOAI22D1BWP12T U1049 ( .A1(n3478), .A2(n3609), .B1(n3477), .B2(n3602), .ZN(
        n915) );
  OAI21D1BWP12T U1050 ( .A1(n1666), .A2(n1665), .B(n1664), .ZN(n1667) );
  TPNR2D1BWP12T U1051 ( .A1(n1666), .A2(n1144), .ZN(n1150) );
  OR2XD1BWP12T U1052 ( .A1(n1666), .A2(n1280), .Z(n1281) );
  NR2XD1BWP12T U1053 ( .A1(n3348), .A2(n1867), .ZN(n1860) );
  XNR2D1BWP12T U1054 ( .A1(n3325), .A2(n3344), .ZN(n1460) );
  TPND2D1BWP12T U1055 ( .A1(n3369), .A2(n3368), .ZN(n3370) );
  INVD2BWP12T U1056 ( .I(n3369), .ZN(n3360) );
  DEL025D1BWP12T U1057 ( .I(write1_in[19]), .Z(n250) );
  ND2XD0BWP12T U1058 ( .A1(n3335), .A2(n3352), .ZN(n816) );
  TPND2D2BWP12T U1059 ( .A1(n3618), .A2(n3617), .ZN(regB_out[19]) );
  OR2D2BWP12T U1060 ( .A1(n270), .A2(n269), .Z(n271) );
  ND2XD4BWP12T U1061 ( .A1(n992), .A2(n991), .ZN(regB_out[0]) );
  TPNR2D3BWP12T U1062 ( .A1(n901), .A2(n900), .ZN(n911) );
  OAI21D2BWP12T U1063 ( .A1(n2038), .A2(n233), .B(n1299), .ZN(n1300) );
  INVD3BWP12T U1064 ( .I(readB_sel[0]), .ZN(n273) );
  INVD3BWP12T U1065 ( .I(readB_sel[0]), .ZN(n290) );
  TPAOI22D2BWP12T U1066 ( .A1(n3580), .A2(immediate2_in[5]), .B1(n295), .B2(
        tmp1[5]), .ZN(n1328) );
  ND3XD1BWP12T U1067 ( .A1(n3343), .A2(n3340), .A3(n3352), .ZN(n3337) );
  CKND0BWP12T U1068 ( .I(n1724), .ZN(n251) );
  INVD2BWP12T U1069 ( .I(r4[1]), .ZN(n1724) );
  TPNR2D3BWP12T U1070 ( .A1(readB_sel[1]), .A2(readB_sel[2]), .ZN(n286) );
  ND2XD4BWP12T U1071 ( .A1(n927), .A2(n926), .ZN(regA_out[19]) );
  NR4D3BWP12T U1072 ( .A1(n917), .A2(n916), .A3(n915), .A4(n914), .ZN(n927) );
  INR2D2BWP12T U1073 ( .A1(r10[3]), .B1(n3479), .ZN(n350) );
  NR4D0BWP12T U1074 ( .A1(n1778), .A2(n1777), .A3(n1776), .A4(n1775), .ZN(
        n1779) );
  TPND2D2BWP12T U1075 ( .A1(n1780), .A2(n1779), .ZN(regB_out[18]) );
  BUFFXD16BWP12T U1076 ( .I(n381), .Z(n3491) );
  AN2XD2BWP12T U1077 ( .A1(n1946), .A2(n[3697]), .Z(n362) );
  NR2D1BWP12T U1078 ( .A1(n800), .A2(n799), .ZN(n803) );
  ND3XD4BWP12T U1079 ( .A1(n1165), .A2(n1164), .A3(n1163), .ZN(regA_out[17])
         );
  NR4D3BWP12T U1080 ( .A1(n1150), .A2(n1149), .A3(n1148), .A4(n1147), .ZN(
        n1165) );
  ND2XD4BWP12T U1081 ( .A1(n320), .A2(readA_sel[0]), .ZN(n1290) );
  BUFFXD6BWP12T U1082 ( .I(n1394), .Z(n1884) );
  CKND2D2BWP12T U1083 ( .A1(n278), .A2(n1685), .ZN(n262) );
  INR2D4BWP12T U1084 ( .A1(n242), .B1(n792), .ZN(n1327) );
  IOA21D1BWP12T U1085 ( .A1(n3474), .A2(r2[26]), .B(n376), .ZN(n377) );
  AOI22D2BWP12T U1086 ( .A1(r9[26]), .A2(n3471), .B1(n3472), .B2(tmp1[26]), 
        .ZN(n376) );
  ND2XD8BWP12T U1087 ( .A1(n911), .A2(n910), .ZN(regA_out[18]) );
  NR4D1BWP12T U1088 ( .A1(n1011), .A2(n1010), .A3(n1009), .A4(n1008), .ZN(
        n1018) );
  OAI22D1BWP12T U1089 ( .A1(n3448), .A2(n3499), .B1(n3476), .B2(n3501), .ZN(
        n1010) );
  ND3D2BWP12T U1090 ( .A1(n446), .A2(n44), .A3(n1867), .ZN(n448) );
  INVD4BWP12T U1091 ( .I(n3668), .ZN(n253) );
  INVD8BWP12T U1092 ( .I(n253), .ZN(regB_out[27]) );
  TPAOI21D1BWP12T U1093 ( .A1(write1_in[30]), .A2(n3381), .B(n1134), .ZN(n3401) );
  INVD2BWP12T U1094 ( .I(readB_sel[4]), .ZN(n292) );
  INVD8BWP12T U1095 ( .I(n1951), .ZN(n3463) );
  ND2D3BWP12T U1096 ( .A1(n964), .A2(n963), .ZN(regA_out[0]) );
  TPND2D2BWP12T U1097 ( .A1(n808), .A2(n807), .ZN(n3668) );
  INR2D1BWP12T U1098 ( .A1(n502), .B1(n526), .ZN(n3248) );
  INVD1BWP12T U1099 ( .I(n3241), .ZN(n575) );
  INR2D1BWP12T U1100 ( .A1(n583), .B1(n550), .ZN(n3241) );
  INR2D1BWP12T U1101 ( .A1(n583), .B1(n582), .ZN(n3622) );
  INR2D1BWP12T U1102 ( .A1(n475), .B1(n526), .ZN(n3229) );
  INR2D1BWP12T U1103 ( .A1(n539), .B1(n582), .ZN(n3623) );
  INR2D1BWP12T U1104 ( .A1(n583), .B1(n497), .ZN(n3289) );
  INR2D1BWP12T U1105 ( .A1(n539), .B1(n497), .ZN(n3284) );
  NR2D1BWP12T U1106 ( .A1(n2914), .A2(reset), .ZN(n3352) );
  INR2D1BWP12T U1107 ( .A1(n521), .B1(n550), .ZN(n3234) );
  INR2D1BWP12T U1108 ( .A1(n502), .B1(n519), .ZN(n3211) );
  INR2D1BWP12T U1109 ( .A1(n551), .B1(n550), .ZN(n3638) );
  INR2D1BWP12T U1110 ( .A1(n521), .B1(n582), .ZN(n3216) );
  INR2D8BWP12T U1111 ( .A1(n294), .B1(n293), .ZN(n295) );
  AN2D1BWP12T U1112 ( .A1(n3471), .A2(r9[10]), .Z(n255) );
  INVD1BWP12T U1113 ( .I(n3352), .ZN(n3394) );
  INVD1BWP12T U1114 ( .I(n3381), .ZN(n3362) );
  INVD2BWP12T U1115 ( .I(r9[9]), .ZN(n2038) );
  INVD2BWP12T U1116 ( .I(r1[3]), .ZN(n2074) );
  INVD2BWP12T U1117 ( .I(r12[1]), .ZN(n2821) );
  INVD2BWP12T U1118 ( .I(r1[12]), .ZN(n2952) );
  INVD1BWP12T U1119 ( .I(reset), .ZN(n3621) );
  TPOAI22D1BWP12T U1120 ( .A1(n3586), .A2(n931), .B1(n3588), .B2(n930), .ZN(
        n932) );
  TPOAI22D1BWP12T U1121 ( .A1(n3612), .A2(n1034), .B1(n3611), .B2(n1033), .ZN(
        n1035) );
  OAI22D1BWP12T U1122 ( .A1(n3438), .A2(n3463), .B1(n3437), .B2(n3436), .ZN(
        n3439) );
  ND2XD4BWP12T U1123 ( .A1(n301), .A2(n286), .ZN(n1901) );
  TPNR3D4BWP12T U1124 ( .A1(readB_sel[4]), .A2(readB_sel[3]), .A3(readB_sel[0]), .ZN(n301) );
  TPNR3D3BWP12T U1125 ( .A1(n291), .A2(n273), .A3(readB_sel[4]), .ZN(n278) );
  INR2D4BWP12T U1126 ( .A1(readB_sel[2]), .B1(readB_sel[1]), .ZN(n280) );
  TPND2D2BWP12T U1127 ( .A1(n278), .A2(n280), .ZN(n1738) );
  INVD1BWP12T U1128 ( .I(n[3696]), .ZN(n260) );
  ND2XD3BWP12T U1129 ( .A1(n257), .A2(readB_sel[3]), .ZN(n276) );
  INVD1P75BWP12T U1130 ( .I(n286), .ZN(n258) );
  OR2XD4BWP12T U1131 ( .A1(n276), .A2(n258), .Z(n3603) );
  INVD1BWP12T U1132 ( .I(r8[4]), .ZN(n259) );
  OAI22D1BWP12T U1133 ( .A1(n1738), .A2(n260), .B1(n3603), .B2(n259), .ZN(n265) );
  ND2D3BWP12T U1134 ( .A1(readB_sel[1]), .A2(readB_sel[2]), .ZN(n261) );
  BUFFXD8BWP12T U1135 ( .I(n262), .Z(n3612) );
  INVD1BWP12T U1136 ( .I(pc_out[4]), .ZN(n2818) );
  TPND2D2BWP12T U1137 ( .A1(n301), .A2(n1685), .ZN(n1915) );
  BUFFD12BWP12T U1138 ( .I(n1915), .Z(n3611) );
  INVD1BWP12T U1139 ( .I(r6[4]), .ZN(n263) );
  OAI22D1BWP12T U1140 ( .A1(n3612), .A2(n2818), .B1(n3611), .B2(n263), .ZN(
        n264) );
  OR2XD2BWP12T U1141 ( .A1(n265), .A2(n264), .Z(n272) );
  INVD1BWP12T U1142 ( .I(r12[4]), .ZN(n1627) );
  INVD4BWP12T U1143 ( .I(n276), .ZN(n1689) );
  ND2XD4BWP12T U1144 ( .A1(n1689), .A2(n280), .ZN(n3600) );
  NR2XD2BWP12T U1145 ( .A1(readB_sel[3]), .A2(readB_sel[4]), .ZN(n299) );
  TPND2D1BWP12T U1146 ( .A1(n299), .A2(n286), .ZN(n266) );
  INR2D2BWP12T U1147 ( .A1(n298), .B1(n266), .ZN(n267) );
  INVD6BWP12T U1148 ( .I(n267), .ZN(n3599) );
  INVD1BWP12T U1149 ( .I(r1[4]), .ZN(n2778) );
  OAI22D1BWP12T U1150 ( .A1(n1627), .A2(n3600), .B1(n3599), .B2(n2778), .ZN(
        n270) );
  INVD1BWP12T U1151 ( .I(lr[4]), .ZN(n2817) );
  ND2D4BWP12T U1152 ( .A1(n1689), .A2(n242), .ZN(n1394) );
  BUFFXD3BWP12T U1153 ( .I(n1394), .Z(n3608) );
  DCCKND4BWP12T U1154 ( .I(readB_sel[1]), .ZN(n268) );
  TPNR2D3BWP12T U1155 ( .A1(n268), .A2(readB_sel[2]), .ZN(n300) );
  INVD1BWP12T U1156 ( .I(r3[4]), .ZN(n1629) );
  TPNR2D3BWP12T U1157 ( .A1(n272), .A2(n271), .ZN(n308) );
  TPNR3D1BWP12T U1158 ( .A1(n273), .A2(readB_sel[4]), .A3(readB_sel[3]), .ZN(
        n274) );
  INR2D2BWP12T U1159 ( .A1(n300), .B1(n276), .ZN(n277) );
  BUFFXD12BWP12T U1160 ( .I(n277), .Z(n3591) );
  ND2D2BWP12T U1161 ( .A1(n278), .A2(n286), .ZN(n279) );
  BUFFXD8BWP12T U1162 ( .I(n279), .Z(n3584) );
  INVD1BWP12T U1163 ( .I(r9[4]), .ZN(n283) );
  INVD1BWP12T U1164 ( .I(r4[4]), .ZN(n282) );
  TPOAI22D1BWP12T U1165 ( .A1(n3584), .A2(n283), .B1(n3582), .B2(n282), .ZN(
        n289) );
  INR3D4BWP12T U1166 ( .A1(readB_sel[3]), .B1(readB_sel[4]), .B2(n290), .ZN(
        n284) );
  ND2D3BWP12T U1167 ( .A1(n284), .A2(n300), .ZN(n285) );
  BUFFXD8BWP12T U1168 ( .I(n285), .Z(n3586) );
  INVD1BWP12T U1169 ( .I(r11[4]), .ZN(n1621) );
  INVD1BWP12T U1170 ( .I(r0[4]), .ZN(n287) );
  TPNR2D1BWP12T U1171 ( .A1(n289), .A2(n288), .ZN(n305) );
  DEL025D1BWP12T U1172 ( .I(n290), .Z(n294) );
  TPNR2D2BWP12T U1173 ( .A1(n292), .A2(n291), .ZN(n297) );
  TPND2D2BWP12T U1174 ( .A1(n297), .A2(n1685), .ZN(n293) );
  ND2XD4BWP12T U1175 ( .A1(n242), .A2(n298), .ZN(n296) );
  INR2D4BWP12T U1176 ( .A1(n242), .B1(n792), .ZN(n3524) );
  INVD4BWP12T U1177 ( .I(n302), .ZN(n1730) );
  AOI22D1BWP12T U1178 ( .A1(n3524), .A2(r7[4]), .B1(n1730), .B2(r2[4]), .ZN(
        n303) );
  AN4D4BWP12T U1179 ( .A1(n306), .A2(n305), .A3(n304), .A4(n303), .Z(n307) );
  ND2XD4BWP12T U1180 ( .A1(n308), .A2(n307), .ZN(regB_out[4]) );
  INVD8BWP12T U1181 ( .I(readA_sel[2]), .ZN(n309) );
  TPNR3D8BWP12T U1182 ( .A1(n1608), .A2(readA_sel[0]), .A3(readA_sel[4]), .ZN(
        n1285) );
  ND2D4BWP12T U1183 ( .A1(n328), .A2(n1285), .ZN(n349) );
  INR2D1BWP12T U1184 ( .A1(r10[10]), .B1(n3422), .ZN(n326) );
  ND2D8BWP12T U1185 ( .A1(readA_sel[2]), .A2(readA_sel[1]), .ZN(n1287) );
  INVD4BWP12T U1186 ( .I(n1287), .ZN(n1275) );
  ND2D3BWP12T U1187 ( .A1(n1275), .A2(n1285), .ZN(n310) );
  INVD6BWP12T U1188 ( .I(n310), .ZN(n1653) );
  INVD8BWP12T U1189 ( .I(readA_sel[1]), .ZN(n1610) );
  ND2D8BWP12T U1190 ( .A1(n1610), .A2(readA_sel[2]), .ZN(n340) );
  INVD8BWP12T U1191 ( .I(n340), .ZN(n317) );
  ND2XD8BWP12T U1192 ( .A1(n335), .A2(n246), .ZN(n315) );
  INVD8BWP12T U1193 ( .I(readA_sel[4]), .ZN(n1613) );
  INVD4BWP12T U1194 ( .I(n1613), .ZN(n314) );
  TPNR2D2BWP12T U1195 ( .A1(n315), .A2(n314), .ZN(n311) );
  INVD6BWP12T U1196 ( .I(n374), .ZN(n3475) );
  OR2XD16BWP12T U1197 ( .A1(n315), .A2(n314), .Z(n339) );
  INVD12BWP12T U1198 ( .I(n339), .ZN(n1934) );
  INVD6BWP12T U1199 ( .I(n316), .ZN(n1933) );
  ND2XD16BWP12T U1200 ( .A1(n1934), .A2(n1933), .ZN(n1666) );
  ND2D8BWP12T U1201 ( .A1(n317), .A2(n1285), .ZN(n1716) );
  INVD12BWP12T U1202 ( .I(n1716), .ZN(n1952) );
  TPNR2D8BWP12T U1203 ( .A1(n339), .A2(n1287), .ZN(n1642) );
  TPND2D2BWP12T U1204 ( .A1(n319), .A2(n318), .ZN(n324) );
  TPNR2D3BWP12T U1205 ( .A1(readA_sel[4]), .A2(readA_sel[3]), .ZN(n320) );
  TPNR2D8BWP12T U1206 ( .A1(readA_sel[1]), .A2(readA_sel[2]), .ZN(n1291) );
  INVD4BWP12T U1207 ( .I(n1291), .ZN(n321) );
  TPNR2D4BWP12T U1208 ( .A1(n1290), .A2(n321), .ZN(n1951) );
  INVD1BWP12T U1209 ( .I(r1[10]), .ZN(n2931) );
  OR2D4BWP12T U1210 ( .A1(n1290), .A2(n1287), .Z(n1414) );
  DCCKND12BWP12T U1211 ( .I(n1414), .ZN(n1950) );
  TPOAI21D2BWP12T U1212 ( .A1(n3463), .A2(n2931), .B(n322), .ZN(n323) );
  TPND2D3BWP12T U1213 ( .A1(n1291), .A2(n1285), .ZN(n327) );
  INVD6BWP12T U1214 ( .I(n327), .ZN(n1633) );
  BUFFXD16BWP12T U1215 ( .I(n1337), .Z(n3490) );
  INR2D2BWP12T U1216 ( .A1(r11[10]), .B1(n3490), .ZN(n333) );
  CKND3BWP12T U1217 ( .I(n1290), .ZN(n329) );
  BUFFXD12BWP12T U1218 ( .I(n1468), .Z(n3488) );
  INVD1BWP12T U1219 ( .I(r3[10]), .ZN(n1031) );
  TPNR2D2BWP12T U1220 ( .A1(n1290), .A2(n340), .ZN(n330) );
  ND2D1BWP12T U1221 ( .A1(n1942), .A2(r5[10]), .ZN(n331) );
  OAI21D1BWP12T U1222 ( .A1(n234), .A2(n1031), .B(n331), .ZN(n332) );
  INR3D2BWP12T U1223 ( .A1(n334), .B1(n333), .B2(n332), .ZN(n347) );
  ND3D2BWP12T U1224 ( .A1(readA_sel[3]), .A2(readA_sel[1]), .A3(readA_sel[4]), 
        .ZN(n337) );
  CKND2D2BWP12T U1225 ( .A1(n335), .A2(readA_sel[2]), .ZN(n336) );
  NR2D3BWP12T U1226 ( .A1(n337), .A2(n336), .ZN(n1156) );
  DCCKND8BWP12T U1227 ( .I(n1156), .ZN(n338) );
  ND2D1BWP12T U1228 ( .A1(n3472), .A2(tmp1[10]), .ZN(n345) );
  CKND2D0BWP12T U1229 ( .A1(n1945), .A2(pc_out[10]), .ZN(n342) );
  INVD4BWP12T U1230 ( .I(n340), .ZN(n1659) );
  ND2D8BWP12T U1231 ( .A1(n1658), .A2(n1659), .ZN(n381) );
  INVD8BWP12T U1232 ( .I(n381), .ZN(n1946) );
  INR3D2BWP12T U1233 ( .A1(n345), .B1(n255), .B2(n344), .ZN(n346) );
  TPAOI21D2BWP12T U1234 ( .A1(r6[3]), .A2(n1926), .B(n350), .ZN(n353) );
  ND2D1BWP12T U1235 ( .A1(n1653), .A2(lr[3]), .ZN(n352) );
  IOA21D2BWP12T U1236 ( .A1(n3475), .A2(r4[3]), .B(n354), .ZN(n359) );
  ND2D1BWP12T U1237 ( .A1(n3471), .A2(r9[3]), .ZN(n357) );
  ND2D1BWP12T U1238 ( .A1(n3472), .A2(tmp1[3]), .ZN(n355) );
  ND3D2BWP12T U1239 ( .A1(n357), .A2(n356), .A3(n355), .ZN(n358) );
  INR2D2BWP12T U1240 ( .A1(r11[3]), .B1(n3490), .ZN(n361) );
  TPNR2D2BWP12T U1241 ( .A1(n362), .A2(n361), .ZN(n370) );
  INVD1BWP12T U1242 ( .I(r3[3]), .ZN(n1393) );
  AN2XD2BWP12T U1243 ( .A1(n1952), .A2(r12[3]), .Z(n364) );
  INR2D2BWP12T U1244 ( .A1(r1[3]), .B1(n3463), .ZN(n363) );
  NR2D2BWP12T U1245 ( .A1(n364), .A2(n363), .ZN(n367) );
  ND2D1BWP12T U1246 ( .A1(n6), .A2(pc_out[3]), .ZN(n366) );
  ND2D1BWP12T U1247 ( .A1(n1950), .A2(r7[3]), .ZN(n365) );
  ND3D2BWP12T U1248 ( .A1(n367), .A2(n366), .A3(n365), .ZN(n368) );
  ND2XD8BWP12T U1249 ( .A1(n371), .A2(n372), .ZN(regA_out[3]) );
  INVD8BWP12T U1250 ( .I(n1642), .ZN(n3481) );
  INVD1BWP12T U1251 ( .I(r6[26]), .ZN(n1200) );
  INVD1BWP12T U1252 ( .I(r10[26]), .ZN(n373) );
  OAI22D0BWP12T U1253 ( .A1(n3481), .A2(n1200), .B1(n373), .B2(n3479), .ZN(
        n380) );
  INVD1BWP12T U1254 ( .I(r4[26]), .ZN(n1185) );
  INVD6BWP12T U1255 ( .I(n375), .ZN(n3476) );
  INVD1BWP12T U1256 ( .I(r0[26]), .ZN(n1187) );
  TPOAI22D1BWP12T U1257 ( .A1(n3448), .A2(n1185), .B1(n3476), .B2(n1187), .ZN(
        n379) );
  INVD9BWP12T U1258 ( .I(n1653), .ZN(n3478) );
  INVD1BWP12T U1259 ( .I(lr[26]), .ZN(n1199) );
  INVD1BWP12T U1260 ( .I(r8[26]), .ZN(n1197) );
  OAI22D0BWP12T U1261 ( .A1(n3478), .A2(n1199), .B1(n3477), .B2(n1197), .ZN(
        n378) );
  INVD1BWP12T U1262 ( .I(n[3674]), .ZN(n1991) );
  INVD1BWP12T U1263 ( .I(r11[26]), .ZN(n1188) );
  OAI22D0BWP12T U1264 ( .A1(n3491), .A2(n1991), .B1(n1188), .B2(n3490), .ZN(
        n387) );
  INVD1BWP12T U1265 ( .I(r5[26]), .ZN(n382) );
  INVD1BWP12T U1266 ( .I(r3[26]), .ZN(n1198) );
  OAI22D1BWP12T U1267 ( .A1(n3489), .A2(n382), .B1(n1198), .B2(n3488), .ZN(
        n386) );
  INVD12BWP12T U1268 ( .I(n1950), .ZN(n3487) );
  INVD1BWP12T U1269 ( .I(r7[26]), .ZN(n383) );
  OAI22D0BWP12T U1270 ( .A1(n3487), .A2(n383), .B1(n3486), .B2(n3646), .ZN(
        n385) );
  INVD1BWP12T U1271 ( .I(r1[26]), .ZN(n1195) );
  INVD1BWP12T U1272 ( .I(r12[26]), .ZN(n1196) );
  NR4D0BWP12T U1273 ( .A1(n387), .A2(n386), .A3(n385), .A4(n384), .ZN(n388) );
  CKND2D2BWP12T U1274 ( .A1(n389), .A2(n388), .ZN(regA_out[26]) );
  INVD1BWP12T U1275 ( .I(write1_sel[1]), .ZN(n390) );
  INR2D1BWP12T U1276 ( .A1(write1_sel[3]), .B1(n457), .ZN(n391) );
  INR2D2BWP12T U1277 ( .A1(n470), .B1(n526), .ZN(n392) );
  BUFFD16BWP12T U1278 ( .I(n392), .Z(n3381) );
  AN2D4BWP12T U1279 ( .A1(write1_in[23]), .A2(n3381), .Z(n394) );
  ND2D1BWP12T U1280 ( .A1(write2_in[24]), .A2(n3379), .ZN(n815) );
  CKND0BWP12T U1281 ( .I(write2_in[23]), .ZN(n1121) );
  TPNR2D0BWP12T U1282 ( .A1(n815), .A2(n1121), .ZN(n393) );
  TPAOI21D2BWP12T U1283 ( .A1(n394), .A2(write1_in[24]), .B(n393), .ZN(n3357)
         );
  TPNR3D1BWP12T U1284 ( .A1(n395), .A2(n256), .A3(n3357), .ZN(n443) );
  CKND2D1BWP12T U1285 ( .A1(write2_in[28]), .A2(n3379), .ZN(n447) );
  INVD1BWP12T U1286 ( .I(write2_in[26]), .ZN(n396) );
  ND2D1BWP12T U1287 ( .A1(write2_sel[2]), .A2(write2_sel[1]), .ZN(n552) );
  OAI21D0BWP12T U1288 ( .A1(write2_in[27]), .A2(n3381), .B(n3352), .ZN(n398)
         );
  INR2XD2BWP12T U1289 ( .A1(n447), .B1(n399), .ZN(n442) );
  INVD8BWP12T U1290 ( .I(write1_in[22]), .ZN(n401) );
  ND2D3BWP12T U1291 ( .A1(write1_in[21]), .A2(n3381), .ZN(n400) );
  NR2XD3BWP12T U1292 ( .A1(n401), .A2(n400), .ZN(n404) );
  CKND0BWP12T U1293 ( .I(write2_in[22]), .ZN(n402) );
  CKND2D1BWP12T U1294 ( .A1(write2_in[25]), .A2(n3379), .ZN(n3320) );
  NR3D1BWP12T U1295 ( .A1(n809), .A2(n402), .A3(n3320), .ZN(n403) );
  TPAOI21D4BWP12T U1296 ( .A1(n404), .A2(write1_in[25]), .B(n403), .ZN(n438)
         );
  TPND2D2BWP12T U1297 ( .A1(write1_in[18]), .A2(n3381), .ZN(n406) );
  TPND2D0BWP12T U1298 ( .A1(write2_in[18]), .A2(n3379), .ZN(n405) );
  TPND2D2BWP12T U1299 ( .A1(n406), .A2(n405), .ZN(n411) );
  INVD1P75BWP12T U1300 ( .I(n3381), .ZN(n3393) );
  IOA21D0BWP12T U1301 ( .A1(write2_in[17]), .A2(write2_in[16]), .B(n3393), 
        .ZN(n407) );
  TPOAI21D2BWP12T U1302 ( .A1(write1_in[16]), .A2(n3393), .B(n407), .ZN(n408)
         );
  NR2XD2BWP12T U1303 ( .A1(n409), .A2(n408), .ZN(n410) );
  TPND2D3BWP12T U1304 ( .A1(n411), .A2(n410), .ZN(n1970) );
  NR2XD2BWP12T U1305 ( .A1(n1970), .A2(n1973), .ZN(n437) );
  INVD1P75BWP12T U1306 ( .I(write1_in[14]), .ZN(n415) );
  INVD1BWP12T U1307 ( .I(n3381), .ZN(n414) );
  ND2D1BWP12T U1308 ( .A1(n2973), .A2(n414), .ZN(n413) );
  TPOAI21D2BWP12T U1309 ( .A1(n415), .A2(n414), .B(n413), .ZN(n664) );
  ND2D1BWP12T U1310 ( .A1(n843), .A2(n3379), .ZN(n416) );
  TPND2D3BWP12T U1311 ( .A1(n417), .A2(n416), .ZN(n544) );
  CKND2D2BWP12T U1312 ( .A1(write1_in[11]), .A2(n3381), .ZN(n419) );
  CKND2D1BWP12T U1313 ( .A1(n2971), .A2(n3379), .ZN(n418) );
  CKND2D2BWP12T U1314 ( .A1(n419), .A2(n418), .ZN(n844) );
  INVD1P75BWP12T U1315 ( .I(write1_in[12]), .ZN(n421) );
  ND2D1BWP12T U1316 ( .A1(n727), .A2(n3379), .ZN(n420) );
  INR2D1BWP12T U1317 ( .A1(n2972), .B1(n1856), .ZN(n422) );
  AO21D4BWP12T U1318 ( .A1(write1_in[13]), .A2(n1856), .B(n422), .Z(n510) );
  INR2D0BWP12T U1319 ( .A1(n3393), .B1(write2_in[19]), .ZN(n423) );
  INVD1BWP12T U1320 ( .I(n423), .ZN(n424) );
  ND2XD3BWP12T U1321 ( .A1(n510), .A2(n424), .ZN(n425) );
  NR2XD2BWP12T U1322 ( .A1(n508), .A2(n425), .ZN(n434) );
  INVD1BWP12T U1323 ( .I(n892), .ZN(n891) );
  ND2D1BWP12T U1324 ( .A1(n3393), .A2(n891), .ZN(n426) );
  TPOAI21D2BWP12T U1325 ( .A1(write1_in[1]), .A2(n3393), .B(n426), .ZN(n2924)
         );
  AN2XD1BWP12T U1326 ( .A1(n2882), .A2(n3393), .Z(n427) );
  TPAOI21D4BWP12T U1327 ( .A1(write1_in[2]), .A2(n1856), .B(n427), .ZN(n2925)
         );
  INVD1BWP12T U1328 ( .I(n3381), .ZN(n429) );
  ND2D1BWP12T U1329 ( .A1(n2913), .A2(n429), .ZN(n428) );
  TPND2D2BWP12T U1330 ( .A1(n2930), .A2(n2929), .ZN(n2944) );
  INR2D1BWP12T U1331 ( .A1(n2887), .B1(n1856), .ZN(n431) );
  TPAOI21D2BWP12T U1332 ( .A1(write1_in[4]), .A2(n1856), .B(n431), .ZN(n2943)
         );
  MUX2D1BWP12T U1333 ( .I0(n2900), .I1(write1_in[5]), .S(n3381), .Z(n732) );
  MUX2XD2BWP12T U1334 ( .I0(write2_in[7]), .I1(write1_in[7]), .S(n3381), .Z(
        n730) );
  CKND2D2BWP12T U1335 ( .A1(n731), .A2(n730), .ZN(n2984) );
  CKAN2D1BWP12T U1336 ( .A1(n2937), .A2(n3393), .Z(n432) );
  TPAOI21D1BWP12T U1337 ( .A1(write1_in[9]), .A2(n1856), .B(n432), .ZN(n2987)
         );
  TPNR2D2BWP12T U1338 ( .A1(n2984), .A2(n2987), .ZN(n433) );
  MUX2XD2BWP12T U1339 ( .I0(n866), .I1(write1_in[8]), .S(n3381), .Z(n2985) );
  TPND2D2BWP12T U1340 ( .A1(n433), .A2(n2985), .ZN(n719) );
  MUX2ND4BWP12T U1341 ( .I0(write1_in[10]), .I1(n2951), .S(n3393), .ZN(n720)
         );
  TPNR2D3BWP12T U1342 ( .A1(n719), .A2(n720), .ZN(n845) );
  NR3XD4BWP12T U1343 ( .A1(n436), .A2(n511), .A3(n435), .ZN(n1971) );
  ND2XD3BWP12T U1344 ( .A1(n437), .A2(n1971), .ZN(n1978) );
  TPNR2D3BWP12T U1345 ( .A1(next_pc_en_BAR), .A2(n439), .ZN(n3398) );
  INVD1BWP12T U1346 ( .I(n439), .ZN(n440) );
  TPAOI31D1BWP12T U1347 ( .A1(n443), .A2(n442), .A3(n44), .B(n441), .ZN(n450)
         );
  NR2D1BWP12T U1348 ( .A1(n3357), .A2(n3340), .ZN(n446) );
  TPND2D0BWP12T U1349 ( .A1(write2_in[27]), .A2(n3379), .ZN(n444) );
  TPND2D3BWP12T U1350 ( .A1(n445), .A2(n444), .ZN(n1867) );
  ND3XD3BWP12T U1351 ( .A1(n448), .A2(n3352), .A3(n3366), .ZN(n449) );
  ND3D1BWP12T U1352 ( .A1(write1_sel[3]), .A2(write1_en), .A3(n457), .ZN(n549)
         );
  TPND2D1BWP12T U1353 ( .A1(n247), .A2(n3216), .ZN(n455) );
  ND2D1BWP12T U1354 ( .A1(n458), .A2(write2_sel[3]), .ZN(n520) );
  INR2D1BWP12T U1355 ( .A1(write2_sel[2]), .B1(write2_sel[1]), .ZN(n584) );
  ND2D1BWP12T U1356 ( .A1(n485), .A2(n584), .ZN(n452) );
  AOI22D0BWP12T U1357 ( .A1(write2_in[26]), .A2(n3218), .B1(n3217), .B2(
        r12[26]), .ZN(n454) );
  BUFFXD6BWP12T U1358 ( .I(write1_in[29]), .Z(n3372) );
  TPND2D1BWP12T U1359 ( .A1(n3372), .A2(n3623), .ZN(n462) );
  INVD1BWP12T U1360 ( .I(write2_sel[3]), .ZN(n464) );
  ND2D1BWP12T U1361 ( .A1(n537), .A2(n584), .ZN(n459) );
  AOI22D0BWP12T U1362 ( .A1(write2_in[29]), .A2(n3281), .B1(n3280), .B2(r4[29]), .ZN(n461) );
  TPND2D1BWP12T U1363 ( .A1(n3372), .A2(n3289), .ZN(n469) );
  ND2D1BWP12T U1364 ( .A1(n585), .A2(n503), .ZN(n466) );
  AOI22D0BWP12T U1365 ( .A1(write2_in[29]), .A2(n3291), .B1(n3290), .B2(r1[29]), .ZN(n468) );
  TPND2D1BWP12T U1366 ( .A1(n247), .A2(n3234), .ZN(n474) );
  INVD1BWP12T U1367 ( .I(n552), .ZN(n480) );
  ND2D1BWP12T U1368 ( .A1(n485), .A2(n480), .ZN(n471) );
  AOI22D0BWP12T U1369 ( .A1(write2_in[26]), .A2(n3236), .B1(n3235), .B2(lr[26]), .ZN(n473) );
  TPND2D1BWP12T U1370 ( .A1(n247), .A2(n3229), .ZN(n479) );
  ND2D1BWP12T U1371 ( .A1(n531), .A2(n584), .ZN(n476) );
  AOI22D0BWP12T U1372 ( .A1(write2_in[26]), .A2(n3231), .B1(n3230), .B2(
        n[3674]), .ZN(n478) );
  TPND2D1BWP12T U1373 ( .A1(n247), .A2(n3241), .ZN(n484) );
  ND2D1BWP12T U1374 ( .A1(n585), .A2(n480), .ZN(n481) );
  ND2D1BWP12T U1375 ( .A1(n575), .A2(n3621), .ZN(n482) );
  AOI22D0BWP12T U1376 ( .A1(write2_in[26]), .A2(n3243), .B1(n3242), .B2(r7[26]), .ZN(n483) );
  TPND2D1BWP12T U1377 ( .A1(n247), .A2(n3211), .ZN(n489) );
  ND2D1BWP12T U1378 ( .A1(n485), .A2(n503), .ZN(n486) );
  AOI22D0BWP12T U1379 ( .A1(write2_in[26]), .A2(n3213), .B1(n3212), .B2(r8[26]), .ZN(n488) );
  TPND2D1BWP12T U1380 ( .A1(n3372), .A2(n3211), .ZN(n491) );
  AOI22D0BWP12T U1381 ( .A1(write2_in[29]), .A2(n3213), .B1(n3212), .B2(r8[29]), .ZN(n490) );
  NR2D1BWP12T U1382 ( .A1(n492), .A2(n552), .ZN(n494) );
  AOI22D0BWP12T U1383 ( .A1(write2_in[26]), .A2(n3263), .B1(n3262), .B2(r6[26]), .ZN(n495) );
  TPND2D1BWP12T U1384 ( .A1(n3372), .A2(n3284), .ZN(n501) );
  ND2D1BWP12T U1385 ( .A1(n537), .A2(n503), .ZN(n498) );
  AOI22D0BWP12T U1386 ( .A1(write2_in[29]), .A2(n3286), .B1(n3285), .B2(r0[29]), .ZN(n500) );
  TPND2D1BWP12T U1387 ( .A1(n247), .A2(n3248), .ZN(n507) );
  ND2D1BWP12T U1388 ( .A1(n531), .A2(n503), .ZN(n504) );
  AOI22D0BWP12T U1389 ( .A1(write2_in[26]), .A2(n3250), .B1(n3249), .B2(r9[26]), .ZN(n506) );
  CKND3BWP12T U1390 ( .I(n510), .ZN(n568) );
  NR2XD2BWP12T U1391 ( .A1(n567), .A2(n568), .ZN(n665) );
  IND2XD1BWP12T U1392 ( .A1(write2_in[16]), .B1(n3393), .ZN(n513) );
  INVD1BWP12T U1393 ( .I(n583), .ZN(n514) );
  CKND2D0BWP12T U1394 ( .A1(write1_in[22]), .A2(n3624), .ZN(n518) );
  INVD1BWP12T U1395 ( .I(write2_sel[1]), .ZN(n529) );
  NR3D1BWP12T U1396 ( .A1(n529), .A2(reset), .A3(write2_sel[2]), .ZN(n536) );
  ND2D1BWP12T U1397 ( .A1(n585), .A2(n536), .ZN(n516) );
  CKND2D1BWP12T U1398 ( .A1(n583), .A2(n538), .ZN(n515) );
  AOI22D0BWP12T U1399 ( .A1(write2_in[22]), .A2(n3028), .B1(n3303), .B2(r3[22]), .ZN(n517) );
  ND2D1BWP12T U1400 ( .A1(n518), .A2(n517), .ZN(n2543) );
  CKND2D0BWP12T U1401 ( .A1(write1_in[22]), .A2(n3627), .ZN(n525) );
  INVD1BWP12T U1402 ( .I(n536), .ZN(n527) );
  CKND2D1BWP12T U1403 ( .A1(n538), .A2(n521), .ZN(n522) );
  AOI22D0BWP12T U1404 ( .A1(write2_in[22]), .A2(n3298), .B1(n3297), .B2(
        r10[22]), .ZN(n524) );
  ND2D1BWP12T U1405 ( .A1(n525), .A2(n524), .ZN(n2319) );
  CKND2D0BWP12T U1406 ( .A1(write1_in[22]), .A2(n3626), .ZN(n533) );
  INR2D1BWP12T U1407 ( .A1(n538), .B1(n526), .ZN(n530) );
  AOI22D0BWP12T U1408 ( .A1(write2_in[22]), .A2(n3307), .B1(n3306), .B2(
        r11[22]), .ZN(n532) );
  ND2D1BWP12T U1409 ( .A1(n533), .A2(n532), .ZN(n2287) );
  INVD1BWP12T U1410 ( .I(n539), .ZN(n535) );
  CKND2D0BWP12T U1411 ( .A1(write1_in[22]), .A2(n3625), .ZN(n543) );
  CKND2D1BWP12T U1412 ( .A1(n537), .A2(n536), .ZN(n541) );
  CKND2D1BWP12T U1413 ( .A1(n539), .A2(n538), .ZN(n540) );
  AOI22D0BWP12T U1414 ( .A1(write2_in[22]), .A2(n3374), .B1(n3373), .B2(r2[22]), .ZN(n542) );
  ND2D1BWP12T U1415 ( .A1(n543), .A2(n542), .ZN(n2575) );
  BUFFD3BWP12T U1416 ( .I(write1_in[20]), .Z(n3051) );
  TPND2D0BWP12T U1417 ( .A1(n3051), .A2(n3234), .ZN(n546) );
  AOI22D0BWP12T U1418 ( .A1(write2_in[20]), .A2(n3236), .B1(n3235), .B2(lr[20]), .ZN(n545) );
  CKND2D1BWP12T U1419 ( .A1(n546), .A2(n545), .ZN(n2221) );
  CKND2D0BWP12T U1420 ( .A1(write1_in[21]), .A2(n3234), .ZN(n548) );
  AOI22D0BWP12T U1421 ( .A1(write2_in[21]), .A2(n3236), .B1(n3235), .B2(lr[21]), .ZN(n547) );
  CKND2D1BWP12T U1422 ( .A1(n548), .A2(n547), .ZN(n2222) );
  INR2XD0BWP12T U1423 ( .A1(write1_sel[4]), .B1(n549), .ZN(n551) );
  CKND2D0BWP12T U1424 ( .A1(write1_in[21]), .A2(n3638), .ZN(n556) );
  AOI22D0BWP12T U1425 ( .A1(write2_in[21]), .A2(n3277), .B1(n3276), .B2(
        tmp1[21]), .ZN(n555) );
  CKND2D1BWP12T U1426 ( .A1(n556), .A2(n555), .ZN(n2158) );
  TPND2D0BWP12T U1427 ( .A1(n3051), .A2(n3638), .ZN(n558) );
  AOI22D0BWP12T U1428 ( .A1(write2_in[20]), .A2(n3277), .B1(n3276), .B2(
        tmp1[20]), .ZN(n557) );
  CKND2D1BWP12T U1429 ( .A1(n558), .A2(n557), .ZN(n2157) );
  TPND2D0BWP12T U1430 ( .A1(n3051), .A2(n3211), .ZN(n560) );
  AOI22D0BWP12T U1431 ( .A1(write2_in[20]), .A2(n3213), .B1(n3212), .B2(r8[20]), .ZN(n559) );
  CKND2D1BWP12T U1432 ( .A1(n560), .A2(n559), .ZN(n2381) );
  CKND2D0BWP12T U1433 ( .A1(write1_in[21]), .A2(n3216), .ZN(n562) );
  AOI22D0BWP12T U1434 ( .A1(write2_in[21]), .A2(n3218), .B1(n3217), .B2(
        r12[21]), .ZN(n561) );
  CKND2D1BWP12T U1435 ( .A1(n562), .A2(n561), .ZN(n2254) );
  CKND2D0BWP12T U1436 ( .A1(write1_in[21]), .A2(n3211), .ZN(n564) );
  AOI22D0BWP12T U1437 ( .A1(write2_in[21]), .A2(n3213), .B1(n3212), .B2(r8[21]), .ZN(n563) );
  CKND2D1BWP12T U1438 ( .A1(n564), .A2(n563), .ZN(n2382) );
  TPND2D0BWP12T U1439 ( .A1(n3051), .A2(n3216), .ZN(n566) );
  AOI22D0BWP12T U1440 ( .A1(write2_in[20]), .A2(n3218), .B1(n3217), .B2(
        r12[20]), .ZN(n565) );
  CKND2D1BWP12T U1441 ( .A1(n566), .A2(n565), .ZN(n2253) );
  CKND2D0BWP12T U1442 ( .A1(write1_in[17]), .A2(n3234), .ZN(n570) );
  AOI22D0BWP12T U1443 ( .A1(write2_in[17]), .A2(n3236), .B1(n3235), .B2(lr[17]), .ZN(n569) );
  ND2D1BWP12T U1444 ( .A1(n570), .A2(n569), .ZN(n2218) );
  CKND2D0BWP12T U1445 ( .A1(write1_in[17]), .A2(n3624), .ZN(n572) );
  AOI22D0BWP12T U1446 ( .A1(write2_in[17]), .A2(n3028), .B1(n3303), .B2(r3[17]), .ZN(n571) );
  ND2D1BWP12T U1447 ( .A1(n572), .A2(n571), .ZN(n2538) );
  CKND2D0BWP12T U1448 ( .A1(write1_in[17]), .A2(n3626), .ZN(n574) );
  AOI22D0BWP12T U1449 ( .A1(write2_in[17]), .A2(n3307), .B1(n3306), .B2(
        r11[17]), .ZN(n573) );
  ND2D1BWP12T U1450 ( .A1(n574), .A2(n573), .ZN(n2282) );
  CKND2D0BWP12T U1451 ( .A1(write1_in[17]), .A2(n3627), .ZN(n577) );
  AOI22D0BWP12T U1452 ( .A1(write2_in[17]), .A2(n3298), .B1(n3297), .B2(
        r10[17]), .ZN(n576) );
  ND2D1BWP12T U1453 ( .A1(n577), .A2(n576), .ZN(n2314) );
  CKND2D0BWP12T U1454 ( .A1(write1_in[17]), .A2(n3625), .ZN(n579) );
  AOI22D0BWP12T U1455 ( .A1(write2_in[17]), .A2(n3374), .B1(n3373), .B2(r2[17]), .ZN(n578) );
  ND2D1BWP12T U1456 ( .A1(n579), .A2(n578), .ZN(n2570) );
  CKND2D0BWP12T U1457 ( .A1(write1_in[17]), .A2(n3211), .ZN(n581) );
  AOI22D0BWP12T U1458 ( .A1(write2_in[17]), .A2(n3213), .B1(n3212), .B2(r8[17]), .ZN(n580) );
  ND2D1BWP12T U1459 ( .A1(n581), .A2(n580), .ZN(n2378) );
  ND2D1BWP12T U1460 ( .A1(n585), .A2(n584), .ZN(n586) );
  CKND2D0BWP12T U1461 ( .A1(write1_in[18]), .A2(n3638), .ZN(n589) );
  AOI22D0BWP12T U1462 ( .A1(write2_in[18]), .A2(n3277), .B1(n3276), .B2(
        tmp1[18]), .ZN(n588) );
  CKND2D1BWP12T U1463 ( .A1(n589), .A2(n588), .ZN(n2155) );
  CKND2D0BWP12T U1464 ( .A1(write1_in[17]), .A2(n3638), .ZN(n591) );
  AOI22D0BWP12T U1465 ( .A1(write2_in[17]), .A2(n3277), .B1(n3276), .B2(
        tmp1[17]), .ZN(n590) );
  ND2D1BWP12T U1466 ( .A1(n591), .A2(n590), .ZN(n2154) );
  CKND2D0BWP12T U1467 ( .A1(write1_in[17]), .A2(n3216), .ZN(n593) );
  AOI22D0BWP12T U1468 ( .A1(write2_in[17]), .A2(n3218), .B1(n3217), .B2(
        r12[17]), .ZN(n592) );
  ND2D1BWP12T U1469 ( .A1(n593), .A2(n592), .ZN(n2250) );
  CKND2D0BWP12T U1470 ( .A1(write1_in[16]), .A2(n3623), .ZN(n595) );
  AOI22D0BWP12T U1471 ( .A1(write2_in[16]), .A2(n3281), .B1(n3280), .B2(r4[16]), .ZN(n594) );
  CKND2D1BWP12T U1472 ( .A1(n595), .A2(n594), .ZN(n2505) );
  CKND2D0BWP12T U1473 ( .A1(write1_in[16]), .A2(n3241), .ZN(n597) );
  AOI22D0BWP12T U1474 ( .A1(write2_in[16]), .A2(n3243), .B1(n3242), .B2(r7[16]), .ZN(n596) );
  CKND2D1BWP12T U1475 ( .A1(n597), .A2(n596), .ZN(n2409) );
  CKND2D0BWP12T U1476 ( .A1(write1_in[16]), .A2(n3622), .ZN(n599) );
  AOI22D0BWP12T U1477 ( .A1(write2_in[16]), .A2(n3273), .B1(n3272), .B2(r5[16]), .ZN(n598) );
  CKND2D1BWP12T U1478 ( .A1(n599), .A2(n598), .ZN(n2473) );
  CKND2D0BWP12T U1479 ( .A1(write1_in[16]), .A2(n3229), .ZN(n601) );
  AOI22D0BWP12T U1480 ( .A1(write2_in[16]), .A2(n3231), .B1(n3230), .B2(
        n[3684]), .ZN(n600) );
  CKND2D1BWP12T U1481 ( .A1(n601), .A2(n600), .ZN(spin[16]) );
  CKND2D0BWP12T U1482 ( .A1(write1_in[16]), .A2(n3248), .ZN(n603) );
  AOI22D0BWP12T U1483 ( .A1(write2_in[16]), .A2(n3250), .B1(n3249), .B2(r9[16]), .ZN(n602) );
  CKND2D1BWP12T U1484 ( .A1(n603), .A2(n602), .ZN(n2345) );
  TPND2D0BWP12T U1485 ( .A1(write1_in[11]), .A2(n3211), .ZN(n605) );
  AOI22D0BWP12T U1486 ( .A1(n2971), .A2(n3213), .B1(n3212), .B2(r8[11]), .ZN(
        n604) );
  CKND2D1BWP12T U1487 ( .A1(n605), .A2(n604), .ZN(n2372) );
  BUFFD4BWP12T U1488 ( .I(write1_in[6]), .Z(n2920) );
  TPND2D0BWP12T U1489 ( .A1(n2920), .A2(n3638), .ZN(n607) );
  AOI22D0BWP12T U1490 ( .A1(n2921), .A2(n3277), .B1(n3276), .B2(tmp1[6]), .ZN(
        n606) );
  CKND2D1BWP12T U1491 ( .A1(n607), .A2(n606), .ZN(n2143) );
  TPND2D0BWP12T U1492 ( .A1(write1_in[4]), .A2(n3241), .ZN(n609) );
  AOI22D0BWP12T U1493 ( .A1(n2887), .A2(n3243), .B1(n3242), .B2(r7[4]), .ZN(
        n608) );
  CKND2D1BWP12T U1494 ( .A1(n609), .A2(n608), .ZN(n2397) );
  TPND2D0BWP12T U1495 ( .A1(write1_in[4]), .A2(n3229), .ZN(n613) );
  INVD0BWP12T U1496 ( .I(n2887), .ZN(n610) );
  NR2D1BWP12T U1497 ( .A1(n610), .A2(n2938), .ZN(n611) );
  RCAOI211D0BWP12T U1498 ( .A1(n3230), .A2(n[3696]), .B(n611), .C(reset), .ZN(
        n612) );
  CKND2D1BWP12T U1499 ( .A1(n613), .A2(n612), .ZN(spin[4]) );
  TPND2D0BWP12T U1500 ( .A1(write1_in[4]), .A2(n3248), .ZN(n615) );
  AOI22D0BWP12T U1501 ( .A1(n2887), .A2(n3250), .B1(n3249), .B2(r9[4]), .ZN(
        n614) );
  CKND2D1BWP12T U1502 ( .A1(n615), .A2(n614), .ZN(n2333) );
  TPND2D0BWP12T U1503 ( .A1(n782), .A2(n3216), .ZN(n617) );
  AOI22D0BWP12T U1504 ( .A1(n3218), .A2(write2_in[0]), .B1(n3217), .B2(r12[0]), 
        .ZN(n616) );
  CKND2D1BWP12T U1505 ( .A1(n617), .A2(n616), .ZN(n2233) );
  TPND2D0BWP12T U1506 ( .A1(n782), .A2(n3241), .ZN(n619) );
  AOI22D0BWP12T U1507 ( .A1(n3243), .A2(write2_in[0]), .B1(n3242), .B2(r7[0]), 
        .ZN(n618) );
  CKND2D1BWP12T U1508 ( .A1(n619), .A2(n618), .ZN(n2393) );
  TPND2D0BWP12T U1509 ( .A1(n782), .A2(n3622), .ZN(n621) );
  AOI22D0BWP12T U1510 ( .A1(n3273), .A2(write2_in[0]), .B1(n3272), .B2(r5[0]), 
        .ZN(n620) );
  CKND2D1BWP12T U1511 ( .A1(n621), .A2(n620), .ZN(n2457) );
  TPND2D0BWP12T U1512 ( .A1(n782), .A2(n3289), .ZN(n623) );
  AOI22D0BWP12T U1513 ( .A1(n3291), .A2(write2_in[0]), .B1(n3290), .B2(r1[0]), 
        .ZN(n622) );
  CKND2D1BWP12T U1514 ( .A1(n623), .A2(n622), .ZN(n2585) );
  TPND2D0BWP12T U1515 ( .A1(n782), .A2(n3229), .ZN(n625) );
  AOI22D0BWP12T U1516 ( .A1(n3231), .A2(write2_in[0]), .B1(n3230), .B2(n[3700]), .ZN(n624) );
  CKND2D1BWP12T U1517 ( .A1(n625), .A2(n624), .ZN(spin[0]) );
  TPND2D0BWP12T U1518 ( .A1(n782), .A2(n3234), .ZN(n627) );
  AOI22D0BWP12T U1519 ( .A1(n3236), .A2(write2_in[0]), .B1(n3235), .B2(lr[0]), 
        .ZN(n626) );
  CKND2D1BWP12T U1520 ( .A1(n627), .A2(n626), .ZN(n2201) );
  TPND2D0BWP12T U1521 ( .A1(n782), .A2(n3248), .ZN(n629) );
  AOI22D0BWP12T U1522 ( .A1(n3250), .A2(write2_in[0]), .B1(n3249), .B2(r9[0]), 
        .ZN(n628) );
  CKND2D1BWP12T U1523 ( .A1(n629), .A2(n628), .ZN(n2329) );
  TPND2D0BWP12T U1524 ( .A1(n782), .A2(n3638), .ZN(n631) );
  AOI22D0BWP12T U1525 ( .A1(write2_in[0]), .A2(n3277), .B1(n3276), .B2(tmp1[0]), .ZN(n630) );
  CKND2D1BWP12T U1526 ( .A1(n631), .A2(n630), .ZN(n2136) );
  TPND2D0BWP12T U1527 ( .A1(n782), .A2(n3211), .ZN(n633) );
  AOI22D0BWP12T U1528 ( .A1(n3213), .A2(write2_in[0]), .B1(n3212), .B2(r8[0]), 
        .ZN(n632) );
  CKND2D1BWP12T U1529 ( .A1(n633), .A2(n632), .ZN(n2361) );
  TPND2D0BWP12T U1530 ( .A1(n782), .A2(n3623), .ZN(n635) );
  AOI22D0BWP12T U1531 ( .A1(n3281), .A2(write2_in[0]), .B1(n3280), .B2(r4[0]), 
        .ZN(n634) );
  CKND2D1BWP12T U1532 ( .A1(n635), .A2(n634), .ZN(n2489) );
  TPND2D1BWP12T U1533 ( .A1(n249), .A2(n3284), .ZN(n637) );
  AOI22D0BWP12T U1534 ( .A1(write2_in[30]), .A2(n3286), .B1(n3285), .B2(r0[30]), .ZN(n636) );
  TPND2D1BWP12T U1535 ( .A1(n249), .A2(n3241), .ZN(n639) );
  AOI22D0BWP12T U1536 ( .A1(write2_in[30]), .A2(n3243), .B1(n3242), .B2(r7[30]), .ZN(n638) );
  TPND2D1BWP12T U1537 ( .A1(n249), .A2(n3289), .ZN(n641) );
  AOI22D0BWP12T U1538 ( .A1(write2_in[30]), .A2(n3291), .B1(n3290), .B2(r1[30]), .ZN(n640) );
  TPND2D1BWP12T U1539 ( .A1(n249), .A2(n3229), .ZN(n643) );
  AOI22D0BWP12T U1540 ( .A1(write2_in[30]), .A2(n3231), .B1(n3230), .B2(
        n[3670]), .ZN(n642) );
  TPND2D1BWP12T U1541 ( .A1(n3372), .A2(n3622), .ZN(n645) );
  AOI22D0BWP12T U1542 ( .A1(write2_in[29]), .A2(n3273), .B1(n3272), .B2(r5[29]), .ZN(n644) );
  TPND2D1BWP12T U1543 ( .A1(n645), .A2(n644), .ZN(n2486) );
  TPND2D1BWP12T U1544 ( .A1(n3372), .A2(n3241), .ZN(n647) );
  AOI22D0BWP12T U1545 ( .A1(write2_in[29]), .A2(n3243), .B1(n3242), .B2(r7[29]), .ZN(n646) );
  TPND2D1BWP12T U1546 ( .A1(n647), .A2(n646), .ZN(n2422) );
  TPND2D1BWP12T U1547 ( .A1(n3372), .A2(n3628), .ZN(n649) );
  AOI22D0BWP12T U1548 ( .A1(write2_in[29]), .A2(n3263), .B1(n3262), .B2(r6[29]), .ZN(n648) );
  TPND2D1BWP12T U1549 ( .A1(n649), .A2(n648), .ZN(n2454) );
  CKND2D0BWP12T U1550 ( .A1(write1_in[22]), .A2(n3623), .ZN(n651) );
  AOI22D0BWP12T U1551 ( .A1(write2_in[22]), .A2(n3281), .B1(n3280), .B2(r4[22]), .ZN(n650) );
  ND2D1BWP12T U1552 ( .A1(n651), .A2(n650), .ZN(n2511) );
  CKND2D0BWP12T U1553 ( .A1(write1_in[22]), .A2(n3248), .ZN(n653) );
  AOI22D0BWP12T U1554 ( .A1(write2_in[22]), .A2(n3250), .B1(n3249), .B2(r9[22]), .ZN(n652) );
  ND2D1BWP12T U1555 ( .A1(n653), .A2(n652), .ZN(n2351) );
  CKND2D0BWP12T U1556 ( .A1(write1_in[22]), .A2(n3229), .ZN(n655) );
  AOI22D0BWP12T U1557 ( .A1(write2_in[22]), .A2(n3231), .B1(n3230), .B2(
        n[3678]), .ZN(n654) );
  ND2D1BWP12T U1558 ( .A1(n655), .A2(n654), .ZN(spin[22]) );
  CKND2D0BWP12T U1559 ( .A1(write1_in[22]), .A2(n3628), .ZN(n657) );
  AOI22D0BWP12T U1560 ( .A1(write2_in[22]), .A2(n3263), .B1(n3262), .B2(r6[22]), .ZN(n656) );
  ND2D1BWP12T U1561 ( .A1(n657), .A2(n656), .ZN(n2447) );
  CKND2D0BWP12T U1562 ( .A1(write1_in[22]), .A2(n3622), .ZN(n659) );
  AOI22D0BWP12T U1563 ( .A1(write2_in[22]), .A2(n3273), .B1(n3272), .B2(r5[22]), .ZN(n658) );
  ND2D1BWP12T U1564 ( .A1(n659), .A2(n658), .ZN(n2479) );
  CKND2D0BWP12T U1565 ( .A1(write1_in[22]), .A2(n3241), .ZN(n661) );
  AOI22D0BWP12T U1566 ( .A1(write2_in[22]), .A2(n3243), .B1(n3242), .B2(r7[22]), .ZN(n660) );
  ND2D1BWP12T U1567 ( .A1(n661), .A2(n660), .ZN(n2415) );
  CKND2D0BWP12T U1568 ( .A1(write1_in[19]), .A2(n3638), .ZN(n663) );
  AOI22D0BWP12T U1569 ( .A1(write2_in[19]), .A2(n3277), .B1(n3276), .B2(
        tmp1[19]), .ZN(n662) );
  CKND2D1BWP12T U1570 ( .A1(n663), .A2(n662), .ZN(n2156) );
  CKND2D0BWP12T U1571 ( .A1(write1_in[19]), .A2(n3216), .ZN(n667) );
  AOI22D0BWP12T U1572 ( .A1(write2_in[19]), .A2(n3218), .B1(n3217), .B2(
        r12[19]), .ZN(n666) );
  CKND2D1BWP12T U1573 ( .A1(n667), .A2(n666), .ZN(n2252) );
  CKND2D0BWP12T U1574 ( .A1(write1_in[19]), .A2(n3211), .ZN(n669) );
  AOI22D0BWP12T U1575 ( .A1(write2_in[19]), .A2(n3213), .B1(n3212), .B2(r8[19]), .ZN(n668) );
  CKND2D1BWP12T U1576 ( .A1(n669), .A2(n668), .ZN(n2380) );
  CKND2D0BWP12T U1577 ( .A1(write1_in[19]), .A2(n3234), .ZN(n671) );
  AOI22D0BWP12T U1578 ( .A1(write2_in[19]), .A2(n3236), .B1(n3235), .B2(lr[19]), .ZN(n670) );
  CKND2D1BWP12T U1579 ( .A1(n671), .A2(n670), .ZN(n2220) );
  CKND2D0BWP12T U1580 ( .A1(write1_in[18]), .A2(n3229), .ZN(n673) );
  AOI22D0BWP12T U1581 ( .A1(write2_in[18]), .A2(n3231), .B1(n3230), .B2(
        n[3682]), .ZN(n672) );
  ND2D1BWP12T U1582 ( .A1(n673), .A2(n672), .ZN(spin[18]) );
  CKND2D0BWP12T U1583 ( .A1(write1_in[18]), .A2(n3234), .ZN(n675) );
  AOI22D0BWP12T U1584 ( .A1(write2_in[18]), .A2(n3236), .B1(n3235), .B2(lr[18]), .ZN(n674) );
  CKND2D1BWP12T U1585 ( .A1(n675), .A2(n674), .ZN(n2219) );
  CKND2D0BWP12T U1586 ( .A1(write1_in[18]), .A2(n3211), .ZN(n677) );
  AOI22D0BWP12T U1587 ( .A1(write2_in[18]), .A2(n3213), .B1(n3212), .B2(r8[18]), .ZN(n676) );
  CKND2D1BWP12T U1588 ( .A1(n677), .A2(n676), .ZN(n2379) );
  CKND2D0BWP12T U1589 ( .A1(write1_in[18]), .A2(n3627), .ZN(n679) );
  AOI22D0BWP12T U1590 ( .A1(write2_in[18]), .A2(n3298), .B1(n3297), .B2(
        r10[18]), .ZN(n678) );
  ND2D1BWP12T U1591 ( .A1(n679), .A2(n678), .ZN(n2315) );
  CKND2D0BWP12T U1592 ( .A1(write1_in[17]), .A2(n3229), .ZN(n681) );
  AOI22D0BWP12T U1593 ( .A1(write2_in[17]), .A2(n3231), .B1(n3230), .B2(
        n[3683]), .ZN(n680) );
  ND2D1BWP12T U1594 ( .A1(n681), .A2(n680), .ZN(spin[17]) );
  CKND2D0BWP12T U1595 ( .A1(write1_in[17]), .A2(n3622), .ZN(n683) );
  AOI22D0BWP12T U1596 ( .A1(write2_in[17]), .A2(n3273), .B1(n3272), .B2(r5[17]), .ZN(n682) );
  ND2D1BWP12T U1597 ( .A1(n683), .A2(n682), .ZN(n2474) );
  CKND2D0BWP12T U1598 ( .A1(write1_in[17]), .A2(n3628), .ZN(n685) );
  AOI22D0BWP12T U1599 ( .A1(write2_in[17]), .A2(n3263), .B1(n3262), .B2(r6[17]), .ZN(n684) );
  ND2D1BWP12T U1600 ( .A1(n685), .A2(n684), .ZN(n2442) );
  CKND2D0BWP12T U1601 ( .A1(write1_in[17]), .A2(n3241), .ZN(n687) );
  AOI22D0BWP12T U1602 ( .A1(write2_in[17]), .A2(n3243), .B1(n3242), .B2(r7[17]), .ZN(n686) );
  ND2D1BWP12T U1603 ( .A1(n687), .A2(n686), .ZN(n2410) );
  CKND2D0BWP12T U1604 ( .A1(write1_in[17]), .A2(n3248), .ZN(n689) );
  AOI22D0BWP12T U1605 ( .A1(write2_in[17]), .A2(n3250), .B1(n3249), .B2(r9[17]), .ZN(n688) );
  ND2D1BWP12T U1606 ( .A1(n689), .A2(n688), .ZN(n2346) );
  CKND2D0BWP12T U1607 ( .A1(write1_in[18]), .A2(n3248), .ZN(n691) );
  AOI22D0BWP12T U1608 ( .A1(write2_in[18]), .A2(n3250), .B1(n3249), .B2(r9[18]), .ZN(n690) );
  ND2D1BWP12T U1609 ( .A1(n691), .A2(n690), .ZN(n2347) );
  CKND2D0BWP12T U1610 ( .A1(write1_in[17]), .A2(n3623), .ZN(n693) );
  AOI22D0BWP12T U1611 ( .A1(write2_in[17]), .A2(n3281), .B1(n3280), .B2(r4[17]), .ZN(n692) );
  ND2D1BWP12T U1612 ( .A1(n693), .A2(n692), .ZN(n2506) );
  CKND2D0BWP12T U1613 ( .A1(write1_in[18]), .A2(n3625), .ZN(n695) );
  AOI22D0BWP12T U1614 ( .A1(write2_in[18]), .A2(n3374), .B1(n3373), .B2(r2[18]), .ZN(n694) );
  ND2D1BWP12T U1615 ( .A1(n695), .A2(n694), .ZN(n2571) );
  CKND2D0BWP12T U1616 ( .A1(write1_in[18]), .A2(n3626), .ZN(n697) );
  AOI22D0BWP12T U1617 ( .A1(write2_in[18]), .A2(n3307), .B1(n3306), .B2(
        r11[18]), .ZN(n696) );
  ND2D1BWP12T U1618 ( .A1(n697), .A2(n696), .ZN(n2283) );
  CKND2D0BWP12T U1619 ( .A1(write1_in[18]), .A2(n3216), .ZN(n699) );
  AOI22D0BWP12T U1620 ( .A1(write2_in[18]), .A2(n3218), .B1(n3217), .B2(
        r12[18]), .ZN(n698) );
  CKND2D1BWP12T U1621 ( .A1(n699), .A2(n698), .ZN(n2251) );
  CKND2D0BWP12T U1622 ( .A1(write1_in[18]), .A2(n3624), .ZN(n702) );
  AOI22D0BWP12T U1623 ( .A1(write2_in[18]), .A2(n3028), .B1(n3303), .B2(r3[18]), .ZN(n701) );
  ND2D1BWP12T U1624 ( .A1(n702), .A2(n701), .ZN(n2539) );
  CKND2D0BWP12T U1625 ( .A1(write1_in[16]), .A2(n3216), .ZN(n704) );
  AOI22D0BWP12T U1626 ( .A1(write2_in[16]), .A2(n3218), .B1(n3217), .B2(
        r12[16]), .ZN(n703) );
  CKND2D1BWP12T U1627 ( .A1(n704), .A2(n703), .ZN(n2249) );
  CKND2D0BWP12T U1628 ( .A1(write1_in[16]), .A2(n3638), .ZN(n706) );
  AOI22D0BWP12T U1629 ( .A1(write2_in[16]), .A2(n3277), .B1(n3276), .B2(
        tmp1[16]), .ZN(n705) );
  CKND2D1BWP12T U1630 ( .A1(n706), .A2(n705), .ZN(n2153) );
  CKND2D0BWP12T U1631 ( .A1(write1_in[16]), .A2(n3626), .ZN(n708) );
  AOI22D0BWP12T U1632 ( .A1(write2_in[16]), .A2(n3307), .B1(n3306), .B2(
        r11[16]), .ZN(n707) );
  ND2D1BWP12T U1633 ( .A1(n708), .A2(n707), .ZN(n2281) );
  CKND2D0BWP12T U1634 ( .A1(write1_in[16]), .A2(n3625), .ZN(n710) );
  AOI22D0BWP12T U1635 ( .A1(write2_in[16]), .A2(n3374), .B1(n3373), .B2(r2[16]), .ZN(n709) );
  ND2D1BWP12T U1636 ( .A1(n710), .A2(n709), .ZN(n2569) );
  CKND2D0BWP12T U1637 ( .A1(write1_in[16]), .A2(n3624), .ZN(n712) );
  AOI22D0BWP12T U1638 ( .A1(write2_in[16]), .A2(n3028), .B1(n3303), .B2(r3[16]), .ZN(n711) );
  ND2D1BWP12T U1639 ( .A1(n712), .A2(n711), .ZN(n2537) );
  CKND2D0BWP12T U1640 ( .A1(write1_in[16]), .A2(n3234), .ZN(n714) );
  AOI22D0BWP12T U1641 ( .A1(write2_in[16]), .A2(n3236), .B1(n3235), .B2(lr[16]), .ZN(n713) );
  CKND2D1BWP12T U1642 ( .A1(n714), .A2(n713), .ZN(n2217) );
  CKND2D0BWP12T U1643 ( .A1(write1_in[16]), .A2(n3211), .ZN(n716) );
  AOI22D0BWP12T U1644 ( .A1(write2_in[16]), .A2(n3213), .B1(n3212), .B2(r8[16]), .ZN(n715) );
  CKND2D1BWP12T U1645 ( .A1(n716), .A2(n715), .ZN(n2377) );
  CKND2D0BWP12T U1646 ( .A1(write1_in[16]), .A2(n3627), .ZN(n718) );
  AOI22D0BWP12T U1647 ( .A1(write2_in[16]), .A2(n3298), .B1(n3297), .B2(
        r10[16]), .ZN(n717) );
  ND2D1BWP12T U1648 ( .A1(n718), .A2(n717), .ZN(n2313) );
  XNR2XD0BWP12T U1649 ( .A1(n720), .A2(n719), .ZN(n722) );
  AOI22D1BWP12T U1650 ( .A1(n2989), .A2(pc_out[10]), .B1(n3398), .B2(
        next_pc_in[10]), .ZN(n721) );
  OAI21D1BWP12T U1651 ( .A1(n722), .A2(n3394), .B(n721), .ZN(n2179) );
  CKND2D0BWP12T U1652 ( .A1(write1_in[12]), .A2(n3625), .ZN(n724) );
  AOI22D0BWP12T U1653 ( .A1(n727), .A2(n3374), .B1(n3373), .B2(r2[12]), .ZN(
        n723) );
  ND2D1BWP12T U1654 ( .A1(n724), .A2(n723), .ZN(n2565) );
  XOR2XD0BWP12T U1655 ( .A1(n2985), .A2(n2984), .Z(n726) );
  AOI22D1BWP12T U1656 ( .A1(n2989), .A2(pc_out[8]), .B1(n3398), .B2(
        next_pc_in[8]), .ZN(n725) );
  OAI21D1BWP12T U1657 ( .A1(n726), .A2(n3394), .B(n725), .ZN(n2177) );
  TPND2D0BWP12T U1658 ( .A1(write1_in[7]), .A2(n3625), .ZN(n735) );
  AOI22D0BWP12T U1659 ( .A1(n3373), .A2(r2[7]), .B1(n3374), .B2(write2_in[7]), 
        .ZN(n734) );
  ND2D1BWP12T U1660 ( .A1(n735), .A2(n734), .ZN(n2560) );
  TPND2D0BWP12T U1661 ( .A1(write1_in[4]), .A2(n3216), .ZN(n737) );
  AOI22D0BWP12T U1662 ( .A1(n2887), .A2(n3218), .B1(n3217), .B2(r12[4]), .ZN(
        n736) );
  CKND2D1BWP12T U1663 ( .A1(n737), .A2(n736), .ZN(n2237) );
  TPND2D0BWP12T U1664 ( .A1(write1_in[7]), .A2(n3627), .ZN(n739) );
  AOI22D0BWP12T U1665 ( .A1(write2_in[7]), .A2(n3298), .B1(n3297), .B2(r10[7]), 
        .ZN(n738) );
  ND2D1BWP12T U1666 ( .A1(n739), .A2(n738), .ZN(n2304) );
  TPND2D0BWP12T U1667 ( .A1(write1_in[7]), .A2(n3628), .ZN(n741) );
  AOI22D0BWP12T U1668 ( .A1(write2_in[7]), .A2(n3263), .B1(n3262), .B2(r6[7]), 
        .ZN(n740) );
  ND2D1BWP12T U1669 ( .A1(n741), .A2(n740), .ZN(n2432) );
  TPND2D0BWP12T U1670 ( .A1(write1_in[4]), .A2(n3638), .ZN(n743) );
  AOI22D0BWP12T U1671 ( .A1(n2887), .A2(n3277), .B1(n3276), .B2(tmp1[4]), .ZN(
        n742) );
  CKND2D1BWP12T U1672 ( .A1(n743), .A2(n742), .ZN(n2141) );
  TPND2D0BWP12T U1673 ( .A1(write1_in[4]), .A2(n3628), .ZN(n745) );
  AOI22D0BWP12T U1674 ( .A1(n2887), .A2(n3263), .B1(n3262), .B2(r6[4]), .ZN(
        n744) );
  ND2D1BWP12T U1675 ( .A1(n745), .A2(n744), .ZN(n2429) );
  TPND2D0BWP12T U1676 ( .A1(write1_in[4]), .A2(n3211), .ZN(n747) );
  AOI22D0BWP12T U1677 ( .A1(n2887), .A2(n3213), .B1(n3212), .B2(r8[4]), .ZN(
        n746) );
  CKND2D1BWP12T U1678 ( .A1(n747), .A2(n746), .ZN(n2365) );
  TPND2D0BWP12T U1679 ( .A1(write1_in[4]), .A2(n3234), .ZN(n749) );
  AOI22D0BWP12T U1680 ( .A1(n2887), .A2(n3236), .B1(n3235), .B2(lr[4]), .ZN(
        n748) );
  CKND2D1BWP12T U1681 ( .A1(n749), .A2(n748), .ZN(n2205) );
  TPND2D0BWP12T U1682 ( .A1(write1_in[7]), .A2(n3626), .ZN(n751) );
  AOI22D0BWP12T U1683 ( .A1(write2_in[7]), .A2(n3307), .B1(n3306), .B2(r11[7]), 
        .ZN(n750) );
  ND2D1BWP12T U1684 ( .A1(n751), .A2(n750), .ZN(n2272) );
  TPND2D0BWP12T U1685 ( .A1(write1_in[7]), .A2(n3624), .ZN(n753) );
  AOI22D0BWP12T U1686 ( .A1(n3303), .A2(r3[7]), .B1(write2_in[7]), .B2(n3028), 
        .ZN(n752) );
  ND2D1BWP12T U1687 ( .A1(n753), .A2(n752), .ZN(n2528) );
  TPND2D0BWP12T U1688 ( .A1(write1_in[3]), .A2(n3229), .ZN(n757) );
  INVD0BWP12T U1689 ( .I(n2913), .ZN(n754) );
  NR2D1BWP12T U1690 ( .A1(n754), .A2(n2938), .ZN(n755) );
  AOI211D0BWP12T U1691 ( .A1(n3230), .A2(n[3697]), .B(n755), .C(reset), .ZN(
        n756) );
  CKND2D1BWP12T U1692 ( .A1(n757), .A2(n756), .ZN(spin[3]) );
  TPND2D0BWP12T U1693 ( .A1(write1_in[5]), .A2(n3229), .ZN(n761) );
  INVD0BWP12T U1694 ( .I(n2900), .ZN(n758) );
  NR2D1BWP12T U1695 ( .A1(n758), .A2(n2938), .ZN(n759) );
  RCAOI211D0BWP12T U1696 ( .A1(n3230), .A2(n[3695]), .B(n759), .C(reset), .ZN(
        n760) );
  CKND2D1BWP12T U1697 ( .A1(n761), .A2(n760), .ZN(spin[5]) );
  TPND2D0BWP12T U1698 ( .A1(write1_in[3]), .A2(n3289), .ZN(n763) );
  AOI22D0BWP12T U1699 ( .A1(n2913), .A2(n3291), .B1(n3290), .B2(r1[3]), .ZN(
        n762) );
  CKND2D1BWP12T U1700 ( .A1(n763), .A2(n762), .ZN(n2588) );
  TPND2D0BWP12T U1701 ( .A1(write1_in[5]), .A2(n3638), .ZN(n765) );
  AOI22D0BWP12T U1702 ( .A1(n2900), .A2(n3277), .B1(n3276), .B2(tmp1[5]), .ZN(
        n764) );
  CKND2D1BWP12T U1703 ( .A1(n765), .A2(n764), .ZN(n2142) );
  TPND2D0BWP12T U1704 ( .A1(n782), .A2(n3624), .ZN(n767) );
  AOI22D0BWP12T U1705 ( .A1(n3303), .A2(r3[0]), .B1(n3028), .B2(write2_in[0]), 
        .ZN(n766) );
  ND2D1BWP12T U1706 ( .A1(n767), .A2(n766), .ZN(n2521) );
  ND2D0BWP12T U1707 ( .A1(n41), .A2(n3624), .ZN(n769) );
  AOI22D0BWP12T U1708 ( .A1(n3303), .A2(r3[2]), .B1(n2882), .B2(n3028), .ZN(
        n768) );
  CKND2D1BWP12T U1709 ( .A1(n769), .A2(n768), .ZN(n2523) );
  TPND2D0BWP12T U1710 ( .A1(n782), .A2(n3627), .ZN(n771) );
  AOI22D0BWP12T U1711 ( .A1(n3298), .A2(write2_in[0]), .B1(n3297), .B2(r10[0]), 
        .ZN(n770) );
  ND2D1BWP12T U1712 ( .A1(n771), .A2(n770), .ZN(n2297) );
  TPND2D0BWP12T U1713 ( .A1(n41), .A2(n3229), .ZN(n775) );
  INVD0BWP12T U1714 ( .I(n2882), .ZN(n772) );
  NR2D1BWP12T U1715 ( .A1(n772), .A2(n2938), .ZN(n773) );
  RCAOI211D0BWP12T U1716 ( .A1(n3230), .A2(n[3698]), .B(n773), .C(reset), .ZN(
        n774) );
  CKND2D1BWP12T U1717 ( .A1(n775), .A2(n774), .ZN(spin[2]) );
  TPND2D0BWP12T U1718 ( .A1(n782), .A2(n3626), .ZN(n777) );
  AOI22D0BWP12T U1719 ( .A1(n3307), .A2(write2_in[0]), .B1(n3306), .B2(r11[0]), 
        .ZN(n776) );
  ND2D1BWP12T U1720 ( .A1(n777), .A2(n776), .ZN(n2265) );
  TPND2D0BWP12T U1721 ( .A1(n782), .A2(n3628), .ZN(n779) );
  AOI22D0BWP12T U1722 ( .A1(n3263), .A2(write2_in[0]), .B1(n3262), .B2(r6[0]), 
        .ZN(n778) );
  ND2D1BWP12T U1723 ( .A1(n779), .A2(n778), .ZN(n2425) );
  MUX2NXD0BWP12T U1724 ( .I0(n782), .I1(write2_in[0]), .S(n3393), .ZN(n781) );
  AOI22D0BWP12T U1725 ( .A1(n2989), .A2(pc_out[0]), .B1(n3398), .B2(
        next_pc_in[0]), .ZN(n780) );
  OAI21D1BWP12T U1726 ( .A1(n781), .A2(n3394), .B(n780), .ZN(n2169) );
  TPND2D0BWP12T U1727 ( .A1(n782), .A2(n3625), .ZN(n784) );
  AOI22D0BWP12T U1728 ( .A1(n3373), .A2(r2[0]), .B1(n3374), .B2(write2_in[0]), 
        .ZN(n783) );
  ND2D1BWP12T U1729 ( .A1(n784), .A2(n783), .ZN(n2553) );
  AOI22D0BWP12T U1730 ( .A1(write2_in[30]), .A2(n3281), .B1(n3280), .B2(r4[30]), .ZN(n3635) );
  AOI22D0BWP12T U1731 ( .A1(write2_in[30]), .A2(n3277), .B1(n3276), .B2(
        tmp1[30]), .ZN(n3639) );
  AOI22D0BWP12T U1732 ( .A1(write2_in[30]), .A2(n3374), .B1(n3373), .B2(r2[30]), .ZN(n3636) );
  AOI22D0BWP12T U1733 ( .A1(write2_in[30]), .A2(n3263), .B1(n3262), .B2(r6[30]), .ZN(n3632) );
  AOI22D0BWP12T U1734 ( .A1(write2_in[29]), .A2(n3028), .B1(n3303), .B2(r3[29]), .ZN(n3629) );
  AOI22D0BWP12T U1735 ( .A1(write2_in[30]), .A2(n3273), .B1(n3272), .B2(r5[30]), .ZN(n3633) );
  INVD1BWP12T U1736 ( .I(r12[15]), .ZN(n1715) );
  INVD1BWP12T U1737 ( .I(r1[15]), .ZN(n1717) );
  OAI22D0BWP12T U1738 ( .A1(n1715), .A2(n3600), .B1(n3599), .B2(n1717), .ZN(
        n789) );
  BUFFXD8BWP12T U1739 ( .I(n1738), .Z(n3605) );
  INVD1BWP12T U1740 ( .I(n[3685]), .ZN(n1711) );
  INVD1BWP12T U1741 ( .I(r8[15]), .ZN(n2699) );
  OAI22D1BWP12T U1742 ( .A1(n3605), .A2(n1711), .B1(n3603), .B2(n2699), .ZN(
        n788) );
  INVD1BWP12T U1743 ( .I(lr[15]), .ZN(n2700) );
  INVD1BWP12T U1744 ( .I(r3[15]), .ZN(n1712) );
  INVD0BWP12T U1745 ( .I(pc_out[15]), .ZN(n785) );
  INVD1BWP12T U1746 ( .I(r6[15]), .ZN(n1705) );
  OAI22D1BWP12T U1747 ( .A1(n3612), .A2(n785), .B1(n3611), .B2(n1705), .ZN(
        n786) );
  INVD1BWP12T U1748 ( .I(r9[15]), .ZN(n1699) );
  INVD1BWP12T U1749 ( .I(r4[15]), .ZN(n1703) );
  INVD1BWP12T U1750 ( .I(r11[15]), .ZN(n1710) );
  BUFFXD12BWP12T U1751 ( .I(n1901), .Z(n3588) );
  INVD1BWP12T U1752 ( .I(r0[15]), .ZN(n1702) );
  BUFFXD8BWP12T U1753 ( .I(n1730), .Z(n1906) );
  AN4D4BWP12T U1754 ( .A1(n796), .A2(n794), .A3(n795), .A4(n793), .Z(n797) );
  AOI22D1BWP12T U1755 ( .A1(tmp1[27]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[27]), .ZN(n804) );
  INVD1BWP12T U1756 ( .I(r11[27]), .ZN(n3434) );
  INVD1BWP12T U1757 ( .I(r0[27]), .ZN(n3420) );
  OAI22D0BWP12T U1758 ( .A1(n3586), .A2(n3434), .B1(n1901), .B2(n3420), .ZN(
        n800) );
  INVD0BWP12T U1759 ( .I(r9[27]), .ZN(n798) );
  INVD1BWP12T U1760 ( .I(r4[27]), .ZN(n3421) );
  OAI22D1BWP12T U1761 ( .A1(n3584), .A2(n798), .B1(n3582), .B2(n3421), .ZN(
        n799) );
  AOI22D1BWP12T U1762 ( .A1(r5[27]), .A2(n3592), .B1(n3591), .B2(r10[27]), 
        .ZN(n802) );
  AOI22D1BWP12T U1763 ( .A1(r7[27]), .A2(n3524), .B1(n3593), .B2(r2[27]), .ZN(
        n801) );
  AN4XD1BWP12T U1764 ( .A1(n804), .A2(n803), .A3(n802), .A4(n801), .Z(n808) );
  INVD1BWP12T U1765 ( .I(r12[27]), .ZN(n3436) );
  INVD1BWP12T U1766 ( .I(r1[27]), .ZN(n3438) );
  OAI22D0BWP12T U1767 ( .A1(n3436), .A2(n3600), .B1(n3599), .B2(n3438), .ZN(
        n806) );
  INVD1BWP12T U1768 ( .I(n[3673]), .ZN(n3435) );
  INVD1BWP12T U1769 ( .I(r8[27]), .ZN(n3425) );
  INVD1BWP12T U1770 ( .I(lr[27]), .ZN(n3426) );
  BUFFD3BWP12T U1771 ( .I(n981), .Z(n3607) );
  INVD1BWP12T U1772 ( .I(r3[27]), .ZN(n3432) );
  TPOAI22D1BWP12T U1773 ( .A1(n3426), .A2(n3571), .B1(n3607), .B2(n3432), .ZN(
        n805) );
  INVD1BWP12T U1774 ( .I(r6[27]), .ZN(n3424) );
  INVD1BWP12T U1775 ( .I(n1973), .ZN(n812) );
  CKND0BWP12T U1776 ( .I(write2_in[21]), .ZN(n809) );
  INR2D1BWP12T U1777 ( .A1(n3393), .B1(n809), .ZN(n810) );
  TPAOI21D2BWP12T U1778 ( .A1(write1_in[21]), .A2(n1856), .B(n810), .ZN(n1977)
         );
  ND2D4BWP12T U1779 ( .A1(write1_in[22]), .A2(n3381), .ZN(n814) );
  CKND2D1BWP12T U1780 ( .A1(write2_in[22]), .A2(n3393), .ZN(n813) );
  ND2D4BWP12T U1781 ( .A1(n814), .A2(n813), .ZN(n1865) );
  TPND2D1BWP12T U1782 ( .A1(n3310), .A2(n3352), .ZN(n3313) );
  OR2D2BWP12T U1783 ( .A1(n3313), .A2(n3335), .Z(n821) );
  TPAOI31D1BWP12T U1784 ( .A1(n3335), .A2(n238), .A3(n3352), .B(n818), .ZN(
        n819) );
  OAI211D1BWP12T U1785 ( .A1(n822), .A2(n821), .B(n820), .C(n819), .ZN(n2193)
         );
  TPND2D1BWP12T U1786 ( .A1(n249), .A2(n3626), .ZN(n824) );
  AOI22D0BWP12T U1787 ( .A1(write2_in[30]), .A2(n3307), .B1(n3306), .B2(
        r11[30]), .ZN(n823) );
  ND2D2BWP12T U1788 ( .A1(n824), .A2(n823), .ZN(n2295) );
  TPND2D1BWP12T U1789 ( .A1(n249), .A2(n3211), .ZN(n826) );
  AOI22D0BWP12T U1790 ( .A1(write2_in[30]), .A2(n3213), .B1(n3212), .B2(r8[30]), .ZN(n825) );
  TPND2D1BWP12T U1791 ( .A1(n249), .A2(n3216), .ZN(n828) );
  AOI22D0BWP12T U1792 ( .A1(write2_in[30]), .A2(n3218), .B1(n3217), .B2(
        r12[30]), .ZN(n827) );
  TPND2D1BWP12T U1793 ( .A1(n249), .A2(n3234), .ZN(n830) );
  AOI22D0BWP12T U1794 ( .A1(write2_in[30]), .A2(n3236), .B1(n3235), .B2(lr[30]), .ZN(n829) );
  TPND2D1BWP12T U1795 ( .A1(n249), .A2(n3248), .ZN(n832) );
  AOI22D0BWP12T U1796 ( .A1(write2_in[30]), .A2(n3250), .B1(n3249), .B2(r9[30]), .ZN(n831) );
  TPND2D1BWP12T U1797 ( .A1(n3372), .A2(n3234), .ZN(n834) );
  AOI22D0BWP12T U1798 ( .A1(write2_in[29]), .A2(n3236), .B1(n3235), .B2(lr[29]), .ZN(n833) );
  ND2D1BWP12T U1799 ( .A1(n834), .A2(n833), .ZN(n2230) );
  TPND2D1BWP12T U1800 ( .A1(n3372), .A2(n3216), .ZN(n836) );
  AOI22D0BWP12T U1801 ( .A1(write2_in[29]), .A2(n3218), .B1(n3217), .B2(
        r12[29]), .ZN(n835) );
  ND2D1BWP12T U1802 ( .A1(n836), .A2(n835), .ZN(n2262) );
  TPND2D1BWP12T U1803 ( .A1(n3372), .A2(n3638), .ZN(n838) );
  AOI22D0BWP12T U1804 ( .A1(write2_in[29]), .A2(n3277), .B1(n3276), .B2(
        tmp1[29]), .ZN(n837) );
  ND2D1BWP12T U1805 ( .A1(n838), .A2(n837), .ZN(n2166) );
  TPND2D1BWP12T U1806 ( .A1(n3372), .A2(n3229), .ZN(n840) );
  AOI22D0BWP12T U1807 ( .A1(write2_in[29]), .A2(n3231), .B1(n3230), .B2(
        n[3671]), .ZN(n839) );
  TPND2D1BWP12T U1808 ( .A1(n840), .A2(n839), .ZN(spin[29]) );
  TPND2D1BWP12T U1809 ( .A1(n3372), .A2(n3248), .ZN(n842) );
  AOI22D0BWP12T U1810 ( .A1(write2_in[29]), .A2(n3250), .B1(n3249), .B2(r9[29]), .ZN(n841) );
  TPND2D1BWP12T U1811 ( .A1(n842), .A2(n841), .ZN(n2358) );
  CKND2D0BWP12T U1812 ( .A1(write1_in[13]), .A2(n3248), .ZN(n847) );
  AOI22D0BWP12T U1813 ( .A1(n2972), .A2(n3250), .B1(n3249), .B2(r9[13]), .ZN(
        n846) );
  CKND2D1BWP12T U1814 ( .A1(n847), .A2(n846), .ZN(n2342) );
  CKND2D0BWP12T U1815 ( .A1(write1_in[13]), .A2(n3626), .ZN(n849) );
  AOI22D0BWP12T U1816 ( .A1(n2972), .A2(n3307), .B1(n3306), .B2(r11[13]), .ZN(
        n848) );
  CKND2D1BWP12T U1817 ( .A1(n849), .A2(n848), .ZN(n2278) );
  CKND2D0BWP12T U1818 ( .A1(n42), .A2(n3627), .ZN(n851) );
  AOI22D0BWP12T U1819 ( .A1(n2972), .A2(n3298), .B1(n3297), .B2(r10[13]), .ZN(
        n850) );
  CKND2D1BWP12T U1820 ( .A1(n851), .A2(n850), .ZN(n2310) );
  CKND2D0BWP12T U1821 ( .A1(write1_in[13]), .A2(n3211), .ZN(n853) );
  AOI22D0BWP12T U1822 ( .A1(n2972), .A2(n3213), .B1(n3212), .B2(r8[13]), .ZN(
        n852) );
  CKND2D1BWP12T U1823 ( .A1(n853), .A2(n852), .ZN(n2374) );
  CKND2D0BWP12T U1824 ( .A1(write1_in[13]), .A2(n3216), .ZN(n855) );
  AOI22D0BWP12T U1825 ( .A1(n2972), .A2(n3218), .B1(n3217), .B2(r12[13]), .ZN(
        n854) );
  CKND2D1BWP12T U1826 ( .A1(n855), .A2(n854), .ZN(n2246) );
  CKND2D0BWP12T U1827 ( .A1(n42), .A2(n3241), .ZN(n857) );
  AOI22D0BWP12T U1828 ( .A1(n2972), .A2(n3243), .B1(n3242), .B2(r7[13]), .ZN(
        n856) );
  CKND2D1BWP12T U1829 ( .A1(n857), .A2(n856), .ZN(n2406) );
  CKND2D0BWP12T U1830 ( .A1(n42), .A2(n3229), .ZN(n859) );
  AOI22D0BWP12T U1831 ( .A1(n2972), .A2(n3231), .B1(n3230), .B2(n[3687]), .ZN(
        n858) );
  CKND2D1BWP12T U1832 ( .A1(n859), .A2(n858), .ZN(spin[13]) );
  CKND2D0BWP12T U1833 ( .A1(write1_in[13]), .A2(n3234), .ZN(n861) );
  AOI22D0BWP12T U1834 ( .A1(n2972), .A2(n3236), .B1(n3235), .B2(lr[13]), .ZN(
        n860) );
  CKND2D1BWP12T U1835 ( .A1(n861), .A2(n860), .ZN(n2214) );
  CKND2D0BWP12T U1836 ( .A1(write1_in[13]), .A2(n3638), .ZN(n863) );
  AOI22D0BWP12T U1837 ( .A1(n2972), .A2(n3277), .B1(n3276), .B2(tmp1[13]), 
        .ZN(n862) );
  CKND2D1BWP12T U1838 ( .A1(n863), .A2(n862), .ZN(n2150) );
  TPND2D0BWP12T U1839 ( .A1(write1_in[8]), .A2(n3638), .ZN(n865) );
  AOI22D0BWP12T U1840 ( .A1(n866), .A2(n3277), .B1(n3276), .B2(tmp1[8]), .ZN(
        n864) );
  CKND2D1BWP12T U1841 ( .A1(n865), .A2(n864), .ZN(n2145) );
  TPND2D0BWP12T U1842 ( .A1(write1_in[7]), .A2(n3229), .ZN(n870) );
  INVD0BWP12T U1843 ( .I(write2_in[7]), .ZN(n867) );
  NR2D1BWP12T U1844 ( .A1(n867), .A2(n2938), .ZN(n868) );
  RCAOI211D0BWP12T U1845 ( .A1(n3230), .A2(n[3693]), .B(n868), .C(reset), .ZN(
        n869) );
  CKND2D1BWP12T U1846 ( .A1(n870), .A2(n869), .ZN(spin[7]) );
  TPND2D0BWP12T U1847 ( .A1(write1_in[7]), .A2(n3248), .ZN(n872) );
  AOI22D0BWP12T U1848 ( .A1(write2_in[7]), .A2(n3250), .B1(n3249), .B2(r9[7]), 
        .ZN(n871) );
  CKND2D1BWP12T U1849 ( .A1(n872), .A2(n871), .ZN(n2336) );
  TPND2D0BWP12T U1850 ( .A1(write1_in[7]), .A2(n3623), .ZN(n874) );
  AOI22D0BWP12T U1851 ( .A1(write2_in[7]), .A2(n3281), .B1(n3280), .B2(r4[7]), 
        .ZN(n873) );
  CKND2D1BWP12T U1852 ( .A1(n874), .A2(n873), .ZN(n2496) );
  TPND2D0BWP12T U1853 ( .A1(write1_in[7]), .A2(n3622), .ZN(n876) );
  AOI22D0BWP12T U1854 ( .A1(write2_in[7]), .A2(n3273), .B1(n3272), .B2(r5[7]), 
        .ZN(n875) );
  CKND2D1BWP12T U1855 ( .A1(n876), .A2(n875), .ZN(n2464) );
  TPND2D0BWP12T U1856 ( .A1(write1_in[7]), .A2(n3234), .ZN(n878) );
  AOI22D0BWP12T U1857 ( .A1(write2_in[7]), .A2(n3236), .B1(n3235), .B2(lr[7]), 
        .ZN(n877) );
  CKND2D1BWP12T U1858 ( .A1(n878), .A2(n877), .ZN(n2208) );
  TPND2D0BWP12T U1859 ( .A1(write1_in[7]), .A2(n3216), .ZN(n880) );
  AOI22D0BWP12T U1860 ( .A1(write2_in[7]), .A2(n3218), .B1(n3217), .B2(r12[7]), 
        .ZN(n879) );
  CKND2D1BWP12T U1861 ( .A1(n880), .A2(n879), .ZN(n2240) );
  TPND2D0BWP12T U1862 ( .A1(write1_in[7]), .A2(n3211), .ZN(n882) );
  AOI22D0BWP12T U1863 ( .A1(write2_in[7]), .A2(n3213), .B1(n3212), .B2(r8[7]), 
        .ZN(n881) );
  CKND2D1BWP12T U1864 ( .A1(n882), .A2(n881), .ZN(n2368) );
  TPND2D0BWP12T U1865 ( .A1(write1_in[7]), .A2(n3241), .ZN(n884) );
  AOI22D0BWP12T U1866 ( .A1(write2_in[7]), .A2(n3243), .B1(n3242), .B2(r7[7]), 
        .ZN(n883) );
  CKND2D1BWP12T U1867 ( .A1(n884), .A2(n883), .ZN(n2400) );
  TPND2D0BWP12T U1868 ( .A1(write1_in[7]), .A2(n3289), .ZN(n886) );
  AOI22D0BWP12T U1869 ( .A1(write2_in[7]), .A2(n3291), .B1(n3290), .B2(r1[7]), 
        .ZN(n885) );
  CKND2D1BWP12T U1870 ( .A1(n886), .A2(n885), .ZN(n2592) );
  TPND2D0BWP12T U1871 ( .A1(write1_in[7]), .A2(n3638), .ZN(n888) );
  AOI22D0BWP12T U1872 ( .A1(write2_in[7]), .A2(n3277), .B1(n3276), .B2(tmp1[7]), .ZN(n887) );
  CKND2D1BWP12T U1873 ( .A1(n888), .A2(n887), .ZN(n2144) );
  TPND2D0BWP12T U1874 ( .A1(write1_in[1]), .A2(n3216), .ZN(n890) );
  AOI22D0BWP12T U1875 ( .A1(n892), .A2(n3218), .B1(n3217), .B2(r12[1]), .ZN(
        n889) );
  CKND2D1BWP12T U1876 ( .A1(n890), .A2(n889), .ZN(n2234) );
  AOI22D0BWP12T U1877 ( .A1(write2_in[29]), .A2(n3307), .B1(n3306), .B2(
        r11[29]), .ZN(n3630) );
  AOI22D0BWP12T U1878 ( .A1(write2_in[30]), .A2(n3028), .B1(n3303), .B2(r3[30]), .ZN(n3634) );
  AOI22D0BWP12T U1879 ( .A1(write2_in[29]), .A2(n3298), .B1(n3297), .B2(
        r10[29]), .ZN(n3631) );
  AOI22D1BWP12T U1880 ( .A1(r9[18]), .A2(n3471), .B1(n3472), .B2(tmp1[18]), 
        .ZN(n893) );
  IOA21D1BWP12T U1881 ( .A1(n3474), .A2(r2[18]), .B(n893), .ZN(n896) );
  INVD1BWP12T U1882 ( .I(r4[18]), .ZN(n1759) );
  INVD1BWP12T U1883 ( .I(r0[18]), .ZN(n1761) );
  OAI22D1BWP12T U1884 ( .A1(n3448), .A2(n1759), .B1(n3476), .B2(n1761), .ZN(
        n894) );
  INVD1BWP12T U1885 ( .I(n894), .ZN(n895) );
  IND2D2BWP12T U1886 ( .A1(n896), .B1(n895), .ZN(n901) );
  INVD1BWP12T U1887 ( .I(lr[18]), .ZN(n1772) );
  INVD1BWP12T U1888 ( .I(r8[18]), .ZN(n2093) );
  OAI22D1BWP12T U1889 ( .A1(n3478), .A2(n1772), .B1(n3477), .B2(n2093), .ZN(
        n899) );
  INVD1BWP12T U1890 ( .I(r6[18]), .ZN(n1773) );
  INVD1BWP12T U1891 ( .I(r10[18]), .ZN(n897) );
  OR2XD2BWP12T U1892 ( .A1(n899), .A2(n898), .Z(n900) );
  INVD1BWP12T U1893 ( .I(n[3682]), .ZN(n1770) );
  INVD1BWP12T U1894 ( .I(r11[18]), .ZN(n1762) );
  TPOAI22D1BWP12T U1895 ( .A1(n3491), .A2(n1770), .B1(n1762), .B2(n3490), .ZN(
        n904) );
  INVD1BWP12T U1896 ( .I(r5[18]), .ZN(n902) );
  INVD1BWP12T U1897 ( .I(r3[18]), .ZN(n1771) );
  INVD1BWP12T U1898 ( .I(r7[18]), .ZN(n905) );
  INVD1BWP12T U1899 ( .I(r1[18]), .ZN(n1769) );
  INVD1BWP12T U1900 ( .I(r12[18]), .ZN(n2094) );
  OAI22D1BWP12T U1901 ( .A1(n1769), .A2(n3463), .B1(n3437), .B2(n2094), .ZN(
        n906) );
  OR2XD2BWP12T U1902 ( .A1(n907), .A2(n906), .Z(n908) );
  AOI22D0BWP12T U1903 ( .A1(write2_in[30]), .A2(n3298), .B1(n3297), .B2(
        r10[30]), .ZN(n3637) );
  AOI22D1BWP12T U1904 ( .A1(r9[19]), .A2(n3471), .B1(n3472), .B2(tmp1[19]), 
        .ZN(n912) );
  INVD1BWP12T U1905 ( .I(r4[19]), .ZN(n3581) );
  INVD1BWP12T U1906 ( .I(r0[19]), .ZN(n3587) );
  TPOAI22D1BWP12T U1907 ( .A1(n3448), .A2(n3581), .B1(n3476), .B2(n3587), .ZN(
        n916) );
  INVD1BWP12T U1908 ( .I(lr[19]), .ZN(n3609) );
  INVD1BWP12T U1909 ( .I(r8[19]), .ZN(n3602) );
  INVD1BWP12T U1910 ( .I(r6[19]), .ZN(n3610) );
  INVD1BWP12T U1911 ( .I(r10[19]), .ZN(n913) );
  INVD1BWP12T U1912 ( .I(r5[19]), .ZN(n918) );
  INVD1BWP12T U1913 ( .I(r3[19]), .ZN(n3606) );
  OAI22D2BWP12T U1914 ( .A1(n3489), .A2(n918), .B1(n3606), .B2(n3488), .ZN(
        n920) );
  INVD1BWP12T U1915 ( .I(n[3681]), .ZN(n3604) );
  INVD1BWP12T U1916 ( .I(r11[19]), .ZN(n3585) );
  TPOAI22D1BWP12T U1917 ( .A1(n3491), .A2(n3604), .B1(n3490), .B2(n3585), .ZN(
        n919) );
  INVD1BWP12T U1918 ( .I(r7[19]), .ZN(n921) );
  OAI22D2BWP12T U1919 ( .A1(n3487), .A2(n921), .B1(n3486), .B2(n3641), .ZN(
        n923) );
  INVD1BWP12T U1920 ( .I(r12[19]), .ZN(n3601) );
  INVD1BWP12T U1921 ( .I(r1[19]), .ZN(n3598) );
  TPOAI22D1BWP12T U1922 ( .A1(n3492), .A2(n3601), .B1(n3463), .B2(n3598), .ZN(
        n922) );
  OR2XD4BWP12T U1923 ( .A1(n923), .A2(n922), .Z(n924) );
  AOI22D1BWP12T U1924 ( .A1(tmp1[11]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[11]), .ZN(n937) );
  AOI22D1BWP12T U1925 ( .A1(n1906), .A2(r2[11]), .B1(n3524), .B2(r7[11]), .ZN(
        n936) );
  INVD0BWP12T U1926 ( .I(r9[11]), .ZN(n929) );
  CKND1BWP12T U1927 ( .I(r4[11]), .ZN(n928) );
  OAI22D1BWP12T U1928 ( .A1(n3584), .A2(n929), .B1(n3582), .B2(n928), .ZN(n933) );
  CKND0BWP12T U1929 ( .I(r11[11]), .ZN(n931) );
  INVD1BWP12T U1930 ( .I(r0[11]), .ZN(n930) );
  TPNR2D1BWP12T U1931 ( .A1(n933), .A2(n932), .ZN(n935) );
  AN4D4BWP12T U1932 ( .A1(n937), .A2(n936), .A3(n935), .A4(n934), .Z(n949) );
  INVD1BWP12T U1933 ( .I(n[3689]), .ZN(n2738) );
  INVD1BWP12T U1934 ( .I(r8[11]), .ZN(n938) );
  INVD0BWP12T U1935 ( .I(lr[11]), .ZN(n939) );
  INVD1BWP12T U1936 ( .I(r3[11]), .ZN(n1652) );
  OAI22D1BWP12T U1937 ( .A1(n939), .A2(n1884), .B1(n1913), .B2(n1652), .ZN(
        n940) );
  OR2XD2BWP12T U1938 ( .A1(n941), .A2(n940), .Z(n947) );
  INVD1BWP12T U1939 ( .I(r12[11]), .ZN(n2737) );
  INVD1BWP12T U1940 ( .I(r1[11]), .ZN(n2969) );
  OAI22D1BWP12T U1941 ( .A1(n2737), .A2(n3600), .B1(n3599), .B2(n2969), .ZN(
        n945) );
  INVD1BWP12T U1942 ( .I(pc_out[11]), .ZN(n943) );
  INVD1BWP12T U1943 ( .I(r6[11]), .ZN(n942) );
  OR2XD2BWP12T U1944 ( .A1(n945), .A2(n944), .Z(n946) );
  TPNR2D2BWP12T U1945 ( .A1(n947), .A2(n946), .ZN(n948) );
  ND2D4BWP12T U1946 ( .A1(n949), .A2(n948), .ZN(regB_out[11]) );
  AOI22D1BWP12T U1947 ( .A1(r9[0]), .A2(n3471), .B1(n3472), .B2(tmp1[0]), .ZN(
        n950) );
  IOA21D1BWP12T U1948 ( .A1(n3474), .A2(r2[0]), .B(n950), .ZN(n955) );
  INVD1P75BWP12T U1949 ( .I(r0[0]), .ZN(n970) );
  ND2D1BWP12T U1950 ( .A1(n3475), .A2(r4[0]), .ZN(n951) );
  OAI21D1BWP12T U1951 ( .A1(n3476), .A2(n970), .B(n951), .ZN(n954) );
  INVD1BWP12T U1952 ( .I(r10[0]), .ZN(n2664) );
  INVD1P75BWP12T U1953 ( .I(r6[0]), .ZN(n986) );
  INVD1BWP12T U1954 ( .I(lr[0]), .ZN(n2665) );
  INVD1P75BWP12T U1955 ( .I(r8[0]), .ZN(n979) );
  TPOAI22D1BWP12T U1956 ( .A1(n3478), .A2(n2665), .B1(n3477), .B2(n979), .ZN(
        n952) );
  NR4D1BWP12T U1957 ( .A1(n955), .A2(n954), .A3(n953), .A4(n952), .ZN(n964) );
  INVD1P75BWP12T U1958 ( .I(n[3700]), .ZN(n978) );
  INVD1P75BWP12T U1959 ( .I(r11[0]), .ZN(n971) );
  TPOAI22D1BWP12T U1960 ( .A1(n3491), .A2(n978), .B1(n971), .B2(n3490), .ZN(
        n962) );
  INVD1BWP12T U1961 ( .I(r5[0]), .ZN(n956) );
  INVD1BWP12T U1962 ( .I(r3[0]), .ZN(n980) );
  INVD1BWP12T U1963 ( .I(r12[0]), .ZN(n984) );
  INVD1BWP12T U1964 ( .I(r1[0]), .ZN(n985) );
  TPOAI22D1BWP12T U1965 ( .A1(n3492), .A2(n984), .B1(n3463), .B2(n985), .ZN(
        n959) );
  NR4D1BWP12T U1966 ( .A1(n962), .A2(n961), .A3(n960), .A4(n959), .ZN(n963) );
  ND2D3BWP12T U1967 ( .A1(n3591), .A2(r10[0]), .ZN(n967) );
  TPAOI22D2BWP12T U1968 ( .A1(n3524), .A2(r7[0]), .B1(n1730), .B2(r2[0]), .ZN(
        n966) );
  ND2D3BWP12T U1969 ( .A1(n295), .A2(tmp1[0]), .ZN(n965) );
  ND3D2BWP12T U1970 ( .A1(n967), .A2(n966), .A3(n965), .ZN(n976) );
  INVD1BWP12T U1971 ( .I(r9[0]), .ZN(n969) );
  INVD1BWP12T U1972 ( .I(r4[0]), .ZN(n968) );
  TPOAI22D4BWP12T U1973 ( .A1(n3586), .A2(n971), .B1(n3588), .B2(n970), .ZN(
        n972) );
  CKND2BWP12T U1974 ( .I(n974), .ZN(n975) );
  INR3XD2BWP12T U1975 ( .A1(n977), .B1(n976), .B2(n975), .ZN(n992) );
  TPOAI22D2BWP12T U1976 ( .A1(n3603), .A2(n979), .B1(n1738), .B2(n978), .ZN(
        n983) );
  OAI22D1BWP12T U1977 ( .A1(n2665), .A2(n1394), .B1(n981), .B2(n980), .ZN(n982) );
  TPOAI22D1BWP12T U1978 ( .A1(n985), .A2(n3599), .B1(n3600), .B2(n984), .ZN(
        n989) );
  INVD1BWP12T U1979 ( .I(pc_out[0]), .ZN(n987) );
  TPOAI22D1BWP12T U1980 ( .A1(n3612), .A2(n987), .B1(n3611), .B2(n986), .ZN(
        n988) );
  TPNR3D4BWP12T U1981 ( .A1(n990), .A2(n989), .A3(n988), .ZN(n991) );
  IOA21D1BWP12T U1982 ( .A1(n3474), .A2(r2[29]), .B(n993), .ZN(n997) );
  INVD1BWP12T U1983 ( .I(r4[29]), .ZN(n3558) );
  INVD1BWP12T U1984 ( .I(r0[29]), .ZN(n3560) );
  OAI22D1BWP12T U1985 ( .A1(n3448), .A2(n3558), .B1(n3476), .B2(n3560), .ZN(
        n996) );
  INVD1BWP12T U1986 ( .I(lr[29]), .ZN(n3572) );
  INVD1BWP12T U1987 ( .I(r8[29]), .ZN(n3569) );
  OAI22D0BWP12T U1988 ( .A1(n3478), .A2(n3572), .B1(n3477), .B2(n3569), .ZN(
        n995) );
  INVD1BWP12T U1989 ( .I(r6[29]), .ZN(n3573) );
  OAI22D1BWP12T U1990 ( .A1(n3481), .A2(n3573), .B1(n3649), .B2(n3422), .ZN(
        n994) );
  NR4D0BWP12T U1991 ( .A1(n997), .A2(n996), .A3(n995), .A4(n994), .ZN(n1005)
         );
  INVD1BWP12T U1992 ( .I(r7[29]), .ZN(n998) );
  OAI22D0BWP12T U1993 ( .A1(n3487), .A2(n998), .B1(n3486), .B2(n3650), .ZN(
        n1003) );
  INVD1BWP12T U1994 ( .I(r5[29]), .ZN(n999) );
  OAI22D1BWP12T U1995 ( .A1(n3489), .A2(n999), .B1(n3651), .B2(n3488), .ZN(
        n1002) );
  INVD1BWP12T U1996 ( .I(n[3671]), .ZN(n3570) );
  OAI22D1BWP12T U1997 ( .A1(n3491), .A2(n3570), .B1(n3652), .B2(n3490), .ZN(
        n1001) );
  INVD1BWP12T U1998 ( .I(r1[29]), .ZN(n3568) );
  INVD1BWP12T U1999 ( .I(r12[29]), .ZN(n3567) );
  OAI22D0BWP12T U2000 ( .A1(n3568), .A2(n3463), .B1(n3437), .B2(n3567), .ZN(
        n1000) );
  NR4D0BWP12T U2001 ( .A1(n1003), .A2(n1002), .A3(n1001), .A4(n1000), .ZN(
        n1004) );
  AOI22D1BWP12T U2002 ( .A1(r9[25]), .A2(n3471), .B1(n3472), .B2(tmp1[25]), 
        .ZN(n1006) );
  IOA21D1BWP12T U2003 ( .A1(n3474), .A2(r2[25]), .B(n1006), .ZN(n1011) );
  INVD1BWP12T U2004 ( .I(r4[25]), .ZN(n3499) );
  INVD1BWP12T U2005 ( .I(r0[25]), .ZN(n3501) );
  INVD1BWP12T U2006 ( .I(lr[25]), .ZN(n3514) );
  INVD1BWP12T U2007 ( .I(r8[25]), .ZN(n3511) );
  OAI22D1BWP12T U2008 ( .A1(n3478), .A2(n3514), .B1(n3477), .B2(n3511), .ZN(
        n1009) );
  INVD1BWP12T U2009 ( .I(r6[25]), .ZN(n3515) );
  INVD1BWP12T U2010 ( .I(r10[25]), .ZN(n1007) );
  TPOAI22D1BWP12T U2011 ( .A1(n3481), .A2(n3515), .B1(n3422), .B2(n1007), .ZN(
        n1008) );
  INVD1BWP12T U2012 ( .I(r5[25]), .ZN(n1012) );
  INVD1BWP12T U2013 ( .I(r3[25]), .ZN(n3513) );
  OAI22D1BWP12T U2014 ( .A1(n3489), .A2(n1012), .B1(n3513), .B2(n3488), .ZN(
        n1015) );
  INVD1BWP12T U2015 ( .I(n[3675]), .ZN(n3512) );
  INVD1BWP12T U2016 ( .I(r11[25]), .ZN(n3502) );
  OAI22D1BWP12T U2017 ( .A1(n3491), .A2(n3512), .B1(n3502), .B2(n3490), .ZN(
        n1014) );
  INVD1BWP12T U2018 ( .I(r1[25]), .ZN(n3509) );
  INVD1BWP12T U2019 ( .I(r12[25]), .ZN(n3510) );
  NR4D1BWP12T U2020 ( .A1(n1016), .A2(n1015), .A3(n1014), .A4(n1013), .ZN(
        n1017) );
  AOI22D1BWP12T U2021 ( .A1(tmp1[10]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[10]), .ZN(n1028) );
  CKND0BWP12T U2022 ( .I(r9[10]), .ZN(n1020) );
  INVD1BWP12T U2023 ( .I(r4[10]), .ZN(n1019) );
  OAI22D1BWP12T U2024 ( .A1(n3584), .A2(n1020), .B1(n3582), .B2(n1019), .ZN(
        n1024) );
  CKND1BWP12T U2025 ( .I(r11[10]), .ZN(n1022) );
  INVD1BWP12T U2026 ( .I(r0[10]), .ZN(n1021) );
  OAI22D1BWP12T U2027 ( .A1(n3586), .A2(n1022), .B1(n3588), .B2(n1021), .ZN(
        n1023) );
  RCAOI22D2BWP12T U2028 ( .A1(r5[10]), .A2(n3592), .B1(n3591), .B2(r10[10]), 
        .ZN(n1026) );
  AOI22D2BWP12T U2029 ( .A1(r7[10]), .A2(n1327), .B1(n1906), .B2(r2[10]), .ZN(
        n1025) );
  AN4XD1BWP12T U2030 ( .A1(n1028), .A2(n1027), .A3(n1026), .A4(n1025), .Z(
        n1040) );
  INVD1BWP12T U2031 ( .I(r12[10]), .ZN(n1029) );
  OAI22D1BWP12T U2032 ( .A1(n1029), .A2(n3600), .B1(n3599), .B2(n2931), .ZN(
        n1038) );
  INVD1BWP12T U2033 ( .I(n[3690]), .ZN(n2118) );
  INVD1BWP12T U2034 ( .I(r8[10]), .ZN(n1030) );
  OAI22D1BWP12T U2035 ( .A1(n3605), .A2(n2118), .B1(n3603), .B2(n1030), .ZN(
        n1037) );
  INVD1BWP12T U2036 ( .I(lr[10]), .ZN(n1032) );
  OAI22D1BWP12T U2037 ( .A1(n1032), .A2(n1884), .B1(n1913), .B2(n1031), .ZN(
        n1036) );
  INVD1BWP12T U2038 ( .I(pc_out[10]), .ZN(n1034) );
  INVD1BWP12T U2039 ( .I(r6[10]), .ZN(n1033) );
  NR4D1BWP12T U2040 ( .A1(n1038), .A2(n1037), .A3(n1036), .A4(n1035), .ZN(
        n1039) );
  INVD1BWP12T U2041 ( .I(r6[22]), .ZN(n1825) );
  OAI22D1BWP12T U2042 ( .A1(n3612), .A2(n3643), .B1(n3611), .B2(n1825), .ZN(
        n1043) );
  INVD1BWP12T U2043 ( .I(r8[22]), .ZN(n2714) );
  OAI22D1BWP12T U2044 ( .A1(n3605), .A2(n2715), .B1(n3603), .B2(n2714), .ZN(
        n1042) );
  INVD1BWP12T U2045 ( .I(r12[22]), .ZN(n1830) );
  INVD1BWP12T U2046 ( .I(r1[22]), .ZN(n1831) );
  OAI22D0BWP12T U2047 ( .A1(n1830), .A2(n3600), .B1(n3599), .B2(n1831), .ZN(
        n1041) );
  OR3XD2BWP12T U2048 ( .A1(n1043), .A2(n1042), .A3(n1041), .Z(n1045) );
  INVD1BWP12T U2049 ( .I(lr[22]), .ZN(n2713) );
  INVD1BWP12T U2050 ( .I(r3[22]), .ZN(n1832) );
  OAI22D0BWP12T U2051 ( .A1(n3571), .A2(n2713), .B1(n1740), .B2(n1832), .ZN(
        n1044) );
  TPNR2D2BWP12T U2052 ( .A1(n1045), .A2(n1044), .ZN(n1054) );
  AOI22D1BWP12T U2053 ( .A1(tmp1[22]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[22]), .ZN(n1052) );
  INVD0BWP12T U2054 ( .I(r9[22]), .ZN(n1046) );
  INVD1BWP12T U2055 ( .I(r4[22]), .ZN(n1823) );
  OAI22D1BWP12T U2056 ( .A1(n3584), .A2(n1046), .B1(n3582), .B2(n1823), .ZN(
        n1048) );
  INVD1BWP12T U2057 ( .I(r11[22]), .ZN(n2712) );
  INVD1BWP12T U2058 ( .I(r0[22]), .ZN(n1822) );
  OAI22D1BWP12T U2059 ( .A1(n3586), .A2(n2712), .B1(n3588), .B2(n1822), .ZN(
        n1047) );
  NR2D1BWP12T U2060 ( .A1(n1048), .A2(n1047), .ZN(n1051) );
  AOI22D1BWP12T U2061 ( .A1(r7[22]), .A2(n3524), .B1(n3593), .B2(r2[22]), .ZN(
        n1050) );
  AOI22D1BWP12T U2062 ( .A1(r5[22]), .A2(n3592), .B1(n3591), .B2(r10[22]), 
        .ZN(n1049) );
  AN4XD1BWP12T U2063 ( .A1(n1052), .A2(n1051), .A3(n1050), .A4(n1049), .Z(
        n1053) );
  TPND2D2BWP12T U2064 ( .A1(n1054), .A2(n1053), .ZN(regB_out[22]) );
  AOI22D1BWP12T U2065 ( .A1(tmp1[16]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[16]), .ZN(n1063) );
  INVD0BWP12T U2066 ( .I(r9[16]), .ZN(n1055) );
  CKND0BWP12T U2067 ( .I(r11[16]), .ZN(n1057) );
  CKND1BWP12T U2068 ( .I(r0[16]), .ZN(n1056) );
  OAI22D1BWP12T U2069 ( .A1(n3586), .A2(n1057), .B1(n3588), .B2(n1056), .ZN(
        n1058) );
  NR2D1BWP12T U2070 ( .A1(n1059), .A2(n1058), .ZN(n1062) );
  AOI22D1BWP12T U2071 ( .A1(r5[16]), .A2(n3592), .B1(n3591), .B2(r10[16]), 
        .ZN(n1061) );
  AOI22D1BWP12T U2072 ( .A1(r7[16]), .A2(n1327), .B1(n1906), .B2(r2[16]), .ZN(
        n1060) );
  AN4XD1BWP12T U2073 ( .A1(n1062), .A2(n1060), .A3(n1061), .A4(n1063), .Z(
        n1070) );
  INVD1BWP12T U2074 ( .I(r12[16]), .ZN(n2866) );
  INVD0BWP12T U2075 ( .I(lr[16]), .ZN(n1064) );
  INVD1BWP12T U2076 ( .I(r3[16]), .ZN(n1226) );
  OAI22D1BWP12T U2077 ( .A1(n1064), .A2(n1884), .B1(n1913), .B2(n1226), .ZN(
        n1066) );
  NR4D0BWP12T U2078 ( .A1(n1068), .A2(n1067), .A3(n1066), .A4(n1065), .ZN(
        n1069) );
  CKND2D2BWP12T U2079 ( .A1(n1070), .A2(n1069), .ZN(regB_out[16]) );
  AOI22D1BWP12T U2080 ( .A1(tmp1[9]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[9]), .ZN(n1077) );
  CKND0BWP12T U2081 ( .I(r11[9]), .ZN(n1073) );
  CKND1BWP12T U2082 ( .I(r0[9]), .ZN(n1072) );
  AOI22D1BWP12T U2083 ( .A1(r5[9]), .A2(n3592), .B1(n3591), .B2(r10[9]), .ZN(
        n1075) );
  AOI22D1BWP12T U2084 ( .A1(r7[9]), .A2(n1327), .B1(n1906), .B2(r2[9]), .ZN(
        n1074) );
  AN4XD1BWP12T U2085 ( .A1(n1074), .A2(n1076), .A3(n1075), .A4(n1077), .Z(
        n1086) );
  INVD1BWP12T U2086 ( .I(r12[9]), .ZN(n1297) );
  INVD1BWP12T U2087 ( .I(r1[9]), .ZN(n2923) );
  OAI22D1BWP12T U2088 ( .A1(n1297), .A2(n3600), .B1(n3599), .B2(n2923), .ZN(
        n1084) );
  INVD1BWP12T U2089 ( .I(n[3691]), .ZN(n1298) );
  INVD1BWP12T U2090 ( .I(r8[9]), .ZN(n2039) );
  OAI22D1BWP12T U2091 ( .A1(n3605), .A2(n1298), .B1(n3603), .B2(n2039), .ZN(
        n1083) );
  INVD1BWP12T U2092 ( .I(lr[9]), .ZN(n1078) );
  INVD1BWP12T U2093 ( .I(r3[9]), .ZN(n1279) );
  OAI22D1BWP12T U2094 ( .A1(n1078), .A2(n1884), .B1(n1913), .B2(n1279), .ZN(
        n1082) );
  INVD1BWP12T U2095 ( .I(pc_out[9]), .ZN(n1080) );
  INVD1BWP12T U2096 ( .I(r6[9]), .ZN(n1079) );
  INVD1BWP12T U2097 ( .I(lr[28]), .ZN(n2677) );
  INVD1BWP12T U2098 ( .I(r8[28]), .ZN(n1804) );
  OAI22D0BWP12T U2099 ( .A1(n3478), .A2(n2677), .B1(n3477), .B2(n1804), .ZN(
        n1089) );
  TPNR2D1BWP12T U2100 ( .A1(n1089), .A2(n1088), .ZN(n1102) );
  INVD1BWP12T U2101 ( .I(r6[28]), .ZN(n1807) );
  INVD1BWP12T U2102 ( .I(r10[28]), .ZN(n1090) );
  INVD1BWP12T U2103 ( .I(r0[28]), .ZN(n1813) );
  ND2D1BWP12T U2104 ( .A1(n3475), .A2(r4[28]), .ZN(n1091) );
  TPOAI21D1BWP12T U2105 ( .A1(n3476), .A2(n1813), .B(n1091), .ZN(n1092) );
  INVD1BWP12T U2106 ( .I(r7[28]), .ZN(n1094) );
  INVD1BWP12T U2107 ( .I(r5[28]), .ZN(n1095) );
  INVD1BWP12T U2108 ( .I(r3[28]), .ZN(n1806) );
  INVD1BWP12T U2109 ( .I(n[3672]), .ZN(n1805) );
  INVD1BWP12T U2110 ( .I(r11[28]), .ZN(n1814) );
  OAI22D1BWP12T U2111 ( .A1(n3491), .A2(n1805), .B1(n1814), .B2(n3490), .ZN(
        n1099) );
  INVD1BWP12T U2112 ( .I(r1[28]), .ZN(n1803) );
  INVD1BWP12T U2113 ( .I(r12[28]), .ZN(n2676) );
  OAI22D1BWP12T U2114 ( .A1(n1803), .A2(n3463), .B1(n3492), .B2(n2676), .ZN(
        n1098) );
  TPNR2D1BWP12T U2115 ( .A1(n1099), .A2(n1098), .ZN(n1100) );
  INVD1BWP12T U2116 ( .I(r5[13]), .ZN(n1103) );
  INVD1BWP12T U2117 ( .I(r3[13]), .ZN(n1537) );
  TPOAI22D1BWP12T U2118 ( .A1(n3489), .A2(n1103), .B1(n1537), .B2(n3488), .ZN(
        n1109) );
  INVD1BWP12T U2119 ( .I(n[3687]), .ZN(n1536) );
  INVD1BWP12T U2120 ( .I(r11[13]), .ZN(n1526) );
  TPOAI22D1BWP12T U2121 ( .A1(n3491), .A2(n1536), .B1(n3490), .B2(n1526), .ZN(
        n1108) );
  INVD1BWP12T U2122 ( .I(r7[13]), .ZN(n1104) );
  INVD1BWP12T U2123 ( .I(pc_out[13]), .ZN(n1539) );
  INVD1BWP12T U2124 ( .I(r1[13]), .ZN(n1533) );
  NR4D2BWP12T U2125 ( .A1(n1109), .A2(n1107), .A3(n1108), .A4(n1106), .ZN(
        n1118) );
  CKND2D2BWP12T U2126 ( .A1(n1111), .A2(n1110), .ZN(n1116) );
  INVD1BWP12T U2127 ( .I(r4[13]), .ZN(n1523) );
  INVD1BWP12T U2128 ( .I(r0[13]), .ZN(n1525) );
  INVD1BWP12T U2129 ( .I(lr[13]), .ZN(n2845) );
  INVD1BWP12T U2130 ( .I(r8[13]), .ZN(n1535) );
  INVD1BWP12T U2131 ( .I(r6[13]), .ZN(n1538) );
  INVD1BWP12T U2132 ( .I(r10[13]), .ZN(n1112) );
  TPOAI22D2BWP12T U2133 ( .A1(n3481), .A2(n1538), .B1(n3479), .B2(n1112), .ZN(
        n1113) );
  NR4D2BWP12T U2134 ( .A1(n1116), .A2(n1115), .A3(n1114), .A4(n1113), .ZN(
        n1117) );
  ND2D1BWP12T U2135 ( .A1(write1_in[23]), .A2(n3381), .ZN(n1125) );
  CKND0BWP12T U2136 ( .I(write2_in[27]), .ZN(n1119) );
  NR2XD0BWP12T U2137 ( .A1(n1119), .A2(n3381), .ZN(n3355) );
  CKND2D0BWP12T U2138 ( .A1(write2_in[26]), .A2(write2_in[24]), .ZN(n1120) );
  TPNR2D0BWP12T U2139 ( .A1(n1121), .A2(n1120), .ZN(n1122) );
  ND2D1BWP12T U2140 ( .A1(n3355), .A2(n1122), .ZN(n1123) );
  TPOAI31D4BWP12T U2141 ( .A1(n1125), .A2(n43), .A3(n1124), .B(n1123), .ZN(
        n3378) );
  TPND2D1BWP12T U2142 ( .A1(n3377), .A2(n3378), .ZN(n1126) );
  INVD1BWP12T U2143 ( .I(n1126), .ZN(n1139) );
  CKND0BWP12T U2144 ( .I(write2_in[30]), .ZN(n1127) );
  NR2D1BWP12T U2145 ( .A1(n1127), .A2(n3381), .ZN(n1134) );
  INVD1P75BWP12T U2146 ( .I(n3401), .ZN(n1130) );
  INVD1BWP12T U2147 ( .I(n3363), .ZN(n3388) );
  AOI21D0BWP12T U2148 ( .A1(n3379), .A2(n3363), .B(n3394), .ZN(n1128) );
  NR2XD1BWP12T U2149 ( .A1(n1130), .A2(n1129), .ZN(n1138) );
  CKND0BWP12T U2150 ( .I(n1134), .ZN(n1132) );
  AOI21D0BWP12T U2151 ( .A1(n3379), .A2(n1132), .B(n3394), .ZN(n1133) );
  TPNR2D0BWP12T U2152 ( .A1(n3399), .A2(n3659), .ZN(n1135) );
  TPAOI21D0BWP12T U2153 ( .A1(next_pc_in[30]), .A2(n3398), .B(n1135), .ZN(
        n1136) );
  TPAOI31D1BWP12T U2154 ( .A1(n1139), .A2(n1138), .A3(n3366), .B(n1137), .ZN(
        n1143) );
  INVD1BWP12T U2155 ( .I(n3366), .ZN(n1141) );
  ND2D1BWP12T U2156 ( .A1(n44), .A2(n3378), .ZN(n3403) );
  ND2D2BWP12T U2157 ( .A1(n1143), .A2(n1142), .ZN(n2199) );
  INVD1BWP12T U2158 ( .I(r2[17]), .ZN(n1144) );
  INVD1BWP12T U2159 ( .I(r4[17]), .ZN(n1873) );
  INR2D2BWP12T U2160 ( .A1(r4[17]), .B1(n3448), .ZN(n1149) );
  INVD1BWP12T U2161 ( .I(r3[17]), .ZN(n1883) );
  TPND2D4BWP12T U2162 ( .A1(n1950), .A2(r7[17]), .ZN(n1145) );
  TPOAI21D1BWP12T U2163 ( .A1(n1883), .A2(n3488), .B(n1145), .ZN(n1148) );
  IOA21D2BWP12T U2164 ( .A1(n1952), .A2(r12[17]), .B(n1146), .ZN(n1147) );
  ND2D1BWP12T U2165 ( .A1(n3471), .A2(r9[17]), .ZN(n1155) );
  INR2D1BWP12T U2166 ( .A1(r11[17]), .B1(n3490), .ZN(n1154) );
  INVD1BWP12T U2167 ( .I(lr[17]), .ZN(n2795) );
  ND2D4BWP12T U2168 ( .A1(n235), .A2(r0[17]), .ZN(n1152) );
  ND2D1BWP12T U2169 ( .A1(n1642), .A2(r6[17]), .ZN(n1162) );
  AN2XD2BWP12T U2170 ( .A1(n1924), .A2(r8[17]), .Z(n1161) );
  INVD1BWP12T U2171 ( .I(r10[17]), .ZN(n1159) );
  AOI22D1BWP12T U2172 ( .A1(n1951), .A2(r1[17]), .B1(n1156), .B2(tmp1[17]), 
        .ZN(n1158) );
  ND2D1BWP12T U2173 ( .A1(n1945), .A2(pc_out[17]), .ZN(n1157) );
  OAI211D1BWP12T U2174 ( .A1(n1159), .A2(n3422), .B(n1158), .C(n1157), .ZN(
        n1160) );
  INR3D2BWP12T U2175 ( .A1(n1162), .B1(n1161), .B2(n1160), .ZN(n1163) );
  AOI22D1BWP12T U2176 ( .A1(tmp1[8]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[8]), .ZN(n1174) );
  AOI22D1BWP12T U2177 ( .A1(r7[8]), .A2(n1327), .B1(n1906), .B2(r2[8]), .ZN(
        n1173) );
  AOI22D1BWP12T U2178 ( .A1(r5[8]), .A2(n3592), .B1(n3591), .B2(r10[8]), .ZN(
        n1172) );
  INVD0BWP12T U2179 ( .I(r9[8]), .ZN(n1166) );
  INVD1BWP12T U2180 ( .I(r4[8]), .ZN(n1369) );
  OAI22D1BWP12T U2181 ( .A1(n3584), .A2(n1166), .B1(n3582), .B2(n1369), .ZN(
        n1170) );
  INVD1BWP12T U2182 ( .I(r11[8]), .ZN(n1168) );
  INVD1BWP12T U2183 ( .I(r0[8]), .ZN(n1167) );
  TPOAI22D1BWP12T U2184 ( .A1(n3586), .A2(n1168), .B1(n3588), .B2(n1167), .ZN(
        n1169) );
  TPNR2D1BWP12T U2185 ( .A1(n1170), .A2(n1169), .ZN(n1171) );
  AN4XD1BWP12T U2186 ( .A1(n1174), .A2(n1173), .A3(n1172), .A4(n1171), .Z(
        n1184) );
  INVD1BWP12T U2187 ( .I(r12[8]), .ZN(n2106) );
  INVD1BWP12T U2188 ( .I(r1[8]), .ZN(n2928) );
  OAI22D0BWP12T U2189 ( .A1(n2106), .A2(n3600), .B1(n3599), .B2(n2928), .ZN(
        n1182) );
  INVD1BWP12T U2190 ( .I(n[3692]), .ZN(n1175) );
  INVD1BWP12T U2191 ( .I(r8[8]), .ZN(n2105) );
  OAI22D1BWP12T U2192 ( .A1(n3605), .A2(n1175), .B1(n3603), .B2(n2105), .ZN(
        n1181) );
  INVD1BWP12T U2193 ( .I(lr[8]), .ZN(n1176) );
  INVD1BWP12T U2194 ( .I(r3[8]), .ZN(n1358) );
  OAI22D1BWP12T U2195 ( .A1(n1176), .A2(n1884), .B1(n1913), .B2(n1358), .ZN(
        n1180) );
  INVD1BWP12T U2196 ( .I(pc_out[8]), .ZN(n1178) );
  INVD1BWP12T U2197 ( .I(r6[8]), .ZN(n1177) );
  OAI22D1BWP12T U2198 ( .A1(n3612), .A2(n1178), .B1(n3611), .B2(n1177), .ZN(
        n1179) );
  NR4D0BWP12T U2199 ( .A1(n1182), .A2(n1181), .A3(n1180), .A4(n1179), .ZN(
        n1183) );
  TPND2D1BWP12T U2200 ( .A1(n1184), .A2(n1183), .ZN(regB_out[8]) );
  AOI22D1BWP12T U2201 ( .A1(tmp1[26]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[26]), .ZN(n1194) );
  INVD1BWP12T U2202 ( .I(r9[26]), .ZN(n1186) );
  OAI22D1BWP12T U2203 ( .A1(n3584), .A2(n1186), .B1(n3582), .B2(n1185), .ZN(
        n1190) );
  OAI22D1BWP12T U2204 ( .A1(n3586), .A2(n1188), .B1(n3588), .B2(n1187), .ZN(
        n1189) );
  NR2D1BWP12T U2205 ( .A1(n1190), .A2(n1189), .ZN(n1193) );
  AOI22D1BWP12T U2206 ( .A1(r5[26]), .A2(n3592), .B1(n3591), .B2(r10[26]), 
        .ZN(n1192) );
  AOI22D1BWP12T U2207 ( .A1(r7[26]), .A2(n3524), .B1(n3593), .B2(r2[26]), .ZN(
        n1191) );
  AN4XD1BWP12T U2208 ( .A1(n1194), .A2(n1193), .A3(n1192), .A4(n1191), .Z(
        n1206) );
  OAI22D0BWP12T U2209 ( .A1(n1196), .A2(n3600), .B1(n3599), .B2(n1195), .ZN(
        n1204) );
  OAI22D1BWP12T U2210 ( .A1(n3605), .A2(n1991), .B1(n3603), .B2(n1197), .ZN(
        n1203) );
  OAI22D1BWP12T U2211 ( .A1(n1199), .A2(n3571), .B1(n3607), .B2(n1198), .ZN(
        n1202) );
  OAI22D1BWP12T U2212 ( .A1(n3612), .A2(n3646), .B1(n3611), .B2(n1200), .ZN(
        n1201) );
  CKND2D2BWP12T U2213 ( .A1(n1206), .A2(n1205), .ZN(regB_out[26]) );
  INVD1BWP12T U2214 ( .I(write1_in[30]), .ZN(n3619) );
  INVD1BWP12T U2215 ( .I(r7[6]), .ZN(n1207) );
  INVD1BWP12T U2216 ( .I(pc_out[6]), .ZN(n1439) );
  TPOAI22D1BWP12T U2217 ( .A1(n3487), .A2(n1207), .B1(n3486), .B2(n1439), .ZN(
        n1212) );
  INVD1BWP12T U2218 ( .I(r5[6]), .ZN(n1208) );
  INVD1BWP12T U2219 ( .I(r3[6]), .ZN(n1436) );
  TPOAI22D1BWP12T U2220 ( .A1(n3489), .A2(n1208), .B1(n3488), .B2(n1436), .ZN(
        n1211) );
  INVD1BWP12T U2221 ( .I(n[3694]), .ZN(n2784) );
  INVD1BWP12T U2222 ( .I(r11[6]), .ZN(n1429) );
  INVD1BWP12T U2223 ( .I(r1[6]), .ZN(n2909) );
  INVD1BWP12T U2224 ( .I(r12[6]), .ZN(n2783) );
  TPOAI22D1BWP12T U2225 ( .A1(n3463), .A2(n2909), .B1(n1716), .B2(n2783), .ZN(
        n1209) );
  NR4D2BWP12T U2226 ( .A1(n1211), .A2(n1212), .A3(n1210), .A4(n1209), .ZN(
        n1221) );
  IOA21D1BWP12T U2227 ( .A1(n3474), .A2(r2[6]), .B(n1213), .ZN(n1215) );
  INVD1BWP12T U2228 ( .I(r4[6]), .ZN(n1426) );
  INVD1BWP12T U2229 ( .I(r0[6]), .ZN(n1428) );
  TPOAI22D1BWP12T U2230 ( .A1(n3448), .A2(n1426), .B1(n3476), .B2(n1428), .ZN(
        n1214) );
  TPNR2D1BWP12T U2231 ( .A1(n1215), .A2(n1214), .ZN(n1220) );
  INVD1BWP12T U2232 ( .I(r6[6]), .ZN(n1438) );
  INVD1BWP12T U2233 ( .I(r10[6]), .ZN(n1216) );
  INVD1BWP12T U2234 ( .I(lr[6]), .ZN(n1437) );
  INVD1BWP12T U2235 ( .I(r8[6]), .ZN(n1435) );
  TPOAI22D1BWP12T U2236 ( .A1(n3478), .A2(n1437), .B1(n3477), .B2(n1435), .ZN(
        n1217) );
  ND3D2BWP12T U2237 ( .A1(n1221), .A2(n1220), .A3(n1219), .ZN(regA_out[6]) );
  ND2D1BWP12T U2238 ( .A1(n1923), .A2(lr[16]), .ZN(n1229) );
  ND2D1BWP12T U2239 ( .A1(n1924), .A2(r8[16]), .ZN(n1224) );
  ND2D1BWP12T U2240 ( .A1(n1950), .A2(r7[16]), .ZN(n1223) );
  ND2D1BWP12T U2241 ( .A1(n1946), .A2(n[3684]), .ZN(n1222) );
  ND3D2BWP12T U2242 ( .A1(n1224), .A2(n1223), .A3(n1222), .ZN(n1228) );
  ND2D1BWP12T U2243 ( .A1(n1942), .A2(r5[16]), .ZN(n1225) );
  OAI21D1BWP12T U2244 ( .A1(n234), .A2(n1226), .B(n1225), .ZN(n1227) );
  INR3D2BWP12T U2245 ( .A1(n1229), .B1(n1228), .B2(n1227), .ZN(n1244) );
  ND2D1BWP12T U2246 ( .A1(n3474), .A2(r2[16]), .ZN(n1232) );
  ND2D1BWP12T U2247 ( .A1(n3471), .A2(r9[16]), .ZN(n1231) );
  ND2D1BWP12T U2248 ( .A1(n3472), .A2(tmp1[16]), .ZN(n1230) );
  ND3D1BWP12T U2249 ( .A1(n1232), .A2(n1231), .A3(n1230), .ZN(n1236) );
  INR2D1BWP12T U2250 ( .A1(r11[16]), .B1(n3490), .ZN(n1234) );
  INR2D1BWP12T U2251 ( .A1(r10[16]), .B1(n3422), .ZN(n1233) );
  OR2D2BWP12T U2252 ( .A1(n1234), .A2(n1233), .Z(n1235) );
  NR2D2BWP12T U2253 ( .A1(n1235), .A2(n1236), .ZN(n1243) );
  AOI22D1BWP12T U2254 ( .A1(n1951), .A2(r1[16]), .B1(n1642), .B2(r6[16]), .ZN(
        n1238) );
  CKND2D0BWP12T U2255 ( .A1(n1945), .A2(pc_out[16]), .ZN(n1237) );
  ND3XD3BWP12T U2256 ( .A1(n1244), .A2(n1243), .A3(n1242), .ZN(regA_out[16])
         );
  TPND2D2BWP12T U2257 ( .A1(n235), .A2(r0[1]), .ZN(n1248) );
  INVD1BWP12T U2258 ( .I(r2[1]), .ZN(n1249) );
  TPND2D2BWP12T U2259 ( .A1(n3471), .A2(r9[1]), .ZN(n1251) );
  ND3D2BWP12T U2260 ( .A1(n1252), .A2(n1251), .A3(n1250), .ZN(n1253) );
  TPNR3D2BWP12T U2261 ( .A1(n1255), .A2(n1254), .A3(n1253), .ZN(n1269) );
  AN2D4BWP12T U2262 ( .A1(n1951), .A2(r1[1]), .Z(n1258) );
  INVD1BWP12T U2263 ( .I(r3[1]), .ZN(n1739) );
  ND2D1BWP12T U2264 ( .A1(n6), .A2(pc_out[1]), .ZN(n1264) );
  ND2XD3BWP12T U2265 ( .A1(n1269), .A2(n1268), .ZN(regA_out[1]) );
  INR2D2BWP12T U2266 ( .A1(r11[9]), .B1(n3490), .ZN(n1270) );
  TPAOI21D2BWP12T U2267 ( .A1(n1924), .A2(r8[9]), .B(n1270), .ZN(n1274) );
  INVD1BWP12T U2268 ( .I(r5[9]), .ZN(n1271) );
  CKND2D0BWP12T U2269 ( .A1(n1275), .A2(lr[9]), .ZN(n1276) );
  INR2D1BWP12T U2270 ( .A1(n1285), .B1(n1276), .ZN(n1277) );
  INVD1BWP12T U2271 ( .I(n1277), .ZN(n1278) );
  TPOAI21D1BWP12T U2272 ( .A1(n3488), .A2(n1279), .B(n1278), .ZN(n1283) );
  INVD1BWP12T U2273 ( .I(r2[9]), .ZN(n1280) );
  CKND2D2BWP12T U2274 ( .A1(n1281), .A2(n248), .ZN(n1282) );
  AN3XD1BWP12T U2275 ( .A1(n1285), .A2(r10[9]), .A3(n1933), .Z(n1289) );
  INR3D0BWP12T U2276 ( .A1(pc_out[9]), .B1(n1287), .B2(n1286), .ZN(n1288) );
  NR2D1BWP12T U2277 ( .A1(n1289), .A2(n1288), .ZN(n1295) );
  INR3D0BWP12T U2278 ( .A1(n1291), .B1(n2923), .B2(n1290), .ZN(n1292) );
  AOI21D1BWP12T U2279 ( .A1(n3472), .A2(tmp1[9]), .B(n1292), .ZN(n1294) );
  ND2D1BWP12T U2280 ( .A1(n1642), .A2(r6[9]), .ZN(n1293) );
  TPND3D1BWP12T U2281 ( .A1(n1295), .A2(n1294), .A3(n1293), .ZN(n1302) );
  TPND2D2BWP12T U2282 ( .A1(n235), .A2(r0[9]), .ZN(n1296) );
  AOI22D1BWP12T U2283 ( .A1(tmp1[21]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[21]), .ZN(n1312) );
  INVD0BWP12T U2284 ( .I(r9[21]), .ZN(n1306) );
  CKND0BWP12T U2285 ( .I(r4[21]), .ZN(n1305) );
  OAI22D1BWP12T U2286 ( .A1(n3584), .A2(n1306), .B1(n3582), .B2(n1305), .ZN(
        n1308) );
  INVD1BWP12T U2287 ( .I(r11[21]), .ZN(n1560) );
  INVD1BWP12T U2288 ( .I(r0[21]), .ZN(n1548) );
  OAI22D1BWP12T U2289 ( .A1(n3586), .A2(n1560), .B1(n3588), .B2(n1548), .ZN(
        n1307) );
  NR2D1BWP12T U2290 ( .A1(n1308), .A2(n1307), .ZN(n1311) );
  AOI22D1BWP12T U2291 ( .A1(r5[21]), .A2(n3592), .B1(n3591), .B2(r10[21]), 
        .ZN(n1310) );
  AOI22D1BWP12T U2292 ( .A1(r7[21]), .A2(n1327), .B1(n3593), .B2(r2[21]), .ZN(
        n1309) );
  AN4XD1BWP12T U2293 ( .A1(n1312), .A2(n1311), .A3(n1310), .A4(n1309), .Z(
        n1319) );
  INVD0BWP12T U2294 ( .I(r12[21]), .ZN(n1313) );
  INVD1BWP12T U2295 ( .I(r1[21]), .ZN(n1562) );
  OAI22D0BWP12T U2296 ( .A1(n1313), .A2(n3600), .B1(n3599), .B2(n1562), .ZN(
        n1317) );
  INVD1BWP12T U2297 ( .I(n[3679]), .ZN(n1561) );
  INVD1BWP12T U2298 ( .I(r8[21]), .ZN(n1551) );
  OAI22D1BWP12T U2299 ( .A1(n3605), .A2(n1561), .B1(n3603), .B2(n1551), .ZN(
        n1316) );
  INVD1BWP12T U2300 ( .I(lr[21]), .ZN(n1552) );
  INVD1BWP12T U2301 ( .I(r3[21]), .ZN(n1557) );
  INVD1BWP12T U2302 ( .I(pc_out[21]), .ZN(n1559) );
  INVD1BWP12T U2303 ( .I(r6[21]), .ZN(n1550) );
  OAI22D1BWP12T U2304 ( .A1(n3612), .A2(n1559), .B1(n3611), .B2(n1550), .ZN(
        n1314) );
  NR4D0BWP12T U2305 ( .A1(n1317), .A2(n1316), .A3(n1315), .A4(n1314), .ZN(
        n1318) );
  CKND2D2BWP12T U2306 ( .A1(n1319), .A2(n1318), .ZN(regB_out[21]) );
  INVD1BWP12T U2307 ( .I(r12[5]), .ZN(n1419) );
  INVD1P75BWP12T U2308 ( .I(r1[5]), .ZN(n2896) );
  OAI22D0BWP12T U2309 ( .A1(n1419), .A2(n3600), .B1(n3599), .B2(n2896), .ZN(
        n1323) );
  INVD1BWP12T U2310 ( .I(r8[5]), .ZN(n1407) );
  OAI22D1BWP12T U2311 ( .A1(n3605), .A2(n1418), .B1(n3603), .B2(n1407), .ZN(
        n1322) );
  INVD1BWP12T U2312 ( .I(r3[5]), .ZN(n1415) );
  OAI22D0BWP12T U2313 ( .A1(n2327), .A2(n1394), .B1(n1740), .B2(n1415), .ZN(
        n1321) );
  INVD1BWP12T U2314 ( .I(pc_out[5]), .ZN(n1412) );
  INVD1BWP12T U2315 ( .I(r6[5]), .ZN(n1404) );
  OAI22D1BWP12T U2316 ( .A1(n3612), .A2(n1412), .B1(n3611), .B2(n1404), .ZN(
        n1320) );
  NR4D0BWP12T U2317 ( .A1(n1323), .A2(n1322), .A3(n1321), .A4(n1320), .ZN(
        n1333) );
  INVD1BWP12T U2318 ( .I(r9[5]), .ZN(n2326) );
  CKND1BWP12T U2319 ( .I(r4[5]), .ZN(n1324) );
  OAI22D1BWP12T U2320 ( .A1(n3584), .A2(n2326), .B1(n3582), .B2(n1324), .ZN(
        n1326) );
  INVD1BWP12T U2321 ( .I(r11[5]), .ZN(n1417) );
  INVD1BWP12T U2322 ( .I(r0[5]), .ZN(n1406) );
  OAI22D1BWP12T U2323 ( .A1(n3586), .A2(n1417), .B1(n1901), .B2(n1406), .ZN(
        n1325) );
  TPNR2D1BWP12T U2324 ( .A1(n1326), .A2(n1325), .ZN(n1331) );
  AOI22D2BWP12T U2325 ( .A1(r5[5]), .A2(n3592), .B1(n3591), .B2(r10[5]), .ZN(
        n1330) );
  AOI22D1BWP12T U2326 ( .A1(n1327), .A2(r7[5]), .B1(n1730), .B2(r2[5]), .ZN(
        n1329) );
  AN4D4BWP12T U2327 ( .A1(n1331), .A2(n1330), .A3(n1329), .A4(n1328), .Z(n1332) );
  TPND2D2BWP12T U2328 ( .A1(n1333), .A2(n1332), .ZN(regB_out[5]) );
  INVD1BWP12T U2329 ( .I(r6[14]), .ZN(n1582) );
  INVD1BWP12T U2330 ( .I(r10[14]), .ZN(n2828) );
  OAI22D1BWP12T U2331 ( .A1(n3481), .A2(n1582), .B1(n2828), .B2(n3422), .ZN(
        n1335) );
  INVD1BWP12T U2332 ( .I(r1[14]), .ZN(n1579) );
  INVD1BWP12T U2333 ( .I(r12[14]), .ZN(n1580) );
  OAI22D1BWP12T U2334 ( .A1(n1579), .A2(n3463), .B1(n3492), .B2(n1580), .ZN(
        n1334) );
  NR2D1BWP12T U2335 ( .A1(n1335), .A2(n1334), .ZN(n1343) );
  INVD1BWP12T U2336 ( .I(r5[14]), .ZN(n1336) );
  INVD1BWP12T U2337 ( .I(r3[14]), .ZN(n1581) );
  OAI22D1BWP12T U2338 ( .A1(n3489), .A2(n1336), .B1(n1581), .B2(n3488), .ZN(
        n1341) );
  INVD1BWP12T U2339 ( .I(r0[14]), .ZN(n1571) );
  INVD1BWP12T U2340 ( .I(r11[14]), .ZN(n1572) );
  OAI22D0BWP12T U2341 ( .A1(n3476), .A2(n1571), .B1(n1572), .B2(n1337), .ZN(
        n1340) );
  INVD1BWP12T U2342 ( .I(r7[14]), .ZN(n1338) );
  MOAI22D1BWP12T U2343 ( .A1(n3487), .A2(n1338), .B1(n6), .B2(pc_out[14]), 
        .ZN(n1339) );
  NR3D1BWP12T U2344 ( .A1(n1341), .A2(n1340), .A3(n1339), .ZN(n1342) );
  CKAN2D2BWP12T U2345 ( .A1(n1343), .A2(n1342), .Z(n1351) );
  INVD1BWP12T U2346 ( .I(lr[14]), .ZN(n2831) );
  INVD1BWP12T U2347 ( .I(r8[14]), .ZN(n2829) );
  OAI22D1BWP12T U2348 ( .A1(n3478), .A2(n2831), .B1(n3477), .B2(n2829), .ZN(
        n1345) );
  INVD1BWP12T U2349 ( .I(r4[14]), .ZN(n1569) );
  INVD1BWP12T U2350 ( .I(n[3686]), .ZN(n2833) );
  OAI22D1BWP12T U2351 ( .A1(n1569), .A2(n3448), .B1(n3491), .B2(n2833), .ZN(
        n1344) );
  NR2D1BWP12T U2352 ( .A1(n1345), .A2(n1344), .ZN(n1349) );
  AOI22D1BWP12T U2353 ( .A1(r9[14]), .A2(n3471), .B1(n3472), .B2(tmp1[14]), 
        .ZN(n1346) );
  IOA21D1BWP12T U2354 ( .A1(n3474), .A2(r2[14]), .B(n1346), .ZN(n1347) );
  INVD1BWP12T U2355 ( .I(n1347), .ZN(n1348) );
  AN2XD2BWP12T U2356 ( .A1(n1349), .A2(n1348), .Z(n1350) );
  INR2D2BWP12T U2357 ( .A1(r11[8]), .B1(n3490), .ZN(n1352) );
  TPAOI21D1BWP12T U2358 ( .A1(n1946), .A2(n[3692]), .B(n1352), .ZN(n1355) );
  ND2D1BWP12T U2359 ( .A1(n1950), .A2(r7[8]), .ZN(n1354) );
  CKND2D0BWP12T U2360 ( .A1(n6), .A2(pc_out[8]), .ZN(n1353) );
  ND3D1BWP12T U2361 ( .A1(n1355), .A2(n1354), .A3(n1353), .ZN(n1363) );
  AN2D1BWP12T U2362 ( .A1(n1952), .A2(r12[8]), .Z(n1362) );
  TPNR2D1BWP12T U2363 ( .A1(n3463), .A2(n2928), .ZN(n1356) );
  INVD1BWP12T U2364 ( .I(n1356), .ZN(n1361) );
  TPOAI21D1BWP12T U2365 ( .A1(n3488), .A2(n1358), .B(n1357), .ZN(n1359) );
  INR2D2BWP12T U2366 ( .A1(r10[8]), .B1(n3479), .ZN(n1364) );
  CKND2D0BWP12T U2367 ( .A1(n1653), .A2(lr[8]), .ZN(n1366) );
  ND2D1BWP12T U2368 ( .A1(n1924), .A2(r8[8]), .ZN(n1365) );
  ND2D3BWP12T U2369 ( .A1(n235), .A2(r0[8]), .ZN(n1368) );
  OAI21D1BWP12T U2370 ( .A1(n3448), .A2(n1369), .B(n1368), .ZN(n1374) );
  ND2D1BWP12T U2371 ( .A1(n3474), .A2(r2[8]), .ZN(n1372) );
  ND2D1BWP12T U2372 ( .A1(n3471), .A2(r9[8]), .ZN(n1371) );
  ND2D1BWP12T U2373 ( .A1(n3472), .A2(tmp1[8]), .ZN(n1370) );
  ND3D2BWP12T U2374 ( .A1(n1372), .A2(n1371), .A3(n1370), .ZN(n1373) );
  TPNR3D2BWP12T U2375 ( .A1(n1375), .A2(n1374), .A3(n1373), .ZN(n1376) );
  INVD1BWP12T U2376 ( .I(r9[3]), .ZN(n1379) );
  INVD1BWP12T U2377 ( .I(r4[3]), .ZN(n1378) );
  INVD1BWP12T U2378 ( .I(r11[3]), .ZN(n1381) );
  INVD1BWP12T U2379 ( .I(r0[3]), .ZN(n1380) );
  AOI22D1BWP12T U2380 ( .A1(tmp1[3]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[3]), .ZN(n1384) );
  AOI22D1BWP12T U2381 ( .A1(n3524), .A2(r7[3]), .B1(n1730), .B2(r2[3]), .ZN(
        n1383) );
  INR2D2BWP12T U2382 ( .A1(n1386), .B1(n1385), .ZN(n1401) );
  INVD1BWP12T U2383 ( .I(r8[3]), .ZN(n1388) );
  INVD1BWP12T U2384 ( .I(n[3697]), .ZN(n1387) );
  TPOAI22D1BWP12T U2385 ( .A1(n3603), .A2(n1388), .B1(n1738), .B2(n1387), .ZN(
        n1391) );
  INVD1BWP12T U2386 ( .I(r12[3]), .ZN(n1389) );
  OR2XD2BWP12T U2387 ( .A1(n1391), .A2(n1390), .Z(n1399) );
  INVD1BWP12T U2388 ( .I(r6[3]), .ZN(n1392) );
  INVD1BWP12T U2389 ( .I(pc_out[3]), .ZN(n2727) );
  INVD1BWP12T U2390 ( .I(lr[3]), .ZN(n1395) );
  OAI22D1BWP12T U2391 ( .A1(n1395), .A2(n1394), .B1(n1740), .B2(n1393), .ZN(
        n1396) );
  OR2XD4BWP12T U2392 ( .A1(n1397), .A2(n1396), .Z(n1398) );
  TPNR2D2BWP12T U2393 ( .A1(n1399), .A2(n1398), .ZN(n1400) );
  TPND2D2BWP12T U2394 ( .A1(n1401), .A2(n1400), .ZN(regB_out[3]) );
  AOI22D2BWP12T U2395 ( .A1(r9[5]), .A2(n3471), .B1(n3472), .B2(tmp1[5]), .ZN(
        n1402) );
  IOA21D2BWP12T U2396 ( .A1(r2[5]), .A2(n3474), .B(n1402), .ZN(n1411) );
  INVD1BWP12T U2397 ( .I(r10[5]), .ZN(n1403) );
  TPND2D2BWP12T U2398 ( .A1(n3475), .A2(r4[5]), .ZN(n1405) );
  TPOAI21D1BWP12T U2399 ( .A1(n3476), .A2(n1406), .B(n1405), .ZN(n1409) );
  TPOAI22D2BWP12T U2400 ( .A1(n3478), .A2(n2327), .B1(n3477), .B2(n1407), .ZN(
        n1408) );
  NR4D2BWP12T U2401 ( .A1(n1411), .A2(n1410), .A3(n1409), .A4(n1408), .ZN(
        n1425) );
  INVD1BWP12T U2402 ( .I(r7[5]), .ZN(n1413) );
  TPOAI22D1BWP12T U2403 ( .A1(n1414), .A2(n1413), .B1(n3486), .B2(n1412), .ZN(
        n1423) );
  INVD1BWP12T U2404 ( .I(r5[5]), .ZN(n1416) );
  TPOAI22D2BWP12T U2405 ( .A1(n3489), .A2(n1416), .B1(n1415), .B2(n3488), .ZN(
        n1422) );
  TPOAI22D2BWP12T U2406 ( .A1(n3491), .A2(n1418), .B1(n3490), .B2(n1417), .ZN(
        n1421) );
  TPOAI22D2BWP12T U2407 ( .A1(n3492), .A2(n1419), .B1(n3463), .B2(n2896), .ZN(
        n1420) );
  NR4D2BWP12T U2408 ( .A1(n1423), .A2(n1422), .A3(n1421), .A4(n1420), .ZN(
        n1424) );
  TPND2D3BWP12T U2409 ( .A1(n1425), .A2(n1424), .ZN(regA_out[5]) );
  AOI22D1BWP12T U2410 ( .A1(tmp1[6]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[6]), .ZN(n1434) );
  AOI22D1BWP12T U2411 ( .A1(r5[6]), .A2(n3592), .B1(n3591), .B2(r10[6]), .ZN(
        n1433) );
  AOI22D1BWP12T U2412 ( .A1(r7[6]), .A2(n1327), .B1(n1906), .B2(r2[6]), .ZN(
        n1432) );
  INVD1BWP12T U2413 ( .I(r9[6]), .ZN(n1427) );
  OAI22D1BWP12T U2414 ( .A1(n3584), .A2(n1427), .B1(n3582), .B2(n1426), .ZN(
        n1431) );
  TPOAI22D1BWP12T U2415 ( .A1(n3586), .A2(n1429), .B1(n3588), .B2(n1428), .ZN(
        n1430) );
  OAI22D1BWP12T U2416 ( .A1(n2783), .A2(n3600), .B1(n3599), .B2(n2909), .ZN(
        n1443) );
  OAI22D1BWP12T U2417 ( .A1(n3605), .A2(n2784), .B1(n3603), .B2(n1435), .ZN(
        n1442) );
  OAI22D1BWP12T U2418 ( .A1(n1437), .A2(n1884), .B1(n1913), .B2(n1436), .ZN(
        n1441) );
  OAI22D1BWP12T U2419 ( .A1(n3612), .A2(n1439), .B1(n3611), .B2(n1438), .ZN(
        n1440) );
  NR4D0BWP12T U2420 ( .A1(n1443), .A2(n1442), .A3(n1441), .A4(n1440), .ZN(
        n1444) );
  TPND2D1BWP12T U2421 ( .A1(n1445), .A2(n1444), .ZN(regB_out[6]) );
  AOI22D1BWP12T U2422 ( .A1(tmp1[23]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[23]), .ZN(n1453) );
  INVD0BWP12T U2423 ( .I(r9[23]), .ZN(n1447) );
  CKND0BWP12T U2424 ( .I(r4[23]), .ZN(n1446) );
  OAI22D1BWP12T U2425 ( .A1(n3584), .A2(n1447), .B1(n3582), .B2(n1446), .ZN(
        n1449) );
  INVD1BWP12T U2426 ( .I(r11[23]), .ZN(n1795) );
  INVD1BWP12T U2427 ( .I(r0[23]), .ZN(n1784) );
  OAI22D1BWP12T U2428 ( .A1(n3586), .A2(n1795), .B1(n3588), .B2(n1784), .ZN(
        n1448) );
  NR2D1BWP12T U2429 ( .A1(n1449), .A2(n1448), .ZN(n1452) );
  AOI22D1BWP12T U2430 ( .A1(r5[23]), .A2(n3592), .B1(n3591), .B2(r10[23]), 
        .ZN(n1451) );
  AOI22D1BWP12T U2431 ( .A1(r7[23]), .A2(n3524), .B1(n3593), .B2(r2[23]), .ZN(
        n1450) );
  AN4XD1BWP12T U2432 ( .A1(n1453), .A2(n1452), .A3(n1451), .A4(n1450), .Z(
        n1458) );
  INVD1BWP12T U2433 ( .I(r8[23]), .ZN(n2689) );
  OAI22D1BWP12T U2434 ( .A1(n3605), .A2(n1796), .B1(n3603), .B2(n2689), .ZN(
        n1455) );
  INVD1BWP12T U2435 ( .I(pc_out[23]), .ZN(n3314) );
  INVD1BWP12T U2436 ( .I(r6[23]), .ZN(n1786) );
  OAI22D1BWP12T U2437 ( .A1(n3612), .A2(n3314), .B1(n3611), .B2(n1786), .ZN(
        n1454) );
  INVD1BWP12T U2438 ( .I(r12[23]), .ZN(n1797) );
  INVD1BWP12T U2439 ( .I(r1[23]), .ZN(n1798) );
  OAI22D0BWP12T U2440 ( .A1(n1797), .A2(n3600), .B1(n3599), .B2(n1798), .ZN(
        n1457) );
  INVD1BWP12T U2441 ( .I(lr[23]), .ZN(n1787) );
  INVD1BWP12T U2442 ( .I(r3[23]), .ZN(n1793) );
  OAI22D1BWP12T U2443 ( .A1(n1787), .A2(n3608), .B1(n3607), .B2(n1793), .ZN(
        n1456) );
  INVD6BWP12T U2444 ( .I(n1865), .ZN(n3325) );
  AOI22D1BWP12T U2445 ( .A1(n2989), .A2(pc_out[22]), .B1(n3398), .B2(
        next_pc_in[22]), .ZN(n1459) );
  TPOAI21D1BWP12T U2446 ( .A1(n1460), .A2(n3394), .B(n1459), .ZN(n2191) );
  INR2D1BWP12T U2447 ( .A1(r11[2]), .B1(n3490), .ZN(n1461) );
  INR2D1BWP12T U2448 ( .A1(r10[2]), .B1(n3422), .ZN(n1465) );
  CKND2D0BWP12T U2449 ( .A1(n6), .A2(pc_out[2]), .ZN(n1464) );
  IND3D2BWP12T U2450 ( .A1(n1465), .B1(n1464), .B2(n1463), .ZN(n1466) );
  INR2D4BWP12T U2451 ( .A1(n1467), .B1(n1466), .ZN(n1485) );
  CKND0BWP12T U2452 ( .I(n1468), .ZN(n1470) );
  INVD1BWP12T U2453 ( .I(r3[2]), .ZN(n1691) );
  ND2D1BWP12T U2454 ( .A1(n1942), .A2(r5[2]), .ZN(n1469) );
  IOA21D1BWP12T U2455 ( .A1(n1470), .A2(r3[2]), .B(n1469), .ZN(n1474) );
  ND2D1BWP12T U2456 ( .A1(n3471), .A2(r9[2]), .ZN(n1476) );
  ND2D1BWP12T U2457 ( .A1(n3472), .A2(tmp1[2]), .ZN(n1475) );
  INVD1BWP12T U2458 ( .I(r1[2]), .ZN(n2088) );
  TPOAI21D2BWP12T U2459 ( .A1(n2088), .A2(n3463), .B(n1479), .ZN(n1482) );
  AN2XD2BWP12T U2460 ( .A1(n1923), .A2(lr[2]), .Z(n1481) );
  TPNR3D2BWP12T U2461 ( .A1(n1482), .A2(n1481), .A3(n1480), .ZN(n1483) );
  ND3XD4BWP12T U2462 ( .A1(n1485), .A2(n1484), .A3(n1483), .ZN(regA_out[2]) );
  INVD1BWP12T U2463 ( .I(r1[20]), .ZN(n1503) );
  INVD1BWP12T U2464 ( .I(r12[20]), .ZN(n1502) );
  TPNR2D1BWP12T U2465 ( .A1(n1488), .A2(n1487), .ZN(n1501) );
  INVD1BWP12T U2466 ( .I(r7[20]), .ZN(n1489) );
  OAI22D1BWP12T U2467 ( .A1(n3487), .A2(n1489), .B1(n3486), .B2(n3642), .ZN(
        n1491) );
  INVD1BWP12T U2468 ( .I(lr[20]), .ZN(n1506) );
  INVD1BWP12T U2469 ( .I(r8[20]), .ZN(n1504) );
  OAI22D1BWP12T U2470 ( .A1(n3478), .A2(n1506), .B1(n3477), .B2(n1504), .ZN(
        n1490) );
  TPNR2D1BWP12T U2471 ( .A1(n1491), .A2(n1490), .ZN(n1500) );
  INVD1BWP12T U2472 ( .I(n[3680]), .ZN(n2027) );
  INVD1BWP12T U2473 ( .I(r11[20]), .ZN(n2026) );
  OAI22D1BWP12T U2474 ( .A1(n3491), .A2(n2027), .B1(n2026), .B2(n3490), .ZN(
        n1494) );
  INVD1BWP12T U2475 ( .I(r6[20]), .ZN(n1507) );
  INVD1BWP12T U2476 ( .I(r10[20]), .ZN(n1492) );
  INVD1BWP12T U2477 ( .I(r5[20]), .ZN(n1495) );
  INVD1BWP12T U2478 ( .I(r3[20]), .ZN(n1505) );
  OAI22D1BWP12T U2479 ( .A1(n3489), .A2(n1495), .B1(n1505), .B2(n3488), .ZN(
        n1497) );
  INVD1BWP12T U2480 ( .I(r4[20]), .ZN(n1512) );
  INVD1BWP12T U2481 ( .I(r0[20]), .ZN(n1514) );
  OAI22D1BWP12T U2482 ( .A1(n3448), .A2(n1512), .B1(n3476), .B2(n1514), .ZN(
        n1496) );
  TPNR2D1BWP12T U2483 ( .A1(n1497), .A2(n1496), .ZN(n1498) );
  OAI22D0BWP12T U2484 ( .A1(n1503), .A2(n3599), .B1(n3600), .B2(n1502), .ZN(
        n1511) );
  OAI22D1BWP12T U2485 ( .A1(n3605), .A2(n2027), .B1(n3603), .B2(n1504), .ZN(
        n1510) );
  OAI22D1BWP12T U2486 ( .A1(n1506), .A2(n3571), .B1(n3607), .B2(n1505), .ZN(
        n1509) );
  OAI22D1BWP12T U2487 ( .A1(n3612), .A2(n3642), .B1(n3611), .B2(n1507), .ZN(
        n1508) );
  NR4D0BWP12T U2488 ( .A1(n1511), .A2(n1510), .A3(n1509), .A4(n1508), .ZN(
        n1522) );
  AOI22D1BWP12T U2489 ( .A1(tmp1[20]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[20]), .ZN(n1520) );
  INVD1BWP12T U2490 ( .I(r9[20]), .ZN(n1513) );
  OAI22D1BWP12T U2491 ( .A1(n3584), .A2(n1513), .B1(n3582), .B2(n1512), .ZN(
        n1516) );
  OAI22D1BWP12T U2492 ( .A1(n3586), .A2(n2026), .B1(n3588), .B2(n1514), .ZN(
        n1515) );
  NR2D1BWP12T U2493 ( .A1(n1516), .A2(n1515), .ZN(n1519) );
  AOI22D1BWP12T U2494 ( .A1(r5[20]), .A2(n3592), .B1(n3591), .B2(r10[20]), 
        .ZN(n1518) );
  AOI22D1BWP12T U2495 ( .A1(r7[20]), .A2(n1327), .B1(n3593), .B2(r2[20]), .ZN(
        n1517) );
  AN4XD1BWP12T U2496 ( .A1(n1520), .A2(n1519), .A3(n1518), .A4(n1517), .Z(
        n1521) );
  TPND2D2BWP12T U2497 ( .A1(n1522), .A2(n1521), .ZN(regB_out[20]) );
  AOI22D1BWP12T U2498 ( .A1(tmp1[13]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[13]), .ZN(n1532) );
  INVD1BWP12T U2499 ( .I(r9[13]), .ZN(n1524) );
  OAI22D1BWP12T U2500 ( .A1(n3584), .A2(n1524), .B1(n3582), .B2(n1523), .ZN(
        n1528) );
  NR2D1BWP12T U2501 ( .A1(n1528), .A2(n1527), .ZN(n1531) );
  AOI22D1BWP12T U2502 ( .A1(r5[13]), .A2(n3592), .B1(n3591), .B2(r10[13]), 
        .ZN(n1530) );
  AOI22D1BWP12T U2503 ( .A1(r7[13]), .A2(n3524), .B1(n1906), .B2(r2[13]), .ZN(
        n1529) );
  AN4XD1BWP12T U2504 ( .A1(n1532), .A2(n1531), .A3(n1530), .A4(n1529), .Z(
        n1545) );
  INVD0BWP12T U2505 ( .I(r12[13]), .ZN(n1534) );
  OAI22D1BWP12T U2506 ( .A1(n1534), .A2(n3600), .B1(n3599), .B2(n1533), .ZN(
        n1543) );
  OAI22D1BWP12T U2507 ( .A1(n1738), .A2(n1536), .B1(n3603), .B2(n1535), .ZN(
        n1542) );
  OAI22D1BWP12T U2508 ( .A1(n2845), .A2(n1884), .B1(n1913), .B2(n1537), .ZN(
        n1541) );
  OAI22D1BWP12T U2509 ( .A1(n3612), .A2(n1539), .B1(n3611), .B2(n1538), .ZN(
        n1540) );
  NR4D0BWP12T U2510 ( .A1(n1543), .A2(n1542), .A3(n1541), .A4(n1540), .ZN(
        n1544) );
  TPND2D2BWP12T U2511 ( .A1(n1545), .A2(n1544), .ZN(regB_out[13]) );
  AOI22D1BWP12T U2512 ( .A1(n3471), .A2(r9[21]), .B1(n3472), .B2(tmp1[21]), 
        .ZN(n1546) );
  IOA21D1BWP12T U2513 ( .A1(n3474), .A2(r2[21]), .B(n1546), .ZN(n1556) );
  ND2D1BWP12T U2514 ( .A1(n3475), .A2(r4[21]), .ZN(n1547) );
  OAI21D1BWP12T U2515 ( .A1(n3476), .A2(n1548), .B(n1547), .ZN(n1555) );
  INVD1BWP12T U2516 ( .I(r10[21]), .ZN(n1549) );
  NR4D0BWP12T U2517 ( .A1(n1556), .A2(n1555), .A3(n1554), .A4(n1553), .ZN(
        n1568) );
  INVD1BWP12T U2518 ( .I(r5[21]), .ZN(n1558) );
  TPOAI22D1BWP12T U2519 ( .A1(n3489), .A2(n1558), .B1(n1557), .B2(n3488), .ZN(
        n1566) );
  MOAI22D1BWP12T U2520 ( .A1(n1562), .A2(n3463), .B1(n1952), .B2(r12[21]), 
        .ZN(n1563) );
  NR4D0BWP12T U2521 ( .A1(n1566), .A2(n1565), .A3(n1564), .A4(n1563), .ZN(
        n1567) );
  TPND2D1BWP12T U2522 ( .A1(n1568), .A2(n1567), .ZN(regA_out[21]) );
  AOI22D1BWP12T U2523 ( .A1(tmp1[14]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[14]), .ZN(n1578) );
  INVD0BWP12T U2524 ( .I(r9[14]), .ZN(n1570) );
  OAI22D1BWP12T U2525 ( .A1(n3584), .A2(n1570), .B1(n3582), .B2(n1569), .ZN(
        n1574) );
  OAI22D1BWP12T U2526 ( .A1(n3586), .A2(n1572), .B1(n3588), .B2(n1571), .ZN(
        n1573) );
  NR2D1BWP12T U2527 ( .A1(n1574), .A2(n1573), .ZN(n1577) );
  AOI22D1BWP12T U2528 ( .A1(r5[14]), .A2(n3592), .B1(n3591), .B2(r10[14]), 
        .ZN(n1576) );
  AOI22D1BWP12T U2529 ( .A1(r7[14]), .A2(n3524), .B1(n1906), .B2(r2[14]), .ZN(
        n1575) );
  AN4XD1BWP12T U2530 ( .A1(n1578), .A2(n1577), .A3(n1576), .A4(n1575), .Z(
        n1589) );
  OAI22D1BWP12T U2531 ( .A1(n1580), .A2(n3600), .B1(n3599), .B2(n1579), .ZN(
        n1587) );
  OAI22D1BWP12T U2532 ( .A1(n3605), .A2(n2833), .B1(n3603), .B2(n2829), .ZN(
        n1586) );
  OAI22D1BWP12T U2533 ( .A1(n2831), .A2(n1884), .B1(n1913), .B2(n1581), .ZN(
        n1585) );
  INVD1BWP12T U2534 ( .I(pc_out[14]), .ZN(n1583) );
  OAI22D1BWP12T U2535 ( .A1(n3612), .A2(n1583), .B1(n3611), .B2(n1582), .ZN(
        n1584) );
  NR4D0BWP12T U2536 ( .A1(n1587), .A2(n1586), .A3(n1585), .A4(n1584), .ZN(
        n1588) );
  TPND2D2BWP12T U2537 ( .A1(n1589), .A2(n1588), .ZN(regB_out[14]) );
  INVD1BWP12T U2538 ( .I(r12[12]), .ZN(n2749) );
  OAI22D0BWP12T U2539 ( .A1(n2749), .A2(n3600), .B1(n3599), .B2(n2952), .ZN(
        n1597) );
  INVD1BWP12T U2540 ( .I(n[3688]), .ZN(n1591) );
  INVD1BWP12T U2541 ( .I(r8[12]), .ZN(n1590) );
  TPOAI22D1BWP12T U2542 ( .A1(n3605), .A2(n1591), .B1(n3603), .B2(n1590), .ZN(
        n1596) );
  INVD1BWP12T U2543 ( .I(lr[12]), .ZN(n1592) );
  INVD1BWP12T U2544 ( .I(r3[12]), .ZN(n1944) );
  OAI22D1BWP12T U2545 ( .A1(n1592), .A2(n1884), .B1(n1913), .B2(n1944), .ZN(
        n1595) );
  INVD1BWP12T U2546 ( .I(pc_out[12]), .ZN(n2750) );
  INVD1BWP12T U2547 ( .I(r6[12]), .ZN(n1593) );
  OAI22D1BWP12T U2548 ( .A1(n3612), .A2(n2750), .B1(n3611), .B2(n1593), .ZN(
        n1594) );
  AOI22D1BWP12T U2549 ( .A1(r7[12]), .A2(n3524), .B1(n1906), .B2(r2[12]), .ZN(
        n1599) );
  AOI22D1BWP12T U2550 ( .A1(r5[12]), .A2(n3592), .B1(n3591), .B2(r10[12]), 
        .ZN(n1598) );
  INVD1BWP12T U2551 ( .I(r9[12]), .ZN(n1600) );
  INVD1BWP12T U2552 ( .I(r4[12]), .ZN(n1932) );
  TPOAI22D1BWP12T U2553 ( .A1(n3584), .A2(n1600), .B1(n3582), .B2(n1932), .ZN(
        n1603) );
  INVD1BWP12T U2554 ( .I(r11[12]), .ZN(n1949) );
  INVD1BWP12T U2555 ( .I(r0[12]), .ZN(n1601) );
  OAI22D1BWP12T U2556 ( .A1(n3586), .A2(n1949), .B1(n1901), .B2(n1601), .ZN(
        n1602) );
  NR2D1BWP12T U2557 ( .A1(n1603), .A2(n1602), .ZN(n1605) );
  AOI22D1BWP12T U2558 ( .A1(tmp1[12]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[12]), .ZN(n1604) );
  CKAN2D2BWP12T U2559 ( .A1(n1605), .A2(n1604), .Z(n1606) );
  OAI21D0BWP12T U2560 ( .A1(r2[4]), .A2(n1610), .B(n1608), .ZN(n1612) );
  CKND0BWP12T U2561 ( .I(readA_sel[2]), .ZN(n1609) );
  AOI21D1BWP12T U2562 ( .A1(n1610), .A2(r4[4]), .B(n1609), .ZN(n1611) );
  NR2D1BWP12T U2563 ( .A1(n1612), .A2(n1611), .ZN(n1617) );
  NR3D1BWP12T U2564 ( .A1(readA_sel[2]), .A2(readA_sel[1]), .A3(r0[4]), .ZN(
        n1615) );
  CKND2D0BWP12T U2565 ( .A1(n335), .A2(n1613), .ZN(n1614) );
  TPNR2D1BWP12T U2566 ( .A1(n1615), .A2(n1614), .ZN(n1616) );
  ND2D1BWP12T U2567 ( .A1(n1642), .A2(r6[4]), .ZN(n1618) );
  TPND2D1BWP12T U2568 ( .A1(n1619), .A2(n1618), .ZN(n1626) );
  TPND2D1BWP12T U2569 ( .A1(n3471), .A2(r9[4]), .ZN(n1620) );
  OAI21D1BWP12T U2570 ( .A1(n3490), .A2(n1621), .B(n1620), .ZN(n1625) );
  ND2D1BWP12T U2571 ( .A1(n1950), .A2(r7[4]), .ZN(n1623) );
  ND2D1BWP12T U2572 ( .A1(n1946), .A2(n[3696]), .ZN(n1622) );
  TPND2D1BWP12T U2573 ( .A1(n1623), .A2(n1622), .ZN(n1624) );
  ND2D1BWP12T U2574 ( .A1(n1942), .A2(r5[4]), .ZN(n1632) );
  NR2D1BWP12T U2575 ( .A1(n3492), .A2(n1627), .ZN(n1631) );
  CKND2D0BWP12T U2576 ( .A1(n1945), .A2(pc_out[4]), .ZN(n1628) );
  OAI21D1BWP12T U2577 ( .A1(n3488), .A2(n1629), .B(n1628), .ZN(n1630) );
  INR3D2BWP12T U2578 ( .A1(n1632), .B1(n1631), .B2(n1630), .ZN(n1640) );
  CKND2D0BWP12T U2579 ( .A1(n1653), .A2(lr[4]), .ZN(n1638) );
  NR2D1BWP12T U2580 ( .A1(n3463), .A2(n2778), .ZN(n1637) );
  INVD1BWP12T U2581 ( .I(r10[4]), .ZN(n1635) );
  CKND2D0BWP12T U2582 ( .A1(n1633), .A2(r8[4]), .ZN(n1634) );
  OAI21D1BWP12T U2583 ( .A1(n3422), .A2(n1635), .B(n1634), .ZN(n1636) );
  INR3D2BWP12T U2584 ( .A1(n1638), .B1(n1637), .B2(n1636), .ZN(n1639) );
  ND3D2BWP12T U2585 ( .A1(n1641), .A2(n1640), .A3(n1639), .ZN(regA_out[4]) );
  AOI22D1BWP12T U2586 ( .A1(n1942), .A2(r5[11]), .B1(n1642), .B2(r6[11]), .ZN(
        n1647) );
  ND2D1BWP12T U2587 ( .A1(n1633), .A2(r8[11]), .ZN(n1646) );
  INR2D2BWP12T U2588 ( .A1(r11[11]), .B1(n3490), .ZN(n1643) );
  INVD1P75BWP12T U2589 ( .I(n1643), .ZN(n1645) );
  ND2D1BWP12T U2590 ( .A1(n1950), .A2(r7[11]), .ZN(n1644) );
  AN4D4BWP12T U2591 ( .A1(n1647), .A2(n1646), .A3(n1645), .A4(n1644), .Z(n1671) );
  ND2D1BWP12T U2592 ( .A1(n3471), .A2(r9[11]), .ZN(n1650) );
  ND2D1BWP12T U2593 ( .A1(n3472), .A2(tmp1[11]), .ZN(n1648) );
  ND2D1BWP12T U2594 ( .A1(n1952), .A2(r12[11]), .ZN(n1651) );
  OAI21D1BWP12T U2595 ( .A1(n1652), .A2(n3488), .B(n1651), .ZN(n1656) );
  ND2D1BWP12T U2596 ( .A1(n1653), .A2(lr[11]), .ZN(n1654) );
  TPNR3D2BWP12T U2597 ( .A1(n1657), .A2(n1656), .A3(n1655), .ZN(n1670) );
  ND2D1BWP12T U2598 ( .A1(n1945), .A2(pc_out[11]), .ZN(n1660) );
  ND2D1BWP12T U2599 ( .A1(n1661), .A2(n1660), .ZN(n1663) );
  OR2XD2BWP12T U2600 ( .A1(n1663), .A2(n1662), .Z(n1668) );
  INVD1BWP12T U2601 ( .I(r2[11]), .ZN(n1665) );
  TPNR2D2BWP12T U2602 ( .A1(n1668), .A2(n1667), .ZN(n1669) );
  ND3XD4BWP12T U2603 ( .A1(n1671), .A2(n1670), .A3(n1669), .ZN(regA_out[11])
         );
  AOI22D1BWP12T U2604 ( .A1(tmp1[2]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[2]), .ZN(n1681) );
  INVD1BWP12T U2605 ( .I(r9[2]), .ZN(n1673) );
  INVD1BWP12T U2606 ( .I(r4[2]), .ZN(n1672) );
  TPOAI22D1BWP12T U2607 ( .A1(n3584), .A2(n1673), .B1(n3582), .B2(n1672), .ZN(
        n1677) );
  INVD1BWP12T U2608 ( .I(r11[2]), .ZN(n1675) );
  INVD1BWP12T U2609 ( .I(r0[2]), .ZN(n1674) );
  OAI22D1BWP12T U2610 ( .A1(n3586), .A2(n1675), .B1(n1901), .B2(n1674), .ZN(
        n1676) );
  TPNR2D1BWP12T U2611 ( .A1(n1677), .A2(n1676), .ZN(n1680) );
  AOI22D2BWP12T U2612 ( .A1(r5[2]), .A2(n3592), .B1(n3591), .B2(r10[2]), .ZN(
        n1679) );
  AOI22D1BWP12T U2613 ( .A1(n3524), .A2(r7[2]), .B1(n1730), .B2(r2[2]), .ZN(
        n1678) );
  AN4D4BWP12T U2614 ( .A1(n1681), .A2(n1680), .A3(n1679), .A4(n1678), .Z(n1698) );
  INVD1BWP12T U2615 ( .I(r12[2]), .ZN(n1682) );
  OAI22D1BWP12T U2616 ( .A1(n1682), .A2(n3600), .B1(n3599), .B2(n2088), .ZN(
        n1696) );
  INVD1BWP12T U2617 ( .I(n[3698]), .ZN(n1684) );
  INVD1BWP12T U2618 ( .I(r8[2]), .ZN(n1683) );
  TPOAI22D1BWP12T U2619 ( .A1(n1738), .A2(n1684), .B1(n3603), .B2(n1683), .ZN(
        n1695) );
  INVD1BWP12T U2620 ( .I(lr[2]), .ZN(n1687) );
  CKND0BWP12T U2621 ( .I(n242), .ZN(n1686) );
  NR2D1BWP12T U2622 ( .A1(n1687), .A2(n1686), .ZN(n1688) );
  CKND2D0BWP12T U2623 ( .A1(n1688), .A2(n1689), .ZN(n1690) );
  OAI21D1BWP12T U2624 ( .A1(n1740), .A2(n1691), .B(n1690), .ZN(n1694) );
  INVD1BWP12T U2625 ( .I(pc_out[2]), .ZN(n2129) );
  INVD1BWP12T U2626 ( .I(r6[2]), .ZN(n1692) );
  TPOAI22D1BWP12T U2627 ( .A1(n3612), .A2(n2129), .B1(n3611), .B2(n1692), .ZN(
        n1693) );
  NR4D2BWP12T U2628 ( .A1(n1696), .A2(n1695), .A3(n1694), .A4(n1693), .ZN(
        n1697) );
  IOA21D1BWP12T U2629 ( .A1(n3474), .A2(r2[15]), .B(n1701), .ZN(n1709) );
  INVD1BWP12T U2630 ( .I(r10[15]), .ZN(n1704) );
  TPOAI22D1BWP12T U2631 ( .A1(n3481), .A2(n1705), .B1(n3479), .B2(n1704), .ZN(
        n1706) );
  NR4D2BWP12T U2632 ( .A1(n1709), .A2(n1708), .A3(n1706), .A4(n1707), .ZN(
        n1723) );
  TPOAI22D1BWP12T U2633 ( .A1(n3491), .A2(n1711), .B1(n1710), .B2(n3490), .ZN(
        n1721) );
  INVD1BWP12T U2634 ( .I(r5[15]), .ZN(n1713) );
  TPOAI22D1BWP12T U2635 ( .A1(n3463), .A2(n1717), .B1(n1716), .B2(n1715), .ZN(
        n1718) );
  NR4D2BWP12T U2636 ( .A1(n1721), .A2(n1720), .A3(n1719), .A4(n1718), .ZN(
        n1722) );
  TPND2D3BWP12T U2637 ( .A1(n1723), .A2(n1722), .ZN(regA_out[15]) );
  INVD1BWP12T U2638 ( .I(r9[1]), .ZN(n1725) );
  TPOAI22D1BWP12T U2639 ( .A1(n3584), .A2(n1725), .B1(n3582), .B2(n1724), .ZN(
        n1729) );
  INVD1BWP12T U2640 ( .I(r11[1]), .ZN(n1727) );
  INVD1BWP12T U2641 ( .I(r0[1]), .ZN(n1726) );
  TPOAI22D1BWP12T U2642 ( .A1(n3586), .A2(n1727), .B1(n3588), .B2(n1726), .ZN(
        n1728) );
  AOI22D1BWP12T U2643 ( .A1(tmp1[1]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[1]), .ZN(n1733) );
  AOI22D1BWP12T U2644 ( .A1(n1327), .A2(r7[1]), .B1(n1730), .B2(r2[1]), .ZN(
        n1732) );
  INR2D2BWP12T U2645 ( .A1(n1735), .B1(n1734), .ZN(n1747) );
  INVD1BWP12T U2646 ( .I(r1[1]), .ZN(n1736) );
  INVD1BWP12T U2647 ( .I(n[3699]), .ZN(n1737) );
  INVD1BWP12T U2648 ( .I(r8[1]), .ZN(n2819) );
  TPOAI22D1BWP12T U2649 ( .A1(n1738), .A2(n1737), .B1(n3603), .B2(n2819), .ZN(
        n1744) );
  INVD1BWP12T U2650 ( .I(lr[1]), .ZN(n2820) );
  TPOAI22D1BWP12T U2651 ( .A1(n2820), .A2(n3608), .B1(n1740), .B2(n1739), .ZN(
        n1743) );
  INVD1BWP12T U2652 ( .I(pc_out[1]), .ZN(n2915) );
  INVD1BWP12T U2653 ( .I(r6[1]), .ZN(n1741) );
  TPOAI22D1BWP12T U2654 ( .A1(n3612), .A2(n2915), .B1(n3611), .B2(n1741), .ZN(
        n1742) );
  NR4D2BWP12T U2655 ( .A1(n1745), .A2(n1744), .A3(n1743), .A4(n1742), .ZN(
        n1746) );
  TPND2D2BWP12T U2656 ( .A1(n1747), .A2(n1746), .ZN(regB_out[1]) );
  AOI22D1BWP12T U2657 ( .A1(tmp1[24]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[24]), .ZN(n1752) );
  INVD1BWP12T U2658 ( .I(r9[24]), .ZN(n1748) );
  INVD1BWP12T U2659 ( .I(r4[24]), .ZN(n3447) );
  INVD1BWP12T U2660 ( .I(r11[24]), .ZN(n3460) );
  INVD1BWP12T U2661 ( .I(r0[24]), .ZN(n3446) );
  AOI22D1BWP12T U2662 ( .A1(r5[24]), .A2(n3592), .B1(n3591), .B2(r10[24]), 
        .ZN(n1750) );
  AOI22D1BWP12T U2663 ( .A1(r7[24]), .A2(n3524), .B1(n3593), .B2(r2[24]), .ZN(
        n1749) );
  AN4XD1BWP12T U2664 ( .A1(n1752), .A2(n1751), .A3(n1750), .A4(n1749), .Z(
        n1758) );
  INVD1BWP12T U2665 ( .I(lr[24]), .ZN(n3450) );
  INVD1BWP12T U2666 ( .I(r3[24]), .ZN(n3458) );
  OAI22D1BWP12T U2667 ( .A1(n3450), .A2(n3571), .B1(n3607), .B2(n3458), .ZN(
        n1756) );
  INVD1BWP12T U2668 ( .I(n[3676]), .ZN(n3461) );
  INVD1BWP12T U2669 ( .I(r8[24]), .ZN(n3449) );
  OAI22D1BWP12T U2670 ( .A1(n3605), .A2(n3461), .B1(n3603), .B2(n3449), .ZN(
        n1755) );
  INVD1BWP12T U2671 ( .I(r12[24]), .ZN(n3462) );
  INVD1BWP12T U2672 ( .I(r1[24]), .ZN(n3464) );
  OAI22D1BWP12T U2673 ( .A1(n3462), .A2(n3600), .B1(n3599), .B2(n3464), .ZN(
        n1754) );
  INVD1BWP12T U2674 ( .I(r6[24]), .ZN(n3452) );
  OAI22D1BWP12T U2675 ( .A1(n3612), .A2(n3644), .B1(n3611), .B2(n3452), .ZN(
        n1753) );
  NR4D0BWP12T U2676 ( .A1(n1756), .A2(n1755), .A3(n1754), .A4(n1753), .ZN(
        n1757) );
  TPND2D2BWP12T U2677 ( .A1(n1758), .A2(n1757), .ZN(regB_out[24]) );
  AOI22D1BWP12T U2678 ( .A1(tmp1[18]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[18]), .ZN(n1768) );
  INVD1BWP12T U2679 ( .I(r9[18]), .ZN(n1760) );
  OAI22D1BWP12T U2680 ( .A1(n3584), .A2(n1760), .B1(n3582), .B2(n1759), .ZN(
        n1764) );
  OAI22D1BWP12T U2681 ( .A1(n3586), .A2(n1762), .B1(n3588), .B2(n1761), .ZN(
        n1763) );
  TPNR2D1BWP12T U2682 ( .A1(n1764), .A2(n1763), .ZN(n1767) );
  AOI22D1BWP12T U2683 ( .A1(r5[18]), .A2(n3592), .B1(n3591), .B2(r10[18]), 
        .ZN(n1766) );
  AOI22D1BWP12T U2684 ( .A1(r7[18]), .A2(n3524), .B1(n1906), .B2(r2[18]), .ZN(
        n1765) );
  AN4XD1BWP12T U2685 ( .A1(n1768), .A2(n1767), .A3(n1766), .A4(n1765), .Z(
        n1780) );
  OAI22D1BWP12T U2686 ( .A1(n1769), .A2(n3599), .B1(n3600), .B2(n2094), .ZN(
        n1778) );
  OAI22D1BWP12T U2687 ( .A1(n3605), .A2(n1770), .B1(n3603), .B2(n2093), .ZN(
        n1777) );
  OAI22D1BWP12T U2688 ( .A1(n1772), .A2(n1884), .B1(n1913), .B2(n1771), .ZN(
        n1776) );
  OAI22D1BWP12T U2689 ( .A1(n3612), .A2(n1774), .B1(n3611), .B2(n1773), .ZN(
        n1775) );
  AOI22D1BWP12T U2690 ( .A1(n3471), .A2(r9[23]), .B1(n3472), .B2(tmp1[23]), 
        .ZN(n1782) );
  TPND2D1BWP12T U2691 ( .A1(n1782), .A2(n1781), .ZN(n1791) );
  ND2D1BWP12T U2692 ( .A1(n3475), .A2(r4[23]), .ZN(n1783) );
  OAI21D1BWP12T U2693 ( .A1(n3476), .A2(n1784), .B(n1783), .ZN(n1790) );
  INVD1BWP12T U2694 ( .I(r10[23]), .ZN(n1785) );
  TPOAI22D1BWP12T U2695 ( .A1(n3481), .A2(n1786), .B1(n3422), .B2(n1785), .ZN(
        n1789) );
  INVD1BWP12T U2696 ( .I(r7[23]), .ZN(n1792) );
  TPOAI22D1BWP12T U2697 ( .A1(n3487), .A2(n1792), .B1(n3486), .B2(n3314), .ZN(
        n1802) );
  INVD1BWP12T U2698 ( .I(r5[23]), .ZN(n1794) );
  TPOAI22D1BWP12T U2699 ( .A1(n3489), .A2(n1794), .B1(n1793), .B2(n3488), .ZN(
        n1801) );
  TPOAI22D2BWP12T U2700 ( .A1(n3491), .A2(n1796), .B1(n1795), .B2(n3490), .ZN(
        n1800) );
  TPOAI22D1BWP12T U2701 ( .A1(n1798), .A2(n3463), .B1(n3492), .B2(n1797), .ZN(
        n1799) );
  OAI22D0BWP12T U2702 ( .A1(n1803), .A2(n3599), .B1(n3600), .B2(n2676), .ZN(
        n1810) );
  OAI22D1BWP12T U2703 ( .A1(n3605), .A2(n1805), .B1(n3603), .B2(n1804), .ZN(
        n1809) );
  OAI22D1BWP12T U2704 ( .A1(n3612), .A2(n3648), .B1(n3611), .B2(n1807), .ZN(
        n1808) );
  AOI22D1BWP12T U2705 ( .A1(tmp1[28]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[28]), .ZN(n1820) );
  INVD1BWP12T U2706 ( .I(r9[28]), .ZN(n1812) );
  INVD0BWP12T U2707 ( .I(r4[28]), .ZN(n1811) );
  OAI22D1BWP12T U2708 ( .A1(n3584), .A2(n1812), .B1(n3582), .B2(n1811), .ZN(
        n1816) );
  OAI22D0BWP12T U2709 ( .A1(n3586), .A2(n1814), .B1(n3588), .B2(n1813), .ZN(
        n1815) );
  NR2D1BWP12T U2710 ( .A1(n1816), .A2(n1815), .ZN(n1819) );
  AOI22D1BWP12T U2711 ( .A1(r5[28]), .A2(n3592), .B1(n3591), .B2(r10[28]), 
        .ZN(n1818) );
  AOI22D1BWP12T U2712 ( .A1(r7[28]), .A2(n3524), .B1(n3593), .B2(r2[28]), .ZN(
        n1817) );
  AOI22D1BWP12T U2713 ( .A1(r9[22]), .A2(n3471), .B1(n3472), .B2(tmp1[22]), 
        .ZN(n1821) );
  TPOAI22D1BWP12T U2714 ( .A1(n3448), .A2(n1823), .B1(n3476), .B2(n1822), .ZN(
        n1828) );
  OAI22D1BWP12T U2715 ( .A1(n3478), .A2(n2713), .B1(n3477), .B2(n2714), .ZN(
        n1827) );
  INVD1BWP12T U2716 ( .I(r10[22]), .ZN(n1824) );
  TPOAI22D1BWP12T U2717 ( .A1(n3481), .A2(n1825), .B1(n3422), .B2(n1824), .ZN(
        n1826) );
  NR4D0BWP12T U2718 ( .A1(n1829), .A2(n1826), .A3(n1827), .A4(n1828), .ZN(
        n1841) );
  OAI22D1BWP12T U2719 ( .A1(n1831), .A2(n3463), .B1(n3492), .B2(n1830), .ZN(
        n1839) );
  INVD1BWP12T U2720 ( .I(r5[22]), .ZN(n1833) );
  TPOAI22D1BWP12T U2721 ( .A1(n3491), .A2(n2715), .B1(n3490), .B2(n2712), .ZN(
        n1837) );
  INVD1BWP12T U2722 ( .I(r7[22]), .ZN(n1835) );
  TPND2D1BWP12T U2723 ( .A1(n1945), .A2(pc_out[22]), .ZN(n1834) );
  TPOAI21D1BWP12T U2724 ( .A1(n3487), .A2(n1835), .B(n1834), .ZN(n1836) );
  NR4D0BWP12T U2725 ( .A1(n1839), .A2(n1838), .A3(n1837), .A4(n1836), .ZN(
        n1840) );
  TPND2D1BWP12T U2726 ( .A1(n1841), .A2(n1840), .ZN(regA_out[22]) );
  INVD1BWP12T U2727 ( .I(r7[7]), .ZN(n1842) );
  INVD1BWP12T U2728 ( .I(pc_out[7]), .ZN(n1916) );
  TPOAI22D1BWP12T U2729 ( .A1(n3487), .A2(n1842), .B1(n3486), .B2(n1916), .ZN(
        n1847) );
  INVD1BWP12T U2730 ( .I(r5[7]), .ZN(n1843) );
  INVD1BWP12T U2731 ( .I(r3[7]), .ZN(n1912) );
  TPOAI22D1BWP12T U2732 ( .A1(n3489), .A2(n1843), .B1(n3488), .B2(n1912), .ZN(
        n1846) );
  INVD1BWP12T U2733 ( .I(n[3693]), .ZN(n1911) );
  INVD1BWP12T U2734 ( .I(r11[7]), .ZN(n1903) );
  TPOAI22D1BWP12T U2735 ( .A1(n3491), .A2(n1911), .B1(n3490), .B2(n1903), .ZN(
        n1845) );
  INVD1P75BWP12T U2736 ( .I(r12[7]), .ZN(n2808) );
  INVD1P75BWP12T U2737 ( .I(r1[7]), .ZN(n2922) );
  TPOAI22D2BWP12T U2738 ( .A1(n3492), .A2(n2808), .B1(n3463), .B2(n2922), .ZN(
        n1844) );
  NR4D2BWP12T U2739 ( .A1(n1847), .A2(n1846), .A3(n1845), .A4(n1844), .ZN(
        n1855) );
  AOI22D2BWP12T U2740 ( .A1(n3471), .A2(r9[7]), .B1(n3472), .B2(tmp1[7]), .ZN(
        n1849) );
  INVD1BWP12T U2741 ( .I(r4[7]), .ZN(n1898) );
  INVD1BWP12T U2742 ( .I(r0[7]), .ZN(n1900) );
  TPOAI22D2BWP12T U2743 ( .A1(n3448), .A2(n1898), .B1(n3476), .B2(n1900), .ZN(
        n1852) );
  INVD1P75BWP12T U2744 ( .I(lr[7]), .ZN(n2810) );
  INVD1P75BWP12T U2745 ( .I(r8[7]), .ZN(n2807) );
  TPOAI22D2BWP12T U2746 ( .A1(n3478), .A2(n2810), .B1(n3477), .B2(n2807), .ZN(
        n1851) );
  INVD1BWP12T U2747 ( .I(r6[7]), .ZN(n1914) );
  INVD1BWP12T U2748 ( .I(r10[7]), .ZN(n2809) );
  TPOAI22D2BWP12T U2749 ( .A1(n3481), .A2(n1914), .B1(n3479), .B2(n2809), .ZN(
        n1850) );
  NR4D3BWP12T U2750 ( .A1(n1853), .A2(n1852), .A3(n1850), .A4(n1851), .ZN(
        n1854) );
  TPND2D3BWP12T U2751 ( .A1(n1855), .A2(n1854), .ZN(regA_out[7]) );
  BUFFD1BWP12T U2752 ( .I(n3381), .Z(n1856) );
  ND3XD1BWP12T U2753 ( .A1(n1860), .A2(n3333), .A3(n1859), .ZN(n1872) );
  INVD1BWP12T U2754 ( .I(n3340), .ZN(n1861) );
  NR2D1BWP12T U2755 ( .A1(n1861), .A2(n3394), .ZN(n1863) );
  INR2D1BWP12T U2756 ( .A1(n1865), .B1(n1864), .ZN(n1866) );
  ND3D1BWP12T U2757 ( .A1(n1866), .A2(n3333), .A3(n3324), .ZN(n1869) );
  TPND2D1BWP12T U2758 ( .A1(n1869), .A2(n1868), .ZN(n1870) );
  ND3D1BWP12T U2759 ( .A1(n1872), .A2(n1871), .A3(n1870), .ZN(n2196) );
  AOI22D1BWP12T U2760 ( .A1(tmp1[17]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[17]), .ZN(n1882) );
  CKND0BWP12T U2761 ( .I(r9[17]), .ZN(n1874) );
  OAI22D1BWP12T U2762 ( .A1(n3584), .A2(n1874), .B1(n3582), .B2(n1873), .ZN(
        n1878) );
  CKND0BWP12T U2763 ( .I(r11[17]), .ZN(n1876) );
  INVD1BWP12T U2764 ( .I(r0[17]), .ZN(n1875) );
  OAI22D1BWP12T U2765 ( .A1(n3586), .A2(n1876), .B1(n3588), .B2(n1875), .ZN(
        n1877) );
  NR2D1BWP12T U2766 ( .A1(n1878), .A2(n1877), .ZN(n1881) );
  AOI22D1BWP12T U2767 ( .A1(r5[17]), .A2(n3592), .B1(n3591), .B2(r10[17]), 
        .ZN(n1880) );
  AOI22D1BWP12T U2768 ( .A1(r7[17]), .A2(n3524), .B1(n1906), .B2(r2[17]), .ZN(
        n1879) );
  AN4XD1BWP12T U2769 ( .A1(n1881), .A2(n1882), .A3(n1880), .A4(n1879), .Z(
        n1890) );
  INVD1BWP12T U2770 ( .I(n[3683]), .ZN(n2796) );
  OAI22D1BWP12T U2771 ( .A1(n2795), .A2(n1884), .B1(n1913), .B2(n1883), .ZN(
        n1886) );
  NR4D0BWP12T U2772 ( .A1(n1888), .A2(n1887), .A3(n1886), .A4(n1885), .ZN(
        n1889) );
  CKND2D2BWP12T U2773 ( .A1(n1890), .A2(n1889), .ZN(regB_out[17]) );
  MUX2XD2BWP12T U2774 ( .I0(write2_in[17]), .I1(write1_in[17]), .S(n3381), .Z(
        n1962) );
  INR2XD0BWP12T U2775 ( .A1(n3393), .B1(write2_in[18]), .ZN(n1892) );
  INVD1BWP12T U2776 ( .I(n1892), .ZN(n1893) );
  MUX2XD2BWP12T U2777 ( .I0(write2_in[19]), .I1(write1_in[19]), .S(n3381), .Z(
        n1894) );
  XNR2D1BWP12T U2778 ( .A1(n1895), .A2(n1894), .ZN(n1897) );
  AOI22D1BWP12T U2779 ( .A1(n2989), .A2(pc_out[19]), .B1(n3398), .B2(
        next_pc_in[19]), .ZN(n1896) );
  TPOAI21D1BWP12T U2780 ( .A1(n1897), .A2(n3394), .B(n1896), .ZN(n2188) );
  INVD1BWP12T U2781 ( .I(r9[7]), .ZN(n1899) );
  OAI22D1BWP12T U2782 ( .A1(n3584), .A2(n1899), .B1(n3582), .B2(n1898), .ZN(
        n1905) );
  NR2D1BWP12T U2783 ( .A1(n1905), .A2(n1904), .ZN(n1910) );
  AOI22D1BWP12T U2784 ( .A1(r5[7]), .A2(n3592), .B1(n3591), .B2(r10[7]), .ZN(
        n1909) );
  AOI22D1BWP12T U2785 ( .A1(tmp1[7]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[7]), .ZN(n1908) );
  AOI22D1BWP12T U2786 ( .A1(n1906), .A2(r2[7]), .B1(n3524), .B2(r7[7]), .ZN(
        n1907) );
  AN4XD1BWP12T U2787 ( .A1(n1910), .A2(n1909), .A3(n1908), .A4(n1907), .Z(
        n1922) );
  OAI22D1BWP12T U2788 ( .A1(n2808), .A2(n3600), .B1(n3599), .B2(n2922), .ZN(
        n1920) );
  OAI22D1BWP12T U2789 ( .A1(n3605), .A2(n1911), .B1(n3603), .B2(n2807), .ZN(
        n1919) );
  OAI22D1BWP12T U2790 ( .A1(n2810), .A2(n3608), .B1(n1913), .B2(n1912), .ZN(
        n1918) );
  OAI22D1BWP12T U2791 ( .A1(n3612), .A2(n1916), .B1(n1915), .B2(n1914), .ZN(
        n1917) );
  NR4D0BWP12T U2792 ( .A1(n1920), .A2(n1919), .A3(n1918), .A4(n1917), .ZN(
        n1921) );
  TPND2D1BWP12T U2793 ( .A1(n1922), .A2(n1921), .ZN(regB_out[7]) );
  INR2D2BWP12T U2794 ( .A1(r10[12]), .B1(n3479), .ZN(n1925) );
  INVD1P75BWP12T U2795 ( .I(n1925), .ZN(n1928) );
  TPND2D2BWP12T U2796 ( .A1(n1926), .A2(r6[12]), .ZN(n1927) );
  ND4D1BWP12T U2797 ( .A1(n1927), .A2(n1929), .A3(n1928), .A4(n1930), .ZN(
        n1941) );
  ND2D3BWP12T U2798 ( .A1(n235), .A2(r0[12]), .ZN(n1931) );
  OAI21D1BWP12T U2799 ( .A1(n3448), .A2(n1932), .B(n1931), .ZN(n1940) );
  AN2XD2BWP12T U2800 ( .A1(n1933), .A2(r2[12]), .Z(n1935) );
  ND2D1BWP12T U2801 ( .A1(n3471), .A2(r9[12]), .ZN(n1937) );
  ND2D1BWP12T U2802 ( .A1(n3472), .A2(tmp1[12]), .ZN(n1936) );
  ND3D1BWP12T U2803 ( .A1(n1938), .A2(n1937), .A3(n1936), .ZN(n1939) );
  TPNR3D1BWP12T U2804 ( .A1(n1941), .A2(n1940), .A3(n1939), .ZN(n1959) );
  ND2D1BWP12T U2805 ( .A1(n1942), .A2(r5[12]), .ZN(n1943) );
  CKND2D0BWP12T U2806 ( .A1(n1945), .A2(pc_out[12]), .ZN(n1948) );
  ND2D1BWP12T U2807 ( .A1(n1946), .A2(n[3688]), .ZN(n1947) );
  OAI211D1BWP12T U2808 ( .A1(n3490), .A2(n1949), .B(n1948), .C(n1947), .ZN(
        n1956) );
  AOI22D0BWP12T U2809 ( .A1(n1952), .A2(r12[12]), .B1(n1951), .B2(r1[12]), 
        .ZN(n1953) );
  TPNR3D1BWP12T U2810 ( .A1(n1957), .A2(n1956), .A3(n1955), .ZN(n1958) );
  TPND2D1BWP12T U2811 ( .A1(n1959), .A2(n1958), .ZN(regA_out[12]) );
  TPNR2D1BWP12T U2812 ( .A1(n1960), .A2(n1961), .ZN(n1963) );
  XNR2D1BWP12T U2813 ( .A1(n1963), .A2(n1962), .ZN(n1965) );
  AOI22D1BWP12T U2814 ( .A1(n2989), .A2(pc_out[17]), .B1(n3398), .B2(
        next_pc_in[17]), .ZN(n1964) );
  XNR2D1BWP12T U2815 ( .A1(n1967), .A2(n1966), .ZN(n1969) );
  AOI22D1BWP12T U2816 ( .A1(n2989), .A2(pc_out[18]), .B1(n3398), .B2(
        next_pc_in[18]), .ZN(n1968) );
  INVD1BWP12T U2817 ( .I(n1970), .ZN(n1972) );
  ND2D1BWP12T U2818 ( .A1(n1972), .A2(n1971), .ZN(n1974) );
  AOI22D1BWP12T U2819 ( .A1(n2989), .A2(pc_out[20]), .B1(n3398), .B2(
        next_pc_in[20]), .ZN(n1975) );
  TPOAI21D1BWP12T U2820 ( .A1(n1976), .A2(n3394), .B(n1975), .ZN(n2189) );
  XNR2XD2BWP12T U2821 ( .A1(n1978), .A2(n1977), .ZN(n1980) );
  AOI22D1BWP12T U2822 ( .A1(n2989), .A2(pc_out[21]), .B1(n3398), .B2(
        next_pc_in[21]), .ZN(n1979) );
  INVD1BWP12T U2823 ( .I(readC_sel[2]), .ZN(n1983) );
  ND3D1BWP12T U2824 ( .A1(readC_sel[3]), .A2(n2864), .A3(n1983), .ZN(n1981) );
  IND2D1BWP12T U2825 ( .A1(readC_sel[1]), .B1(readC_sel[0]), .ZN(n1990) );
  IND2D1BWP12T U2826 ( .A1(readC_sel[0]), .B1(readC_sel[1]), .ZN(n1984) );
  ND3D1BWP12T U2827 ( .A1(readC_sel[2]), .A2(readC_sel[3]), .A3(n2864), .ZN(
        n1989) );
  ND2D1BWP12T U2828 ( .A1(readC_sel[1]), .A2(readC_sel[0]), .ZN(n1988) );
  CKND1BWP12T U2829 ( .I(readC_sel[3]), .ZN(n1982) );
  ND2D1BWP12T U2830 ( .A1(readC_sel[2]), .A2(n1982), .ZN(n1985) );
  ND2D1BWP12T U2831 ( .A1(n1983), .A2(n1982), .ZN(n1987) );
  TPNR2D0BWP12T U2832 ( .A1(n1990), .A2(n1985), .ZN(n2757) );
  NR2D1BWP12T U2833 ( .A1(n1987), .A2(n1988), .ZN(n2858) );
  INVD1BWP12T U2834 ( .I(n2875), .ZN(n2832) );
  AOI22D0BWP12T U2835 ( .A1(r12[31]), .A2(n2848), .B1(n2874), .B2(pc_out[31]), 
        .ZN(n2001) );
  AOI22D0BWP12T U2836 ( .A1(lr[31]), .A2(n2869), .B1(n2875), .B2(n[3669]), 
        .ZN(n2000) );
  AOI22D0BWP12T U2837 ( .A1(r8[31]), .A2(n2873), .B1(n2870), .B2(r11[31]), 
        .ZN(n1999) );
  AOI22D0BWP12T U2838 ( .A1(r7[31]), .A2(n2854), .B1(n2853), .B2(r4[31]), .ZN(
        n1995) );
  AOI22D0BWP12T U2839 ( .A1(r2[31]), .A2(n2856), .B1(n2855), .B2(r6[31]), .ZN(
        n1994) );
  AOI22D0BWP12T U2840 ( .A1(r5[31]), .A2(n2757), .B1(n2857), .B2(r1[31]), .ZN(
        n1993) );
  AOI22D0BWP12T U2841 ( .A1(r0[31]), .A2(n2859), .B1(n2858), .B2(r3[31]), .ZN(
        n1992) );
  ND4D1BWP12T U2842 ( .A1(n1995), .A2(n1994), .A3(n1993), .A4(n1992), .ZN(
        n1997) );
  CKND1BWP12T U2843 ( .I(r9[31]), .ZN(n3536) );
  INVD1BWP12T U2844 ( .I(r10[31]), .ZN(n3480) );
  OAI22D0BWP12T U2845 ( .A1(n2653), .A2(n3536), .B1(n3480), .B2(n2827), .ZN(
        n1996) );
  AOI21D1BWP12T U2846 ( .A1(n1997), .A2(n2864), .B(n1996), .ZN(n1998) );
  ND4D1BWP12T U2847 ( .A1(n2001), .A2(n2000), .A3(n1999), .A4(n1998), .ZN(
        regC_out[31]) );
  AOI22D0BWP12T U2848 ( .A1(pc_out[29]), .A2(n2874), .B1(n2873), .B2(r8[29]), 
        .ZN(n2011) );
  AOI22D0BWP12T U2849 ( .A1(lr[29]), .A2(n2869), .B1(n2848), .B2(r12[29]), 
        .ZN(n2010) );
  AOI22D0BWP12T U2850 ( .A1(r10[29]), .A2(n2872), .B1(n2870), .B2(r11[29]), 
        .ZN(n2009) );
  AOI22D0BWP12T U2851 ( .A1(r7[29]), .A2(n2854), .B1(n2853), .B2(r4[29]), .ZN(
        n2005) );
  AOI22D0BWP12T U2852 ( .A1(r2[29]), .A2(n2856), .B1(n2855), .B2(r6[29]), .ZN(
        n2004) );
  AOI22D0BWP12T U2853 ( .A1(r5[29]), .A2(n2757), .B1(n2857), .B2(r1[29]), .ZN(
        n2003) );
  AOI22D0BWP12T U2854 ( .A1(r0[29]), .A2(n2859), .B1(n2858), .B2(r3[29]), .ZN(
        n2002) );
  ND4D1BWP12T U2855 ( .A1(n2005), .A2(n2004), .A3(n2003), .A4(n2002), .ZN(
        n2007) );
  INVD1BWP12T U2856 ( .I(r9[29]), .ZN(n3559) );
  OAI22D0BWP12T U2857 ( .A1(n3570), .A2(n2832), .B1(n2653), .B2(n3559), .ZN(
        n2006) );
  AOI21D1BWP12T U2858 ( .A1(n2007), .A2(n2864), .B(n2006), .ZN(n2008) );
  ND4D1BWP12T U2859 ( .A1(n2011), .A2(n2010), .A3(n2009), .A4(n2008), .ZN(
        regC_out[29]) );
  AOI22D0BWP12T U2860 ( .A1(pc_out[27]), .A2(n2874), .B1(n2873), .B2(r8[27]), 
        .ZN(n2021) );
  AOI22D0BWP12T U2861 ( .A1(lr[27]), .A2(n2869), .B1(n2848), .B2(r12[27]), 
        .ZN(n2020) );
  AOI22D0BWP12T U2862 ( .A1(r9[27]), .A2(n2871), .B1(n2872), .B2(r10[27]), 
        .ZN(n2019) );
  AOI22D0BWP12T U2863 ( .A1(r7[27]), .A2(n2854), .B1(n2853), .B2(r4[27]), .ZN(
        n2015) );
  AOI22D0BWP12T U2864 ( .A1(r2[27]), .A2(n2856), .B1(n2855), .B2(r6[27]), .ZN(
        n2014) );
  AOI22D0BWP12T U2865 ( .A1(r5[27]), .A2(n2757), .B1(n2857), .B2(r1[27]), .ZN(
        n2013) );
  AOI22D0BWP12T U2866 ( .A1(r0[27]), .A2(n2859), .B1(n2858), .B2(r3[27]), .ZN(
        n2012) );
  ND4D1BWP12T U2867 ( .A1(n2015), .A2(n2014), .A3(n2013), .A4(n2012), .ZN(
        n2017) );
  OAI22D0BWP12T U2868 ( .A1(n3435), .A2(n2832), .B1(n2711), .B2(n3434), .ZN(
        n2016) );
  AOI21D1BWP12T U2869 ( .A1(n2017), .A2(n2864), .B(n2016), .ZN(n2018) );
  ND4D1BWP12T U2870 ( .A1(n2021), .A2(n2020), .A3(n2019), .A4(n2018), .ZN(
        regC_out[27]) );
  AOI22D0BWP12T U2871 ( .A1(pc_out[20]), .A2(n2874), .B1(n2873), .B2(r8[20]), 
        .ZN(n2033) );
  AOI22D0BWP12T U2872 ( .A1(lr[20]), .A2(n2869), .B1(n2848), .B2(r12[20]), 
        .ZN(n2032) );
  AOI22D0BWP12T U2873 ( .A1(r9[20]), .A2(n2871), .B1(n2872), .B2(r10[20]), 
        .ZN(n2031) );
  AOI22D0BWP12T U2874 ( .A1(r7[20]), .A2(n2854), .B1(n2853), .B2(r4[20]), .ZN(
        n2025) );
  AOI22D0BWP12T U2875 ( .A1(r2[20]), .A2(n2856), .B1(n2855), .B2(r6[20]), .ZN(
        n2024) );
  AOI22D0BWP12T U2876 ( .A1(r5[20]), .A2(n2757), .B1(n2857), .B2(r1[20]), .ZN(
        n2023) );
  AOI22D0BWP12T U2877 ( .A1(r0[20]), .A2(n2859), .B1(n2858), .B2(r3[20]), .ZN(
        n2022) );
  ND4D1BWP12T U2878 ( .A1(n2025), .A2(n2024), .A3(n2023), .A4(n2022), .ZN(
        n2029) );
  OAI22D0BWP12T U2879 ( .A1(n2027), .A2(n2832), .B1(n2711), .B2(n2026), .ZN(
        n2028) );
  AOI21D1BWP12T U2880 ( .A1(n2029), .A2(n2864), .B(n2028), .ZN(n2030) );
  ND4D1BWP12T U2881 ( .A1(n2033), .A2(n2032), .A3(n2031), .A4(n2030), .ZN(
        regC_out[20]) );
  AOI22D0BWP12T U2882 ( .A1(r12[9]), .A2(n2848), .B1(n2874), .B2(pc_out[9]), 
        .ZN(n2045) );
  AOI22D0BWP12T U2883 ( .A1(lr[9]), .A2(n2869), .B1(n2875), .B2(n[3691]), .ZN(
        n2044) );
  AOI22D0BWP12T U2884 ( .A1(r10[9]), .A2(n2872), .B1(n2870), .B2(r11[9]), .ZN(
        n2043) );
  AOI22D0BWP12T U2885 ( .A1(r7[9]), .A2(n2854), .B1(n2853), .B2(r4[9]), .ZN(
        n2037) );
  AOI22D0BWP12T U2886 ( .A1(r2[9]), .A2(n2856), .B1(n2855), .B2(r6[9]), .ZN(
        n2036) );
  AOI22D0BWP12T U2887 ( .A1(r5[9]), .A2(n2757), .B1(n2857), .B2(r1[9]), .ZN(
        n2035) );
  AOI22D0BWP12T U2888 ( .A1(r0[9]), .A2(n2859), .B1(n2858), .B2(r3[9]), .ZN(
        n2034) );
  ND4D1BWP12T U2889 ( .A1(n2037), .A2(n2036), .A3(n2035), .A4(n2034), .ZN(
        n2041) );
  INVD1BWP12T U2890 ( .I(n2873), .ZN(n2830) );
  OAI22D0BWP12T U2891 ( .A1(n2830), .A2(n2039), .B1(n2038), .B2(n2653), .ZN(
        n2040) );
  AOI21D1BWP12T U2892 ( .A1(n2041), .A2(n2864), .B(n2040), .ZN(n2042) );
  ND4D1BWP12T U2893 ( .A1(n2045), .A2(n2044), .A3(n2043), .A4(n2042), .ZN(
        regC_out[9]) );
  AOI22D0BWP12T U2894 ( .A1(r12[25]), .A2(n2848), .B1(n2871), .B2(r9[25]), 
        .ZN(n2055) );
  AOI22D0BWP12T U2895 ( .A1(lr[25]), .A2(n2869), .B1(n2875), .B2(n[3675]), 
        .ZN(n2054) );
  AOI22D0BWP12T U2896 ( .A1(r10[25]), .A2(n2872), .B1(n2870), .B2(r11[25]), 
        .ZN(n2053) );
  AOI22D0BWP12T U2897 ( .A1(r7[25]), .A2(n2854), .B1(n2853), .B2(r4[25]), .ZN(
        n2049) );
  AOI22D0BWP12T U2898 ( .A1(r2[25]), .A2(n2856), .B1(n2855), .B2(r6[25]), .ZN(
        n2048) );
  AOI22D0BWP12T U2899 ( .A1(r5[25]), .A2(n2757), .B1(n2857), .B2(r1[25]), .ZN(
        n2047) );
  AOI22D0BWP12T U2900 ( .A1(r0[25]), .A2(n2859), .B1(n2858), .B2(r3[25]), .ZN(
        n2046) );
  ND4D1BWP12T U2901 ( .A1(n2049), .A2(n2048), .A3(n2047), .A4(n2046), .ZN(
        n2051) );
  OAI22D0BWP12T U2902 ( .A1(n3645), .A2(n2822), .B1(n2830), .B2(n3511), .ZN(
        n2050) );
  AOI21D1BWP12T U2903 ( .A1(n2051), .A2(n2864), .B(n2050), .ZN(n2052) );
  ND4D1BWP12T U2904 ( .A1(n2055), .A2(n2054), .A3(n2053), .A4(n2052), .ZN(
        regC_out[25]) );
  NR2XD0BWP12T U2905 ( .A1(readD_sel[1]), .A2(readD_sel[0]), .ZN(n2069) );
  INVD1BWP12T U2906 ( .I(n2069), .ZN(n2060) );
  IND2D1BWP12T U2907 ( .A1(readD_sel[2]), .B1(readD_sel[3]), .ZN(n2059) );
  NR2D1BWP12T U2908 ( .A1(n2060), .A2(n2059), .ZN(n2954) );
  IND2D1BWP12T U2909 ( .A1(readD_sel[3]), .B1(readD_sel[2]), .ZN(n2058) );
  NR2D1BWP12T U2910 ( .A1(n2060), .A2(n2058), .ZN(n2953) );
  AOI22D0BWP12T U2911 ( .A1(r8[3]), .A2(n2954), .B1(n2953), .B2(r4[3]), .ZN(
        n2057) );
  ND2D1BWP12T U2912 ( .A1(readD_sel[3]), .A2(readD_sel[2]), .ZN(n2071) );
  IND2D1BWP12T U2913 ( .A1(readD_sel[1]), .B1(readD_sel[0]), .ZN(n2065) );
  NR2D1BWP12T U2914 ( .A1(n2071), .A2(n2065), .ZN(n2956) );
  IND2D1BWP12T U2915 ( .A1(readD_sel[0]), .B1(readD_sel[1]), .ZN(n2067) );
  NR2D1BWP12T U2916 ( .A1(n2059), .A2(n2067), .ZN(n2955) );
  AOI22D0BWP12T U2917 ( .A1(n[3697]), .A2(n2956), .B1(n2955), .B2(r10[3]), 
        .ZN(n2056) );
  CKND2D1BWP12T U2918 ( .A1(n2057), .A2(n2056), .ZN(n2077) );
  CKND2D1BWP12T U2919 ( .A1(readD_sel[1]), .A2(readD_sel[0]), .ZN(n2070) );
  NR2D1BWP12T U2920 ( .A1(n2070), .A2(n2058), .ZN(n2958) );
  NR2D1BWP12T U2921 ( .A1(n2065), .A2(n2058), .ZN(n2957) );
  AOI22D0BWP12T U2922 ( .A1(r7[3]), .A2(n2958), .B1(n2957), .B2(r5[3]), .ZN(
        n2064) );
  NR2D1BWP12T U2923 ( .A1(n2071), .A2(n2067), .ZN(n2960) );
  NR2D1BWP12T U2924 ( .A1(n2059), .A2(n2065), .ZN(n2959) );
  AOI22D0BWP12T U2925 ( .A1(lr[3]), .A2(n2960), .B1(n2959), .B2(r9[3]), .ZN(
        n2063) );
  NR2D1BWP12T U2926 ( .A1(n2067), .A2(n2058), .ZN(n2962) );
  NR2D1BWP12T U2927 ( .A1(n2059), .A2(n2070), .ZN(n2961) );
  AOI22D0BWP12T U2928 ( .A1(r6[3]), .A2(n2962), .B1(n2961), .B2(r11[3]), .ZN(
        n2062) );
  NR2D1BWP12T U2929 ( .A1(n2071), .A2(n2060), .ZN(n2963) );
  CKND2D0BWP12T U2930 ( .A1(n2963), .A2(r12[3]), .ZN(n2061) );
  ND4D1BWP12T U2931 ( .A1(n2064), .A2(n2063), .A3(n2062), .A4(n2061), .ZN(
        n2076) );
  NR2D1BWP12T U2932 ( .A1(readD_sel[3]), .A2(readD_sel[2]), .ZN(n2068) );
  INVD1BWP12T U2933 ( .I(n2068), .ZN(n2066) );
  OR2XD1BWP12T U2934 ( .A1(n2065), .A2(n2066), .Z(n2968) );
  NR2D1BWP12T U2935 ( .A1(n2070), .A2(n2066), .ZN(n2965) );
  NR2D1BWP12T U2936 ( .A1(n2067), .A2(n2066), .ZN(n2964) );
  AOI22D0BWP12T U2937 ( .A1(r3[3]), .A2(n2965), .B1(n2964), .B2(r2[3]), .ZN(
        n2073) );
  AN2XD1BWP12T U2938 ( .A1(n2069), .A2(n2068), .Z(n2967) );
  NR2D1BWP12T U2939 ( .A1(n2071), .A2(n2070), .ZN(n2966) );
  AOI22D0BWP12T U2940 ( .A1(n2967), .A2(r0[3]), .B1(pc_out[3]), .B2(n2966), 
        .ZN(n2072) );
  OAI211D0BWP12T U2941 ( .A1(n2074), .A2(n2968), .B(n2073), .C(n2072), .ZN(
        n2075) );
  OA31D1BWP12T U2942 ( .A1(n2077), .A2(n2076), .A3(n2075), .B(n2970), .Z(
        regD_out[3]) );
  AOI22D0BWP12T U2943 ( .A1(lr[30]), .A2(n2869), .B1(n2875), .B2(n[3670]), 
        .ZN(n2087) );
  AOI22D0BWP12T U2944 ( .A1(r9[30]), .A2(n2871), .B1(n2872), .B2(r10[30]), 
        .ZN(n2086) );
  AOI22D0BWP12T U2945 ( .A1(r7[30]), .A2(n2854), .B1(n2853), .B2(r4[30]), .ZN(
        n2081) );
  AOI22D0BWP12T U2946 ( .A1(r2[30]), .A2(n2856), .B1(n2855), .B2(r6[30]), .ZN(
        n2080) );
  AOI22D0BWP12T U2947 ( .A1(r5[30]), .A2(n2757), .B1(n2857), .B2(r1[30]), .ZN(
        n2079) );
  AOI22D0BWP12T U2948 ( .A1(r0[30]), .A2(n2859), .B1(n2858), .B2(r3[30]), .ZN(
        n2078) );
  ND4D1BWP12T U2949 ( .A1(n2081), .A2(n2080), .A3(n2079), .A4(n2078), .ZN(
        n2084) );
  INVD1BWP12T U2950 ( .I(n2848), .ZN(n2867) );
  OAI22D0BWP12T U2951 ( .A1(n2867), .A2(n3665), .B1(n3663), .B2(n2711), .ZN(
        n2083) );
  OAI22D0BWP12T U2952 ( .A1(n3659), .A2(n2822), .B1(n2830), .B2(n3655), .ZN(
        n2082) );
  AOI211D1BWP12T U2953 ( .A1(n2084), .A2(n2864), .B(n2083), .C(n2082), .ZN(
        n2085) );
  ND3D1BWP12T U2954 ( .A1(n2087), .A2(n2086), .A3(n2085), .ZN(regC_out[30]) );
  AOI22D0BWP12T U2955 ( .A1(pc_out[18]), .A2(n2874), .B1(n2871), .B2(r9[18]), 
        .ZN(n2100) );
  AOI22D0BWP12T U2956 ( .A1(lr[18]), .A2(n2869), .B1(n2875), .B2(n[3682]), 
        .ZN(n2099) );
  AOI22D0BWP12T U2957 ( .A1(r10[18]), .A2(n2872), .B1(n2870), .B2(r11[18]), 
        .ZN(n2098) );
  AOI22D0BWP12T U2958 ( .A1(r7[18]), .A2(n2854), .B1(n2853), .B2(r4[18]), .ZN(
        n2092) );
  AOI22D0BWP12T U2959 ( .A1(r2[18]), .A2(n2856), .B1(n2855), .B2(r6[18]), .ZN(
        n2091) );
  AOI22D0BWP12T U2960 ( .A1(r5[18]), .A2(n2757), .B1(n2857), .B2(r1[18]), .ZN(
        n2090) );
  AOI22D0BWP12T U2961 ( .A1(r0[18]), .A2(n2859), .B1(n2858), .B2(r3[18]), .ZN(
        n2089) );
  ND4D1BWP12T U2962 ( .A1(n2092), .A2(n2091), .A3(n2090), .A4(n2089), .ZN(
        n2096) );
  OAI22D0BWP12T U2963 ( .A1(n2867), .A2(n2094), .B1(n2093), .B2(n2830), .ZN(
        n2095) );
  AOI21D1BWP12T U2964 ( .A1(n2096), .A2(n2864), .B(n2095), .ZN(n2097) );
  ND4D1BWP12T U2965 ( .A1(n2100), .A2(n2099), .A3(n2098), .A4(n2097), .ZN(
        regC_out[18]) );
  AOI22D0BWP12T U2966 ( .A1(pc_out[8]), .A2(n2874), .B1(n2871), .B2(r9[8]), 
        .ZN(n2112) );
  AOI22D0BWP12T U2967 ( .A1(lr[8]), .A2(n2869), .B1(n2875), .B2(n[3692]), .ZN(
        n2111) );
  AOI22D0BWP12T U2968 ( .A1(r10[8]), .A2(n2872), .B1(n2870), .B2(r11[8]), .ZN(
        n2110) );
  AOI22D0BWP12T U2969 ( .A1(r7[8]), .A2(n2854), .B1(n2853), .B2(r4[8]), .ZN(
        n2104) );
  AOI22D0BWP12T U2970 ( .A1(r2[8]), .A2(n2856), .B1(n2855), .B2(r6[8]), .ZN(
        n2103) );
  AOI22D0BWP12T U2971 ( .A1(r5[8]), .A2(n2757), .B1(n2857), .B2(r1[8]), .ZN(
        n2102) );
  AOI22D0BWP12T U2972 ( .A1(r0[8]), .A2(n2859), .B1(n2858), .B2(r3[8]), .ZN(
        n2101) );
  ND4D1BWP12T U2973 ( .A1(n2104), .A2(n2103), .A3(n2102), .A4(n2101), .ZN(
        n2108) );
  OAI22D0BWP12T U2974 ( .A1(n2867), .A2(n2106), .B1(n2105), .B2(n2830), .ZN(
        n2107) );
  AOI21D1BWP12T U2975 ( .A1(n2108), .A2(n2864), .B(n2107), .ZN(n2109) );
  ND4D1BWP12T U2976 ( .A1(n2112), .A2(n2111), .A3(n2110), .A4(n2109), .ZN(
        regC_out[8]) );
  AOI22D0BWP12T U2977 ( .A1(r7[10]), .A2(n2854), .B1(n2853), .B2(r4[10]), .ZN(
        n2116) );
  AOI22D0BWP12T U2978 ( .A1(r2[10]), .A2(n2856), .B1(n2855), .B2(r6[10]), .ZN(
        n2115) );
  AOI22D0BWP12T U2979 ( .A1(r5[10]), .A2(n2757), .B1(n2857), .B2(r1[10]), .ZN(
        n2114) );
  AOI22D0BWP12T U2980 ( .A1(r0[10]), .A2(n2859), .B1(n2858), .B2(r3[10]), .ZN(
        n2113) );
  ND4D1BWP12T U2981 ( .A1(n2116), .A2(n2115), .A3(n2114), .A4(n2113), .ZN(
        n2117) );
  MOAI22D0BWP12T U2982 ( .A1(n2832), .A2(n2118), .B1(n2117), .B2(n2864), .ZN(
        n2119) );
  AOI21D0BWP12T U2983 ( .A1(lr[10]), .A2(n2869), .B(n2119), .ZN(n2123) );
  AOI22D0BWP12T U2984 ( .A1(r9[10]), .A2(n2871), .B1(n2870), .B2(r11[10]), 
        .ZN(n2122) );
  AOI22D0BWP12T U2985 ( .A1(r8[10]), .A2(n2873), .B1(n2872), .B2(r10[10]), 
        .ZN(n2121) );
  AOI22D0BWP12T U2986 ( .A1(r12[10]), .A2(n2848), .B1(n2874), .B2(pc_out[10]), 
        .ZN(n2120) );
  ND4D1BWP12T U2987 ( .A1(n2123), .A2(n2122), .A3(n2121), .A4(n2120), .ZN(
        regC_out[10]) );
  AOI22D0BWP12T U2988 ( .A1(r7[2]), .A2(n2854), .B1(n2853), .B2(r4[2]), .ZN(
        n2127) );
  AOI22D0BWP12T U2989 ( .A1(r2[2]), .A2(n2856), .B1(n2855), .B2(r6[2]), .ZN(
        n2126) );
  AOI22D0BWP12T U2990 ( .A1(r5[2]), .A2(n2757), .B1(n2857), .B2(r1[2]), .ZN(
        n2125) );
  AOI22D0BWP12T U2991 ( .A1(r0[2]), .A2(n2859), .B1(n2858), .B2(r3[2]), .ZN(
        n2124) );
  ND4D1BWP12T U2992 ( .A1(n2127), .A2(n2126), .A3(n2125), .A4(n2124), .ZN(
        n2128) );
  MOAI22D0BWP12T U2993 ( .A1(n2822), .A2(n2129), .B1(n2128), .B2(n2864), .ZN(
        n2130) );
  AOI21D0BWP12T U2994 ( .A1(lr[2]), .A2(n2869), .B(n2130), .ZN(n2134) );
  AOI22D0BWP12T U2995 ( .A1(r9[2]), .A2(n2871), .B1(n2870), .B2(r11[2]), .ZN(
        n2133) );
  AOI22D0BWP12T U2996 ( .A1(r8[2]), .A2(n2873), .B1(n2872), .B2(r10[2]), .ZN(
        n2132) );
  AOI22D0BWP12T U2997 ( .A1(r12[2]), .A2(n2848), .B1(n2875), .B2(n[3698]), 
        .ZN(n2131) );
  ND4D1BWP12T U2998 ( .A1(n2134), .A2(n2133), .A3(n2132), .A4(n2131), .ZN(
        regC_out[2]) );
  AOI22D0BWP12T U2999 ( .A1(pc_out[5]), .A2(n2874), .B1(n2873), .B2(r8[5]), 
        .ZN(n2583) );
  AOI22D0BWP12T U3000 ( .A1(r12[5]), .A2(n2848), .B1(n2875), .B2(n[3695]), 
        .ZN(n2551) );
  AOI22D0BWP12T U3001 ( .A1(r10[5]), .A2(n2872), .B1(n2870), .B2(r11[5]), .ZN(
        n2550) );
  AOI22D0BWP12T U3002 ( .A1(r7[5]), .A2(n2854), .B1(n2853), .B2(r4[5]), .ZN(
        n2294) );
  AOI22D0BWP12T U3003 ( .A1(r2[5]), .A2(n2856), .B1(n2855), .B2(r6[5]), .ZN(
        n2167) );
  AOI22D0BWP12T U3004 ( .A1(r5[5]), .A2(n2757), .B1(n2857), .B2(r1[5]), .ZN(
        n2137) );
  AOI22D0BWP12T U3005 ( .A1(r0[5]), .A2(n2859), .B1(n2858), .B2(r3[5]), .ZN(
        n2135) );
  ND4D1BWP12T U3006 ( .A1(n2294), .A2(n2167), .A3(n2137), .A4(n2135), .ZN(
        n2487) );
  INVD1BWP12T U3007 ( .I(n2869), .ZN(n2846) );
  OAI22D0BWP12T U3008 ( .A1(n2846), .A2(n2327), .B1(n2326), .B2(n2653), .ZN(
        n2455) );
  AOI21D0BWP12T U3009 ( .A1(n2487), .A2(n2864), .B(n2455), .ZN(n2519) );
  ND4D1BWP12T U3010 ( .A1(n2583), .A2(n2551), .A3(n2550), .A4(n2519), .ZN(
        regC_out[5]) );
  AOI22D0BWP12T U3011 ( .A1(pc_out[19]), .A2(n2874), .B1(n2873), .B2(r8[19]), 
        .ZN(n2659) );
  AOI22D0BWP12T U3012 ( .A1(n[3681]), .A2(n2875), .B1(n2848), .B2(r12[19]), 
        .ZN(n2658) );
  AOI22D0BWP12T U3013 ( .A1(r10[19]), .A2(n2872), .B1(n2870), .B2(r11[19]), 
        .ZN(n2657) );
  AOI22D0BWP12T U3014 ( .A1(r7[19]), .A2(n2854), .B1(n2853), .B2(r4[19]), .ZN(
        n2652) );
  AOI22D0BWP12T U3015 ( .A1(r2[19]), .A2(n2856), .B1(n2855), .B2(r6[19]), .ZN(
        n2651) );
  AOI22D0BWP12T U3016 ( .A1(r5[19]), .A2(n2757), .B1(n2857), .B2(r1[19]), .ZN(
        n2650) );
  AOI22D0BWP12T U3017 ( .A1(r0[19]), .A2(n2859), .B1(n2858), .B2(r3[19]), .ZN(
        n2649) );
  ND4D1BWP12T U3018 ( .A1(n2652), .A2(n2651), .A3(n2650), .A4(n2649), .ZN(
        n2655) );
  INVD1BWP12T U3019 ( .I(r9[19]), .ZN(n3583) );
  OAI22D0BWP12T U3020 ( .A1(n2846), .A2(n3609), .B1(n3583), .B2(n2653), .ZN(
        n2654) );
  AOI21D1BWP12T U3021 ( .A1(n2655), .A2(n2864), .B(n2654), .ZN(n2656) );
  ND4D1BWP12T U3022 ( .A1(n2659), .A2(n2658), .A3(n2657), .A4(n2656), .ZN(
        regC_out[19]) );
  AOI22D0BWP12T U3023 ( .A1(pc_out[0]), .A2(n2874), .B1(n2873), .B2(r8[0]), 
        .ZN(n2671) );
  AOI22D0BWP12T U3024 ( .A1(n[3700]), .A2(n2875), .B1(n2848), .B2(r12[0]), 
        .ZN(n2670) );
  AOI22D0BWP12T U3025 ( .A1(r9[0]), .A2(n2871), .B1(n2870), .B2(r11[0]), .ZN(
        n2669) );
  AOI22D0BWP12T U3026 ( .A1(r7[0]), .A2(n2854), .B1(n2853), .B2(r4[0]), .ZN(
        n2663) );
  AOI22D0BWP12T U3027 ( .A1(r2[0]), .A2(n2856), .B1(n2855), .B2(r6[0]), .ZN(
        n2662) );
  AOI22D0BWP12T U3028 ( .A1(r5[0]), .A2(n2757), .B1(n2857), .B2(r1[0]), .ZN(
        n2661) );
  AOI22D0BWP12T U3029 ( .A1(r0[0]), .A2(n2859), .B1(n2858), .B2(r3[0]), .ZN(
        n2660) );
  ND4D1BWP12T U3030 ( .A1(n2663), .A2(n2662), .A3(n2661), .A4(n2660), .ZN(
        n2667) );
  OAI22D0BWP12T U3031 ( .A1(n2846), .A2(n2665), .B1(n2664), .B2(n2827), .ZN(
        n2666) );
  AOI21D1BWP12T U3032 ( .A1(n2667), .A2(n2864), .B(n2666), .ZN(n2668) );
  ND4D1BWP12T U3033 ( .A1(n2671), .A2(n2670), .A3(n2669), .A4(n2668), .ZN(
        regC_out[0]) );
  AOI22D0BWP12T U3034 ( .A1(r8[28]), .A2(n2873), .B1(n2872), .B2(r10[28]), 
        .ZN(n2683) );
  AOI22D0BWP12T U3035 ( .A1(n[3672]), .A2(n2875), .B1(n2874), .B2(pc_out[28]), 
        .ZN(n2682) );
  AOI22D0BWP12T U3036 ( .A1(r9[28]), .A2(n2871), .B1(n2870), .B2(r11[28]), 
        .ZN(n2681) );
  AOI22D0BWP12T U3037 ( .A1(r7[28]), .A2(n2854), .B1(n2853), .B2(r4[28]), .ZN(
        n2675) );
  AOI22D0BWP12T U3038 ( .A1(r2[28]), .A2(n2856), .B1(n2855), .B2(r6[28]), .ZN(
        n2674) );
  AOI22D0BWP12T U3039 ( .A1(r5[28]), .A2(n2757), .B1(n2857), .B2(r1[28]), .ZN(
        n2673) );
  AOI22D0BWP12T U3040 ( .A1(r0[28]), .A2(n2859), .B1(n2858), .B2(r3[28]), .ZN(
        n2672) );
  ND4D1BWP12T U3041 ( .A1(n2675), .A2(n2674), .A3(n2673), .A4(n2672), .ZN(
        n2679) );
  OAI22D0BWP12T U3042 ( .A1(n2846), .A2(n2677), .B1(n2676), .B2(n2867), .ZN(
        n2678) );
  AOI21D1BWP12T U3043 ( .A1(n2679), .A2(n2864), .B(n2678), .ZN(n2680) );
  ND4D1BWP12T U3044 ( .A1(n2683), .A2(n2682), .A3(n2681), .A4(n2680), .ZN(
        regC_out[28]) );
  AOI22D0BWP12T U3045 ( .A1(r7[23]), .A2(n2854), .B1(n2853), .B2(r4[23]), .ZN(
        n2687) );
  AOI22D0BWP12T U3046 ( .A1(r2[23]), .A2(n2856), .B1(n2855), .B2(r6[23]), .ZN(
        n2686) );
  AOI22D0BWP12T U3047 ( .A1(r5[23]), .A2(n2757), .B1(n2857), .B2(r1[23]), .ZN(
        n2685) );
  AOI22D0BWP12T U3048 ( .A1(r0[23]), .A2(n2859), .B1(n2858), .B2(r3[23]), .ZN(
        n2684) );
  ND4D1BWP12T U3049 ( .A1(n2687), .A2(n2686), .A3(n2685), .A4(n2684), .ZN(
        n2688) );
  MOAI22D0BWP12T U3050 ( .A1(n2830), .A2(n2689), .B1(n2688), .B2(n2864), .ZN(
        n2690) );
  AOI21D0BWP12T U3051 ( .A1(lr[23]), .A2(n2869), .B(n2690), .ZN(n2694) );
  AOI22D0BWP12T U3052 ( .A1(r9[23]), .A2(n2871), .B1(n2870), .B2(r11[23]), 
        .ZN(n2693) );
  AOI22D0BWP12T U3053 ( .A1(pc_out[23]), .A2(n2874), .B1(n2872), .B2(r10[23]), 
        .ZN(n2692) );
  AOI22D0BWP12T U3054 ( .A1(n[3677]), .A2(n2875), .B1(n2848), .B2(r12[23]), 
        .ZN(n2691) );
  ND4D1BWP12T U3055 ( .A1(n2694), .A2(n2693), .A3(n2692), .A4(n2691), .ZN(
        regC_out[23]) );
  AOI22D0BWP12T U3056 ( .A1(pc_out[15]), .A2(n2874), .B1(n2872), .B2(r10[15]), 
        .ZN(n2706) );
  AOI22D0BWP12T U3057 ( .A1(n[3685]), .A2(n2875), .B1(n2848), .B2(r12[15]), 
        .ZN(n2705) );
  AOI22D0BWP12T U3058 ( .A1(r9[15]), .A2(n2871), .B1(n2870), .B2(r11[15]), 
        .ZN(n2704) );
  AOI22D0BWP12T U3059 ( .A1(r7[15]), .A2(n2854), .B1(n2853), .B2(r4[15]), .ZN(
        n2698) );
  AOI22D0BWP12T U3060 ( .A1(r2[15]), .A2(n2856), .B1(n2855), .B2(r6[15]), .ZN(
        n2697) );
  AOI22D0BWP12T U3061 ( .A1(r5[15]), .A2(n2757), .B1(n2857), .B2(r1[15]), .ZN(
        n2696) );
  AOI22D0BWP12T U3062 ( .A1(r0[15]), .A2(n2859), .B1(n2858), .B2(r3[15]), .ZN(
        n2695) );
  ND4D1BWP12T U3063 ( .A1(n2698), .A2(n2697), .A3(n2696), .A4(n2695), .ZN(
        n2702) );
  OAI22D0BWP12T U3064 ( .A1(n2846), .A2(n2700), .B1(n2699), .B2(n2830), .ZN(
        n2701) );
  AOI21D1BWP12T U3065 ( .A1(n2702), .A2(n2864), .B(n2701), .ZN(n2703) );
  ND4D1BWP12T U3066 ( .A1(n2706), .A2(n2705), .A3(n2704), .A4(n2703), .ZN(
        regC_out[15]) );
  AOI22D0BWP12T U3067 ( .A1(r12[22]), .A2(n2848), .B1(n2874), .B2(pc_out[22]), 
        .ZN(n2721) );
  AOI22D0BWP12T U3068 ( .A1(r9[22]), .A2(n2871), .B1(n2872), .B2(r10[22]), 
        .ZN(n2720) );
  AOI22D0BWP12T U3069 ( .A1(r7[22]), .A2(n2854), .B1(n2853), .B2(r4[22]), .ZN(
        n2710) );
  AOI22D0BWP12T U3070 ( .A1(r2[22]), .A2(n2856), .B1(n2855), .B2(r6[22]), .ZN(
        n2709) );
  AOI22D0BWP12T U3071 ( .A1(r5[22]), .A2(n2757), .B1(n2857), .B2(r1[22]), .ZN(
        n2708) );
  AOI22D0BWP12T U3072 ( .A1(r0[22]), .A2(n2859), .B1(n2858), .B2(r3[22]), .ZN(
        n2707) );
  ND4D1BWP12T U3073 ( .A1(n2710), .A2(n2709), .A3(n2708), .A4(n2707), .ZN(
        n2718) );
  OAI22D0BWP12T U3074 ( .A1(n2846), .A2(n2713), .B1(n2712), .B2(n2711), .ZN(
        n2717) );
  OAI22D0BWP12T U3075 ( .A1(n2715), .A2(n2832), .B1(n2830), .B2(n2714), .ZN(
        n2716) );
  AOI211D1BWP12T U3076 ( .A1(n2718), .A2(n2864), .B(n2717), .C(n2716), .ZN(
        n2719) );
  ND3D1BWP12T U3077 ( .A1(n2721), .A2(n2720), .A3(n2719), .ZN(regC_out[22]) );
  AOI22D0BWP12T U3078 ( .A1(r7[3]), .A2(n2854), .B1(n2853), .B2(r4[3]), .ZN(
        n2725) );
  AOI22D0BWP12T U3079 ( .A1(r2[3]), .A2(n2856), .B1(n2855), .B2(r6[3]), .ZN(
        n2724) );
  AOI22D0BWP12T U3080 ( .A1(r5[3]), .A2(n2757), .B1(n2857), .B2(r1[3]), .ZN(
        n2723) );
  AOI22D0BWP12T U3081 ( .A1(r0[3]), .A2(n2859), .B1(n2858), .B2(r3[3]), .ZN(
        n2722) );
  ND4D1BWP12T U3082 ( .A1(n2725), .A2(n2724), .A3(n2723), .A4(n2722), .ZN(
        n2726) );
  MOAI22D0BWP12T U3083 ( .A1(n2822), .A2(n2727), .B1(n2726), .B2(n2864), .ZN(
        n2728) );
  AOI21D0BWP12T U3084 ( .A1(lr[3]), .A2(n2869), .B(n2728), .ZN(n2732) );
  AOI22D0BWP12T U3085 ( .A1(r9[3]), .A2(n2871), .B1(n2870), .B2(r11[3]), .ZN(
        n2731) );
  AOI22D0BWP12T U3086 ( .A1(r8[3]), .A2(n2873), .B1(n2872), .B2(r10[3]), .ZN(
        n2730) );
  AOI22D0BWP12T U3087 ( .A1(r12[3]), .A2(n2848), .B1(n2875), .B2(n[3697]), 
        .ZN(n2729) );
  ND4D1BWP12T U3088 ( .A1(n2732), .A2(n2731), .A3(n2730), .A4(n2729), .ZN(
        regC_out[3]) );
  AOI22D0BWP12T U3089 ( .A1(r8[11]), .A2(n2873), .B1(n2871), .B2(r9[11]), .ZN(
        n2744) );
  AOI22D0BWP12T U3090 ( .A1(lr[11]), .A2(n2869), .B1(n2874), .B2(pc_out[11]), 
        .ZN(n2743) );
  AOI22D0BWP12T U3091 ( .A1(r10[11]), .A2(n2872), .B1(n2870), .B2(r11[11]), 
        .ZN(n2742) );
  AOI22D0BWP12T U3092 ( .A1(r7[11]), .A2(n2854), .B1(n2853), .B2(r4[11]), .ZN(
        n2736) );
  AOI22D0BWP12T U3093 ( .A1(r2[11]), .A2(n2856), .B1(n2855), .B2(r6[11]), .ZN(
        n2735) );
  AOI22D0BWP12T U3094 ( .A1(r5[11]), .A2(n2757), .B1(n2857), .B2(r1[11]), .ZN(
        n2734) );
  AOI22D0BWP12T U3095 ( .A1(r0[11]), .A2(n2859), .B1(n2858), .B2(r3[11]), .ZN(
        n2733) );
  ND4D1BWP12T U3096 ( .A1(n2736), .A2(n2735), .A3(n2734), .A4(n2733), .ZN(
        n2740) );
  OAI22D0BWP12T U3097 ( .A1(n2738), .A2(n2832), .B1(n2867), .B2(n2737), .ZN(
        n2739) );
  AOI21D1BWP12T U3098 ( .A1(n2740), .A2(n2864), .B(n2739), .ZN(n2741) );
  ND4D1BWP12T U3099 ( .A1(n2744), .A2(n2743), .A3(n2742), .A4(n2741), .ZN(
        regC_out[11]) );
  AOI22D0BWP12T U3100 ( .A1(r8[12]), .A2(n2873), .B1(n2871), .B2(r9[12]), .ZN(
        n2756) );
  AOI22D0BWP12T U3101 ( .A1(lr[12]), .A2(n2869), .B1(n2875), .B2(n[3688]), 
        .ZN(n2755) );
  AOI22D0BWP12T U3102 ( .A1(r10[12]), .A2(n2872), .B1(n2870), .B2(r11[12]), 
        .ZN(n2754) );
  AOI22D0BWP12T U3103 ( .A1(r7[12]), .A2(n2854), .B1(n2853), .B2(r4[12]), .ZN(
        n2748) );
  AOI22D0BWP12T U3104 ( .A1(r2[12]), .A2(n2856), .B1(n2855), .B2(r6[12]), .ZN(
        n2747) );
  AOI22D0BWP12T U3105 ( .A1(r5[12]), .A2(n2757), .B1(n2857), .B2(r1[12]), .ZN(
        n2746) );
  AOI22D0BWP12T U3106 ( .A1(r0[12]), .A2(n2859), .B1(n2858), .B2(r3[12]), .ZN(
        n2745) );
  ND4D1BWP12T U3107 ( .A1(n2748), .A2(n2747), .A3(n2746), .A4(n2745), .ZN(
        n2752) );
  OAI22D0BWP12T U3108 ( .A1(n2750), .A2(n2822), .B1(n2867), .B2(n2749), .ZN(
        n2751) );
  AOI21D1BWP12T U3109 ( .A1(n2752), .A2(n2864), .B(n2751), .ZN(n2753) );
  ND4D1BWP12T U3110 ( .A1(n2756), .A2(n2755), .A3(n2754), .A4(n2753), .ZN(
        regC_out[12]) );
  AOI22D0BWP12T U3111 ( .A1(r7[21]), .A2(n2854), .B1(n2853), .B2(r4[21]), .ZN(
        n2761) );
  AOI22D0BWP12T U3112 ( .A1(r2[21]), .A2(n2856), .B1(n2855), .B2(r6[21]), .ZN(
        n2760) );
  AOI22D0BWP12T U3113 ( .A1(r5[21]), .A2(n2757), .B1(n2857), .B2(r1[21]), .ZN(
        n2759) );
  AOI22D0BWP12T U3114 ( .A1(r0[21]), .A2(n2859), .B1(n2858), .B2(r3[21]), .ZN(
        n2758) );
  ND4D1BWP12T U3115 ( .A1(n2761), .A2(n2760), .A3(n2759), .A4(n2758), .ZN(
        n2767) );
  AOI22D0BWP12T U3116 ( .A1(r8[21]), .A2(n2873), .B1(n2871), .B2(r9[21]), .ZN(
        n2765) );
  AOI22D0BWP12T U3117 ( .A1(lr[21]), .A2(n2869), .B1(n2875), .B2(n[3679]), 
        .ZN(n2764) );
  AOI22D0BWP12T U3118 ( .A1(r12[21]), .A2(n2848), .B1(n2874), .B2(pc_out[21]), 
        .ZN(n2763) );
  AOI22D0BWP12T U3119 ( .A1(r10[21]), .A2(n2872), .B1(n2870), .B2(r11[21]), 
        .ZN(n2762) );
  ND4D1BWP12T U3120 ( .A1(n2765), .A2(n2764), .A3(n2763), .A4(n2762), .ZN(
        n2766) );
  AO21D1BWP12T U3121 ( .A1(n2864), .A2(n2767), .B(n2766), .Z(regC_out[21]) );
  AOI22D0BWP12T U3122 ( .A1(pc_out[24]), .A2(n2874), .B1(n2873), .B2(r8[24]), 
        .ZN(n2777) );
  AOI22D0BWP12T U3123 ( .A1(r9[24]), .A2(n2871), .B1(n2870), .B2(r11[24]), 
        .ZN(n2776) );
  AOI22D0BWP12T U3124 ( .A1(r7[24]), .A2(n2854), .B1(n2853), .B2(r4[24]), .ZN(
        n2771) );
  AOI22D0BWP12T U3125 ( .A1(r2[24]), .A2(n2856), .B1(n2855), .B2(r6[24]), .ZN(
        n2770) );
  AOI22D0BWP12T U3126 ( .A1(r5[24]), .A2(n2757), .B1(n2857), .B2(r1[24]), .ZN(
        n2769) );
  AOI22D0BWP12T U3127 ( .A1(r0[24]), .A2(n2859), .B1(n2858), .B2(r3[24]), .ZN(
        n2768) );
  ND4D1BWP12T U3128 ( .A1(n2771), .A2(n2770), .A3(n2769), .A4(n2768), .ZN(
        n2774) );
  INVD1BWP12T U3129 ( .I(r10[24]), .ZN(n3451) );
  OAI22D0BWP12T U3130 ( .A1(n2867), .A2(n3462), .B1(n3451), .B2(n2827), .ZN(
        n2773) );
  OAI22D0BWP12T U3131 ( .A1(n3461), .A2(n2832), .B1(n2846), .B2(n3450), .ZN(
        n2772) );
  AOI211D1BWP12T U3132 ( .A1(n2774), .A2(n2864), .B(n2773), .C(n2772), .ZN(
        n2775) );
  ND3D1BWP12T U3133 ( .A1(n2777), .A2(n2776), .A3(n2775), .ZN(regC_out[24]) );
  AOI22D0BWP12T U3134 ( .A1(r8[6]), .A2(n2873), .B1(n2871), .B2(r9[6]), .ZN(
        n2790) );
  AOI22D0BWP12T U3135 ( .A1(lr[6]), .A2(n2869), .B1(n2874), .B2(pc_out[6]), 
        .ZN(n2789) );
  AOI22D0BWP12T U3136 ( .A1(r10[6]), .A2(n2872), .B1(n2870), .B2(r11[6]), .ZN(
        n2788) );
  AOI22D0BWP12T U3137 ( .A1(r7[6]), .A2(n2854), .B1(n2853), .B2(r4[6]), .ZN(
        n2782) );
  AOI22D0BWP12T U3138 ( .A1(r2[6]), .A2(n2856), .B1(n2855), .B2(r6[6]), .ZN(
        n2781) );
  AOI22D0BWP12T U3139 ( .A1(r5[6]), .A2(n2757), .B1(n2857), .B2(r1[6]), .ZN(
        n2780) );
  AOI22D0BWP12T U3140 ( .A1(r0[6]), .A2(n2859), .B1(n2858), .B2(r3[6]), .ZN(
        n2779) );
  ND4D1BWP12T U3141 ( .A1(n2782), .A2(n2781), .A3(n2780), .A4(n2779), .ZN(
        n2786) );
  OAI22D0BWP12T U3142 ( .A1(n2784), .A2(n2832), .B1(n2867), .B2(n2783), .ZN(
        n2785) );
  AOI21D1BWP12T U3143 ( .A1(n2786), .A2(n2864), .B(n2785), .ZN(n2787) );
  ND4D1BWP12T U3144 ( .A1(n2790), .A2(n2789), .A3(n2788), .A4(n2787), .ZN(
        regC_out[6]) );
  AOI22D0BWP12T U3145 ( .A1(r8[17]), .A2(n2873), .B1(n2872), .B2(r10[17]), 
        .ZN(n2802) );
  AOI22D0BWP12T U3146 ( .A1(r12[17]), .A2(n2848), .B1(n2874), .B2(pc_out[17]), 
        .ZN(n2801) );
  AOI22D0BWP12T U3147 ( .A1(r9[17]), .A2(n2871), .B1(n2870), .B2(r11[17]), 
        .ZN(n2800) );
  AOI22D0BWP12T U3148 ( .A1(r7[17]), .A2(n2854), .B1(n2853), .B2(r4[17]), .ZN(
        n2794) );
  AOI22D0BWP12T U3149 ( .A1(r2[17]), .A2(n2856), .B1(n2855), .B2(r6[17]), .ZN(
        n2793) );
  AOI22D0BWP12T U3150 ( .A1(r5[17]), .A2(n2757), .B1(n2857), .B2(r1[17]), .ZN(
        n2792) );
  AOI22D0BWP12T U3151 ( .A1(r0[17]), .A2(n2859), .B1(n2858), .B2(r3[17]), .ZN(
        n2791) );
  ND4D1BWP12T U3152 ( .A1(n2794), .A2(n2793), .A3(n2792), .A4(n2791), .ZN(
        n2798) );
  OAI22D0BWP12T U3153 ( .A1(n2796), .A2(n2832), .B1(n2846), .B2(n2795), .ZN(
        n2797) );
  AOI21D1BWP12T U3154 ( .A1(n2798), .A2(n2864), .B(n2797), .ZN(n2799) );
  ND4D1BWP12T U3155 ( .A1(n2802), .A2(n2801), .A3(n2800), .A4(n2799), .ZN(
        regC_out[17]) );
  AOI22D0BWP12T U3156 ( .A1(n[3693]), .A2(n2875), .B1(n2874), .B2(pc_out[7]), 
        .ZN(n2816) );
  AOI22D0BWP12T U3157 ( .A1(r9[7]), .A2(n2871), .B1(n2870), .B2(r11[7]), .ZN(
        n2815) );
  AOI22D0BWP12T U3158 ( .A1(r7[7]), .A2(n2854), .B1(n2853), .B2(r4[7]), .ZN(
        n2806) );
  AOI22D0BWP12T U3159 ( .A1(r2[7]), .A2(n2856), .B1(n2855), .B2(r6[7]), .ZN(
        n2805) );
  AOI22D0BWP12T U3160 ( .A1(r5[7]), .A2(n2757), .B1(n2857), .B2(r1[7]), .ZN(
        n2804) );
  AOI22D0BWP12T U3161 ( .A1(r0[7]), .A2(n2859), .B1(n2858), .B2(r3[7]), .ZN(
        n2803) );
  ND4D1BWP12T U3162 ( .A1(n2806), .A2(n2805), .A3(n2804), .A4(n2803), .ZN(
        n2813) );
  OAI22D0BWP12T U3163 ( .A1(n2867), .A2(n2808), .B1(n2807), .B2(n2830), .ZN(
        n2812) );
  OAI22D0BWP12T U3164 ( .A1(n2846), .A2(n2810), .B1(n2809), .B2(n2827), .ZN(
        n2811) );
  AOI211D1BWP12T U3165 ( .A1(n2813), .A2(n2864), .B(n2812), .C(n2811), .ZN(
        n2814) );
  ND3D1BWP12T U3166 ( .A1(n2816), .A2(n2815), .A3(n2814), .ZN(regC_out[7]) );
  AOI22D0BWP12T U3167 ( .A1(r12[14]), .A2(n2848), .B1(n2874), .B2(pc_out[14]), 
        .ZN(n2839) );
  AOI22D0BWP12T U3168 ( .A1(r9[14]), .A2(n2871), .B1(n2870), .B2(r11[14]), 
        .ZN(n2838) );
  AOI22D0BWP12T U3169 ( .A1(r7[14]), .A2(n2854), .B1(n2853), .B2(r4[14]), .ZN(
        n2826) );
  AOI22D0BWP12T U3170 ( .A1(r2[14]), .A2(n2856), .B1(n2855), .B2(r6[14]), .ZN(
        n2825) );
  AOI22D0BWP12T U3171 ( .A1(r5[14]), .A2(n2757), .B1(n2857), .B2(r1[14]), .ZN(
        n2824) );
  AOI22D0BWP12T U3172 ( .A1(r0[14]), .A2(n2859), .B1(n2858), .B2(r3[14]), .ZN(
        n2823) );
  ND4D1BWP12T U3173 ( .A1(n2826), .A2(n2825), .A3(n2824), .A4(n2823), .ZN(
        n2836) );
  OAI22D0BWP12T U3174 ( .A1(n2830), .A2(n2829), .B1(n2828), .B2(n2827), .ZN(
        n2835) );
  OAI22D0BWP12T U3175 ( .A1(n2833), .A2(n2832), .B1(n2846), .B2(n2831), .ZN(
        n2834) );
  AOI211D1BWP12T U3176 ( .A1(n2836), .A2(n2864), .B(n2835), .C(n2834), .ZN(
        n2837) );
  ND3D1BWP12T U3177 ( .A1(n2839), .A2(n2838), .A3(n2837), .ZN(regC_out[14]) );
  AOI22D0BWP12T U3178 ( .A1(r7[13]), .A2(n2854), .B1(n2853), .B2(r4[13]), .ZN(
        n2843) );
  AOI22D0BWP12T U3179 ( .A1(r2[13]), .A2(n2856), .B1(n2855), .B2(r6[13]), .ZN(
        n2842) );
  AOI22D0BWP12T U3180 ( .A1(r5[13]), .A2(n2757), .B1(n2857), .B2(r1[13]), .ZN(
        n2841) );
  AOI22D0BWP12T U3181 ( .A1(r0[13]), .A2(n2859), .B1(n2858), .B2(r3[13]), .ZN(
        n2840) );
  ND4D1BWP12T U3182 ( .A1(n2843), .A2(n2842), .A3(n2841), .A4(n2840), .ZN(
        n2844) );
  MOAI22D0BWP12T U3183 ( .A1(n2846), .A2(n2845), .B1(n2844), .B2(n2864), .ZN(
        n2847) );
  AOI21D0BWP12T U3184 ( .A1(n[3687]), .A2(n2875), .B(n2847), .ZN(n2852) );
  AOI22D0BWP12T U3185 ( .A1(r10[13]), .A2(n2872), .B1(n2870), .B2(r11[13]), 
        .ZN(n2851) );
  AOI22D0BWP12T U3186 ( .A1(r8[13]), .A2(n2873), .B1(n2871), .B2(r9[13]), .ZN(
        n2850) );
  AOI22D0BWP12T U3187 ( .A1(r12[13]), .A2(n2848), .B1(n2874), .B2(pc_out[13]), 
        .ZN(n2849) );
  ND4D1BWP12T U3188 ( .A1(n2852), .A2(n2851), .A3(n2850), .A4(n2849), .ZN(
        regC_out[13]) );
  AOI22D0BWP12T U3189 ( .A1(r7[16]), .A2(n2854), .B1(n2853), .B2(r4[16]), .ZN(
        n2863) );
  AOI22D0BWP12T U3190 ( .A1(r2[16]), .A2(n2856), .B1(n2855), .B2(r6[16]), .ZN(
        n2862) );
  AOI22D0BWP12T U3191 ( .A1(r5[16]), .A2(n2757), .B1(n2857), .B2(r1[16]), .ZN(
        n2861) );
  AOI22D0BWP12T U3192 ( .A1(r0[16]), .A2(n2859), .B1(n2858), .B2(r3[16]), .ZN(
        n2860) );
  ND4D1BWP12T U3193 ( .A1(n2863), .A2(n2862), .A3(n2861), .A4(n2860), .ZN(
        n2865) );
  MOAI22D0BWP12T U3194 ( .A1(n2867), .A2(n2866), .B1(n2865), .B2(n2864), .ZN(
        n2868) );
  AOI21D0BWP12T U3195 ( .A1(lr[16]), .A2(n2869), .B(n2868), .ZN(n2879) );
  AOI22D0BWP12T U3196 ( .A1(r9[16]), .A2(n2871), .B1(n2870), .B2(r11[16]), 
        .ZN(n2878) );
  AOI22D0BWP12T U3197 ( .A1(r8[16]), .A2(n2873), .B1(n2872), .B2(r10[16]), 
        .ZN(n2877) );
  AOI22D0BWP12T U3198 ( .A1(n[3684]), .A2(n2875), .B1(n2874), .B2(pc_out[16]), 
        .ZN(n2876) );
  ND4D1BWP12T U3199 ( .A1(n2879), .A2(n2878), .A3(n2877), .A4(n2876), .ZN(
        regC_out[16]) );
  CKND2D1BWP12T U3200 ( .A1(n41), .A2(n3638), .ZN(n2881) );
  AOI22D0BWP12T U3201 ( .A1(n2882), .A2(n3277), .B1(n3276), .B2(tmp1[2]), .ZN(
        n2880) );
  ND2D1BWP12T U3202 ( .A1(n2881), .A2(n2880), .ZN(n2139) );
  TPND2D0BWP12T U3203 ( .A1(write1_in[4]), .A2(n3626), .ZN(n2884) );
  AOI22D0BWP12T U3204 ( .A1(n2887), .A2(n3307), .B1(n3306), .B2(r11[4]), .ZN(
        n2883) );
  ND2D1BWP12T U3205 ( .A1(n2884), .A2(n2883), .ZN(n2269) );
  TPND2D0BWP12T U3206 ( .A1(write1_in[4]), .A2(n3627), .ZN(n2886) );
  AOI22D0BWP12T U3207 ( .A1(n2887), .A2(n3298), .B1(n3297), .B2(r10[4]), .ZN(
        n2885) );
  ND2D1BWP12T U3208 ( .A1(n2886), .A2(n2885), .ZN(n2301) );
  AOI22D0BWP12T U3209 ( .A1(r8[5]), .A2(n2954), .B1(n2953), .B2(r4[5]), .ZN(
        n2889) );
  AOI22D0BWP12T U3210 ( .A1(n[3695]), .A2(n2956), .B1(n2955), .B2(r10[5]), 
        .ZN(n2888) );
  CKND2D1BWP12T U3211 ( .A1(n2889), .A2(n2888), .ZN(n2899) );
  AOI22D0BWP12T U3212 ( .A1(r7[5]), .A2(n2958), .B1(n2957), .B2(r5[5]), .ZN(
        n2893) );
  AOI22D0BWP12T U3213 ( .A1(lr[5]), .A2(n2960), .B1(n2959), .B2(r9[5]), .ZN(
        n2892) );
  AOI22D0BWP12T U3214 ( .A1(r6[5]), .A2(n2962), .B1(n2961), .B2(r11[5]), .ZN(
        n2891) );
  CKND2D0BWP12T U3215 ( .A1(n2963), .A2(r12[5]), .ZN(n2890) );
  ND4D1BWP12T U3216 ( .A1(n2893), .A2(n2892), .A3(n2891), .A4(n2890), .ZN(
        n2898) );
  AOI22D0BWP12T U3217 ( .A1(r3[5]), .A2(n2965), .B1(n2964), .B2(r2[5]), .ZN(
        n2895) );
  AOI22D0BWP12T U3218 ( .A1(n2967), .A2(r0[5]), .B1(pc_out[5]), .B2(n2966), 
        .ZN(n2894) );
  OAI211D0BWP12T U3219 ( .A1(n2896), .A2(n2968), .B(n2895), .C(n2894), .ZN(
        n2897) );
  OA31D1BWP12T U3220 ( .A1(n2899), .A2(n2898), .A3(n2897), .B(n2970), .Z(
        regD_out[5]) );
  AOI22D0BWP12T U3221 ( .A1(r8[6]), .A2(n2954), .B1(n2953), .B2(r4[6]), .ZN(
        n2902) );
  AOI22D0BWP12T U3222 ( .A1(n[3694]), .A2(n2956), .B1(n2955), .B2(r10[6]), 
        .ZN(n2901) );
  CKND2D1BWP12T U3223 ( .A1(n2902), .A2(n2901), .ZN(n2912) );
  AOI22D0BWP12T U3224 ( .A1(r7[6]), .A2(n2958), .B1(n2957), .B2(r5[6]), .ZN(
        n2906) );
  AOI22D0BWP12T U3225 ( .A1(lr[6]), .A2(n2960), .B1(n2959), .B2(r9[6]), .ZN(
        n2905) );
  AOI22D0BWP12T U3226 ( .A1(r6[6]), .A2(n2962), .B1(n2961), .B2(r11[6]), .ZN(
        n2904) );
  CKND2D0BWP12T U3227 ( .A1(n2963), .A2(r12[6]), .ZN(n2903) );
  ND4D1BWP12T U3228 ( .A1(n2906), .A2(n2905), .A3(n2904), .A4(n2903), .ZN(
        n2911) );
  AOI22D0BWP12T U3229 ( .A1(r3[6]), .A2(n2965), .B1(n2964), .B2(r2[6]), .ZN(
        n2908) );
  AOI22D0BWP12T U3230 ( .A1(n2967), .A2(r0[6]), .B1(pc_out[6]), .B2(n2966), 
        .ZN(n2907) );
  OAI211D0BWP12T U3231 ( .A1(n2909), .A2(n2968), .B(n2908), .C(n2907), .ZN(
        n2910) );
  OA31D1BWP12T U3232 ( .A1(n2912), .A2(n2911), .A3(n2910), .B(n2970), .Z(
        regD_out[6]) );
  TPND2D0BWP12T U3233 ( .A1(n2920), .A2(n3229), .ZN(n2919) );
  INVD0BWP12T U3234 ( .I(n2921), .ZN(n2916) );
  NR2D1BWP12T U3235 ( .A1(n2916), .A2(n2938), .ZN(n2917) );
  RCAOI211D0BWP12T U3236 ( .A1(n3230), .A2(n[3694]), .B(n2917), .C(reset), 
        .ZN(n2918) );
  ND2D1BWP12T U3237 ( .A1(n2919), .A2(n2918), .ZN(spin[6]) );
  AOI22D0BWP12T U3238 ( .A1(n2989), .A2(pc_out[2]), .B1(n3398), .B2(
        next_pc_in[2]), .ZN(n2926) );
  OAI21D1BWP12T U3239 ( .A1(n2927), .A2(n3394), .B(n2926), .ZN(n2171) );
  BUFFXD4BWP12T U3240 ( .I(write1_in[9]), .Z(n2936) );
  TPND2D0BWP12T U3241 ( .A1(n2936), .A2(n3229), .ZN(n2935) );
  CKND0BWP12T U3242 ( .I(n2937), .ZN(n2932) );
  NR2XD0BWP12T U3243 ( .A1(n2932), .A2(n2938), .ZN(n2933) );
  RCAOI211D0BWP12T U3244 ( .A1(n3230), .A2(n[3691]), .B(n2933), .C(reset), 
        .ZN(n2934) );
  ND2D1BWP12T U3245 ( .A1(n2935), .A2(n2934), .ZN(spin[9]) );
  CKND2D1BWP12T U3246 ( .A1(write1_in[10]), .A2(n3229), .ZN(n2942) );
  CKND0BWP12T U3247 ( .I(n2951), .ZN(n2939) );
  NR2XD0BWP12T U3248 ( .A1(n2939), .A2(n2938), .ZN(n2940) );
  RCAOI211D0BWP12T U3249 ( .A1(n3230), .A2(n[3690]), .B(n2940), .C(reset), 
        .ZN(n2941) );
  ND2D1BWP12T U3250 ( .A1(n2942), .A2(n2941), .ZN(spin[10]) );
  CKND2D1BWP12T U3251 ( .A1(write1_in[10]), .A2(n3638), .ZN(n2946) );
  AOI22D0BWP12T U3252 ( .A1(n2951), .A2(n3277), .B1(n3276), .B2(tmp1[10]), 
        .ZN(n2945) );
  ND2D1BWP12T U3253 ( .A1(n2946), .A2(n2945), .ZN(n2147) );
  CKND2D1BWP12T U3254 ( .A1(write1_in[10]), .A2(n3216), .ZN(n2948) );
  AOI22D0BWP12T U3255 ( .A1(n2951), .A2(n3218), .B1(n3217), .B2(r12[10]), .ZN(
        n2947) );
  ND2D1BWP12T U3256 ( .A1(n2948), .A2(n2947), .ZN(n2243) );
  CKND2D1BWP12T U3257 ( .A1(write1_in[10]), .A2(n3234), .ZN(n2950) );
  AOI22D0BWP12T U3258 ( .A1(n2951), .A2(n3236), .B1(n3235), .B2(lr[10]), .ZN(
        n2949) );
  ND2D1BWP12T U3259 ( .A1(n2950), .A2(n2949), .ZN(n2211) );
  CKND2D0BWP12T U3260 ( .A1(write1_in[16]), .A2(n3628), .ZN(n2975) );
  AOI22D0BWP12T U3261 ( .A1(write2_in[16]), .A2(n3263), .B1(n3262), .B2(r6[16]), .ZN(n2974) );
  ND2D1BWP12T U3262 ( .A1(n2975), .A2(n2974), .ZN(n2441) );
  CKND2D0BWP12T U3263 ( .A1(write1_in[18]), .A2(n3622), .ZN(n2977) );
  AOI22D0BWP12T U3264 ( .A1(write2_in[18]), .A2(n3273), .B1(n3272), .B2(r5[18]), .ZN(n2976) );
  ND2D1BWP12T U3265 ( .A1(n2977), .A2(n2976), .ZN(n2475) );
  CKND2D0BWP12T U3266 ( .A1(write1_in[18]), .A2(n3241), .ZN(n2979) );
  AOI22D0BWP12T U3267 ( .A1(write2_in[18]), .A2(n3243), .B1(n3242), .B2(r7[18]), .ZN(n2978) );
  ND2D1BWP12T U3268 ( .A1(n2979), .A2(n2978), .ZN(n2411) );
  CKND2D0BWP12T U3269 ( .A1(write1_in[18]), .A2(n3623), .ZN(n2981) );
  AOI22D0BWP12T U3270 ( .A1(write2_in[18]), .A2(n3281), .B1(n3280), .B2(r4[18]), .ZN(n2980) );
  ND2D1BWP12T U3271 ( .A1(n2981), .A2(n2980), .ZN(n2507) );
  CKND2D0BWP12T U3272 ( .A1(write1_in[18]), .A2(n3628), .ZN(n2983) );
  AOI22D0BWP12T U3273 ( .A1(write2_in[18]), .A2(n3263), .B1(n3262), .B2(r6[18]), .ZN(n2982) );
  ND2D1BWP12T U3274 ( .A1(n2983), .A2(n2982), .ZN(n2443) );
  CKND0BWP12T U3275 ( .I(n2984), .ZN(n2986) );
  ND2D1BWP12T U3276 ( .A1(n2986), .A2(n2985), .ZN(n2988) );
  XNR2D1BWP12T U3277 ( .A1(n2988), .A2(n2987), .ZN(n2991) );
  AOI22D1BWP12T U3278 ( .A1(n2989), .A2(pc_out[9]), .B1(n3398), .B2(
        next_pc_in[9]), .ZN(n2990) );
  OAI21D1BWP12T U3279 ( .A1(n2991), .A2(n3394), .B(n2990), .ZN(n2178) );
  CKND2D0BWP12T U3280 ( .A1(write1_in[19]), .A2(n3241), .ZN(n2993) );
  AOI22D0BWP12T U3281 ( .A1(write2_in[19]), .A2(n3243), .B1(n3242), .B2(r7[19]), .ZN(n2992) );
  ND2D1BWP12T U3282 ( .A1(n2993), .A2(n2992), .ZN(n2412) );
  CKND2D0BWP12T U3283 ( .A1(write1_in[19]), .A2(n3622), .ZN(n2995) );
  AOI22D0BWP12T U3284 ( .A1(write2_in[19]), .A2(n3273), .B1(n3272), .B2(r5[19]), .ZN(n2994) );
  ND2D1BWP12T U3285 ( .A1(n2995), .A2(n2994), .ZN(n2476) );
  CKND2D0BWP12T U3286 ( .A1(write1_in[19]), .A2(n3623), .ZN(n2997) );
  AOI22D0BWP12T U3287 ( .A1(write2_in[19]), .A2(n3281), .B1(n3280), .B2(r4[19]), .ZN(n2996) );
  ND2D1BWP12T U3288 ( .A1(n2997), .A2(n2996), .ZN(n2508) );
  CKND2D0BWP12T U3289 ( .A1(n250), .A2(n3628), .ZN(n2999) );
  AOI22D0BWP12T U3290 ( .A1(write2_in[19]), .A2(n3263), .B1(n3262), .B2(r6[19]), .ZN(n2998) );
  ND2D1BWP12T U3291 ( .A1(n2999), .A2(n2998), .ZN(n2444) );
  CKND2D0BWP12T U3292 ( .A1(write1_in[19]), .A2(n3248), .ZN(n3001) );
  AOI22D0BWP12T U3293 ( .A1(write2_in[19]), .A2(n3250), .B1(n3249), .B2(r9[19]), .ZN(n3000) );
  ND2D1BWP12T U3294 ( .A1(n3001), .A2(n3000), .ZN(n2348) );
  CKND2D0BWP12T U3295 ( .A1(n250), .A2(n3229), .ZN(n3003) );
  AOI22D0BWP12T U3296 ( .A1(write2_in[19]), .A2(n3231), .B1(n3230), .B2(
        n[3681]), .ZN(n3002) );
  ND2D1BWP12T U3297 ( .A1(n3003), .A2(n3002), .ZN(spin[19]) );
  CKND2D0BWP12T U3298 ( .A1(n250), .A2(n3625), .ZN(n3005) );
  AOI22D0BWP12T U3299 ( .A1(write2_in[19]), .A2(n3374), .B1(n3373), .B2(r2[19]), .ZN(n3004) );
  ND2D1BWP12T U3300 ( .A1(n3005), .A2(n3004), .ZN(n2572) );
  CKND2D0BWP12T U3301 ( .A1(n250), .A2(n3624), .ZN(n3007) );
  AOI22D0BWP12T U3302 ( .A1(write2_in[19]), .A2(n3028), .B1(n3303), .B2(r3[19]), .ZN(n3006) );
  ND2D1BWP12T U3303 ( .A1(n3007), .A2(n3006), .ZN(n2540) );
  CKND2D0BWP12T U3304 ( .A1(n250), .A2(n3626), .ZN(n3009) );
  AOI22D0BWP12T U3305 ( .A1(write2_in[19]), .A2(n3307), .B1(n3306), .B2(
        r11[19]), .ZN(n3008) );
  ND2D1BWP12T U3306 ( .A1(n3009), .A2(n3008), .ZN(n2284) );
  CKND2D0BWP12T U3307 ( .A1(n250), .A2(n3627), .ZN(n3011) );
  AOI22D0BWP12T U3308 ( .A1(write2_in[19]), .A2(n3298), .B1(n3297), .B2(
        r10[19]), .ZN(n3010) );
  ND2D1BWP12T U3309 ( .A1(n3011), .A2(n3010), .ZN(n2316) );
  CKND2D0BWP12T U3310 ( .A1(write1_in[21]), .A2(n3241), .ZN(n3013) );
  AOI22D0BWP12T U3311 ( .A1(write2_in[21]), .A2(n3243), .B1(n3242), .B2(r7[21]), .ZN(n3012) );
  ND2D1BWP12T U3312 ( .A1(n3013), .A2(n3012), .ZN(n2414) );
  CKND2D0BWP12T U3313 ( .A1(write1_in[21]), .A2(n3622), .ZN(n3015) );
  AOI22D0BWP12T U3314 ( .A1(write2_in[21]), .A2(n3273), .B1(n3272), .B2(r5[21]), .ZN(n3014) );
  ND2D1BWP12T U3315 ( .A1(n3015), .A2(n3014), .ZN(n2478) );
  CKND2D0BWP12T U3316 ( .A1(write1_in[21]), .A2(n3623), .ZN(n3017) );
  AOI22D0BWP12T U3317 ( .A1(write2_in[21]), .A2(n3281), .B1(n3280), .B2(r4[21]), .ZN(n3016) );
  ND2D1BWP12T U3318 ( .A1(n3017), .A2(n3016), .ZN(n2510) );
  CKND2D0BWP12T U3319 ( .A1(write1_in[21]), .A2(n3628), .ZN(n3019) );
  AOI22D0BWP12T U3320 ( .A1(write2_in[21]), .A2(n3263), .B1(n3262), .B2(r6[21]), .ZN(n3018) );
  ND2D1BWP12T U3321 ( .A1(n3019), .A2(n3018), .ZN(n2446) );
  CKND2D0BWP12T U3322 ( .A1(write1_in[21]), .A2(n3248), .ZN(n3021) );
  AOI22D0BWP12T U3323 ( .A1(write2_in[21]), .A2(n3250), .B1(n3249), .B2(r9[21]), .ZN(n3020) );
  ND2D1BWP12T U3324 ( .A1(n3021), .A2(n3020), .ZN(n2350) );
  CKND2D0BWP12T U3325 ( .A1(write1_in[21]), .A2(n3229), .ZN(n3023) );
  AOI22D0BWP12T U3326 ( .A1(write2_in[21]), .A2(n3231), .B1(n3230), .B2(
        n[3679]), .ZN(n3022) );
  ND2D1BWP12T U3327 ( .A1(n3023), .A2(n3022), .ZN(spin[21]) );
  CKND2D0BWP12T U3328 ( .A1(write1_in[21]), .A2(n3627), .ZN(n3025) );
  AOI22D0BWP12T U3329 ( .A1(write2_in[21]), .A2(n3298), .B1(n3297), .B2(
        r10[21]), .ZN(n3024) );
  ND2D1BWP12T U3330 ( .A1(n3025), .A2(n3024), .ZN(n2318) );
  CKND2D0BWP12T U3331 ( .A1(write1_in[21]), .A2(n3625), .ZN(n3027) );
  AOI22D0BWP12T U3332 ( .A1(write2_in[21]), .A2(n3374), .B1(n3373), .B2(r2[21]), .ZN(n3026) );
  ND2D1BWP12T U3333 ( .A1(n3027), .A2(n3026), .ZN(n2574) );
  CKND2D0BWP12T U3334 ( .A1(write1_in[21]), .A2(n3624), .ZN(n3030) );
  AOI22D0BWP12T U3335 ( .A1(write2_in[21]), .A2(n3028), .B1(n3303), .B2(r3[21]), .ZN(n3029) );
  ND2D1BWP12T U3336 ( .A1(n3030), .A2(n3029), .ZN(n2542) );
  CKND2D0BWP12T U3337 ( .A1(write1_in[21]), .A2(n3626), .ZN(n3032) );
  AOI22D0BWP12T U3338 ( .A1(write2_in[21]), .A2(n3307), .B1(n3306), .B2(
        r11[21]), .ZN(n3031) );
  ND2D1BWP12T U3339 ( .A1(n3032), .A2(n3031), .ZN(n2286) );
  TPND2D0BWP12T U3340 ( .A1(n3051), .A2(n3623), .ZN(n3034) );
  AOI22D0BWP12T U3341 ( .A1(write2_in[20]), .A2(n3281), .B1(n3280), .B2(r4[20]), .ZN(n3033) );
  ND2D1BWP12T U3342 ( .A1(n3034), .A2(n3033), .ZN(n2509) );
  TPND2D0BWP12T U3343 ( .A1(n3051), .A2(n3229), .ZN(n3036) );
  AOI22D0BWP12T U3344 ( .A1(write2_in[20]), .A2(n3231), .B1(n3230), .B2(
        n[3680]), .ZN(n3035) );
  ND2D1BWP12T U3345 ( .A1(n3036), .A2(n3035), .ZN(spin[20]) );
  TPND2D0BWP12T U3346 ( .A1(n3051), .A2(n3241), .ZN(n3038) );
  AOI22D0BWP12T U3347 ( .A1(write2_in[20]), .A2(n3243), .B1(n3242), .B2(r7[20]), .ZN(n3037) );
  ND2D1BWP12T U3348 ( .A1(n3038), .A2(n3037), .ZN(n2413) );
  TPND2D0BWP12T U3349 ( .A1(n3051), .A2(n3628), .ZN(n3040) );
  AOI22D0BWP12T U3350 ( .A1(write2_in[20]), .A2(n3263), .B1(n3262), .B2(r6[20]), .ZN(n3039) );
  ND2D1BWP12T U3351 ( .A1(n3040), .A2(n3039), .ZN(n2445) );
  TPND2D0BWP12T U3352 ( .A1(n3051), .A2(n3627), .ZN(n3042) );
  AOI22D0BWP12T U3353 ( .A1(write2_in[20]), .A2(n3298), .B1(n3297), .B2(
        r10[20]), .ZN(n3041) );
  ND2D1BWP12T U3354 ( .A1(n3042), .A2(n3041), .ZN(n2317) );
  TPND2D0BWP12T U3355 ( .A1(n3051), .A2(n3624), .ZN(n3044) );
  AOI22D0BWP12T U3356 ( .A1(write2_in[20]), .A2(n3028), .B1(n3303), .B2(r3[20]), .ZN(n3043) );
  ND2D1BWP12T U3357 ( .A1(n3044), .A2(n3043), .ZN(n2541) );
  TPND2D0BWP12T U3358 ( .A1(n3051), .A2(n3622), .ZN(n3046) );
  AOI22D0BWP12T U3359 ( .A1(write2_in[20]), .A2(n3273), .B1(n3272), .B2(r5[20]), .ZN(n3045) );
  ND2D1BWP12T U3360 ( .A1(n3046), .A2(n3045), .ZN(n2477) );
  TPND2D0BWP12T U3361 ( .A1(n3051), .A2(n3248), .ZN(n3048) );
  AOI22D0BWP12T U3362 ( .A1(write2_in[20]), .A2(n3250), .B1(n3249), .B2(r9[20]), .ZN(n3047) );
  ND2D1BWP12T U3363 ( .A1(n3048), .A2(n3047), .ZN(n2349) );
  TPND2D0BWP12T U3364 ( .A1(n3051), .A2(n3626), .ZN(n3050) );
  AOI22D0BWP12T U3365 ( .A1(write2_in[20]), .A2(n3307), .B1(n3306), .B2(
        r11[20]), .ZN(n3049) );
  ND2D1BWP12T U3366 ( .A1(n3050), .A2(n3049), .ZN(n2285) );
  TPND2D0BWP12T U3367 ( .A1(n3051), .A2(n3625), .ZN(n3053) );
  AOI22D0BWP12T U3368 ( .A1(write2_in[20]), .A2(n3374), .B1(n3373), .B2(r2[20]), .ZN(n3052) );
  ND2D1BWP12T U3369 ( .A1(n3053), .A2(n3052), .ZN(n2573) );
  CKND2D0BWP12T U3370 ( .A1(write1_in[22]), .A2(n3216), .ZN(n3055) );
  AOI22D0BWP12T U3371 ( .A1(write2_in[22]), .A2(n3218), .B1(n3217), .B2(
        r12[22]), .ZN(n3054) );
  ND2D1BWP12T U3372 ( .A1(n3055), .A2(n3054), .ZN(n2255) );
  CKND2D0BWP12T U3373 ( .A1(write1_in[22]), .A2(n3638), .ZN(n3057) );
  AOI22D0BWP12T U3374 ( .A1(write2_in[22]), .A2(n3277), .B1(n3276), .B2(
        tmp1[22]), .ZN(n3056) );
  ND2D1BWP12T U3375 ( .A1(n3057), .A2(n3056), .ZN(n2159) );
  CKND2D0BWP12T U3376 ( .A1(write1_in[22]), .A2(n3211), .ZN(n3059) );
  AOI22D0BWP12T U3377 ( .A1(write2_in[22]), .A2(n3213), .B1(n3212), .B2(r8[22]), .ZN(n3058) );
  ND2D1BWP12T U3378 ( .A1(n3059), .A2(n3058), .ZN(n2383) );
  CKND2D0BWP12T U3379 ( .A1(write1_in[22]), .A2(n3234), .ZN(n3061) );
  AOI22D0BWP12T U3380 ( .A1(write2_in[22]), .A2(n3236), .B1(n3235), .B2(lr[22]), .ZN(n3060) );
  ND2D1BWP12T U3381 ( .A1(n3061), .A2(n3060), .ZN(n2223) );
  ND2D1BWP12T U3382 ( .A1(write1_in[24]), .A2(n3229), .ZN(n3063) );
  AOI22D0BWP12T U3383 ( .A1(write2_in[24]), .A2(n3231), .B1(n3230), .B2(
        n[3676]), .ZN(n3062) );
  ND2D1BWP12T U3384 ( .A1(n3063), .A2(n3062), .ZN(spin[24]) );
  ND2D1BWP12T U3385 ( .A1(write1_in[24]), .A2(n3211), .ZN(n3065) );
  AOI22D0BWP12T U3386 ( .A1(write2_in[24]), .A2(n3213), .B1(n3212), .B2(r8[24]), .ZN(n3064) );
  ND2D1BWP12T U3387 ( .A1(n3065), .A2(n3064), .ZN(n2385) );
  ND2D1BWP12T U3388 ( .A1(write1_in[24]), .A2(n3216), .ZN(n3067) );
  AOI22D0BWP12T U3389 ( .A1(write2_in[24]), .A2(n3218), .B1(n3217), .B2(
        r12[24]), .ZN(n3066) );
  ND2D1BWP12T U3390 ( .A1(n3067), .A2(n3066), .ZN(n2257) );
  ND2D1BWP12T U3391 ( .A1(write1_in[24]), .A2(n3623), .ZN(n3069) );
  AOI22D0BWP12T U3392 ( .A1(write2_in[24]), .A2(n3281), .B1(n3280), .B2(r4[24]), .ZN(n3068) );
  ND2D1BWP12T U3393 ( .A1(n3069), .A2(n3068), .ZN(n2513) );
  ND2D1BWP12T U3394 ( .A1(write1_in[24]), .A2(n3622), .ZN(n3071) );
  AOI22D0BWP12T U3395 ( .A1(write2_in[24]), .A2(n3273), .B1(n3272), .B2(r5[24]), .ZN(n3070) );
  ND2D1BWP12T U3396 ( .A1(n3071), .A2(n3070), .ZN(n2481) );
  ND2D1BWP12T U3397 ( .A1(write1_in[24]), .A2(n3234), .ZN(n3073) );
  AOI22D0BWP12T U3398 ( .A1(write2_in[24]), .A2(n3236), .B1(n3235), .B2(lr[24]), .ZN(n3072) );
  ND2D1BWP12T U3399 ( .A1(n3073), .A2(n3072), .ZN(n2225) );
  ND2D1BWP12T U3400 ( .A1(write1_in[24]), .A2(n3638), .ZN(n3075) );
  AOI22D0BWP12T U3401 ( .A1(write2_in[24]), .A2(n3277), .B1(n3276), .B2(
        tmp1[24]), .ZN(n3074) );
  ND2D1BWP12T U3402 ( .A1(n3075), .A2(n3074), .ZN(n2161) );
  ND2D1BWP12T U3403 ( .A1(write1_in[24]), .A2(n3241), .ZN(n3077) );
  AOI22D0BWP12T U3404 ( .A1(write2_in[24]), .A2(n3243), .B1(n3242), .B2(r7[24]), .ZN(n3076) );
  ND2D1BWP12T U3405 ( .A1(n3077), .A2(n3076), .ZN(n2417) );
  ND2D1BWP12T U3406 ( .A1(write1_in[24]), .A2(n3248), .ZN(n3079) );
  AOI22D0BWP12T U3407 ( .A1(write2_in[24]), .A2(n3250), .B1(n3249), .B2(r9[24]), .ZN(n3078) );
  ND2D1BWP12T U3408 ( .A1(n3079), .A2(n3078), .ZN(n2353) );
  ND2D1BWP12T U3409 ( .A1(write1_in[24]), .A2(n3628), .ZN(n3081) );
  AOI22D0BWP12T U3410 ( .A1(write2_in[24]), .A2(n3263), .B1(n3262), .B2(r6[24]), .ZN(n3080) );
  ND2D1BWP12T U3411 ( .A1(n3081), .A2(n3080), .ZN(n2449) );
  ND2D1BWP12T U3412 ( .A1(write1_in[24]), .A2(n3625), .ZN(n3083) );
  AOI22D0BWP12T U3413 ( .A1(write2_in[24]), .A2(n3374), .B1(n3373), .B2(r2[24]), .ZN(n3082) );
  ND2D1BWP12T U3414 ( .A1(n3083), .A2(n3082), .ZN(n2577) );
  ND2D1BWP12T U3415 ( .A1(write1_in[24]), .A2(n3624), .ZN(n3085) );
  AOI22D0BWP12T U3416 ( .A1(write2_in[24]), .A2(n3028), .B1(n3303), .B2(r3[24]), .ZN(n3084) );
  ND2D1BWP12T U3417 ( .A1(n3085), .A2(n3084), .ZN(n2545) );
  ND2D1BWP12T U3418 ( .A1(write1_in[24]), .A2(n3627), .ZN(n3087) );
  AOI22D0BWP12T U3419 ( .A1(write2_in[24]), .A2(n3298), .B1(n3297), .B2(
        r10[24]), .ZN(n3086) );
  ND2D1BWP12T U3420 ( .A1(n3087), .A2(n3086), .ZN(n2321) );
  ND2D1BWP12T U3421 ( .A1(write1_in[24]), .A2(n3626), .ZN(n3089) );
  AOI22D0BWP12T U3422 ( .A1(write2_in[24]), .A2(n3307), .B1(n3306), .B2(
        r11[24]), .ZN(n3088) );
  ND2D1BWP12T U3423 ( .A1(n3089), .A2(n3088), .ZN(n2289) );
  BUFFXD4BWP12T U3424 ( .I(write1_in[23]), .Z(n3124) );
  CKND2D1BWP12T U3425 ( .A1(n3124), .A2(n3234), .ZN(n3091) );
  AOI22D0BWP12T U3426 ( .A1(write2_in[23]), .A2(n3236), .B1(n3235), .B2(lr[23]), .ZN(n3090) );
  ND2D1BWP12T U3427 ( .A1(n3091), .A2(n3090), .ZN(n2224) );
  CKND2D1BWP12T U3428 ( .A1(n3124), .A2(n3216), .ZN(n3093) );
  AOI22D0BWP12T U3429 ( .A1(write2_in[23]), .A2(n3218), .B1(n3217), .B2(
        r12[23]), .ZN(n3092) );
  ND2D1BWP12T U3430 ( .A1(n3093), .A2(n3092), .ZN(n2256) );
  CKND2D1BWP12T U3431 ( .A1(n3124), .A2(n3638), .ZN(n3095) );
  AOI22D0BWP12T U3432 ( .A1(write2_in[23]), .A2(n3277), .B1(n3276), .B2(
        tmp1[23]), .ZN(n3094) );
  ND2D1BWP12T U3433 ( .A1(n3095), .A2(n3094), .ZN(n2160) );
  CKND2D1BWP12T U3434 ( .A1(n3124), .A2(n3229), .ZN(n3097) );
  AOI22D0BWP12T U3435 ( .A1(write2_in[23]), .A2(n3231), .B1(n3230), .B2(
        n[3677]), .ZN(n3096) );
  ND2D1BWP12T U3436 ( .A1(n3097), .A2(n3096), .ZN(spin[23]) );
  CKND2D1BWP12T U3437 ( .A1(n3124), .A2(n3627), .ZN(n3099) );
  AOI22D0BWP12T U3438 ( .A1(write2_in[23]), .A2(n3298), .B1(n3297), .B2(
        r10[23]), .ZN(n3098) );
  ND2D1BWP12T U3439 ( .A1(n3099), .A2(n3098), .ZN(n2320) );
  CKND2D1BWP12T U3440 ( .A1(n3124), .A2(n3622), .ZN(n3101) );
  AOI22D0BWP12T U3441 ( .A1(write2_in[23]), .A2(n3273), .B1(n3272), .B2(r5[23]), .ZN(n3100) );
  ND2D1BWP12T U3442 ( .A1(n3101), .A2(n3100), .ZN(n2480) );
  CKND2D1BWP12T U3443 ( .A1(n3124), .A2(n3241), .ZN(n3103) );
  AOI22D0BWP12T U3444 ( .A1(write2_in[23]), .A2(n3243), .B1(n3242), .B2(r7[23]), .ZN(n3102) );
  ND2D1BWP12T U3445 ( .A1(n3103), .A2(n3102), .ZN(n2416) );
  CKND2D1BWP12T U3446 ( .A1(n3124), .A2(n3211), .ZN(n3105) );
  AOI22D0BWP12T U3447 ( .A1(write2_in[23]), .A2(n3213), .B1(n3212), .B2(r8[23]), .ZN(n3104) );
  ND2D1BWP12T U3448 ( .A1(n3105), .A2(n3104), .ZN(n2384) );
  CKND2D1BWP12T U3449 ( .A1(n3124), .A2(n3289), .ZN(n3107) );
  AOI22D0BWP12T U3450 ( .A1(write2_in[23]), .A2(n3291), .B1(n3290), .B2(r1[23]), .ZN(n3106) );
  ND2D1BWP12T U3451 ( .A1(n3107), .A2(n3106), .ZN(n2608) );
  CKND2D1BWP12T U3452 ( .A1(n3124), .A2(n3284), .ZN(n3109) );
  AOI22D0BWP12T U3453 ( .A1(write2_in[23]), .A2(n3286), .B1(n3285), .B2(r0[23]), .ZN(n3108) );
  ND2D1BWP12T U3454 ( .A1(n3109), .A2(n3108), .ZN(n2640) );
  CKND2D1BWP12T U3455 ( .A1(n3124), .A2(n3623), .ZN(n3111) );
  AOI22D0BWP12T U3456 ( .A1(write2_in[23]), .A2(n3281), .B1(n3280), .B2(r4[23]), .ZN(n3110) );
  ND2D1BWP12T U3457 ( .A1(n3111), .A2(n3110), .ZN(n2512) );
  CKND2D1BWP12T U3458 ( .A1(n3124), .A2(n3248), .ZN(n3113) );
  AOI22D0BWP12T U3459 ( .A1(write2_in[23]), .A2(n3250), .B1(n3249), .B2(r9[23]), .ZN(n3112) );
  ND2D1BWP12T U3460 ( .A1(n3113), .A2(n3112), .ZN(n2352) );
  CKND2D1BWP12T U3461 ( .A1(n3124), .A2(n3628), .ZN(n3115) );
  AOI22D0BWP12T U3462 ( .A1(write2_in[23]), .A2(n3263), .B1(n3262), .B2(r6[23]), .ZN(n3114) );
  ND2D1BWP12T U3463 ( .A1(n3115), .A2(n3114), .ZN(n2448) );
  BUFFD3BWP12T U3464 ( .I(write1_in[27]), .Z(n3175) );
  AOI22D0BWP12T U3465 ( .A1(write2_in[27]), .A2(n3231), .B1(n3230), .B2(
        n[3673]), .ZN(n3116) );
  CKND2D1BWP12T U3466 ( .A1(n3124), .A2(n3624), .ZN(n3119) );
  AOI22D0BWP12T U3467 ( .A1(write2_in[23]), .A2(n3028), .B1(n3303), .B2(r3[23]), .ZN(n3118) );
  ND2D1BWP12T U3468 ( .A1(n3119), .A2(n3118), .ZN(n2544) );
  CKND2D1BWP12T U3469 ( .A1(n3124), .A2(n3625), .ZN(n3121) );
  AOI22D0BWP12T U3470 ( .A1(write2_in[23]), .A2(n3374), .B1(n3373), .B2(r2[23]), .ZN(n3120) );
  ND2D1BWP12T U3471 ( .A1(n3121), .A2(n3120), .ZN(n2576) );
  AOI22D0BWP12T U3472 ( .A1(write2_in[27]), .A2(n3213), .B1(n3212), .B2(r8[27]), .ZN(n3122) );
  CKND2D1BWP12T U3473 ( .A1(n3124), .A2(n3626), .ZN(n3126) );
  AOI22D0BWP12T U3474 ( .A1(write2_in[23]), .A2(n3307), .B1(n3306), .B2(
        r11[23]), .ZN(n3125) );
  ND2D1BWP12T U3475 ( .A1(n3126), .A2(n3125), .ZN(n2288) );
  AOI22D0BWP12T U3476 ( .A1(write2_in[27]), .A2(n3218), .B1(n3217), .B2(
        r12[27]), .ZN(n3127) );
  AOI22D0BWP12T U3477 ( .A1(write2_in[27]), .A2(n3291), .B1(n3290), .B2(r1[27]), .ZN(n3129) );
  AOI22D0BWP12T U3478 ( .A1(write2_in[27]), .A2(n3286), .B1(n3285), .B2(r0[27]), .ZN(n3131) );
  AOI22D0BWP12T U3479 ( .A1(write2_in[27]), .A2(n3281), .B1(n3280), .B2(r4[27]), .ZN(n3133) );
  AOI22D0BWP12T U3480 ( .A1(write2_in[27]), .A2(n3273), .B1(n3272), .B2(r5[27]), .ZN(n3135) );
  AOI22D0BWP12T U3481 ( .A1(write2_in[27]), .A2(n3277), .B1(n3276), .B2(
        tmp1[27]), .ZN(n3137) );
  AOI22D0BWP12T U3482 ( .A1(write2_in[27]), .A2(n3236), .B1(n3235), .B2(lr[27]), .ZN(n3139) );
  AOI22D0BWP12T U3483 ( .A1(write2_in[27]), .A2(n3243), .B1(n3242), .B2(r7[27]), .ZN(n3141) );
  AOI22D0BWP12T U3484 ( .A1(write2_in[27]), .A2(n3250), .B1(n3249), .B2(r9[27]), .ZN(n3143) );
  AOI22D0BWP12T U3485 ( .A1(write2_in[25]), .A2(n3213), .B1(n3212), .B2(r8[25]), .ZN(n3145) );
  AOI22D0BWP12T U3486 ( .A1(write2_in[25]), .A2(n3218), .B1(n3217), .B2(
        r12[25]), .ZN(n3147) );
  ND2D1BWP12T U3487 ( .A1(n3148), .A2(n3147), .ZN(n2258) );
  AOI22D0BWP12T U3488 ( .A1(write2_in[25]), .A2(n3291), .B1(n3290), .B2(r1[25]), .ZN(n3149) );
  AOI22D0BWP12T U3489 ( .A1(write2_in[25]), .A2(n3281), .B1(n3280), .B2(r4[25]), .ZN(n3151) );
  ND2D1BWP12T U3490 ( .A1(n3152), .A2(n3151), .ZN(n2514) );
  AOI22D0BWP12T U3491 ( .A1(write2_in[25]), .A2(n3286), .B1(n3285), .B2(r0[25]), .ZN(n3153) );
  ND2D1BWP12T U3492 ( .A1(n3154), .A2(n3153), .ZN(n2642) );
  AOI22D0BWP12T U3493 ( .A1(write2_in[25]), .A2(n3273), .B1(n3272), .B2(r5[25]), .ZN(n3155) );
  ND2D1BWP12T U3494 ( .A1(n3156), .A2(n3155), .ZN(n2482) );
  AOI22D0BWP12T U3495 ( .A1(write2_in[25]), .A2(n3231), .B1(n3230), .B2(
        n[3675]), .ZN(n3157) );
  ND2D1BWP12T U3496 ( .A1(n3158), .A2(n3157), .ZN(spin[25]) );
  AOI22D0BWP12T U3497 ( .A1(write2_in[25]), .A2(n3277), .B1(n3276), .B2(
        tmp1[25]), .ZN(n3159) );
  AOI22D0BWP12T U3498 ( .A1(write2_in[25]), .A2(n3236), .B1(n3235), .B2(lr[25]), .ZN(n3161) );
  ND2D1BWP12T U3499 ( .A1(write1_in[25]), .A2(n3241), .ZN(n3164) );
  AOI22D0BWP12T U3500 ( .A1(write2_in[25]), .A2(n3243), .B1(n3242), .B2(r7[25]), .ZN(n3163) );
  ND2D1BWP12T U3501 ( .A1(n3164), .A2(n3163), .ZN(n2418) );
  AOI22D0BWP12T U3502 ( .A1(write2_in[27]), .A2(n3263), .B1(n3262), .B2(r6[27]), .ZN(n3165) );
  AOI22D0BWP12T U3503 ( .A1(write2_in[27]), .A2(n3307), .B1(n3306), .B2(
        r11[27]), .ZN(n3167) );
  AOI22D0BWP12T U3504 ( .A1(write2_in[27]), .A2(n3028), .B1(n3303), .B2(r3[27]), .ZN(n3169) );
  AOI22D0BWP12T U3505 ( .A1(write2_in[27]), .A2(n3374), .B1(n3373), .B2(r2[27]), .ZN(n3171) );
  AOI22D0BWP12T U3506 ( .A1(write2_in[25]), .A2(n3250), .B1(n3249), .B2(r9[25]), .ZN(n3173) );
  ND2D1BWP12T U3507 ( .A1(n3174), .A2(n3173), .ZN(n2354) );
  AOI22D0BWP12T U3508 ( .A1(write2_in[27]), .A2(n3298), .B1(n3297), .B2(
        r10[27]), .ZN(n3176) );
  ND2D1BWP12T U3509 ( .A1(write1_in[25]), .A2(n3628), .ZN(n3179) );
  AOI22D0BWP12T U3510 ( .A1(write2_in[25]), .A2(n3263), .B1(n3262), .B2(r6[25]), .ZN(n3178) );
  ND2D1BWP12T U3511 ( .A1(n3179), .A2(n3178), .ZN(n2450) );
  ND2D1BWP12T U3512 ( .A1(write1_in[25]), .A2(n3627), .ZN(n3181) );
  AOI22D0BWP12T U3513 ( .A1(write2_in[25]), .A2(n3298), .B1(n3297), .B2(
        r10[25]), .ZN(n3180) );
  ND2D1BWP12T U3514 ( .A1(n3181), .A2(n3180), .ZN(n2322) );
  ND2D1BWP12T U3515 ( .A1(write1_in[25]), .A2(n3625), .ZN(n3183) );
  AOI22D0BWP12T U3516 ( .A1(write2_in[25]), .A2(n3374), .B1(n3373), .B2(r2[25]), .ZN(n3182) );
  ND2D1BWP12T U3517 ( .A1(n3183), .A2(n3182), .ZN(n2578) );
  AOI22D0BWP12T U3518 ( .A1(write2_in[25]), .A2(n3028), .B1(n3303), .B2(r3[25]), .ZN(n3185) );
  ND2D1BWP12T U3519 ( .A1(n3186), .A2(n3185), .ZN(n2546) );
  ND2D1BWP12T U3520 ( .A1(write1_in[25]), .A2(n3626), .ZN(n3188) );
  AOI22D0BWP12T U3521 ( .A1(write2_in[25]), .A2(n3307), .B1(n3306), .B2(
        r11[25]), .ZN(n3187) );
  ND2D1BWP12T U3522 ( .A1(n3188), .A2(n3187), .ZN(n2290) );
  TPND2D1BWP12T U3523 ( .A1(n3259), .A2(n3211), .ZN(n3190) );
  AOI22D0BWP12T U3524 ( .A1(write2_in[31]), .A2(n3213), .B1(n3212), .B2(r8[31]), .ZN(n3189) );
  ND2D1BWP12T U3525 ( .A1(n3190), .A2(n3189), .ZN(n2392) );
  TPND2D1BWP12T U3526 ( .A1(n3259), .A2(n3216), .ZN(n3192) );
  AOI22D0BWP12T U3527 ( .A1(write2_in[31]), .A2(n3218), .B1(n3217), .B2(
        r12[31]), .ZN(n3191) );
  ND2D1BWP12T U3528 ( .A1(n3192), .A2(n3191), .ZN(n2264) );
  TPND2D1BWP12T U3529 ( .A1(n3259), .A2(n3623), .ZN(n3194) );
  AOI22D0BWP12T U3530 ( .A1(write2_in[31]), .A2(n3281), .B1(n3280), .B2(r4[31]), .ZN(n3193) );
  ND2D1BWP12T U3531 ( .A1(n3194), .A2(n3193), .ZN(n2520) );
  TPND2D1BWP12T U3532 ( .A1(n3259), .A2(n3284), .ZN(n3196) );
  AOI22D0BWP12T U3533 ( .A1(write2_in[31]), .A2(n3286), .B1(n3285), .B2(r0[31]), .ZN(n3195) );
  ND2D1BWP12T U3534 ( .A1(n3196), .A2(n3195), .ZN(n2648) );
  TPND2D1BWP12T U3535 ( .A1(n3259), .A2(n3622), .ZN(n3198) );
  AOI22D0BWP12T U3536 ( .A1(write2_in[31]), .A2(n3273), .B1(n3272), .B2(r5[31]), .ZN(n3197) );
  ND2D1BWP12T U3537 ( .A1(n3198), .A2(n3197), .ZN(n2488) );
  TPND2D1BWP12T U3538 ( .A1(n3259), .A2(n3289), .ZN(n3200) );
  AOI22D0BWP12T U3539 ( .A1(write2_in[31]), .A2(n3291), .B1(n3290), .B2(r1[31]), .ZN(n3199) );
  ND2D1BWP12T U3540 ( .A1(n3200), .A2(n3199), .ZN(n2616) );
  CKND2D1BWP12T U3541 ( .A1(n3259), .A2(n3229), .ZN(n3202) );
  AOI22D0BWP12T U3542 ( .A1(write2_in[31]), .A2(n3231), .B1(n3230), .B2(
        n[3669]), .ZN(n3201) );
  TPND2D1BWP12T U3543 ( .A1(n3259), .A2(n3234), .ZN(n3204) );
  AOI22D0BWP12T U3544 ( .A1(write2_in[31]), .A2(n3236), .B1(n3235), .B2(lr[31]), .ZN(n3203) );
  ND2D1BWP12T U3545 ( .A1(n3204), .A2(n3203), .ZN(n2232) );
  TPND2D1BWP12T U3546 ( .A1(n3259), .A2(n3638), .ZN(n3206) );
  AOI22D0BWP12T U3547 ( .A1(write2_in[31]), .A2(n3277), .B1(n3276), .B2(
        tmp1[31]), .ZN(n3205) );
  ND2D1BWP12T U3548 ( .A1(n3206), .A2(n3205), .ZN(n2168) );
  AOI22D0BWP12T U3549 ( .A1(write2_in[31]), .A2(n3243), .B1(n3242), .B2(r7[31]), .ZN(n3207) );
  ND2D1BWP12T U3550 ( .A1(n3259), .A2(n3248), .ZN(n3210) );
  AOI22D0BWP12T U3551 ( .A1(write2_in[31]), .A2(n3250), .B1(n3249), .B2(r9[31]), .ZN(n3209) );
  TPND2D1BWP12T U3552 ( .A1(n3294), .A2(n3211), .ZN(n3215) );
  AOI22D0BWP12T U3553 ( .A1(write2_in[28]), .A2(n3213), .B1(r8[28]), .B2(n3212), .ZN(n3214) );
  ND2D1BWP12T U3554 ( .A1(n3215), .A2(n3214), .ZN(n2389) );
  TPND2D1BWP12T U3555 ( .A1(n3294), .A2(n3216), .ZN(n3220) );
  AOI22D0BWP12T U3556 ( .A1(write2_in[28]), .A2(n3218), .B1(r12[28]), .B2(
        n3217), .ZN(n3219) );
  ND2D1BWP12T U3557 ( .A1(n3220), .A2(n3219), .ZN(n2261) );
  TPND2D1BWP12T U3558 ( .A1(n3294), .A2(n3622), .ZN(n3222) );
  AOI22D0BWP12T U3559 ( .A1(write2_in[28]), .A2(n3273), .B1(r5[28]), .B2(n3272), .ZN(n3221) );
  ND2D1BWP12T U3560 ( .A1(n3222), .A2(n3221), .ZN(n2485) );
  TPND2D1BWP12T U3561 ( .A1(n3294), .A2(n3289), .ZN(n3224) );
  AOI22D0BWP12T U3562 ( .A1(write2_in[28]), .A2(n3291), .B1(r1[28]), .B2(n3290), .ZN(n3223) );
  ND2D1BWP12T U3563 ( .A1(n3224), .A2(n3223), .ZN(n2613) );
  TPND2D1BWP12T U3564 ( .A1(n3294), .A2(n3623), .ZN(n3226) );
  AOI22D0BWP12T U3565 ( .A1(write2_in[28]), .A2(n3281), .B1(r4[28]), .B2(n3280), .ZN(n3225) );
  ND2D1BWP12T U3566 ( .A1(n3226), .A2(n3225), .ZN(n2517) );
  TPND2D1BWP12T U3567 ( .A1(n3294), .A2(n3284), .ZN(n3228) );
  AOI22D0BWP12T U3568 ( .A1(write2_in[28]), .A2(n3286), .B1(r0[28]), .B2(n3285), .ZN(n3227) );
  ND2D1BWP12T U3569 ( .A1(n3228), .A2(n3227), .ZN(n2645) );
  TPND2D1BWP12T U3570 ( .A1(n3294), .A2(n3229), .ZN(n3233) );
  AOI22D0BWP12T U3571 ( .A1(write2_in[28]), .A2(n3231), .B1(n[3672]), .B2(
        n3230), .ZN(n3232) );
  ND2D1BWP12T U3572 ( .A1(n3233), .A2(n3232), .ZN(spin[28]) );
  TPND2D1BWP12T U3573 ( .A1(n3294), .A2(n3234), .ZN(n3238) );
  AOI22D0BWP12T U3574 ( .A1(write2_in[28]), .A2(n3236), .B1(lr[28]), .B2(n3235), .ZN(n3237) );
  TPND2D1BWP12T U3575 ( .A1(n3294), .A2(n3638), .ZN(n3240) );
  AOI22D0BWP12T U3576 ( .A1(write2_in[28]), .A2(n3277), .B1(tmp1[28]), .B2(
        n3276), .ZN(n3239) );
  ND2D1BWP12T U3577 ( .A1(n3240), .A2(n3239), .ZN(n2165) );
  TPND2D1BWP12T U3578 ( .A1(n3294), .A2(n3241), .ZN(n3245) );
  AOI22D0BWP12T U3579 ( .A1(write2_in[28]), .A2(n3243), .B1(r7[28]), .B2(n3242), .ZN(n3244) );
  ND2D1BWP12T U3580 ( .A1(n3245), .A2(n3244), .ZN(n2421) );
  AOI22D0BWP12T U3581 ( .A1(write2_in[31]), .A2(n3263), .B1(n3262), .B2(r6[31]), .ZN(n3246) );
  TPND2D1BWP12T U3582 ( .A1(n3294), .A2(n3248), .ZN(n3252) );
  AOI22D0BWP12T U3583 ( .A1(write2_in[28]), .A2(n3250), .B1(r9[28]), .B2(n3249), .ZN(n3251) );
  ND2D1BWP12T U3584 ( .A1(n3252), .A2(n3251), .ZN(n2357) );
  CKND2D1BWP12T U3585 ( .A1(n3259), .A2(n3627), .ZN(n3254) );
  AOI22D0BWP12T U3586 ( .A1(write2_in[31]), .A2(n3298), .B1(n3297), .B2(
        r10[31]), .ZN(n3253) );
  CKND2D1BWP12T U3587 ( .A1(n3259), .A2(n3624), .ZN(n3256) );
  AOI22D0BWP12T U3588 ( .A1(write2_in[31]), .A2(n3028), .B1(n3303), .B2(r3[31]), .ZN(n3255) );
  CKND2D1BWP12T U3589 ( .A1(n3259), .A2(n3625), .ZN(n3258) );
  AOI22D0BWP12T U3590 ( .A1(write2_in[31]), .A2(n3374), .B1(n3373), .B2(r2[31]), .ZN(n3257) );
  CKND2D1BWP12T U3591 ( .A1(n3259), .A2(n3626), .ZN(n3261) );
  AOI22D0BWP12T U3592 ( .A1(write2_in[31]), .A2(n3307), .B1(n3306), .B2(
        r11[31]), .ZN(n3260) );
  TPND2D1BWP12T U3593 ( .A1(n3294), .A2(n3628), .ZN(n3265) );
  AOI22D0BWP12T U3594 ( .A1(write2_in[28]), .A2(n3263), .B1(r6[28]), .B2(n3262), .ZN(n3264) );
  ND2D1BWP12T U3595 ( .A1(n3265), .A2(n3264), .ZN(n2453) );
  TPND2D1BWP12T U3596 ( .A1(n3294), .A2(n3627), .ZN(n3267) );
  AOI22D0BWP12T U3597 ( .A1(write2_in[28]), .A2(n3298), .B1(r10[28]), .B2(
        n3297), .ZN(n3266) );
  ND2D1BWP12T U3598 ( .A1(n3267), .A2(n3266), .ZN(n2325) );
  TPND2D1BWP12T U3599 ( .A1(n3294), .A2(n3625), .ZN(n3269) );
  AOI22D0BWP12T U3600 ( .A1(write2_in[28]), .A2(n3374), .B1(r2[28]), .B2(n3373), .ZN(n3268) );
  ND2D1BWP12T U3601 ( .A1(n3269), .A2(n3268), .ZN(n2581) );
  TPND2D1BWP12T U3602 ( .A1(n3294), .A2(n3624), .ZN(n3271) );
  AOI22D0BWP12T U3603 ( .A1(write2_in[28]), .A2(n3028), .B1(r3[28]), .B2(n3303), .ZN(n3270) );
  ND2D1BWP12T U3604 ( .A1(n3271), .A2(n3270), .ZN(n2549) );
  TPND2D1BWP12T U3605 ( .A1(n247), .A2(n3622), .ZN(n3275) );
  AOI22D0BWP12T U3606 ( .A1(write2_in[26]), .A2(n3273), .B1(n3272), .B2(r5[26]), .ZN(n3274) );
  TPND2D1BWP12T U3607 ( .A1(n247), .A2(n3638), .ZN(n3279) );
  AOI22D0BWP12T U3608 ( .A1(write2_in[26]), .A2(n3277), .B1(n3276), .B2(
        tmp1[26]), .ZN(n3278) );
  TPND2D1BWP12T U3609 ( .A1(n247), .A2(n3623), .ZN(n3283) );
  AOI22D0BWP12T U3610 ( .A1(write2_in[26]), .A2(n3281), .B1(n3280), .B2(r4[26]), .ZN(n3282) );
  TPND2D1BWP12T U3611 ( .A1(n247), .A2(n3284), .ZN(n3288) );
  AOI22D0BWP12T U3612 ( .A1(write2_in[26]), .A2(n3286), .B1(n3285), .B2(r0[26]), .ZN(n3287) );
  TPND2D1BWP12T U3613 ( .A1(n247), .A2(n3289), .ZN(n3293) );
  AOI22D0BWP12T U3614 ( .A1(write2_in[26]), .A2(n3291), .B1(n3290), .B2(r1[26]), .ZN(n3292) );
  TPND2D1BWP12T U3615 ( .A1(n3294), .A2(n3626), .ZN(n3296) );
  AOI22D0BWP12T U3616 ( .A1(write2_in[28]), .A2(n3307), .B1(r11[28]), .B2(
        n3306), .ZN(n3295) );
  ND2D1BWP12T U3617 ( .A1(n3296), .A2(n3295), .ZN(n2293) );
  TPND2D1BWP12T U3618 ( .A1(n247), .A2(n3627), .ZN(n3300) );
  AOI22D0BWP12T U3619 ( .A1(write2_in[26]), .A2(n3298), .B1(n3297), .B2(
        r10[26]), .ZN(n3299) );
  TPND2D1BWP12T U3620 ( .A1(n247), .A2(n3625), .ZN(n3302) );
  AOI22D0BWP12T U3621 ( .A1(write2_in[26]), .A2(n3374), .B1(n3373), .B2(r2[26]), .ZN(n3301) );
  TPND2D1BWP12T U3622 ( .A1(n247), .A2(n3624), .ZN(n3305) );
  AOI22D0BWP12T U3623 ( .A1(write2_in[26]), .A2(n3028), .B1(n3303), .B2(r3[26]), .ZN(n3304) );
  TPND2D1BWP12T U3624 ( .A1(n247), .A2(n3626), .ZN(n3309) );
  AOI22D0BWP12T U3625 ( .A1(write2_in[26]), .A2(n3307), .B1(n3306), .B2(
        r11[26]), .ZN(n3308) );
  TPNR3D1BWP12T U3626 ( .A1(n3310), .A2(n3394), .A3(n3325), .ZN(n3311) );
  TPND2D1BWP12T U3627 ( .A1(n3333), .A2(n3311), .ZN(n3319) );
  INR2D1BWP12T U3628 ( .A1(n3352), .B1(n238), .ZN(n3312) );
  INVD1BWP12T U3629 ( .I(n3313), .ZN(n3316) );
  ND3D1BWP12T U3630 ( .A1(n3319), .A2(n3318), .A3(n3317), .ZN(n2192) );
  AN2XD2BWP12T U3631 ( .A1(next_cpsr_in[3]), .A2(n3621), .Z(cpsrin[3]) );
  AN2XD2BWP12T U3632 ( .A1(next_cpsr_in[2]), .A2(n3621), .Z(cpsrin[2]) );
  CKAN2D1BWP12T U3633 ( .A1(n3320), .A2(n3352), .Z(n3321) );
  TPND2D2BWP12T U3634 ( .A1(n3324), .A2(n3352), .ZN(n3329) );
  ND2D1BWP12T U3635 ( .A1(n3328), .A2(n3327), .ZN(n3332) );
  NR2XD1BWP12T U3636 ( .A1(n3329), .A2(n45), .ZN(n3331) );
  INVD4BWP12T U3637 ( .I(n3335), .ZN(n3336) );
  NR2XD2BWP12T U3638 ( .A1(n3336), .A2(n238), .ZN(n3343) );
  TPND2D1BWP12T U3639 ( .A1(n3338), .A2(n3339), .ZN(n3351) );
  TPOAI21D1BWP12T U3640 ( .A1(n3343), .A2(n3342), .B(n3341), .ZN(n3346) );
  AN2XD2BWP12T U3641 ( .A1(n3347), .A2(n3344), .Z(n3345) );
  TPNR2D1BWP12T U3642 ( .A1(n3346), .A2(n3345), .ZN(n3350) );
  ND2D1BWP12T U3643 ( .A1(n3348), .A2(n3347), .ZN(n3349) );
  ND3D1BWP12T U3644 ( .A1(n3351), .A2(n3350), .A3(n3349), .ZN(n2195) );
  OA21XD0BWP12T U3645 ( .A1(write2_in[28]), .A2(n3381), .B(n3352), .Z(n3354)
         );
  INR2D1BWP12T U3646 ( .A1(n3381), .B1(write1_in[28]), .ZN(n3353) );
  AN2XD0BWP12T U3647 ( .A1(n3355), .A2(write2_in[26]), .Z(n3356) );
  TPNR2D1BWP12T U3648 ( .A1(n3358), .A2(n3357), .ZN(n3359) );
  TPND2D1BWP12T U3649 ( .A1(n3359), .A2(n3377), .ZN(n3369) );
  TPND2D1BWP12T U3650 ( .A1(n3360), .A2(n3361), .ZN(n3371) );
  AN2XD1BWP12T U3651 ( .A1(n3352), .A2(n3364), .Z(n3365) );
  INVD1BWP12T U3652 ( .I(n3367), .ZN(n3368) );
  TPND2D1BWP12T U3653 ( .A1(n3372), .A2(n3625), .ZN(n3376) );
  AOI22D0BWP12T U3654 ( .A1(write2_in[29]), .A2(n3374), .B1(n3373), .B2(r2[29]), .ZN(n3375) );
  ND2D1BWP12T U3655 ( .A1(n3376), .A2(n3375), .ZN(n2582) );
  TPND2D1BWP12T U3656 ( .A1(n3378), .A2(n3377), .ZN(n3387) );
  TPNR2D1BWP12T U3657 ( .A1(write1_in[30]), .A2(n3362), .ZN(n3383) );
  AOI21D0BWP12T U3658 ( .A1(n3379), .A2(write2_in[31]), .B(n3394), .ZN(n3380)
         );
  OAI21D0BWP12T U3659 ( .A1(write2_in[30]), .A2(n3381), .B(n3380), .ZN(n3382)
         );
  TPND2D1BWP12T U3660 ( .A1(n3385), .A2(n3384), .ZN(n3386) );
  CKND2D0BWP12T U3661 ( .A1(n3388), .A2(write2_in[28]), .ZN(n3389) );
  TPOAI21D2BWP12T U3662 ( .A1(n3620), .A2(n3390), .B(n3389), .ZN(n3392) );
  TPND2D1BWP12T U3663 ( .A1(n3391), .A2(n3392), .ZN(n3407) );
  OAI21D1BWP12T U3664 ( .A1(write2_in[31]), .A2(n1856), .B(n3352), .ZN(n3395)
         );
  TPAOI21D4BWP12T U3665 ( .A1(n3396), .A2(n1856), .B(n3395), .ZN(n3402) );
  AOI21D1BWP12T U3666 ( .A1(n3402), .A2(n3401), .B(n3400), .ZN(n3405) );
  TPND2D1BWP12T U3667 ( .A1(n3403), .A2(n3402), .ZN(n3404) );
  ND4D1BWP12T U3668 ( .A1(n3407), .A2(n3406), .A3(n3405), .A4(n3404), .ZN(
        n2200) );
  AOI22D0BWP12T U3669 ( .A1(n3472), .A2(tmp1[30]), .B1(n3471), .B2(r9[30]), 
        .ZN(n3408) );
  IOA21D1BWP12T U3670 ( .A1(n3474), .A2(r2[30]), .B(n3408), .ZN(n3412) );
  OAI22D0BWP12T U3671 ( .A1(n3448), .A2(n3654), .B1(n3476), .B2(n3653), .ZN(
        n3411) );
  OAI22D0BWP12T U3672 ( .A1(n3478), .A2(n3656), .B1(n3477), .B2(n3655), .ZN(
        n3410) );
  OAI22D1BWP12T U3673 ( .A1(n3481), .A2(n3658), .B1(n3657), .B2(n3422), .ZN(
        n3409) );
  NR4D0BWP12T U3674 ( .A1(n3412), .A2(n3411), .A3(n3410), .A4(n3409), .ZN(
        n3418) );
  OAI22D0BWP12T U3675 ( .A1(n3487), .A2(n3660), .B1(n3486), .B2(n3659), .ZN(
        n3416) );
  OAI22D0BWP12T U3676 ( .A1(n3489), .A2(n3662), .B1(n3661), .B2(n3488), .ZN(
        n3415) );
  OAI22D0BWP12T U3677 ( .A1(n3491), .A2(n3664), .B1(n3663), .B2(n3490), .ZN(
        n3414) );
  OAI22D0BWP12T U3678 ( .A1(n3666), .A2(n3463), .B1(n3492), .B2(n3665), .ZN(
        n3413) );
  NR4D0BWP12T U3679 ( .A1(n3416), .A2(n3415), .A3(n3414), .A4(n3413), .ZN(
        n3417) );
  ND2D1BWP12T U3680 ( .A1(n3418), .A2(n3417), .ZN(regA_out[30]) );
  AOI22D1BWP12T U3681 ( .A1(r9[27]), .A2(n3471), .B1(n3472), .B2(tmp1[27]), 
        .ZN(n3419) );
  OAI22D1BWP12T U3682 ( .A1(n3448), .A2(n3421), .B1(n3476), .B2(n3420), .ZN(
        n3429) );
  INVD1BWP12T U3683 ( .I(r10[27]), .ZN(n3423) );
  OAI22D1BWP12T U3684 ( .A1(n3481), .A2(n3424), .B1(n3423), .B2(n3422), .ZN(
        n3428) );
  OAI22D1BWP12T U3685 ( .A1(n3478), .A2(n3426), .B1(n3477), .B2(n3425), .ZN(
        n3427) );
  NR4D0BWP12T U3686 ( .A1(n3430), .A2(n3429), .A3(n3428), .A4(n3427), .ZN(
        n3444) );
  INVD1BWP12T U3687 ( .I(r7[27]), .ZN(n3431) );
  OAI22D1BWP12T U3688 ( .A1(n3487), .A2(n3431), .B1(n3486), .B2(n3647), .ZN(
        n3442) );
  INVD1BWP12T U3689 ( .I(r5[27]), .ZN(n3433) );
  OAI22D1BWP12T U3690 ( .A1(n3489), .A2(n3433), .B1(n3432), .B2(n3488), .ZN(
        n3441) );
  OAI22D1BWP12T U3691 ( .A1(n3491), .A2(n3435), .B1(n3434), .B2(n3490), .ZN(
        n3440) );
  NR4D0BWP12T U3692 ( .A1(n3442), .A2(n3441), .A3(n3440), .A4(n3439), .ZN(
        n3443) );
  AOI22D0BWP12T U3693 ( .A1(r9[24]), .A2(n3471), .B1(n3472), .B2(tmp1[24]), 
        .ZN(n3445) );
  IOA21D1BWP12T U3694 ( .A1(n3474), .A2(r2[24]), .B(n3445), .ZN(n3456) );
  OAI22D1BWP12T U3695 ( .A1(n3448), .A2(n3447), .B1(n3476), .B2(n3446), .ZN(
        n3455) );
  OAI22D1BWP12T U3696 ( .A1(n3478), .A2(n3450), .B1(n3477), .B2(n3449), .ZN(
        n3454) );
  OAI22D1BWP12T U3697 ( .A1(n3481), .A2(n3452), .B1(n3451), .B2(n3422), .ZN(
        n3453) );
  NR4D0BWP12T U3698 ( .A1(n3456), .A2(n3455), .A3(n3454), .A4(n3453), .ZN(
        n3470) );
  INVD1BWP12T U3699 ( .I(r7[24]), .ZN(n3457) );
  OAI22D1BWP12T U3700 ( .A1(n3487), .A2(n3457), .B1(n3486), .B2(n3644), .ZN(
        n3468) );
  INVD1BWP12T U3701 ( .I(r5[24]), .ZN(n3459) );
  OAI22D1BWP12T U3702 ( .A1(n3489), .A2(n3459), .B1(n3458), .B2(n3488), .ZN(
        n3467) );
  OAI22D1BWP12T U3703 ( .A1(n3491), .A2(n3461), .B1(n3460), .B2(n3490), .ZN(
        n3466) );
  OAI22D1BWP12T U3704 ( .A1(n3464), .A2(n3463), .B1(n3492), .B2(n3462), .ZN(
        n3465) );
  NR4D0BWP12T U3705 ( .A1(n3468), .A2(n3467), .A3(n3466), .A4(n3465), .ZN(
        n3469) );
  AOI22D0BWP12T U3706 ( .A1(n3472), .A2(tmp1[31]), .B1(n3471), .B2(r9[31]), 
        .ZN(n3473) );
  IOA21D1BWP12T U3707 ( .A1(n3474), .A2(r2[31]), .B(n3473), .ZN(n3485) );
  INVD1BWP12T U3708 ( .I(r0[31]), .ZN(n3537) );
  INVD1BWP12T U3709 ( .I(lr[31]), .ZN(n3550) );
  INVD1BWP12T U3710 ( .I(r8[31]), .ZN(n3547) );
  OAI22D0BWP12T U3711 ( .A1(n3478), .A2(n3550), .B1(n3477), .B2(n3547), .ZN(
        n3483) );
  INVD1BWP12T U3712 ( .I(r6[31]), .ZN(n3551) );
  OAI22D0BWP12T U3713 ( .A1(n3481), .A2(n3551), .B1(n3480), .B2(n3479), .ZN(
        n3482) );
  NR4D0BWP12T U3714 ( .A1(n3485), .A2(n3484), .A3(n3483), .A4(n3482), .ZN(
        n3498) );
  INVD1BWP12T U3715 ( .I(r3[31]), .ZN(n3549) );
  INVD1BWP12T U3716 ( .I(n[3669]), .ZN(n3548) );
  INVD1BWP12T U3717 ( .I(r11[31]), .ZN(n3538) );
  OAI22D0BWP12T U3718 ( .A1(n3491), .A2(n3548), .B1(n3538), .B2(n3490), .ZN(
        n3494) );
  INVD1BWP12T U3719 ( .I(r1[31]), .ZN(n3545) );
  INVD1BWP12T U3720 ( .I(r12[31]), .ZN(n3546) );
  OAI22D0BWP12T U3721 ( .A1(n3545), .A2(n3463), .B1(n3492), .B2(n3546), .ZN(
        n3493) );
  NR4D0BWP12T U3722 ( .A1(n3496), .A2(n3495), .A3(n3494), .A4(n3493), .ZN(
        n3497) );
  AOI22D1BWP12T U3723 ( .A1(tmp1[25]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[25]), .ZN(n3508) );
  INVD0BWP12T U3724 ( .I(r9[25]), .ZN(n3500) );
  OAI22D1BWP12T U3725 ( .A1(n3584), .A2(n3500), .B1(n3582), .B2(n3499), .ZN(
        n3504) );
  OAI22D1BWP12T U3726 ( .A1(n3586), .A2(n3502), .B1(n3588), .B2(n3501), .ZN(
        n3503) );
  NR2D1BWP12T U3727 ( .A1(n3504), .A2(n3503), .ZN(n3507) );
  AOI22D1BWP12T U3728 ( .A1(r5[25]), .A2(n3592), .B1(n3591), .B2(r10[25]), 
        .ZN(n3506) );
  AOI22D1BWP12T U3729 ( .A1(r7[25]), .A2(n1327), .B1(n3593), .B2(r2[25]), .ZN(
        n3505) );
  AN4XD1BWP12T U3730 ( .A1(n3508), .A2(n3507), .A3(n3506), .A4(n3505), .Z(
        n3521) );
  OAI22D0BWP12T U3731 ( .A1(n3510), .A2(n3600), .B1(n3599), .B2(n3509), .ZN(
        n3519) );
  OAI22D1BWP12T U3732 ( .A1(n3605), .A2(n3512), .B1(n3603), .B2(n3511), .ZN(
        n3518) );
  OAI22D1BWP12T U3733 ( .A1(n3514), .A2(n3571), .B1(n3607), .B2(n3513), .ZN(
        n3517) );
  OAI22D1BWP12T U3734 ( .A1(n3612), .A2(n3645), .B1(n3611), .B2(n3515), .ZN(
        n3516) );
  NR4D0BWP12T U3735 ( .A1(n3519), .A2(n3518), .A3(n3517), .A4(n3516), .ZN(
        n3520) );
  ND2D1BWP12T U3736 ( .A1(n3521), .A2(n3520), .ZN(regB_out[25]) );
  OAI22D1BWP12T U3737 ( .A1(n3584), .A2(n3640), .B1(n3582), .B2(n3654), .ZN(
        n3523) );
  OAI22D1BWP12T U3738 ( .A1(n3586), .A2(n3663), .B1(n3588), .B2(n3653), .ZN(
        n3522) );
  NR2D1BWP12T U3739 ( .A1(n3523), .A2(n3522), .ZN(n3527) );
  AOI22D1BWP12T U3740 ( .A1(r5[30]), .A2(n3592), .B1(n3591), .B2(r10[30]), 
        .ZN(n3526) );
  AOI22D1BWP12T U3741 ( .A1(r7[30]), .A2(n3524), .B1(n3593), .B2(r2[30]), .ZN(
        n3525) );
  AN4XD1BWP12T U3742 ( .A1(n3528), .A2(n3527), .A3(n3525), .A4(n3526), .Z(
        n3534) );
  OAI22D0BWP12T U3743 ( .A1(n3666), .A2(n3599), .B1(n3600), .B2(n3665), .ZN(
        n3532) );
  OAI22D1BWP12T U3744 ( .A1(n3605), .A2(n3664), .B1(n3603), .B2(n3655), .ZN(
        n3531) );
  OAI22D1BWP12T U3745 ( .A1(n3612), .A2(n3659), .B1(n3611), .B2(n3658), .ZN(
        n3529) );
  NR4D0BWP12T U3746 ( .A1(n3532), .A2(n3531), .A3(n3530), .A4(n3529), .ZN(
        n3533) );
  AOI22D1BWP12T U3747 ( .A1(tmp1[31]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[31]), .ZN(n3544) );
  CKND0BWP12T U3748 ( .I(r4[31]), .ZN(n3535) );
  OAI22D1BWP12T U3749 ( .A1(n3584), .A2(n3536), .B1(n3582), .B2(n3535), .ZN(
        n3540) );
  OAI22D1BWP12T U3750 ( .A1(n3586), .A2(n3538), .B1(n3588), .B2(n3537), .ZN(
        n3539) );
  NR2D1BWP12T U3751 ( .A1(n3540), .A2(n3539), .ZN(n3543) );
  AOI22D1BWP12T U3752 ( .A1(r5[31]), .A2(n3592), .B1(n3591), .B2(r10[31]), 
        .ZN(n3542) );
  AOI22D1BWP12T U3753 ( .A1(r7[31]), .A2(n3524), .B1(n3593), .B2(r2[31]), .ZN(
        n3541) );
  AN4XD1BWP12T U3754 ( .A1(n3544), .A2(n3543), .A3(n3542), .A4(n3541), .Z(
        n3557) );
  OAI22D0BWP12T U3755 ( .A1(n3546), .A2(n3600), .B1(n3599), .B2(n3545), .ZN(
        n3555) );
  OAI22D1BWP12T U3756 ( .A1(n3605), .A2(n3548), .B1(n3603), .B2(n3547), .ZN(
        n3554) );
  OAI22D1BWP12T U3757 ( .A1(n3550), .A2(n3571), .B1(n3607), .B2(n3549), .ZN(
        n3553) );
  OAI22D1BWP12T U3758 ( .A1(n3612), .A2(n3667), .B1(n3611), .B2(n3551), .ZN(
        n3552) );
  NR4D0BWP12T U3759 ( .A1(n3555), .A2(n3554), .A3(n3553), .A4(n3552), .ZN(
        n3556) );
  ND2D1BWP12T U3760 ( .A1(n3557), .A2(n3556), .ZN(regB_out[31]) );
  AOI22D1BWP12T U3761 ( .A1(tmp1[29]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[29]), .ZN(n3566) );
  OAI22D1BWP12T U3762 ( .A1(n3584), .A2(n3559), .B1(n3582), .B2(n3558), .ZN(
        n3562) );
  OAI22D1BWP12T U3763 ( .A1(n3586), .A2(n3652), .B1(n3588), .B2(n3560), .ZN(
        n3561) );
  AOI22D1BWP12T U3764 ( .A1(r5[29]), .A2(n3592), .B1(n3591), .B2(r10[29]), 
        .ZN(n3564) );
  AOI22D1BWP12T U3765 ( .A1(r7[29]), .A2(n1327), .B1(n3593), .B2(r2[29]), .ZN(
        n3563) );
  OAI22D0BWP12T U3766 ( .A1(n3568), .A2(n3599), .B1(n3600), .B2(n3567), .ZN(
        n3577) );
  OAI22D1BWP12T U3767 ( .A1(n3605), .A2(n3570), .B1(n3603), .B2(n3569), .ZN(
        n3576) );
  OAI22D1BWP12T U3768 ( .A1(n3572), .A2(n3571), .B1(n3607), .B2(n3651), .ZN(
        n3575) );
  OAI22D1BWP12T U3769 ( .A1(n3612), .A2(n3650), .B1(n3611), .B2(n3573), .ZN(
        n3574) );
  NR4D0BWP12T U3770 ( .A1(n3577), .A2(n3576), .A3(n3575), .A4(n3574), .ZN(
        n3578) );
  AOI22D1BWP12T U3771 ( .A1(tmp1[19]), .A2(n295), .B1(n3580), .B2(
        immediate2_in[19]), .ZN(n3597) );
  OAI22D1BWP12T U3772 ( .A1(n3584), .A2(n3583), .B1(n3582), .B2(n3581), .ZN(
        n3590) );
  OAI22D1BWP12T U3773 ( .A1(n3588), .A2(n3587), .B1(n3586), .B2(n3585), .ZN(
        n3589) );
  NR2D1BWP12T U3774 ( .A1(n3590), .A2(n3589), .ZN(n3596) );
  AOI22D1BWP12T U3775 ( .A1(r5[19]), .A2(n3592), .B1(n3591), .B2(r10[19]), 
        .ZN(n3595) );
  AOI22D1BWP12T U3776 ( .A1(r7[19]), .A2(n1327), .B1(n3593), .B2(r2[19]), .ZN(
        n3594) );
  AN4XD1BWP12T U3777 ( .A1(n3597), .A2(n3596), .A3(n3595), .A4(n3594), .Z(
        n3618) );
  OAI22D0BWP12T U3778 ( .A1(n3601), .A2(n3600), .B1(n3599), .B2(n3598), .ZN(
        n3616) );
  OAI22D1BWP12T U3779 ( .A1(n3605), .A2(n3604), .B1(n3603), .B2(n3602), .ZN(
        n3615) );
  OAI22D1BWP12T U3780 ( .A1(n3609), .A2(n3608), .B1(n3607), .B2(n3606), .ZN(
        n3614) );
  OAI22D1BWP12T U3781 ( .A1(n3612), .A2(n3641), .B1(n3611), .B2(n3610), .ZN(
        n3613) );
  NR4D0BWP12T U3782 ( .A1(n3616), .A2(n3615), .A3(n3614), .A4(n3613), .ZN(
        n3617) );
endmodule


module ALU_VARIABLE ( a, b, op, c_in, result, c_out, z, n, v );
  input [31:0] a;
  input [31:0] b;
  input [3:0] op;
  output [31:0] result;
  input c_in;
  output c_out, z, n, v;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328;

  DEL100D1BWP12T U3 ( .I(n4609), .Z(n1) );
  IOA21D2BWP12T U4 ( .A1(n746), .A2(n745), .B(n573), .ZN(n718) );
  CKND6BWP12T U5 ( .I(n513), .ZN(n514) );
  INVD2BWP12T U6 ( .I(n2135), .ZN(n2460) );
  ND2XD8BWP12T U7 ( .A1(n3103), .A2(n5292), .ZN(n5) );
  ND2D8BWP12T U8 ( .A1(n5), .A2(n24), .ZN(result[27]) );
  BUFFXD8BWP12T U9 ( .I(n2527), .Z(n2) );
  NR2D3BWP12T U10 ( .A1(a[4]), .A2(n515), .ZN(n516) );
  DCCKND4BWP12T U11 ( .I(n847), .ZN(n33) );
  INVD1BWP12T U12 ( .I(n2458), .ZN(n2459) );
  ND2XD4BWP12T U13 ( .A1(n1525), .A2(n1499), .ZN(n1560) );
  BUFFXD3BWP12T U14 ( .I(n521), .Z(n2303) );
  INVD3BWP12T U15 ( .I(n1765), .ZN(n1762) );
  TPND2D2BWP12T U16 ( .A1(n1753), .A2(n1752), .ZN(n1765) );
  IND2XD2BWP12T U17 ( .A1(n707), .B1(n709), .ZN(n673) );
  TPOAI21D2BWP12T U18 ( .A1(n1309), .A2(n3050), .B(n3051), .ZN(n1310) );
  NR2XD2BWP12T U19 ( .A1(n4), .A2(n3), .ZN(n2993) );
  CKND3BWP12T U20 ( .I(n1415), .ZN(n3) );
  XNR3XD4BWP12T U21 ( .A1(n1419), .A2(n1418), .A3(n1417), .ZN(n4) );
  INVD2BWP12T U22 ( .I(n1602), .ZN(n837) );
  CKND2D2BWP12T U23 ( .A1(n837), .A2(n836), .ZN(n841) );
  CKND0BWP12T U24 ( .I(n3939), .ZN(n2232) );
  INVD4BWP12T U25 ( .I(b[10]), .ZN(n3652) );
  DCCKND8BWP12T U26 ( .I(n4909), .ZN(n4935) );
  XOR3XD4BWP12T U27 ( .A1(n1335), .A2(n1334), .A3(n1333), .Z(n1350) );
  TPOAI22D2BWP12T U28 ( .A1(n2523), .A2(n1327), .B1(n1377), .B2(n2521), .ZN(
        n1333) );
  NR2D3BWP12T U29 ( .A1(n1576), .A2(n1575), .ZN(n1578) );
  OAI21D2BWP12T U30 ( .A1(n1579), .A2(n1578), .B(n1577), .ZN(n444) );
  INVD2BWP12T U31 ( .I(n550), .ZN(n490) );
  TPND2D4BWP12T U32 ( .A1(n431), .A2(n432), .ZN(n434) );
  ND2D8BWP12T U33 ( .A1(n433), .A2(n434), .ZN(n525) );
  TPND2D2BWP12T U34 ( .A1(n483), .A2(n550), .ZN(n489) );
  DCCKND12BWP12T U35 ( .I(n3915), .ZN(n4568) );
  XOR3XD4BWP12T U36 ( .A1(n2560), .A2(n2561), .A3(n2562), .Z(n2492) );
  TPND2D2BWP12T U37 ( .A1(n602), .A2(n738), .ZN(n604) );
  TPOAI21D1BWP12T U38 ( .A1(n903), .A2(n904), .B(n901), .ZN(n730) );
  INVD4BWP12T U39 ( .I(n1945), .ZN(n1941) );
  INVD8BWP12T U40 ( .I(n3590), .ZN(n2123) );
  NR3XD0BWP12T U41 ( .A1(n3102), .A2(n4597), .A3(n5145), .ZN(n9) );
  TPNR2D2BWP12T U42 ( .A1(n2462), .A2(n3334), .ZN(n1743) );
  TPOAI21D4BWP12T U43 ( .A1(n427), .A2(n1650), .B(n1648), .ZN(n768) );
  TPNR2D2BWP12T U44 ( .A1(n629), .A2(a[3]), .ZN(n515) );
  BUFFXD8BWP12T U45 ( .I(n1858), .Z(n6) );
  BUFFD8BWP12T U46 ( .I(n3913), .Z(n7) );
  ND2D4BWP12T U47 ( .A1(n484), .A2(n2220), .ZN(n488) );
  INVD8BWP12T U48 ( .I(n512), .ZN(n2185) );
  ND3XD1BWP12T U49 ( .A1(n9), .A2(n3166), .A3(n8), .ZN(n4596) );
  TPNR2D1BWP12T U50 ( .A1(n4988), .A2(n5100), .ZN(n8) );
  NR2XD3BWP12T U51 ( .A1(n1971), .A2(n10), .ZN(n2095) );
  TPNR2D3BWP12T U52 ( .A1(n1970), .A2(n1969), .ZN(n10) );
  TPND2D2BWP12T U53 ( .A1(n1720), .A2(n1722), .ZN(n457) );
  ND3XD4BWP12T U54 ( .A1(n455), .A2(n456), .A3(n457), .ZN(n1770) );
  XOR3XD4BWP12T U55 ( .A1(n1494), .A2(n11), .A3(n1383), .Z(n1472) );
  TPOAI21D2BWP12T U56 ( .A1(n1492), .A2(n2518), .B(n1491), .ZN(n11) );
  TPOAI22D1BWP12T U57 ( .A1(n52), .A2(n1856), .B1(n2477), .B2(n2006), .ZN(
        n1959) );
  OAI22D2BWP12T U58 ( .A1(n2535), .A2(n1432), .B1(n2533), .B2(n1504), .ZN(
        n1470) );
  CKND2D2BWP12T U59 ( .A1(n1733), .A2(n12), .ZN(n2464) );
  CKND2D2BWP12T U60 ( .A1(n1731), .A2(n3914), .ZN(n12) );
  TPND2D3BWP12T U61 ( .A1(n4943), .A2(n4568), .ZN(n1731) );
  IOA21D2BWP12T U62 ( .A1(n55), .A2(n1335), .B(n1328), .ZN(n1478) );
  INVD3BWP12T U63 ( .I(n3590), .ZN(n71) );
  TPND2D2BWP12T U64 ( .A1(n1281), .A2(n1280), .ZN(n1282) );
  TPND2D2BWP12T U65 ( .A1(n1610), .A2(n1633), .ZN(n1617) );
  TPOAI22D1BWP12T U66 ( .A1(n2016), .A2(n587), .B1(n586), .B2(n2519), .ZN(n633) );
  OAI21D1BWP12T U67 ( .A1(n633), .A2(n634), .B(n635), .ZN(n593) );
  ND2XD8BWP12T U68 ( .A1(n543), .A2(n2527), .ZN(n2529) );
  XNR2XD2BWP12T U69 ( .A1(n5033), .A2(n4500), .ZN(n707) );
  INVD2BWP12T U70 ( .I(n707), .ZN(n708) );
  RCOAI21D2BWP12T U71 ( .A1(n1572), .A2(n875), .B(n1573), .ZN(n877) );
  XNR3XD4BWP12T U72 ( .A1(n909), .A2(n908), .A3(n13), .ZN(n1572) );
  CKND3BWP12T U73 ( .I(n905), .ZN(n13) );
  BUFFXD8BWP12T U74 ( .I(n1384), .Z(n14) );
  INVD2BWP12T U75 ( .I(n740), .ZN(n599) );
  XNR2XD4BWP12T U76 ( .A1(n4914), .A2(n4896), .ZN(n1870) );
  TPND2D2BWP12T U77 ( .A1(n625), .A2(n628), .ZN(n609) );
  TPOAI22D2BWP12T U78 ( .A1(n2020), .A2(n667), .B1(n14), .B2(n666), .ZN(n696)
         );
  IOA21D2BWP12T U79 ( .A1(n688), .A2(n687), .B(n686), .ZN(n1722) );
  XOR3XD4BWP12T U80 ( .A1(n1609), .A2(n1607), .A3(n15), .Z(n1633) );
  CKND3BWP12T U81 ( .I(n1608), .ZN(n15) );
  TPND2D2BWP12T U82 ( .A1(n4596), .A2(n4595), .ZN(z) );
  OAI22D2BWP12T U83 ( .A1(n631), .A2(n2530), .B1(n2532), .B2(n754), .ZN(n803)
         );
  ND2D8BWP12T U84 ( .A1(n3913), .A2(n691), .ZN(n1679) );
  RCOAI21D2BWP12T U85 ( .A1(n2471), .A2(n600), .B(n467), .ZN(n618) );
  TPNR2D3BWP12T U86 ( .A1(n1706), .A2(n1756), .ZN(n1708) );
  TPOAI22D4BWP12T U87 ( .A1(n1709), .A2(n1708), .B1(n49), .B2(n1707), .ZN(
        n1897) );
  CKND2D2BWP12T U88 ( .A1(n2001), .A2(n2000), .ZN(n2002) );
  INVD2BWP12T U89 ( .I(n1973), .ZN(n1978) );
  XNR2XD2BWP12T U90 ( .A1(n436), .A2(n4944), .ZN(n1928) );
  BUFFD8BWP12T U91 ( .I(n4700), .Z(n16) );
  TPOAI22D2BWP12T U92 ( .A1(n601), .A2(n1872), .B1(n2469), .B2(n600), .ZN(n738) );
  TPOAI21D1BWP12T U93 ( .A1(n1777), .A2(n1776), .B(n1775), .ZN(n1779) );
  TPND2D2BWP12T U94 ( .A1(n1779), .A2(n1778), .ZN(n1882) );
  TPOAI22D2BWP12T U95 ( .A1(n705), .A2(n57), .B1(n704), .B2(n703), .ZN(n1724)
         );
  CKND3BWP12T U96 ( .I(n701), .ZN(n704) );
  TPOAI21D2BWP12T U97 ( .A1(n674), .A2(n2532), .B(n673), .ZN(n701) );
  TPND2D3BWP12T U98 ( .A1(n1769), .A2(n1768), .ZN(n1886) );
  BUFFD8BWP12T U99 ( .I(n4676), .Z(n17) );
  CKND2D2BWP12T U100 ( .A1(n18), .A2(n1884), .ZN(n1943) );
  ND2D3BWP12T U101 ( .A1(n1881), .A2(n19), .ZN(n18) );
  CKND3BWP12T U102 ( .I(n20), .ZN(n19) );
  NR2XD2BWP12T U103 ( .A1(n1882), .A2(n1883), .ZN(n20) );
  BUFFD8BWP12T U104 ( .I(b[27]), .Z(n21) );
  BUFFD8BWP12T U105 ( .I(n4610), .Z(n22) );
  TPOAI22D2BWP12T U106 ( .A1(n1689), .A2(n670), .B1(n671), .B2(n2481), .ZN(
        n700) );
  BUFFXD12BWP12T U107 ( .I(a[15]), .Z(n1906) );
  XNR3XD4BWP12T U108 ( .A1(n1852), .A2(n1855), .A3(n1851), .ZN(n1862) );
  ND2D3BWP12T U109 ( .A1(n1798), .A2(n1797), .ZN(n1851) );
  TPOAI22D1BWP12T U110 ( .A1(n52), .A2(n2093), .B1(n2477), .B2(n2478), .ZN(
        n2569) );
  BUFFD3BWP12T U111 ( .I(n2527), .Z(n23) );
  INVD12BWP12T U112 ( .I(n629), .ZN(n3911) );
  INVD1BWP12T U113 ( .I(n4672), .ZN(n445) );
  INVD8BWP12T U114 ( .I(n4500), .ZN(n3887) );
  XNR3XD4BWP12T U115 ( .A1(n1974), .A2(n1975), .A3(n1973), .ZN(n2028) );
  XNR3XD4BWP12T U116 ( .A1(n766), .A2(n765), .A3(n764), .ZN(n1648) );
  CKND3BWP12T U117 ( .I(n2799), .ZN(n24) );
  XNR2XD4BWP12T U118 ( .A1(n3157), .A2(n2738), .ZN(n3103) );
  TPOAI21D2BWP12T U119 ( .A1(n1747), .A2(n1748), .B(n1745), .ZN(n1746) );
  INVD18BWP12T U120 ( .I(n5112), .ZN(n5292) );
  TPNR2D2BWP12T U121 ( .A1(n1525), .A2(n1499), .ZN(n1561) );
  TPOAI22D2BWP12T U122 ( .A1(n2479), .A2(n1386), .B1(n2005), .B2(n1486), .ZN(
        n1456) );
  BUFFD8BWP12T U123 ( .I(n4732), .Z(n25) );
  TPND2D3BWP12T U124 ( .A1(n499), .A2(a[14]), .ZN(n502) );
  BUFFD8BWP12T U125 ( .I(b[14]), .Z(n5264) );
  XNR2XD4BWP12T U126 ( .A1(n3911), .A2(n5264), .ZN(n1485) );
  TPOAI22D4BWP12T U127 ( .A1(n1426), .A2(n3015), .B1(n439), .B2(n2476), .ZN(
        n1439) );
  TPND2D3BWP12T U128 ( .A1(n1207), .A2(n1208), .ZN(n1210) );
  OR2D2BWP12T U129 ( .A1(n1652), .A2(n925), .Z(n923) );
  BUFFD8BWP12T U130 ( .I(n5122), .Z(n26) );
  TPND2D1BWP12T U131 ( .A1(n1374), .A2(n1373), .ZN(n1375) );
  INVD8BWP12T U132 ( .I(n473), .ZN(n3938) );
  TPOAI22D1BWP12T U133 ( .A1(n1689), .A2(n1688), .B1(n2115), .B2(n1801), .ZN(
        n1780) );
  XNR3XD4BWP12T U134 ( .A1(n27), .A2(n2592), .A3(n2591), .ZN(n2598) );
  XOR3XD4BWP12T U135 ( .A1(n2503), .A2(n2502), .A3(n28), .Z(n27) );
  CKND3BWP12T U136 ( .I(n2501), .ZN(n28) );
  INVD8BWP12T U137 ( .I(n4565), .ZN(n450) );
  CKBD1BWP12T U138 ( .I(n2535), .Z(n29) );
  ND2D8BWP12T U139 ( .A1(n2351), .A2(n2139), .ZN(n5112) );
  TPND2D3BWP12T U140 ( .A1(n768), .A2(n767), .ZN(n846) );
  TPND2D2BWP12T U141 ( .A1(n3158), .A2(n3159), .ZN(n3148) );
  INR2D4BWP12T U142 ( .A1(n3152), .B1(n30), .ZN(n3158) );
  CKND3BWP12T U143 ( .I(n3144), .ZN(n30) );
  INVD3BWP12T U144 ( .I(n1377), .ZN(n1379) );
  INVD8BWP12T U145 ( .I(n4943), .ZN(n3913) );
  ND2XD4BWP12T U146 ( .A1(n4644), .A2(n5292), .ZN(n4667) );
  ND2D8BWP12T U147 ( .A1(n4667), .A2(n4666), .ZN(result[24]) );
  BUFFD8BWP12T U148 ( .I(n4991), .Z(n31) );
  BUFFXD12BWP12T U149 ( .I(n4770), .Z(n32) );
  INVD6BWP12T U150 ( .I(n629), .ZN(n513) );
  INVD3BWP12T U151 ( .I(n1153), .ZN(n1154) );
  RCOAI21D2BWP12T U152 ( .A1(n1767), .A2(n1766), .B(n1765), .ZN(n1769) );
  TPOAI22D2BWP12T U153 ( .A1(n2573), .A2(n693), .B1(n2571), .B2(n1693), .ZN(
        n1728) );
  IOA21D2BWP12T U154 ( .A1(n2010), .A2(n2009), .B(n2008), .ZN(n2011) );
  TPND2D2BWP12T U155 ( .A1(n33), .A2(n743), .ZN(n769) );
  XOR3XD4BWP12T U156 ( .A1(n720), .A2(n719), .A3(n718), .Z(n847) );
  TPOAI22D4BWP12T U157 ( .A1(n1872), .A2(n824), .B1(n757), .B2(n2469), .ZN(
        n899) );
  TPND2D1BWP12T U158 ( .A1(n898), .A2(n899), .ZN(n758) );
  INVD8BWP12T U159 ( .I(n3652), .ZN(n3939) );
  TPOAI22D2BWP12T U160 ( .A1(n1484), .A2(n2575), .B1(n1907), .B2(n34), .ZN(
        n1509) );
  TPOAI22D2BWP12T U161 ( .A1(n1907), .A2(n1502), .B1(n2575), .B2(n34), .ZN(
        n1542) );
  XNR2XD4BWP12T U162 ( .A1(n4301), .A2(n1906), .ZN(n34) );
  OAI21D1BWP12T U163 ( .A1(n1232), .A2(n1231), .B(n35), .ZN(n1230) );
  XOR3XD4BWP12T U164 ( .A1(n1232), .A2(n1188), .A3(n35), .Z(n1207) );
  OAI22D4BWP12T U165 ( .A1(n1872), .A2(n1187), .B1(n1234), .B2(n2469), .ZN(n35) );
  CKND3BWP12T U166 ( .I(b[8]), .ZN(n474) );
  TPOAI22D2BWP12T U167 ( .A1(n1689), .A2(n1354), .B1(n2115), .B2(n36), .ZN(
        n1372) );
  OAI22D2BWP12T U168 ( .A1(n1689), .A2(n36), .B1(n1487), .B2(n2481), .ZN(n1464) );
  XNR2XD2BWP12T U169 ( .A1(n4511), .A2(n3899), .ZN(n36) );
  TPOAI22D2BWP12T U170 ( .A1(n2518), .A2(n37), .B1(n865), .B2(n2516), .ZN(
        n1444) );
  OAI22D2BWP12T U171 ( .A1(n2518), .A2(n1445), .B1(n2516), .B2(n37), .ZN(n1489) );
  XNR2XD1BWP12T U172 ( .A1(n5196), .A2(a[17]), .ZN(n37) );
  BUFFD12BWP12T U173 ( .I(n1106), .Z(n5081) );
  OR2D2BWP12T U174 ( .A1(n601), .A2(n1384), .Z(n565) );
  XOR2XD4BWP12T U175 ( .A1(n4916), .A2(n5033), .Z(n1740) );
  BUFFD6BWP12T U176 ( .I(a[20]), .Z(n2141) );
  TPNR2D2BWP12T U177 ( .A1(n547), .A2(n1969), .ZN(n482) );
  XNR2D2BWP12T U178 ( .A1(n3948), .A2(n4568), .ZN(n1711) );
  TPNR2D1BWP12T U179 ( .A1(n625), .A2(n628), .ZN(n611) );
  INVD3BWP12T U180 ( .I(n1313), .ZN(n1362) );
  XNR2XD4BWP12T U181 ( .A1(n2123), .A2(n4700), .ZN(n666) );
  OR2D4BWP12T U182 ( .A1(n2020), .A2(n757), .Z(n564) );
  TPNR2D3BWP12T U183 ( .A1(n2469), .A2(n1385), .ZN(n1313) );
  TPND2D1BWP12T U184 ( .A1(n1457), .A2(n1456), .ZN(n1458) );
  TPND2D2BWP12T U185 ( .A1(n5145), .A2(n5292), .ZN(n5179) );
  CKAN2D2BWP12T U186 ( .A1(n38), .A2(n695), .Z(n1726) );
  XOR2D2BWP12T U187 ( .A1(n38), .A2(n695), .Z(n584) );
  TPOAI22D2BWP12T U188 ( .A1(n2518), .A2(n494), .B1(n535), .B2(n2022), .ZN(n38) );
  ND2D3BWP12T U189 ( .A1(n39), .A2(n2042), .ZN(n3146) );
  TPNR2D3BWP12T U190 ( .A1(n39), .A2(n2042), .ZN(n3145) );
  XNR3XD4BWP12T U191 ( .A1(n2129), .A2(n2128), .A3(n2131), .ZN(n39) );
  ND2XD3BWP12T U192 ( .A1(n41), .A2(n40), .ZN(n1518) );
  ND2D3BWP12T U193 ( .A1(n1473), .A2(n1472), .ZN(n40) );
  TPOAI21D2BWP12T U194 ( .A1(n1473), .A2(n1472), .B(n1471), .ZN(n41) );
  XNR3XD4BWP12T U195 ( .A1(n1456), .A2(n1455), .A3(n42), .ZN(n1473) );
  CKND3BWP12T U196 ( .I(n1518), .ZN(n45) );
  CKND3BWP12T U197 ( .I(n1457), .ZN(n42) );
  ND2XD8BWP12T U198 ( .A1(n43), .A2(n809), .ZN(n2532) );
  XOR2XD4BWP12T U199 ( .A1(n4500), .A2(n2141), .Z(n43) );
  ND2D3BWP12T U200 ( .A1(n708), .A2(n43), .ZN(n710) );
  ND2XD3BWP12T U201 ( .A1(n3131), .A2(n404), .ZN(n1675) );
  TPND2D3BWP12T U202 ( .A1(n1674), .A2(n1673), .ZN(n404) );
  TPND2D2BWP12T U203 ( .A1(n1584), .A2(n1583), .ZN(n1516) );
  ND2D3BWP12T U204 ( .A1(n44), .A2(n1517), .ZN(n1584) );
  XNR3XD4BWP12T U205 ( .A1(n1482), .A2(n1483), .A3(n424), .ZN(n1517) );
  ND2D3BWP12T U206 ( .A1(n45), .A2(n46), .ZN(n44) );
  DCCKND4BWP12T U207 ( .I(n419), .ZN(n46) );
  XOR3XD4BWP12T U208 ( .A1(n1433), .A2(n1469), .A3(n1468), .Z(n424) );
  ND2D3BWP12T U209 ( .A1(n1467), .A2(n1466), .ZN(n1483) );
  TPOAI22D2BWP12T U210 ( .A1(n1799), .A2(n728), .B1(n2467), .B2(n47), .ZN(n904) );
  TPOAI22D2BWP12T U211 ( .A1(n870), .A2(n2467), .B1(n1799), .B2(n47), .ZN(n880) );
  XNR2XD4BWP12T U212 ( .A1(n3939), .A2(n5079), .ZN(n47) );
  TPAOI21D1BWP12T U213 ( .A1(n4282), .A2(n4281), .B(n5240), .ZN(n5227) );
  TPOAI22D1BWP12T U214 ( .A1(n3591), .A2(n4635), .B1(n3588), .B2(n3888), .ZN(
        n239) );
  TPOAI22D2BWP12T U215 ( .A1(n3557), .A2(n3948), .B1(n3618), .B2(n2394), .ZN(
        n5127) );
  TPND2D2BWP12T U216 ( .A1(n2391), .A2(n2390), .ZN(n3557) );
  OAI222D0BWP12T U217 ( .A1(n4815), .A2(n4307), .B1(n4817), .B2(n4319), .C1(
        n5183), .C2(n4306), .ZN(n5130) );
  OAI22D0BWP12T U218 ( .A1(n3620), .A2(n3609), .B1(n3608), .B2(n3618), .ZN(
        n3602) );
  NR2D1BWP12T U219 ( .A1(n3620), .A2(n3730), .ZN(n3621) );
  TPNR2D1BWP12T U220 ( .A1(n2903), .A2(n2902), .ZN(n3620) );
  TPNR2D1BWP12T U221 ( .A1(n4891), .A2(n4892), .ZN(n225) );
  AO31XD2BWP12T U222 ( .A1(n4421), .A2(n226), .A3(n4413), .B(n228), .Z(n2635)
         );
  DCCKND4BWP12T U223 ( .I(n4311), .ZN(n4242) );
  XOR2XD4BWP12T U224 ( .A1(n3040), .A2(n3039), .Z(n5250) );
  TPNR2D1BWP12T U225 ( .A1(n2270), .A2(n2190), .ZN(n4046) );
  TPOAI21D1BWP12T U226 ( .A1(n4046), .A2(n4043), .B(n4416), .ZN(n4048) );
  CKND2D2BWP12T U227 ( .A1(n2270), .A2(n2190), .ZN(n4416) );
  XNR2D2BWP12T U228 ( .A1(n3948), .A2(n5079), .ZN(n1235) );
  ND2D4BWP12T U229 ( .A1(n4810), .A2(n4809), .ZN(result[17]) );
  TPOAI21D1BWP12T U230 ( .A1(n3084), .A2(n3076), .B(n412), .ZN(n3081) );
  ND2D4BWP12T U231 ( .A1(n4724), .A2(n4723), .ZN(result[19]) );
  TPND2D1BWP12T U232 ( .A1(n5070), .A2(n3060), .ZN(n3069) );
  XNR2D2BWP12T U233 ( .A1(n3063), .A2(n3055), .ZN(n5070) );
  TPND2D4BWP12T U234 ( .A1(n403), .A2(n436), .ZN(n486) );
  TPND2D2BWP12T U235 ( .A1(n1006), .A2(n2626), .ZN(n2943) );
  INVD3BWP12T U236 ( .I(n3895), .ZN(n48) );
  INVD2BWP12T U237 ( .I(a[15]), .ZN(n3895) );
  XNR2XD2BWP12T U238 ( .A1(n1812), .A2(n1277), .ZN(n1326) );
  ND2D3BWP12T U239 ( .A1(n1679), .A2(n2773), .ZN(n1733) );
  DCCKBD4BWP12T U240 ( .I(n1906), .Z(n4508) );
  XNR2XD2BWP12T U241 ( .A1(n48), .A2(n3939), .ZN(n546) );
  BUFFD2BWP12T U242 ( .I(n1755), .Z(n49) );
  DEL025D1BWP12T U243 ( .I(n3115), .Z(n50) );
  TPNR2D2BWP12T U244 ( .A1(n3109), .A2(n2991), .ZN(n3115) );
  XNR2XD2BWP12T U245 ( .A1(a[14]), .A2(n6), .ZN(n51) );
  INVD16BWP12T U246 ( .I(n507), .ZN(n1858) );
  TPND2D2BWP12T U247 ( .A1(n4785), .A2(n5292), .ZN(n4810) );
  TPND2D3BWP12T U248 ( .A1(n5100), .A2(n5292), .ZN(n2384) );
  XNR2D1BWP12T U249 ( .A1(n3016), .A2(n2123), .ZN(n990) );
  TPOAI22D2BWP12T U250 ( .A1(n2518), .A2(n1925), .B1(n2023), .B2(n2516), .ZN(
        n1994) );
  CKND2D2BWP12T U251 ( .A1(n1703), .A2(n1702), .ZN(n1704) );
  OR3D2BWP12T U252 ( .A1(n3042), .A2(n3041), .A3(n5250), .Z(n3070) );
  XOR3D2BWP12T U253 ( .A1(n2552), .A2(n2553), .A3(n2550), .Z(n2512) );
  TPOAI21D1BWP12T U254 ( .A1(n1703), .A2(n1702), .B(n1701), .ZN(n1705) );
  INVD1P25BWP12T U255 ( .I(n2005), .ZN(n63) );
  TPNR2D1BWP12T U256 ( .A1(n2643), .A2(n2642), .ZN(n3575) );
  INVD3BWP12T U257 ( .I(n2635), .ZN(n4408) );
  DCCKBD4BWP12T U258 ( .I(n2479), .Z(n52) );
  XOR3XD4BWP12T U259 ( .A1(n1043), .A2(n1044), .A3(n1046), .Z(n1003) );
  OAI22D4BWP12T U260 ( .A1(n1049), .A2(n2005), .B1(n2479), .B2(n1022), .ZN(
        n1057) );
  XNR2D2BWP12T U261 ( .A1(n3948), .A2(n3911), .ZN(n1009) );
  IND2XD8BWP12T U262 ( .A1(a[0]), .B1(a[1]), .ZN(n2476) );
  TPAOI31D1BWP12T U263 ( .A1(n966), .A2(n965), .A3(n3024), .B(n964), .ZN(n53)
         );
  TPAOI31D1BWP12T U264 ( .A1(n966), .A2(n965), .A3(n3024), .B(n964), .ZN(n3011) );
  AN2D1BWP12T U265 ( .A1(n2041), .A2(n2040), .Z(n54) );
  ND2XD4BWP12T U266 ( .A1(n1940), .A2(n1939), .ZN(n2040) );
  INVD9BWP12T U267 ( .I(n468), .ZN(n2014) );
  TPOAI22D4BWP12T U268 ( .A1(n710), .A2(n709), .B1(n2530), .B2(n1691), .ZN(
        n1685) );
  DCCKND4BWP12T U269 ( .I(n1550), .ZN(n1454) );
  TPOAI22D1BWP12T U270 ( .A1(n1329), .A2(n3015), .B1(n1326), .B2(n1969), .ZN(
        n55) );
  TPOAI22D1BWP12T U271 ( .A1(n1329), .A2(n3015), .B1(n1326), .B2(n1969), .ZN(
        n1334) );
  INVD2BWP12T U272 ( .I(n618), .ZN(n477) );
  INVD4BWP12T U273 ( .I(a[7]), .ZN(n3590) );
  XNR2D2BWP12T U274 ( .A1(a[17]), .A2(n3948), .ZN(n865) );
  XNR2D2BWP12T U275 ( .A1(b[1]), .A2(n1906), .ZN(n1355) );
  INVD2BWP12T U276 ( .I(n2910), .ZN(n56) );
  DCCKND8BWP12T U277 ( .I(a[9]), .ZN(n2910) );
  XNR2XD2BWP12T U278 ( .A1(n48), .A2(n3938), .ZN(n795) );
  XNR2XD2BWP12T U279 ( .A1(n1906), .A2(n4770), .ZN(n2007) );
  XNR2XD2BWP12T U280 ( .A1(n1906), .A2(n5085), .ZN(n694) );
  XNR2D2BWP12T U281 ( .A1(n3930), .A2(n48), .ZN(n555) );
  XNR2D2BWP12T U282 ( .A1(n3948), .A2(n1906), .ZN(n1484) );
  TPND2D3BWP12T U283 ( .A1(n3653), .A2(n4509), .ZN(n2961) );
  DCCKND4BWP12T U284 ( .I(n3899), .ZN(n3653) );
  XNR2D2BWP12T U285 ( .A1(n4676), .A2(n513), .ZN(n706) );
  OA22D1BWP12T U286 ( .A1(n2481), .A2(n671), .B1(n1689), .B2(n670), .Z(n57) );
  XNR2XD2BWP12T U287 ( .A1(n4511), .A2(n4794), .ZN(n671) );
  XNR2XD2BWP12T U288 ( .A1(n4511), .A2(n4826), .ZN(n670) );
  TPND2D2BWP12T U289 ( .A1(n1990), .A2(n1989), .ZN(n1991) );
  ND2D4BWP12T U290 ( .A1(n1675), .A2(n3134), .ZN(n3123) );
  DEL025D1BWP12T U291 ( .I(n696), .Z(n58) );
  HA1D2BWP12T U292 ( .A(n1810), .B(n1809), .CO(n1877), .S(n1806) );
  TPOAI22D4BWP12T U293 ( .A1(n397), .A2(n1741), .B1(n1740), .B2(n2519), .ZN(
        n1809) );
  TPAOI21D4BWP12T U294 ( .A1(n1699), .A2(n1700), .B(n1698), .ZN(n1755) );
  INVD2BWP12T U295 ( .I(n627), .ZN(n610) );
  TPND2D2BWP12T U296 ( .A1(n1926), .A2(n2017), .ZN(n2545) );
  XNR2D2BWP12T U297 ( .A1(a[17]), .A2(n3930), .ZN(n535) );
  TPOAI22D1BWP12T U298 ( .A1(n2545), .A2(n2018), .B1(n2085), .B2(n413), .ZN(
        n2103) );
  INVD4BWP12T U299 ( .I(a[2]), .ZN(n2220) );
  INVD4BWP12T U300 ( .I(a[1]), .ZN(n484) );
  OR2XD1BWP12T U301 ( .A1(n964), .A2(n3023), .Z(n3029) );
  TPNR2D3BWP12T U302 ( .A1(n60), .A2(n59), .ZN(n964) );
  INVD2P3BWP12T U303 ( .I(n962), .ZN(n59) );
  DCCKND4BWP12T U304 ( .I(n963), .ZN(n60) );
  TPND2D2BWP12T U305 ( .A1(n62), .A2(n61), .ZN(n1898) );
  ND2D3BWP12T U306 ( .A1(n1759), .A2(n1757), .ZN(n61) );
  TPOAI21D2BWP12T U307 ( .A1(n1759), .A2(n1757), .B(n1760), .ZN(n62) );
  XOR3XD4BWP12T U308 ( .A1(n1782), .A2(n1780), .A3(n1783), .Z(n1760) );
  OAI22D2BWP12T U309 ( .A1(n1687), .A2(n2479), .B1(n2005), .B2(n1710), .ZN(
        n1782) );
  XOR3XD4BWP12T U310 ( .A1(n1818), .A2(n1815), .A3(n1817), .Z(n1757) );
  TPOAI21D2BWP12T U311 ( .A1(n2464), .A2(n1682), .B(n1681), .ZN(n1817) );
  XNR2D2BWP12T U312 ( .A1(n1812), .A2(n689), .ZN(n1739) );
  TPOAI22D4BWP12T U313 ( .A1(n1969), .A2(n1813), .B1(n1910), .B2(n3015), .ZN(
        n1905) );
  OAI21D0BWP12T U314 ( .A1(n1562), .A2(n1561), .B(n1560), .ZN(n1568) );
  IND2D4BWP12T U315 ( .A1(n1559), .B1(n1560), .ZN(n1501) );
  TPOAI21D1BWP12T U316 ( .A1(n781), .A2(n647), .B(n779), .ZN(n649) );
  XNR3XD4BWP12T U317 ( .A1(n777), .A2(n778), .A3(n776), .ZN(n647) );
  TPOAI22D1BWP12T U318 ( .A1(n2479), .A2(n2006), .B1(n2093), .B2(n2005), .ZN(
        n2090) );
  CKND2D2BWP12T U319 ( .A1(n969), .A2(n65), .ZN(n66) );
  TPND2D2BWP12T U320 ( .A1(n64), .A2(n970), .ZN(n67) );
  TPND2D3BWP12T U321 ( .A1(n66), .A2(n67), .ZN(n974) );
  INVD2BWP12T U322 ( .I(n969), .ZN(n64) );
  INVD2BWP12T U323 ( .I(n970), .ZN(n65) );
  IOA21D2BWP12T U324 ( .A1(n976), .A2(n975), .B(n974), .ZN(n977) );
  TPNR2D1BWP12T U325 ( .A1(n791), .A2(n790), .ZN(n645) );
  XNR2XD2BWP12T U326 ( .A1(n4565), .A2(n4896), .ZN(n511) );
  OR2D2BWP12T U327 ( .A1(n1264), .A2(n1263), .Z(n1267) );
  XNR2D2BWP12T U328 ( .A1(a[1]), .A2(b[18]), .ZN(n1426) );
  XNR2D2BWP12T U329 ( .A1(n4511), .A2(n4732), .ZN(n1688) );
  OAI21D1BWP12T U330 ( .A1(n424), .A2(n1564), .B(n1563), .ZN(n1569) );
  TPND2D2BWP12T U331 ( .A1(n1220), .A2(n1219), .ZN(n1292) );
  TPND2D2BWP12T U332 ( .A1(n1215), .A2(n1214), .ZN(n1220) );
  TPND2D2BWP12T U333 ( .A1(n1213), .A2(n1212), .ZN(n1215) );
  INVD4BWP12T U334 ( .I(n1213), .ZN(n1218) );
  TPND2D1BWP12T U335 ( .A1(n3063), .A2(n3047), .ZN(n3049) );
  ND2D4BWP12T U336 ( .A1(n1663), .A2(n1662), .ZN(n3106) );
  XOR3XD4BWP12T U337 ( .A1(n1582), .A2(n1581), .A3(n1580), .Z(n1626) );
  DCCKND4BWP12T U338 ( .I(n2516), .ZN(n68) );
  INVD2BWP12T U339 ( .I(n1253), .ZN(n1255) );
  IOA21D1BWP12T U340 ( .A1(n1252), .A2(n1253), .B(n1251), .ZN(n1257) );
  XNR2XD2BWP12T U341 ( .A1(n3016), .A2(n436), .ZN(n928) );
  DEL025D1BWP12T U342 ( .I(n1542), .Z(n69) );
  DCCKND4BWP12T U343 ( .I(a[2]), .ZN(n70) );
  DCCKBD12BWP12T U344 ( .I(b[1]), .Z(n3908) );
  BUFFXD12BWP12T U345 ( .I(b[1]), .Z(n4849) );
  XNR2XD2BWP12T U346 ( .A1(b[1]), .A2(n4503), .ZN(n1794) );
  XNR2D2BWP12T U347 ( .A1(n5079), .A2(b[1]), .ZN(n1142) );
  XNR2XD2BWP12T U348 ( .A1(b[1]), .A2(n4565), .ZN(n882) );
  XNR2D2BWP12T U349 ( .A1(n2014), .A2(b[1]), .ZN(n586) );
  INVD4BWP12T U350 ( .I(n521), .ZN(n1007) );
  BUFFXD0BWP12T U351 ( .I(a[14]), .Z(n5256) );
  CKND2D2BWP12T U352 ( .A1(n3165), .A2(n3164), .ZN(n5145) );
  NR2XD1BWP12T U353 ( .A1(n1350), .A2(n1349), .ZN(n1352) );
  TPNR2D1BWP12T U354 ( .A1(n889), .A2(n1581), .ZN(n891) );
  INVD2BWP12T U355 ( .I(n1582), .ZN(n889) );
  BUFFXD3BWP12T U356 ( .I(b[30]), .Z(n5153) );
  MUX2ND0BWP12T U357 ( .I0(n5295), .I1(n5294), .S(n5153), .ZN(n5147) );
  OAI21D2BWP12T U358 ( .A1(n1718), .A2(n1717), .B(n1715), .ZN(n1716) );
  CKND2D2BWP12T U359 ( .A1(n3649), .A2(n4508), .ZN(n3447) );
  XNR2D2BWP12T U360 ( .A1(n4301), .A2(n2123), .ZN(n1102) );
  OAI22D2BWP12T U361 ( .A1(n1689), .A2(n3898), .B1(n2481), .B2(n1017), .ZN(
        n1063) );
  BUFFD2BWP12T U362 ( .I(n786), .Z(n440) );
  ND2XD8BWP12T U363 ( .A1(n486), .A2(n485), .ZN(n2523) );
  XNR2D2BWP12T U364 ( .A1(n3016), .A2(n3911), .ZN(n948) );
  ND2D4BWP12T U365 ( .A1(n1738), .A2(n1737), .ZN(n1805) );
  CKND2D2BWP12T U366 ( .A1(n430), .A2(n1805), .ZN(n1807) );
  TPND2D2BWP12T U367 ( .A1(n3098), .A2(n3097), .ZN(n3149) );
  ND2D3BWP12T U368 ( .A1(n2041), .A2(n2040), .ZN(n3141) );
  TPND2D2BWP12T U369 ( .A1(n416), .A2(n417), .ZN(n1910) );
  TPNR2D1BWP12T U370 ( .A1(n1892), .A2(n1891), .ZN(n1895) );
  XNR2D2BWP12T U371 ( .A1(n3948), .A2(n2014), .ZN(n680) );
  TPOAI21D2BWP12T U372 ( .A1(n477), .A2(n476), .B(n475), .ZN(n583) );
  INVD1BWP12T U373 ( .I(n1293), .ZN(n1289) );
  DEL025D1BWP12T U374 ( .I(n3123), .Z(n72) );
  TPOAI22D2BWP12T U375 ( .A1(n2523), .A2(n591), .B1(n2521), .B2(n590), .ZN(
        n635) );
  TPOAI21D1BWP12T U376 ( .A1(n534), .A2(n533), .B(n531), .ZN(n532) );
  CKND2D2BWP12T U377 ( .A1(n766), .A2(n763), .ZN(n641) );
  XNR2XD4BWP12T U378 ( .A1(n3911), .A2(n4301), .ZN(n1022) );
  OAI22D2BWP12T U379 ( .A1(n2529), .A2(n1690), .B1(n1711), .B2(n2527), .ZN(
        n1783) );
  TPND2D1BWP12T U380 ( .A1(n1125), .A2(n1124), .ZN(n1126) );
  AN3XD2BWP12T U381 ( .A1(n4933), .A2(n4932), .A3(n4931), .Z(n4934) );
  INVD1BWP12T U382 ( .I(n1812), .ZN(n414) );
  XNR2D1BWP12T U383 ( .A1(n5079), .A2(n4794), .ZN(n1800) );
  XNR2D1BWP12T U384 ( .A1(n5196), .A2(n4503), .ZN(n1867) );
  XNR2D1BWP12T U385 ( .A1(n4503), .A2(n3948), .ZN(n2021) );
  CKND2D2BWP12T U386 ( .A1(n1905), .A2(n1904), .ZN(n399) );
  CKND0BWP12T U387 ( .I(n2012), .ZN(n2010) );
  BUFFXD3BWP12T U388 ( .I(n1799), .Z(n2465) );
  TPOAI22D1BWP12T U389 ( .A1(n2535), .A2(n510), .B1(n2533), .B2(n711), .ZN(
        n531) );
  OAI22D1BWP12T U390 ( .A1(n2479), .A2(n706), .B1(n1687), .B2(n2005), .ZN(
        n1686) );
  ND2D1BWP12T U391 ( .A1(n1178), .A2(n1177), .ZN(n1179) );
  TPNR2D2BWP12T U392 ( .A1(n1206), .A2(n1205), .ZN(n1211) );
  TPND2D2BWP12T U393 ( .A1(n1320), .A2(n1319), .ZN(n1365) );
  TPOAI22D1BWP12T U394 ( .A1(n2573), .A2(n3890), .B1(n2571), .B2(n881), .ZN(
        n1425) );
  OAI21D1BWP12T U395 ( .A1(n1546), .A2(n1545), .B(n1544), .ZN(n1612) );
  INVD1BWP12T U396 ( .I(n1623), .ZN(n916) );
  CKND2D0BWP12T U397 ( .A1(n1035), .A2(n1036), .ZN(n1027) );
  OAI22D1BWP12T U398 ( .A1(n1689), .A2(n1018), .B1(n2115), .B2(n1050), .ZN(
        n1062) );
  XNR2XD2BWP12T U399 ( .A1(n4501), .A2(n3938), .ZN(n1024) );
  XNR2D2BWP12T U400 ( .A1(n4501), .A2(n4896), .ZN(n982) );
  INVD1BWP12T U401 ( .I(n856), .ZN(n850) );
  IND2D1BWP12T U402 ( .A1(n623), .B1(n526), .ZN(n528) );
  TPOAI21D1BWP12T U403 ( .A1(n520), .A2(n519), .B(n518), .ZN(n660) );
  INVD1BWP12T U404 ( .I(n607), .ZN(n520) );
  TPNR2D1BWP12T U405 ( .A1(n1520), .A2(n1521), .ZN(n1523) );
  AN2D1BWP12T U406 ( .A1(n1569), .A2(n1568), .Z(n1570) );
  NR2D2BWP12T U407 ( .A1(n1567), .A2(n1566), .ZN(n1571) );
  CKND2D2BWP12T U408 ( .A1(n1618), .A2(n1634), .ZN(n1619) );
  TPND2D2BWP12T U409 ( .A1(n1401), .A2(n1400), .ZN(n1418) );
  TPOAI21D1BWP12T U410 ( .A1(n1397), .A2(n1398), .B(n1396), .ZN(n1401) );
  NR2D2BWP12T U411 ( .A1(n3076), .A2(n418), .ZN(n1600) );
  CKND2D0BWP12T U412 ( .A1(n4801), .A2(n4301), .ZN(n3603) );
  AOI21D1BWP12T U413 ( .A1(n3882), .A2(n4861), .B(n3838), .ZN(n4870) );
  CKND2D2BWP12T U414 ( .A1(n936), .A2(n3019), .ZN(n937) );
  TPNR2D3BWP12T U415 ( .A1(n981), .A2(n980), .ZN(n3008) );
  BUFFXD6BWP12T U416 ( .I(b[24]), .Z(n4655) );
  INVD1BWP12T U417 ( .I(n570), .ZN(n556) );
  ND2D1BWP12T U418 ( .A1(n722), .A2(n723), .ZN(n562) );
  IOA21D1BWP12T U419 ( .A1(n5141), .A2(n5305), .B(n5140), .ZN(n5142) );
  INR2D1BWP12T U420 ( .A1(n2725), .B1(n2724), .ZN(n2726) );
  ND2D1BWP12T U421 ( .A1(n2412), .A2(n2348), .ZN(n5105) );
  INVD1BWP12T U422 ( .I(n1794), .ZN(n1795) );
  IND2D1BWP12T U423 ( .A1(n3016), .B1(n4990), .ZN(n1911) );
  ND2D1BWP12T U424 ( .A1(n1812), .A2(n1811), .ZN(n416) );
  INVD1BWP12T U425 ( .I(n1790), .ZN(n1787) );
  INVD2BWP12T U426 ( .I(n1697), .ZN(n1695) );
  OR2XD2BWP12T U427 ( .A1(n2575), .A2(n1736), .Z(n1737) );
  TPOAI22D2BWP12T U428 ( .A1(n2530), .A2(n1786), .B1(n2532), .B2(n1691), .ZN(
        n1717) );
  ND2D1BWP12T U429 ( .A1(n1852), .A2(n1851), .ZN(n1853) );
  OAI22D1BWP12T U430 ( .A1(n2481), .A2(n2024), .B1(n1689), .B2(n1931), .ZN(
        n1949) );
  TPOAI22D1BWP12T U431 ( .A1(n2529), .A2(n1930), .B1(n2), .B2(n1954), .ZN(
        n1950) );
  CKND2D0BWP12T U432 ( .A1(n1883), .A2(n1882), .ZN(n1884) );
  TPOAI22D1BWP12T U433 ( .A1(n2120), .A2(n2519), .B1(n2016), .B2(n2015), .ZN(
        n2104) );
  XOR2D2BWP12T U434 ( .A1(n1812), .A2(b[16]), .Z(n1329) );
  ND2D1BWP12T U435 ( .A1(n1461), .A2(n1460), .ZN(n1462) );
  OAI22D1BWP12T U436 ( .A1(n2523), .A2(n1427), .B1(n2521), .B2(n872), .ZN(
        n1512) );
  INVD1BWP12T U437 ( .I(n908), .ZN(n910) );
  INVD2BWP12T U438 ( .I(n821), .ZN(n799) );
  INVD1BWP12T U439 ( .I(n2518), .ZN(n537) );
  ND2D1BWP12T U440 ( .A1(n1751), .A2(n1750), .ZN(n1752) );
  TPOAI21D1BWP12T U441 ( .A1(n1751), .A2(n1750), .B(n1749), .ZN(n1753) );
  INVD2BWP12T U442 ( .I(n1960), .ZN(n1965) );
  INVD2BWP12T U443 ( .I(n1216), .ZN(n1212) );
  TPND2D1BWP12T U444 ( .A1(n1434), .A2(n1433), .ZN(n1435) );
  INVD1BWP12T U445 ( .I(n1469), .ZN(n1434) );
  ND2D1BWP12T U446 ( .A1(n1440), .A2(n1439), .ZN(n1441) );
  TPND2D1BWP12T U447 ( .A1(n731), .A2(n730), .ZN(n834) );
  ND2D1BWP12T U448 ( .A1(n880), .A2(n879), .ZN(n826) );
  ND2D1BWP12T U449 ( .A1(n868), .A2(n869), .ZN(n814) );
  INVD2BWP12T U450 ( .I(n655), .ZN(n657) );
  INVD2BWP12T U451 ( .I(n1981), .ZN(n1934) );
  ND2D1BWP12T U452 ( .A1(n2562), .A2(n2561), .ZN(n2563) );
  IOA21D1BWP12T U453 ( .A1(n2061), .A2(n2060), .B(n2059), .ZN(n2509) );
  OAI21D0BWP12T U454 ( .A1(n2061), .A2(n2060), .B(n2058), .ZN(n2059) );
  INVD1BWP12T U455 ( .I(n1162), .ZN(n1158) );
  TPNR2D1BWP12T U456 ( .A1(n1239), .A2(n1238), .ZN(n1241) );
  TPND2D1BWP12T U457 ( .A1(n1287), .A2(n1286), .ZN(n1393) );
  ND2D1BWP12T U458 ( .A1(n1283), .A2(n1282), .ZN(n1287) );
  RCOAI21D1BWP12T U459 ( .A1(n1345), .A2(n1344), .B(n1343), .ZN(n1389) );
  ND2D1BWP12T U460 ( .A1(n1366), .A2(n1365), .ZN(n1323) );
  OAI22D1BWP12T U461 ( .A1(n1689), .A2(n1487), .B1(n2481), .B2(n1506), .ZN(
        n1507) );
  TPNR2D1BWP12T U462 ( .A1(n1568), .A2(n1569), .ZN(n1566) );
  INVD2BWP12T U463 ( .I(n1634), .ZN(n1610) );
  INVD2BWP12T U464 ( .I(n1633), .ZN(n1618) );
  CKND2D2BWP12T U465 ( .A1(n896), .A2(n895), .ZN(n761) );
  INVD1BWP12T U466 ( .I(n3518), .ZN(n3487) );
  NR2D1BWP12T U467 ( .A1(n1024), .A2(n3015), .ZN(n984) );
  TPNR2D1BWP12T U468 ( .A1(n982), .A2(n1969), .ZN(n983) );
  XNR2XD2BWP12T U469 ( .A1(n5196), .A2(n436), .ZN(n949) );
  IOA21D1BWP12T U470 ( .A1(n699), .A2(n698), .B(n697), .ZN(n1725) );
  NR3D1BWP12T U471 ( .A1(n3021), .A2(n5221), .A3(n3020), .ZN(n3022) );
  TPND2D1BWP12T U472 ( .A1(n1986), .A2(n1985), .ZN(n1987) );
  INVD2BWP12T U473 ( .I(n1521), .ZN(n1388) );
  INVD2BWP12T U474 ( .I(n25), .ZN(n3641) );
  TPND2D3BWP12T U475 ( .A1(n1660), .A2(n1659), .ZN(n1666) );
  CKND2D2BWP12T U476 ( .A1(n1621), .A2(n917), .ZN(n919) );
  ND2D1BWP12T U477 ( .A1(n1840), .A2(n1836), .ZN(n1837) );
  XNR2XD2BWP12T U478 ( .A1(b[1]), .A2(n4501), .ZN(n933) );
  CKND2D0BWP12T U479 ( .A1(n1054), .A2(n1053), .ZN(n1055) );
  TPOAI22D1BWP12T U480 ( .A1(n3588), .A2(n3889), .B1(n3887), .B2(n3587), .ZN(
        n3518) );
  INVD1BWP12T U481 ( .I(n3782), .ZN(n2845) );
  INVD1BWP12T U482 ( .I(n1062), .ZN(n1019) );
  TPOAI22D2BWP12T U483 ( .A1(n1024), .A2(n1969), .B1(n1023), .B2(n3015), .ZN(
        n1035) );
  TPNR2D4BWP12T U484 ( .A1(n943), .A2(n2005), .ZN(n955) );
  ND2D1BWP12T U485 ( .A1(n2320), .A2(n2319), .ZN(n2324) );
  TPND2D2BWP12T U486 ( .A1(n853), .A2(n852), .ZN(n1673) );
  ND2D1BWP12T U487 ( .A1(n663), .A2(n660), .ZN(n530) );
  OAI21D1BWP12T U488 ( .A1(n663), .A2(n660), .B(n661), .ZN(n529) );
  AOI21D0BWP12T U489 ( .A1(n5153), .A2(n5148), .B(n5255), .ZN(n3916) );
  MUX2ND0BWP12T U490 ( .I0(n4943), .I1(n4568), .S(b[0]), .ZN(n4312) );
  OR2XD1BWP12T U491 ( .A1(n4990), .A2(n3668), .Z(n3294) );
  TPND2D3BWP12T U492 ( .A1(n1250), .A2(n1249), .ZN(n3064) );
  INVD2BWP12T U493 ( .I(n1304), .ZN(n1249) );
  TPND2D1BWP12T U494 ( .A1(n3062), .A2(n3064), .ZN(n3046) );
  ND2D1BWP12T U495 ( .A1(n1418), .A2(n1419), .ZN(n1407) );
  OAI22D0BWP12T U496 ( .A1(n3619), .A2(n3607), .B1(n3614), .B2(n3730), .ZN(
        n3695) );
  INVD1BWP12T U497 ( .I(n2242), .ZN(n3308) );
  ND2D1BWP12T U498 ( .A1(n1642), .A2(n1641), .ZN(n1647) );
  INVD1BWP12T U499 ( .I(b[22]), .ZN(n3637) );
  BUFFD2BWP12T U500 ( .I(n4500), .Z(n4672) );
  ND2D3BWP12T U501 ( .A1(n1667), .A2(n1666), .ZN(n3117) );
  CKND0BWP12T U502 ( .I(n3936), .ZN(n2355) );
  NR2D1BWP12T U503 ( .A1(n2975), .A2(n3779), .ZN(n3782) );
  TPND2D1BWP12T U504 ( .A1(n3710), .A2(n3709), .ZN(n5009) );
  TPOAI22D1BWP12T U505 ( .A1(n1969), .A2(n933), .B1(n930), .B2(n3015), .ZN(
        n932) );
  ND2D1BWP12T U506 ( .A1(n1079), .A2(n1073), .ZN(n447) );
  NR2D0BWP12T U507 ( .A1(n4920), .A2(b[22]), .ZN(n2326) );
  TPNR2D1BWP12T U508 ( .A1(n3160), .A2(n3159), .ZN(n3161) );
  NR3D1BWP12T U509 ( .A1(n3602), .A2(n3601), .A3(n3600), .ZN(n4861) );
  AOI31D0BWP12T U510 ( .A1(n3599), .A2(n3598), .A3(n3597), .B(n3948), .ZN(
        n3600) );
  AOI22D0BWP12T U511 ( .A1(n3596), .A2(n436), .B1(n3595), .B2(n4541), .ZN(
        n3597) );
  INVD3BWP12T U512 ( .I(n3082), .ZN(n3002) );
  TPND2D2BWP12T U513 ( .A1(n1665), .A2(n1664), .ZN(n3110) );
  INR3D0BWP12T U514 ( .A1(n2719), .B1(n2718), .B2(n2717), .ZN(n2725) );
  TPNR2D3BWP12T U515 ( .A1(n942), .A2(n941), .ZN(n2730) );
  TPND2D2BWP12T U516 ( .A1(n2943), .A2(n1048), .ZN(n2801) );
  TPNR2D2BWP12T U517 ( .A1(n2871), .A2(n2869), .ZN(n1048) );
  CKND2D0BWP12T U518 ( .A1(n1079), .A2(n1073), .ZN(n2802) );
  CKND2D2BWP12T U519 ( .A1(n507), .A2(n1906), .ZN(n500) );
  TPNR2D2BWP12T U520 ( .A1(n495), .A2(n3015), .ZN(n481) );
  XOR3D2BWP12T U521 ( .A1(n623), .A2(n622), .A3(n621), .Z(n653) );
  OAI22D1BWP12T U522 ( .A1(n2479), .A2(n756), .B1(n630), .B2(n2005), .ZN(n804)
         );
  CKND2D2BWP12T U523 ( .A1(n3134), .A2(n3130), .ZN(n3124) );
  INR2D1BWP12T U524 ( .A1(n3062), .B1(n3061), .ZN(n3055) );
  OAI21D1BWP12T U525 ( .A1(n53), .A2(n3008), .B(n3009), .ZN(n2628) );
  XOR2XD4BWP12T U526 ( .A1(n4565), .A2(a[18]), .Z(n508) );
  TPND2D1BWP12T U527 ( .A1(n559), .A2(n558), .ZN(n720) );
  ND2D1BWP12T U528 ( .A1(n569), .A2(n570), .ZN(n558) );
  INVD1BWP12T U529 ( .I(n746), .ZN(n572) );
  TPND2D2BWP12T U530 ( .A1(n484), .A2(n2220), .ZN(n403) );
  IND2D1BWP12T U531 ( .A1(b[0]), .B1(n5079), .ZN(n1107) );
  TPND2D1BWP12T U532 ( .A1(n2412), .A2(n2266), .ZN(n4965) );
  NR2D2BWP12T U533 ( .A1(n4873), .A2(n4872), .ZN(n4874) );
  TPND2D1BWP12T U534 ( .A1(n3021), .A2(n5292), .ZN(n2733) );
  IND3D4BWP12T U535 ( .A1(n5224), .B1(n5223), .B2(n5222), .ZN(result[2]) );
  ND2D1BWP12T U536 ( .A1(n5221), .A2(n5292), .ZN(n5222) );
  TPND2D1BWP12T U537 ( .A1(n5220), .A2(n5322), .ZN(n5223) );
  TPND2D1BWP12T U538 ( .A1(n5248), .A2(n5247), .ZN(n5249) );
  AOI211D1BWP12T U539 ( .A1(n5305), .A2(n3235), .B(n2938), .C(n2937), .ZN(
        n2939) );
  TPND2D1BWP12T U540 ( .A1(n3034), .A2(n5292), .ZN(n2989) );
  OAI22D1BWP12T U541 ( .A1(n2523), .A2(n692), .B1(n2521), .B2(n1683), .ZN(
        n1742) );
  OAI22D2BWP12T U542 ( .A1(n2523), .A2(n872), .B1(n2521), .B2(n812), .ZN(n867)
         );
  OAI22D1BWP12T U543 ( .A1(n2479), .A2(n1113), .B1(n1141), .B2(n2005), .ZN(
        n1130) );
  OAI21D2BWP12T U544 ( .A1(n420), .A2(n1112), .B(n1111), .ZN(n1129) );
  INVD3BWP12T U545 ( .I(n4970), .ZN(n5303) );
  TPND2D2BWP12T U546 ( .A1(n2412), .A2(n2345), .ZN(n5312) );
  INVD1BWP12T U547 ( .I(n5212), .ZN(n5327) );
  TPOAI22D1BWP12T U548 ( .A1(n397), .A2(n681), .B1(n680), .B2(n2519), .ZN(n688) );
  NR2D2BWP12T U549 ( .A1(n1799), .A2(n675), .ZN(n676) );
  TPOAI21D1BWP12T U550 ( .A1(n1125), .A2(n1124), .B(n1123), .ZN(n1127) );
  CKND2D0BWP12T U551 ( .A1(n3336), .A2(n3671), .ZN(n73) );
  MAOI22D1BWP12T U552 ( .A1(n3337), .A2(n73), .B1(n3337), .B2(n73), .ZN(n4854)
         );
  CKND0BWP12T U553 ( .I(n4826), .ZN(n74) );
  AOI221D0BWP12T U554 ( .A1(n5257), .A2(n4826), .B1(n5258), .B2(n74), .C(n5296), .ZN(n4823) );
  OAI22D0BWP12T U555 ( .A1(n3575), .A2(n3609), .B1(n3577), .B2(n3607), .ZN(n75) );
  IAO21D0BWP12T U556 ( .A1(n3574), .A2(n3618), .B(n75), .ZN(n76) );
  OAI211D1BWP12T U557 ( .A1(n3576), .A2(n3730), .B(n3882), .C(n76), .ZN(n3723)
         );
  OAI22D0BWP12T U558 ( .A1(n3589), .A2(n3895), .B1(n3591), .B2(n4578), .ZN(n77) );
  OAI22D1BWP12T U559 ( .A1(n3588), .A2(n5260), .B1(n3587), .B2(n4790), .ZN(n78) );
  NR2D1BWP12T U560 ( .A1(n77), .A2(n78), .ZN(n3513) );
  NR2D0BWP12T U561 ( .A1(n4313), .A2(n4308), .ZN(n79) );
  OAI22D0BWP12T U562 ( .A1(n4311), .A2(n4312), .B1(n4315), .B2(n4310), .ZN(n80) );
  AOI211D0BWP12T U563 ( .A1(n4990), .A2(n2839), .B(n79), .C(n80), .ZN(n81) );
  OAI222D0BWP12T U564 ( .A1(n5183), .A2(n81), .B1(n4271), .B2(n4817), .C1(
        n4815), .C2(n4238), .ZN(n5165) );
  NR2D0BWP12T U565 ( .A1(n5146), .A2(n4557), .ZN(n82) );
  IND4D1BWP12T U566 ( .A1(n4571), .B1(n4582), .B2(n82), .B3(n4559), .ZN(n83)
         );
  MAOI22D0BWP12T U567 ( .A1(n2615), .A2(n83), .B1(n2615), .B2(n83), .ZN(n5102)
         );
  MUX2ND0BWP12T U568 ( .I0(n4899), .I1(n3843), .S(n3905), .ZN(n84) );
  NR2D0BWP12T U569 ( .A1(n3844), .A2(n84), .ZN(n5253) );
  AOI21D0BWP12T U570 ( .A1(n4330), .A2(n4491), .B(n4332), .ZN(n85) );
  CKND2D0BWP12T U571 ( .A1(n4329), .A2(n4333), .ZN(n86) );
  MAOI22D0BWP12T U572 ( .A1(n85), .A2(n86), .B1(n85), .B2(n86), .ZN(n4787) );
  CKND2D0BWP12T U573 ( .A1(n3265), .A2(n3414), .ZN(n87) );
  IND2D1BWP12T U574 ( .A1(n3409), .B1(n3483), .ZN(n88) );
  AOI32D0BWP12T U575 ( .A1(n3412), .A2(n3410), .A3(n88), .B1(n3411), .B2(n3410), .ZN(n89) );
  MOAI22D0BWP12T U576 ( .A1(n87), .A2(n89), .B1(n87), .B2(n89), .ZN(n4629) );
  INVD1BWP12T U577 ( .I(n4096), .ZN(n90) );
  AOI21D0BWP12T U578 ( .A1(n4084), .A2(n90), .B(n4088), .ZN(n91) );
  MAOI22D0BWP12T U579 ( .A1(n91), .A2(n2866), .B1(n91), .B2(n2866), .ZN(n4098)
         );
  AOI21D0BWP12T U580 ( .A1(n3221), .A2(n3222), .B(n3220), .ZN(n92) );
  OAI21D1BWP12T U581 ( .A1(n3223), .A2(n92), .B(n3224), .ZN(n93) );
  CKND2D0BWP12T U582 ( .A1(n2633), .A2(n2632), .ZN(n94) );
  MOAI22D0BWP12T U583 ( .A1(n93), .A2(n94), .B1(n93), .B2(n94), .ZN(n3212) );
  OAI22D0BWP12T U584 ( .A1(n4997), .A2(n5271), .B1(n4996), .B2(n5232), .ZN(n95) );
  CKND0BWP12T U585 ( .I(n407), .ZN(n96) );
  AOI22D0BWP12T U586 ( .A1(n4989), .A2(n5297), .B1(n4998), .B2(n5281), .ZN(n97) );
  IOA22D0BWP12T U587 ( .B1(n407), .B2(n4994), .A1(n5161), .A2(n4995), .ZN(n98)
         );
  NR2D0BWP12T U588 ( .A1(n4990), .A2(n5255), .ZN(n99) );
  OAI32D0BWP12T U589 ( .A1(n98), .A2(n5296), .A3(n99), .B1(n31), .B2(n98), 
        .ZN(n100) );
  OAI211D1BWP12T U590 ( .A1(n5299), .A2(n96), .B(n97), .C(n100), .ZN(n101) );
  RCAOI211D1BWP12T U591 ( .A1(n5313), .A2(n4999), .B(n95), .C(n101), .ZN(n102)
         );
  IOA21D1BWP12T U592 ( .A1(n5000), .A2(n5303), .B(n102), .ZN(n103) );
  TPAOI21D1BWP12T U593 ( .A1(n5308), .A2(n5001), .B(n103), .ZN(n5004) );
  CKND2D0BWP12T U594 ( .A1(n4433), .A2(n4434), .ZN(n104) );
  MAOI22D0BWP12T U595 ( .A1(n4435), .A2(n104), .B1(n4435), .B2(n104), .ZN(
        n4843) );
  INR2D0BWP12T U596 ( .A1(n3596), .B1(n4541), .ZN(n3503) );
  CKND0BWP12T U597 ( .I(n3938), .ZN(n105) );
  AOI221D0BWP12T U598 ( .A1(n5257), .A2(n3938), .B1(n5258), .B2(n105), .C(
        n5296), .ZN(n2637) );
  CKND0BWP12T U599 ( .I(n4488), .ZN(n106) );
  AN3XD0BWP12T U600 ( .A1(n107), .A2(n4491), .A3(n4453), .Z(n108) );
  AOI211D1BWP12T U601 ( .A1(n4453), .A2(n106), .B(n4456), .C(n108), .ZN(n109)
         );
  CKND2D0BWP12T U602 ( .A1(n4455), .A2(n4454), .ZN(n110) );
  MAOI22D1BWP12T U603 ( .A1(n109), .A2(n110), .B1(n109), .B2(n110), .ZN(n4981)
         );
  CKND0BWP12T U604 ( .I(n4478), .ZN(n107) );
  INR3D0BWP12T U605 ( .A1(n4577), .B1(n4576), .B2(n5234), .ZN(n111) );
  MOAI22D0BWP12T U606 ( .A1(n5049), .A2(n111), .B1(n5049), .B2(n111), .ZN(
        n5059) );
  CKND0BWP12T U607 ( .I(n5163), .ZN(n112) );
  MAOI22D0BWP12T U608 ( .A1(n4297), .A2(n112), .B1(n4297), .B2(n4271), .ZN(
        n113) );
  OAI21D1BWP12T U609 ( .A1(n4299), .A2(n113), .B(n5276), .ZN(n5280) );
  CKND2D0BWP12T U610 ( .A1(n4013), .A2(n4103), .ZN(n114) );
  CKND2D0BWP12T U611 ( .A1(n4013), .A2(n4112), .ZN(n115) );
  OAI211D1BWP12T U612 ( .A1(n4116), .A2(n114), .B(n4012), .C(n115), .ZN(n116)
         );
  MOAI22D0BWP12T U613 ( .A1(n4353), .A2(n116), .B1(n4353), .B2(n116), .ZN(
        n4686) );
  CKND0BWP12T U614 ( .I(n3578), .ZN(n117) );
  OAI21D0BWP12T U615 ( .A1(n3838), .A2(n117), .B(n3844), .ZN(n118) );
  AOI21D1BWP12T U616 ( .A1(n3723), .A2(n118), .B(n5323), .ZN(n5078) );
  MOAI22D0BWP12T U617 ( .A1(n4508), .A2(n25), .B1(n4508), .B2(n25), .ZN(n119)
         );
  OAI22D1BWP12T U618 ( .A1(n51), .A2(n119), .B1(n2575), .B2(n2574), .ZN(n120)
         );
  MOAI22D0BWP12T U619 ( .A1(n4565), .A2(n5264), .B1(n4565), .B2(n5264), .ZN(
        n121) );
  OAI22D0BWP12T U620 ( .A1(n2573), .A2(n2572), .B1(n2571), .B2(n121), .ZN(n122) );
  MAOI22D0BWP12T U621 ( .A1(n120), .A2(n122), .B1(n120), .B2(n122), .ZN(n123)
         );
  MAOI22D0BWP12T U622 ( .A1(n2578), .A2(n123), .B1(n2578), .B2(n123), .ZN(
        n2579) );
  IND2D0BWP12T U623 ( .A1(n4061), .B1(n4062), .ZN(n4396) );
  OAI22D0BWP12T U624 ( .A1(n4225), .A2(n3871), .B1(n4182), .B2(n3872), .ZN(
        n124) );
  OAI22D1BWP12T U625 ( .A1(n3818), .A2(n3869), .B1(n4219), .B2(n3870), .ZN(
        n125) );
  NR2D1BWP12T U626 ( .A1(n124), .A2(n125), .ZN(n3862) );
  CKND0BWP12T U627 ( .I(n3579), .ZN(n126) );
  AOI21D0BWP12T U628 ( .A1(n3580), .A2(n126), .B(n4940), .ZN(n4614) );
  INR3D0BWP12T U629 ( .A1(n4577), .B1(n4576), .B2(n4575), .ZN(n127) );
  MOAI22D0BWP12T U630 ( .A1(n5256), .A2(n127), .B1(n5256), .B2(n127), .ZN(
        n5268) );
  CKND0BWP12T U631 ( .I(n32), .ZN(n128) );
  OAI221D0BWP12T U632 ( .A1(n32), .A2(n5295), .B1(n128), .B2(n5294), .C(n5254), 
        .ZN(n4767) );
  CKND0BWP12T U633 ( .I(n3723), .ZN(n129) );
  AOI21D0BWP12T U634 ( .A1(n3724), .A2(n4301), .B(n129), .ZN(n5073) );
  CKND2D0BWP12T U635 ( .A1(n4045), .A2(n4043), .ZN(n130) );
  MOAI22D0BWP12T U636 ( .A1(n4050), .A2(n130), .B1(n4050), .B2(n130), .ZN(
        n4055) );
  OAI211D0BWP12T U637 ( .A1(n4801), .A2(n5155), .B(n4800), .C(n4799), .ZN(n131) );
  OAI22D0BWP12T U638 ( .A1(n4804), .A2(n5104), .B1(n4803), .B2(n5312), .ZN(
        n132) );
  AOI211D1BWP12T U639 ( .A1(n4805), .A2(n5303), .B(n131), .C(n132), .ZN(n133)
         );
  IOA21D1BWP12T U640 ( .A1(n4787), .A2(n5313), .B(n133), .ZN(n4806) );
  OAI21D0BWP12T U641 ( .A1(n3996), .A2(n4333), .B(n3999), .ZN(n134) );
  AOI21D1BWP12T U642 ( .A1(n2281), .A2(n4332), .B(n134), .ZN(n4344) );
  OAI22D0BWP12T U643 ( .A1(n4311), .A2(n4227), .B1(n4309), .B2(n4234), .ZN(
        n135) );
  OAI22D0BWP12T U644 ( .A1(n4313), .A2(n4221), .B1(n4315), .B2(n4226), .ZN(
        n136) );
  NR2D1BWP12T U645 ( .A1(n135), .A2(n136), .ZN(n4813) );
  NR2D0BWP12T U646 ( .A1(n3780), .A2(n3872), .ZN(n137) );
  OAI22D1BWP12T U647 ( .A1(n3779), .A2(n3869), .B1(n3871), .B2(n3781), .ZN(
        n138) );
  AOI211D0BWP12T U648 ( .A1(n3782), .A2(n5196), .B(n137), .C(n138), .ZN(n4899)
         );
  ND2D1BWP12T U649 ( .A1(n2815), .A2(n2811), .ZN(n139) );
  OAI211D1BWP12T U650 ( .A1(n2154), .A2(n2961), .B(n2819), .C(n139), .ZN(n3243) );
  CKND0BWP12T U651 ( .I(n4944), .ZN(n140) );
  OAI32D0BWP12T U652 ( .A1(n140), .A2(n4943), .A3(n5255), .B1(n5254), .B2(n140), .ZN(n141) );
  AOI221D0BWP12T U653 ( .A1(n5257), .A2(n4944), .B1(n5258), .B2(n140), .C(
        n5296), .ZN(n142) );
  CKND0BWP12T U654 ( .I(n4943), .ZN(n143) );
  AOI22D0BWP12T U655 ( .A1(n4943), .A2(n142), .B1(n5299), .B2(n143), .ZN(n144)
         );
  AOI211D1BWP12T U656 ( .A1(n4945), .A2(n4974), .B(n141), .C(n144), .ZN(n4946)
         );
  NR4D0BWP12T U657 ( .A1(n5001), .A2(n5174), .A3(n4777), .A4(n4622), .ZN(n145)
         );
  AN4D0BWP12T U658 ( .A1(n3431), .A2(n3430), .A3(n3429), .A4(n3428), .Z(n146)
         );
  NR4D0BWP12T U659 ( .A1(n4963), .A2(n3446), .A3(n4645), .A4(n4983), .ZN(n147)
         );
  ND2D1BWP12T U660 ( .A1(n4127), .A2(n4126), .ZN(n148) );
  NR3D1BWP12T U661 ( .A1(n148), .A2(n4128), .A3(n4592), .ZN(n149) );
  MUX2ND0BWP12T U662 ( .I0(n4591), .I1(n4590), .S(n3015), .ZN(n150) );
  OAI211D1BWP12T U663 ( .A1(n4499), .A2(n4498), .B(n149), .C(n150), .ZN(n151)
         );
  AO31D1BWP12T U664 ( .A1(n145), .A2(n146), .A3(n147), .B(n151), .Z(n4593) );
  MOAI22D0BWP12T U665 ( .A1(n3887), .A2(n3650), .B1(n445), .B2(n3650), .ZN(
        n152) );
  OAI22D0BWP12T U666 ( .A1(n2530), .A2(n152), .B1(n2532), .B2(n2531), .ZN(
        n2537) );
  MOAI22D0BWP12T U667 ( .A1(n5108), .A2(n5196), .B1(n5108), .B2(n5196), .ZN(
        n153) );
  OAI22D1BWP12T U668 ( .A1(n2549), .A2(n2548), .B1(n2547), .B2(n153), .ZN(n154) );
  MOAI22D0BWP12T U669 ( .A1(n4990), .A2(n4301), .B1(n4990), .B2(n4301), .ZN(
        n155) );
  OAI22D0BWP12T U670 ( .A1(n155), .A2(n2017), .B1(n2545), .B2(n2546), .ZN(n156) );
  MOAI22D0BWP12T U671 ( .A1(n154), .A2(n156), .B1(n154), .B2(n156), .ZN(n2559)
         );
  CKND0BWP12T U672 ( .I(n3553), .ZN(n157) );
  INVD1BWP12T U673 ( .I(n2678), .ZN(n158) );
  AOI221D1BWP12T U674 ( .A1(n2779), .A2(n3553), .B1(n3564), .B2(n157), .C(n158), .ZN(n2772) );
  CKND0BWP12T U675 ( .I(n4309), .ZN(n159) );
  AOI22D0BWP12T U676 ( .A1(n2888), .A2(n4228), .B1(n4226), .B2(n159), .ZN(n160) );
  AOI22D0BWP12T U677 ( .A1(n4242), .A2(n4216), .B1(n4199), .B2(n4244), .ZN(
        n161) );
  ND2D1BWP12T U678 ( .A1(n160), .A2(n161), .ZN(n4296) );
  OAI22D0BWP12T U679 ( .A1(n3589), .A2(n5079), .B1(n5234), .B2(n3591), .ZN(
        n162) );
  OAI22D1BWP12T U680 ( .A1(n3588), .A2(n2848), .B1(n4502), .B2(n3587), .ZN(
        n163) );
  TPNR2D1BWP12T U681 ( .A1(n162), .A2(n163), .ZN(n3515) );
  CKND0BWP12T U682 ( .I(n4977), .ZN(n164) );
  AOI221D0BWP12T U683 ( .A1(n5257), .A2(n4977), .B1(n5258), .B2(n164), .C(
        n5296), .ZN(n4976) );
  CKND2D0BWP12T U684 ( .A1(n4301), .A2(n5156), .ZN(n165) );
  AOI31D1BWP12T U685 ( .A1(n3875), .A2(n3729), .A3(n165), .B(n5323), .ZN(n5272) );
  CKND0BWP12T U686 ( .I(n4266), .ZN(n166) );
  AOI22D0BWP12T U687 ( .A1(n4208), .A2(n166), .B1(n4268), .B2(n4267), .ZN(
        n4766) );
  IIND4D0BWP12T U688 ( .A1(n4576), .A2(n4575), .B1(n4577), .B2(n5260), .ZN(
        n167) );
  MAOI22D0BWP12T U689 ( .A1(n4508), .A2(n167), .B1(n4508), .B2(n167), .ZN(
        n4758) );
  AOI21D1BWP12T U690 ( .A1(n3401), .A2(n3483), .B(n3404), .ZN(n168) );
  CKND2D0BWP12T U691 ( .A1(n3392), .A2(n3390), .ZN(n169) );
  MAOI22D0BWP12T U692 ( .A1(n168), .A2(n169), .B1(n168), .B2(n169), .ZN(n4720)
         );
  CKND0BWP12T U693 ( .I(n4491), .ZN(n170) );
  OAI21D1BWP12T U694 ( .A1(n4354), .A2(n170), .B(n4357), .ZN(n171) );
  MOAI22D0BWP12T U695 ( .A1(n4353), .A2(n171), .B1(n4353), .B2(n171), .ZN(
        n4670) );
  INR2D0BWP12T U696 ( .A1(n3875), .B1(n4925), .ZN(n172) );
  OA21XD0BWP12T U697 ( .A1(n172), .A2(n5214), .B(n4285), .Z(n3720) );
  NR4D0BWP12T U698 ( .A1(n5061), .A2(n4752), .A3(n5251), .A4(n5141), .ZN(n173)
         );
  OR4XD1BWP12T U699 ( .A1(n3214), .A2(n3213), .A3(n3212), .A4(n4910), .Z(n174)
         );
  OR4XD1BWP12T U700 ( .A1(n4853), .A2(n5306), .A3(n5203), .A4(n174), .Z(n175)
         );
  NR4D0BWP12T U701 ( .A1(n3234), .A2(n4884), .A3(n5021), .A4(n175), .ZN(n176)
         );
  NR3D0BWP12T U702 ( .A1(n3235), .A2(n4665), .A3(n4984), .ZN(n177) );
  NR4D0BWP12T U703 ( .A1(n3253), .A2(n5226), .A3(n5097), .A4(n4779), .ZN(n178)
         );
  ND4D1BWP12T U704 ( .A1(n5204), .A2(n176), .A3(n177), .A4(n178), .ZN(n179) );
  OR4D0BWP12T U705 ( .A1(n4624), .A2(n5002), .A3(n4938), .A4(n3291), .Z(n180)
         );
  NR4D0BWP12T U706 ( .A1(n4641), .A2(n4669), .A3(n179), .A4(n180), .ZN(n181)
         );
  NR4D0BWP12T U707 ( .A1(n4808), .A2(n4839), .A3(n5175), .A4(n3315), .ZN(n182)
         );
  IND4D1BWP12T U708 ( .A1(n4693), .B1(n173), .B2(n181), .B3(n182), .ZN(n4594)
         );
  OAI21D0BWP12T U709 ( .A1(n2825), .A2(n5255), .B(n5254), .ZN(n183) );
  AOI211D0BWP12T U710 ( .A1(b[22]), .A2(n183), .B(n4636), .C(n5151), .ZN(n184)
         );
  OAI22D0BWP12T U711 ( .A1(n4890), .A2(n4924), .B1(n4634), .B2(n5155), .ZN(
        n185) );
  AOI21D0BWP12T U712 ( .A1(n5252), .A2(n4632), .B(n185), .ZN(n186) );
  AOI22D1BWP12T U713 ( .A1(n4631), .A2(n5313), .B1(n4630), .B2(n5303), .ZN(
        n187) );
  AOI22D0BWP12T U714 ( .A1(n4638), .A2(n5297), .B1(n5281), .B2(n4637), .ZN(
        n188) );
  ND4D1BWP12T U715 ( .A1(n184), .A2(n186), .A3(n187), .A4(n188), .ZN(n4639) );
  MOAI22D0BWP12T U716 ( .A1(n4914), .A2(n3939), .B1(n4914), .B2(n3939), .ZN(
        n189) );
  OAI22D0BWP12T U717 ( .A1(n2519), .A2(n189), .B1(n397), .B2(n2520), .ZN(n2525) );
  INR3D0BWP12T U718 ( .A1(n3539), .B1(n3517), .B2(n3948), .ZN(n3488) );
  AOI22D0BWP12T U719 ( .A1(n4139), .A2(n4242), .B1(n4137), .B2(n2888), .ZN(
        n190) );
  AOI22D0BWP12T U720 ( .A1(n4138), .A2(n2839), .B1(n3761), .B2(n4244), .ZN(
        n191) );
  TPND2D1BWP12T U721 ( .A1(n190), .A2(n191), .ZN(n4189) );
  OAI22D0BWP12T U722 ( .A1(n4215), .A2(n3872), .B1(n3780), .B2(n3871), .ZN(
        n192) );
  OAI22D0BWP12T U723 ( .A1(n3781), .A2(n3870), .B1(n2975), .B2(n3869), .ZN(
        n193) );
  NR2D1BWP12T U724 ( .A1(n192), .A2(n193), .ZN(n3860) );
  AOI21D1BWP12T U725 ( .A1(n3380), .A2(n3483), .B(n3382), .ZN(n194) );
  CKND2D0BWP12T U726 ( .A1(n3379), .A2(n3383), .ZN(n195) );
  MAOI22D0BWP12T U727 ( .A1(n194), .A2(n195), .B1(n194), .B2(n195), .ZN(n4786)
         );
  AOI21D0BWP12T U728 ( .A1(n4349), .A2(n4491), .B(n4352), .ZN(n196) );
  MAOI22D0BWP12T U729 ( .A1(n196), .A2(n4340), .B1(n196), .B2(n4340), .ZN(
        n4694) );
  CKND0BWP12T U730 ( .I(n4208), .ZN(n197) );
  AOI22D0BWP12T U731 ( .A1(n4299), .A2(n4275), .B1(n4297), .B2(n4278), .ZN(
        n198) );
  CKND0BWP12T U732 ( .I(n4298), .ZN(n199) );
  OAI211D1BWP12T U733 ( .A1(n4239), .A2(n197), .B(n198), .C(n199), .ZN(n4684)
         );
  CKND0BWP12T U734 ( .I(n4892), .ZN(n200) );
  OAI221D0BWP12T U735 ( .A1(n4892), .A2(n5295), .B1(n200), .B2(n5294), .C(
        n5254), .ZN(n4893) );
  AOI21D0BWP12T U736 ( .A1(n4660), .A2(n3875), .B(n5214), .ZN(n201) );
  NR2D1BWP12T U737 ( .A1(n2981), .A2(n201), .ZN(n3713) );
  INR3D0BWP12T U738 ( .A1(n3910), .B1(n4543), .B2(n4542), .ZN(n202) );
  MOAI22D0BWP12T U739 ( .A1(n3679), .A2(n202), .B1(n3679), .B2(n202), .ZN(
        n4535) );
  CKND0BWP12T U740 ( .I(n4116), .ZN(n203) );
  AOI21D1BWP12T U741 ( .A1(n3985), .A2(n203), .B(n3988), .ZN(n204) );
  MAOI22D0BWP12T U742 ( .A1(n204), .A2(n4457), .B1(n204), .B2(n4457), .ZN(
        n4952) );
  MOAI22D0BWP12T U743 ( .A1(n4568), .A2(n3937), .B1(n4568), .B2(n3937), .ZN(
        n205) );
  OAI22D0BWP12T U744 ( .A1(n2529), .A2(n2528), .B1(n23), .B2(n205), .ZN(n2538)
         );
  IND2D0BWP12T U745 ( .A1(n3973), .B1(n3980), .ZN(n206) );
  OAI211D1BWP12T U746 ( .A1(n3975), .A2(n2210), .B(n4480), .C(n206), .ZN(n3986) );
  IAO21D0BWP12T U747 ( .A1(n3549), .A2(n3905), .B(n3708), .ZN(n4678) );
  CKND2D0BWP12T U748 ( .A1(n3483), .A2(n3433), .ZN(n207) );
  AOI32D1BWP12T U749 ( .A1(n3480), .A2(n3432), .A3(n207), .B1(n3434), .B2(
        n3432), .ZN(n208) );
  MOAI22D0BWP12T U750 ( .A1(n3435), .A2(n208), .B1(n3435), .B2(n208), .ZN(
        n4645) );
  TPND2D1BWP12T U751 ( .A1(n5186), .A2(n5185), .ZN(n209) );
  NR3D1BWP12T U752 ( .A1(n209), .A2(n5211), .A3(n5312), .ZN(n5187) );
  OAI21D0BWP12T U753 ( .A1(n4096), .A2(n4095), .B(n4094), .ZN(n210) );
  CKND2D0BWP12T U754 ( .A1(n4388), .A2(n4097), .ZN(n211) );
  MOAI22D0BWP12T U755 ( .A1(n210), .A2(n211), .B1(n210), .B2(n211), .ZN(n5242)
         );
  CKND2D0BWP12T U756 ( .A1(n2945), .A2(n2636), .ZN(n212) );
  MAOI22D1BWP12T U757 ( .A1(n4408), .A2(n212), .B1(n4408), .B2(n212), .ZN(
        n4443) );
  CKND2D0BWP12T U758 ( .A1(n3217), .A2(n3215), .ZN(n213) );
  MOAI22D0BWP12T U759 ( .A1(n3222), .A2(n213), .B1(n3222), .B2(n213), .ZN(
        n3213) );
  CKND2D0BWP12T U760 ( .A1(n3875), .A2(n5127), .ZN(n214) );
  AO21D1BWP12T U761 ( .A1(n3844), .A2(n214), .B(n4288), .Z(n3737) );
  INR3D0BWP12T U762 ( .A1(n4582), .B1(n4571), .B2(n4570), .ZN(n215) );
  MOAI22D0BWP12T U763 ( .A1(n4943), .A2(n215), .B1(n4943), .B2(n215), .ZN(
        n4951) );
  CKND2D0BWP12T U764 ( .A1(n4455), .A2(n4453), .ZN(n216) );
  CKND0BWP12T U765 ( .I(n4491), .ZN(n217) );
  OAI32D0BWP12T U766 ( .A1(n216), .A2(n4478), .A3(n217), .B1(n4488), .B2(n216), 
        .ZN(n218) );
  AOI211D1BWP12T U767 ( .A1(n4455), .A2(n4456), .B(n218), .C(n2203), .ZN(n219)
         );
  MAOI22D0BWP12T U768 ( .A1(n4457), .A2(n219), .B1(n4457), .B2(n219), .ZN(
        n4937) );
  INR2D2BWP12T U769 ( .A1(n3013), .B1(n3014), .ZN(n220) );
  MAOI22D0BWP12T U770 ( .A1(n3019), .A2(n220), .B1(n3019), .B2(n220), .ZN(
        n5221) );
  AOI22D0BWP12T U771 ( .A1(n3545), .A2(n5322), .B1(n3253), .B2(n5305), .ZN(
        n221) );
  ND2D1BWP12T U772 ( .A1(n2867), .A2(n221), .ZN(n222) );
  AO211D4BWP12T U773 ( .A1(n3042), .A2(n5292), .B(n2868), .C(n222), .Z(
        result[10]) );
  OAI22D1BWP12T U774 ( .A1(n2545), .A2(n2085), .B1(n2546), .B2(n413), .ZN(
        n2552) );
  OAI21D0BWP12T U775 ( .A1(n4005), .A2(n3999), .B(n4342), .ZN(n223) );
  AOI21D1BWP12T U776 ( .A1(n4002), .A2(n2202), .B(n223), .ZN(n4011) );
  IOA21D1BWP12T U777 ( .A1(n5160), .A2(n3707), .B(n3698), .ZN(n3717) );
  OAI21D0BWP12T U778 ( .A1(n4091), .A2(n4085), .B(n4382), .ZN(n224) );
  RCAOI21D1BWP12T U779 ( .A1(n2196), .A2(n4088), .B(n224), .ZN(n4094) );
  NR2D1BWP12T U780 ( .A1(n4417), .A2(n225), .ZN(n226) );
  ND2D1BWP12T U781 ( .A1(n226), .A2(n4415), .ZN(n227) );
  OAI211D1BWP12T U782 ( .A1(n4416), .A2(n225), .B(n4422), .C(n227), .ZN(n228)
         );
  CKND0BWP12T U783 ( .I(n4175), .ZN(n229) );
  CKND2D0BWP12T U784 ( .A1(n5108), .A2(n3853), .ZN(n230) );
  OAI221D1BWP12T U785 ( .A1(n4175), .A2(n3537), .B1(n229), .B2(n4176), .C(n230), .ZN(n3547) );
  OAI22D0BWP12T U786 ( .A1(n4311), .A2(n3762), .B1(n4309), .B2(n4139), .ZN(
        n231) );
  OAI22D0BWP12T U787 ( .A1(n4313), .A2(n3761), .B1(n4315), .B2(n3760), .ZN(
        n232) );
  NR2D1BWP12T U788 ( .A1(n231), .A2(n232), .ZN(n4203) );
  AN3XD0BWP12T U789 ( .A1(n2612), .A2(n5105), .A3(n5203), .Z(n233) );
  CKND0BWP12T U790 ( .I(n5106), .ZN(n234) );
  AOI211D0BWP12T U791 ( .A1(n5107), .A2(n5108), .B(n233), .C(n234), .ZN(n5109)
         );
  CKND0BWP12T U792 ( .I(n3314), .ZN(n235) );
  AOI21D0BWP12T U793 ( .A1(n3311), .A2(n235), .B(n3313), .ZN(n236) );
  OAI21D1BWP12T U794 ( .A1(n236), .A2(n3310), .B(n3312), .ZN(n237) );
  CKND2D0BWP12T U795 ( .A1(n3379), .A2(n3383), .ZN(n238) );
  MOAI22D0BWP12T U796 ( .A1(n237), .A2(n238), .B1(n237), .B2(n238), .ZN(n4808)
         );
  OAI22D0BWP12T U797 ( .A1(n3587), .A2(n4916), .B1(n3589), .B2(n3887), .ZN(
        n240) );
  NR2D1BWP12T U798 ( .A1(n239), .A2(n240), .ZN(n3535) );
  CKND2D0BWP12T U799 ( .A1(n3890), .A2(n3889), .ZN(n241) );
  TPNR2D2BWP12T U800 ( .A1(n4580), .A2(n241), .ZN(n4572) );
  OAI21D0BWP12T U801 ( .A1(n4029), .A2(n4026), .B(n4393), .ZN(n242) );
  AOI21D1BWP12T U802 ( .A1(n2197), .A2(n4025), .B(n242), .ZN(n2198) );
  CKND0BWP12T U803 ( .I(n3279), .ZN(n243) );
  AOI21D1BWP12T U804 ( .A1(n3280), .A2(n3452), .B(n243), .ZN(n3283) );
  ND2D1BWP12T U805 ( .A1(n4434), .A2(n4433), .ZN(n244) );
  MAOI22D0BWP12T U806 ( .A1(n4059), .A2(n244), .B1(n4059), .B2(n244), .ZN(
        n4844) );
  AOI22D0BWP12T U807 ( .A1(n4301), .A2(n3831), .B1(n3795), .B2(n4178), .ZN(
        n245) );
  CKND2D0BWP12T U808 ( .A1(n3832), .A2(n3948), .ZN(n246) );
  ND3D0BWP12T U809 ( .A1(n246), .A2(n245), .A3(n3817), .ZN(n4680) );
  INVD1BWP12T U810 ( .I(n4366), .ZN(n247) );
  OA21D1BWP12T U811 ( .A1(n4361), .A2(n247), .B(n4080), .Z(n4104) );
  MOAI22D0BWP12T U812 ( .A1(n2418), .A2(n2703), .B1(n4541), .B2(n2272), .ZN(
        n4415) );
  AOI22D0BWP12T U813 ( .A1(n3853), .A2(n3762), .B1(n3852), .B2(n3761), .ZN(
        n248) );
  AOI22D0BWP12T U814 ( .A1(n3854), .A2(n4139), .B1(n3855), .B2(n4137), .ZN(
        n249) );
  ND2D1BWP12T U815 ( .A1(n248), .A2(n249), .ZN(n3768) );
  OA222D1BWP12T U816 ( .A1(n3619), .A2(n3609), .B1(n3620), .B2(n3607), .C1(
        n3618), .C2(n3614), .Z(n250) );
  OA211D1BWP12T U817 ( .A1(n3608), .A2(n3730), .B(n3882), .C(n250), .Z(n2920)
         );
  CKND0BWP12T U818 ( .I(n5235), .ZN(n251) );
  CKND0BWP12T U819 ( .I(n5237), .ZN(n252) );
  OAI221D0BWP12T U820 ( .A1(n5237), .A2(n5295), .B1(n252), .B2(n5294), .C(
        n5254), .ZN(n253) );
  OAI32D0BWP12T U821 ( .A1(n252), .A2(n5234), .A3(n5255), .B1(n5254), .B2(n252), .ZN(n254) );
  AO221D0BWP12T U822 ( .A1(n5235), .A2(n5236), .B1(n251), .B2(n253), .C(n254), 
        .Z(n5238) );
  OAI21D1BWP12T U823 ( .A1(n2863), .A2(n2927), .B(n4085), .ZN(n255) );
  TPAOI21D1BWP12T U824 ( .A1(n2274), .A2(n2924), .B(n255), .ZN(n4381) );
  CKND2D0BWP12T U825 ( .A1(n3848), .A2(n5181), .ZN(n256) );
  TPND3D1BWP12T U826 ( .A1(n256), .A2(n2666), .A3(n2665), .ZN(n257) );
  RCAOI211D1BWP12T U827 ( .A1(n5313), .A2(n4443), .B(n2667), .C(n257), .ZN(
        n2672) );
  NR2D0BWP12T U828 ( .A1(n4311), .A2(n4225), .ZN(n258) );
  OAI22D0BWP12T U829 ( .A1(n4315), .A2(n4219), .B1(n4313), .B2(n4182), .ZN(
        n259) );
  AOI211D0BWP12T U830 ( .A1(n2839), .A2(n4232), .B(n258), .C(n259), .ZN(n4294)
         );
  AO222D0BWP12T U831 ( .A1(n3855), .A2(n3794), .B1(n4165), .B2(n3852), .C1(
        n3853), .C2(n4164), .Z(n260) );
  AOI21D0BWP12T U832 ( .A1(n3854), .A2(n3793), .B(n260), .ZN(n261) );
  AOI21D0BWP12T U833 ( .A1(n3795), .A2(n3880), .B(n3838), .ZN(n262) );
  AOI22D1BWP12T U834 ( .A1(n3831), .A2(n4260), .B1(n3832), .B2(n4262), .ZN(
        n263) );
  OAI211D1BWP12T U835 ( .A1(n261), .A2(n4953), .B(n262), .C(n263), .ZN(n4996)
         );
  OAI222D0BWP12T U836 ( .A1(n4817), .A2(n4816), .B1(n5183), .B2(n4813), .C1(
        n4815), .C2(n4814), .ZN(n264) );
  AOI22D1BWP12T U837 ( .A1(n4818), .A2(n5303), .B1(n5281), .B2(n264), .ZN(
        n4834) );
  IND3D1BWP12T U838 ( .A1(n3298), .B1(n2605), .B2(n2603), .ZN(n265) );
  CKND0BWP12T U839 ( .I(n2604), .ZN(n266) );
  AOI21D0BWP12T U840 ( .A1(n2606), .A2(n2605), .B(n266), .ZN(n267) );
  ND2D1BWP12T U841 ( .A1(n2609), .A2(n2608), .ZN(n268) );
  AOI33D1BWP12T U842 ( .A1(n265), .A2(n5305), .A3(n267), .B1(n2607), .B2(n5308), .B3(n268), .ZN(n5107) );
  CKND0BWP12T U843 ( .I(n5033), .ZN(n269) );
  OAI32D0BWP12T U844 ( .A1(n269), .A2(n5030), .A3(n5255), .B1(n5254), .B2(n269), .ZN(n270) );
  AOI21D0BWP12T U845 ( .A1(n5031), .A2(n5254), .B(n5032), .ZN(n271) );
  AOI211D0BWP12T U846 ( .A1(n5032), .A2(n5236), .B(n270), .C(n271), .ZN(n272)
         );
  OAI21D0BWP12T U847 ( .A1(n5029), .A2(n5271), .B(n272), .ZN(n5038) );
  IOA21D1BWP12T U848 ( .A1(n3588), .A2(n5108), .B(n3727), .ZN(n3509) );
  OAI222D0BWP12T U849 ( .A1(n4311), .A2(n4137), .B1(n4313), .B2(n4138), .C1(
        n4315), .C2(n4139), .ZN(n273) );
  AO21D1BWP12T U850 ( .A1(n2839), .A2(n4140), .B(n273), .Z(n4253) );
  IAO21D0BWP12T U851 ( .A1(n2773), .A2(n21), .B(n3974), .ZN(n4475) );
  IOA21D0BWP12T U852 ( .A1(n3273), .A2(n3267), .B(n3272), .ZN(n274) );
  AOI21D1BWP12T U853 ( .A1(n2176), .A2(n3269), .B(n274), .ZN(n3285) );
  IND2D0BWP12T U854 ( .A1(n3594), .B1(n4501), .ZN(n3599) );
  IAO21D0BWP12T U855 ( .A1(n3649), .A2(n4508), .B(n2242), .ZN(n3380) );
  CKND0BWP12T U856 ( .I(n3595), .ZN(n275) );
  OAI22D0BWP12T U857 ( .A1(n3806), .A2(n436), .B1(n5030), .B2(n275), .ZN(n3502) );
  CKND2D0BWP12T U858 ( .A1(n5081), .A2(n3897), .ZN(n276) );
  NR2D1BWP12T U859 ( .A1(n4519), .A2(n276), .ZN(n4574) );
  CKND0BWP12T U860 ( .I(n4024), .ZN(n277) );
  CKND0BWP12T U861 ( .I(n4027), .ZN(n278) );
  CKND2D0BWP12T U862 ( .A1(n4023), .A2(n278), .ZN(n279) );
  IOA21D0BWP12T U863 ( .A1(n278), .A2(n4025), .B(n4026), .ZN(n280) );
  AOI31D0BWP12T U864 ( .A1(n4028), .A2(n4023), .A3(n278), .B(n280), .ZN(n281)
         );
  OAI31D0BWP12T U865 ( .A1(n4096), .A2(n277), .A3(n279), .B(n281), .ZN(n282)
         );
  MOAI22D0BWP12T U866 ( .A1(n4449), .A2(n282), .B1(n4449), .B2(n282), .ZN(
        n4761) );
  NR2D1BWP12T U867 ( .A1(n4541), .A2(n4543), .ZN(n283) );
  MOAI22D0BWP12T U868 ( .A1(n5030), .A2(n283), .B1(n5030), .B2(n283), .ZN(
        n5020) );
  OAI21D0BWP12T U869 ( .A1(n3579), .A2(n3882), .B(n3875), .ZN(n284) );
  OAI21D1BWP12T U870 ( .A1(n3732), .A2(n284), .B(n3565), .ZN(n5230) );
  OAI21D0BWP12T U871 ( .A1(n2818), .A2(n2885), .B(n2819), .ZN(n285) );
  AOI21D1BWP12T U872 ( .A1(n2233), .A2(n2882), .B(n285), .ZN(n3419) );
  CKND0BWP12T U873 ( .I(n4971), .ZN(n286) );
  CKND0BWP12T U874 ( .I(n4978), .ZN(n287) );
  CKND0BWP12T U875 ( .I(n4977), .ZN(n288) );
  OAI32D0BWP12T U876 ( .A1(n288), .A2(a[25]), .A3(n5255), .B1(n5254), .B2(n288), .ZN(n289) );
  MUX2ND0BWP12T U877 ( .I0(n4976), .I1(n5299), .S(n4975), .ZN(n290) );
  AO211D0BWP12T U878 ( .A1(n4974), .A2(n287), .B(n289), .C(n290), .Z(n291) );
  AOI22D1BWP12T U879 ( .A1(n5297), .A2(n4973), .B1(n4979), .B2(n4980), .ZN(
        n292) );
  IOA21D1BWP12T U880 ( .A1(n4972), .A2(n5252), .B(n292), .ZN(n293) );
  AOI211D1BWP12T U881 ( .A1(n5313), .A2(n4981), .B(n291), .C(n293), .ZN(n294)
         );
  AOI22D0BWP12T U882 ( .A1(n4982), .A2(n5281), .B1(n5308), .B2(n4983), .ZN(
        n295) );
  OAI211D1BWP12T U883 ( .A1(n4970), .A2(n286), .B(n294), .C(n295), .ZN(n296)
         );
  AO21D1BWP12T U884 ( .A1(n5305), .A2(n4984), .B(n296), .Z(n4985) );
  IND3D1BWP12T U885 ( .A1(op[3]), .B1(op[0]), .B2(n2353), .ZN(n2423) );
  IND2D0BWP12T U886 ( .A1(n3016), .B1(n4503), .ZN(n297) );
  TPOAI22D1BWP12T U887 ( .A1(n1868), .A2(n3914), .B1(n2462), .B2(n297), .ZN(
        n1776) );
  IND2D1BWP12T U888 ( .A1(n4356), .B1(n4355), .ZN(n4353) );
  RCIAO21D1BWP12T U889 ( .A1(n3527), .A2(n3618), .B(n4300), .ZN(n3704) );
  AOI21D0BWP12T U890 ( .A1(n3617), .A2(n5108), .B(n3625), .ZN(n298) );
  OAI21D1BWP12T U891 ( .A1(n2779), .A2(n3730), .B(n298), .ZN(n3578) );
  IOA21D1BWP12T U892 ( .A1(n3496), .A2(n5108), .B(n3537), .ZN(n4995) );
  OAI22D1BWP12T U893 ( .A1(n4311), .A2(n4198), .B1(n4309), .B2(n4216), .ZN(
        n299) );
  OAI22D0BWP12T U894 ( .A1(n4313), .A2(n4199), .B1(n4201), .B2(n4200), .ZN(
        n300) );
  NR2D1BWP12T U895 ( .A1(n299), .A2(n300), .ZN(n5163) );
  CKND2D0BWP12T U896 ( .A1(n4678), .A2(n4301), .ZN(n301) );
  AOI21D1BWP12T U897 ( .A1(n301), .A2(n5035), .B(n5323), .ZN(n5029) );
  ND2D1BWP12T U898 ( .A1(n4577), .A2(n4574), .ZN(n302) );
  MAOI22D0BWP12T U899 ( .A1(n5234), .A2(n302), .B1(n5234), .B2(n302), .ZN(
        n5231) );
  OAI32D0BWP12T U900 ( .A1(n3658), .A2(n4511), .A3(n5255), .B1(n5254), .B2(
        n3658), .ZN(n303) );
  INVD1BWP12T U901 ( .I(n2909), .ZN(n304) );
  AOI221D0BWP12T U902 ( .A1(n5257), .A2(n2909), .B1(n5258), .B2(n304), .C(
        n5296), .ZN(n305) );
  MUX2ND0BWP12T U903 ( .I0(n305), .I1(n5299), .S(n2910), .ZN(n306) );
  NR2D1BWP12T U904 ( .A1(n303), .A2(n306), .ZN(n2911) );
  CKND0BWP12T U905 ( .I(n3905), .ZN(n307) );
  OAI221D0BWP12T U906 ( .A1(n3905), .A2(n4144), .B1(n307), .B2(n3860), .C(
        n5214), .ZN(n3842) );
  NR2D0BWP12T U907 ( .A1(n4925), .A2(n5312), .ZN(n308) );
  OAI21D1BWP12T U908 ( .A1(n308), .A2(n5321), .B(n4285), .ZN(n2666) );
  NR2D0BWP12T U909 ( .A1(n4849), .A2(n2314), .ZN(n309) );
  TPND2D1BWP12T U910 ( .A1(n309), .A2(n3539), .ZN(n3806) );
  CKND2D0BWP12T U911 ( .A1(n3268), .A2(n3442), .ZN(n310) );
  CKND0BWP12T U912 ( .I(n3483), .ZN(n311) );
  OAI32D0BWP12T U913 ( .A1(n310), .A2(n3470), .A3(n311), .B1(n3480), .B2(n310), 
        .ZN(n312) );
  AOI211D1BWP12T U914 ( .A1(n3268), .A2(n3444), .B(n312), .C(n3267), .ZN(n313)
         );
  MAOI22D0BWP12T U915 ( .A1(n3445), .A2(n313), .B1(n3445), .B2(n313), .ZN(
        n4963) );
  CKND0BWP12T U916 ( .I(n4116), .ZN(n314) );
  AOI21D0BWP12T U917 ( .A1(n3985), .A2(n314), .B(n3988), .ZN(n315) );
  OAI32D1BWP12T U918 ( .A1(n2618), .A2(n2616), .A3(n315), .B1(n2619), .B2(
        n2618), .ZN(n316) );
  INR2D1BWP12T U919 ( .A1(n2617), .B1(n316), .ZN(n317) );
  IOA21D0BWP12T U920 ( .A1(n2622), .A2(n2621), .B(n2620), .ZN(n318) );
  AOI22D0BWP12T U921 ( .A1(n5303), .A2(n317), .B1(n5313), .B2(n318), .ZN(n2623) );
  NR2D0BWP12T U922 ( .A1(n3648), .A2(n4788), .ZN(n319) );
  NR2D0BWP12T U923 ( .A1(n3310), .A2(n319), .ZN(n320) );
  CKND0BWP12T U924 ( .I(n3314), .ZN(n321) );
  ND2D1BWP12T U925 ( .A1(n3313), .A2(n320), .ZN(n322) );
  OAI211D1BWP12T U926 ( .A1(n3312), .A2(n319), .B(n3383), .C(n322), .ZN(n323)
         );
  AOI31D1BWP12T U927 ( .A1(n3311), .A2(n320), .A3(n321), .B(n323), .ZN(n324)
         );
  MAOI22D0BWP12T U928 ( .A1(n324), .A2(n3388), .B1(n324), .B2(n3388), .ZN(
        n4752) );
  AOI21D1BWP12T U929 ( .A1(n4659), .A2(n5252), .B(n4658), .ZN(n325) );
  AOI22D1BWP12T U930 ( .A1(n4821), .A2(n4660), .B1(n5303), .B2(n4662), .ZN(
        n326) );
  CKND2D0BWP12T U931 ( .A1(n5313), .A2(n4663), .ZN(n327) );
  ND4D1BWP12T U932 ( .A1(n325), .A2(n4661), .A3(n326), .A4(n327), .ZN(n328) );
  AO21D1BWP12T U933 ( .A1(n4645), .A2(n5308), .B(n328), .Z(n4664) );
  OAI22D1BWP12T U934 ( .A1(n2464), .A2(n2114), .B1(n2462), .B2(n2463), .ZN(
        n2555) );
  CKND2D0BWP12T U935 ( .A1(n2703), .A2(n2691), .ZN(n329) );
  MOAI22D0BWP12T U936 ( .A1(n4421), .A2(n329), .B1(n4421), .B2(n329), .ZN(
        n4426) );
  IND2D0BWP12T U937 ( .A1(n2947), .B1(n2948), .ZN(n2953) );
  IAO21D0BWP12T U938 ( .A1(b[0]), .A2(n4501), .B(n5290), .ZN(n4133) );
  IND2D1BWP12T U939 ( .A1(n4990), .B1(n4607), .ZN(n4557) );
  AO211D0BWP12T U940 ( .A1(n4301), .A2(n4890), .B(n3838), .C(n4287), .Z(n4882)
         );
  AOI21D1BWP12T U941 ( .A1(n4045), .A2(n4050), .B(n4044), .ZN(n330) );
  CKND2D0BWP12T U942 ( .A1(n4047), .A2(n4416), .ZN(n331) );
  MAOI22D0BWP12T U943 ( .A1(n330), .A2(n331), .B1(n330), .B2(n331), .ZN(n5011)
         );
  IOA21D0BWP12T U944 ( .A1(n3492), .A2(n3703), .B(n3704), .ZN(n3544) );
  AOI21D0BWP12T U945 ( .A1(n4978), .A2(n4301), .B(n2920), .ZN(n332) );
  AOI21D1BWP12T U946 ( .A1(n4174), .A2(n4281), .B(n332), .ZN(n4323) );
  CKND0BWP12T U947 ( .I(n3311), .ZN(n333) );
  NR3D0BWP12T U948 ( .A1(n3260), .A2(n334), .A3(n3259), .ZN(n335) );
  CKND0BWP12T U949 ( .I(n335), .ZN(n336) );
  CKND0BWP12T U950 ( .I(n3263), .ZN(n334) );
  OAI32D0BWP12T U951 ( .A1(n334), .A2(n3259), .A3(n3264), .B1(n3261), .B2(n334), .ZN(n337) );
  AOI211D0BWP12T U952 ( .A1(n335), .A2(n3313), .B(n3262), .C(n337), .ZN(n338)
         );
  OAI31D0BWP12T U953 ( .A1(n3314), .A2(n333), .A3(n336), .B(n338), .ZN(n339)
         );
  CKND2D0BWP12T U954 ( .A1(n3265), .A2(n3414), .ZN(n340) );
  MOAI22D0BWP12T U955 ( .A1(n339), .A2(n340), .B1(n339), .B2(n340), .ZN(n4641)
         );
  CKND2D0BWP12T U956 ( .A1(n2958), .A2(n2633), .ZN(n341) );
  MAOI22D0BWP12T U957 ( .A1(n3421), .A2(n341), .B1(n3421), .B2(n341), .ZN(
        n3355) );
  AN3XD0BWP12T U958 ( .A1(op[1]), .A2(op[2]), .A3(n2351), .Z(n5236) );
  MOAI22D0BWP12T U959 ( .A1(n5030), .A2(n22), .B1(n5030), .B2(n22), .ZN(n342)
         );
  OAI22D0BWP12T U960 ( .A1(n52), .A2(n2478), .B1(n2477), .B2(n342), .ZN(n2484)
         );
  MOAI22D0BWP12T U961 ( .A1(n4788), .A2(n4826), .B1(n4788), .B2(n4826), .ZN(
        n343) );
  OAI22D0BWP12T U962 ( .A1(n2516), .A2(n343), .B1(n2518), .B2(n2517), .ZN(
        n2526) );
  OAI22D0BWP12T U963 ( .A1(n4315), .A2(n4131), .B1(n4313), .B2(n4130), .ZN(
        n344) );
  OAI22D0BWP12T U964 ( .A1(n4311), .A2(n4153), .B1(n4309), .B2(n4129), .ZN(
        n345) );
  NR2D1BWP12T U965 ( .A1(n344), .A2(n345), .ZN(n4239) );
  OAI21D0BWP12T U966 ( .A1(b[0]), .A2(n1812), .B(n1969), .ZN(n3017) );
  CKND2D0BWP12T U967 ( .A1(n4430), .A2(n4429), .ZN(n346) );
  MAOI22D0BWP12T U968 ( .A1(n4057), .A2(n346), .B1(n4057), .B2(n346), .ZN(
        n5198) );
  OAI21D0BWP12T U969 ( .A1(n5196), .A2(n4200), .B(n3872), .ZN(n347) );
  ND2D1BWP12T U970 ( .A1(n347), .A2(n2845), .ZN(n3821) );
  INR3D0BWP12T U971 ( .A1(n7), .B1(n2773), .B2(n4570), .ZN(n4559) );
  MAOI22D0BWP12T U972 ( .A1(n3293), .A2(n3300), .B1(n2177), .B2(n3283), .ZN(
        n348) );
  OAI211D1BWP12T U973 ( .A1(n3285), .A2(n2178), .B(n348), .C(n3299), .ZN(n2606) );
  CKND0BWP12T U974 ( .I(n4403), .ZN(n349) );
  CKND0BWP12T U975 ( .I(n4406), .ZN(n350) );
  CKND2D0BWP12T U976 ( .A1(n4402), .A2(n350), .ZN(n351) );
  IOA21D0BWP12T U977 ( .A1(n350), .A2(n4404), .B(n4405), .ZN(n352) );
  AOI31D1BWP12T U978 ( .A1(n4402), .A2(n4407), .A3(n350), .B(n352), .ZN(n353)
         );
  OAI31D1BWP12T U979 ( .A1(n4408), .A2(n349), .A3(n351), .B(n353), .ZN(n354)
         );
  MOAI22D0BWP12T U980 ( .A1(n4409), .A2(n354), .B1(n4409), .B2(n354), .ZN(
        n5270) );
  CKND0BWP12T U981 ( .I(b[22]), .ZN(n355) );
  AOI221D0BWP12T U982 ( .A1(n5257), .A2(b[22]), .B1(n5258), .B2(n355), .C(
        n5296), .ZN(n356) );
  MUX2ND0BWP12T U983 ( .I0(n356), .I1(n5299), .S(n4635), .ZN(n4636) );
  AOI21D0BWP12T U984 ( .A1(n3342), .A2(n3350), .B(n3344), .ZN(n357) );
  RCIAO22D1BWP12T U985 ( .B1(n357), .B2(n3341), .A1(n357), .A2(n3341), .ZN(
        n5014) );
  CKND2D0BWP12T U986 ( .A1(n4577), .A2(n3900), .ZN(n358) );
  MAOI22D0BWP12T U987 ( .A1(n2153), .A2(n358), .B1(n2153), .B2(n358), .ZN(
        n4524) );
  CKND0BWP12T U988 ( .I(n3778), .ZN(n359) );
  MAOI22D0BWP12T U989 ( .A1(n5181), .A2(n359), .B1(n4202), .B2(n5017), .ZN(
        n461) );
  NR2D0BWP12T U990 ( .A1(n3535), .A2(n3607), .ZN(n360) );
  OAI22D1BWP12T U991 ( .A1(n3558), .A2(n3730), .B1(n3731), .B2(n3609), .ZN(
        n361) );
  AOI211D0BWP12T U992 ( .A1(n3707), .A2(n3536), .B(n360), .C(n361), .ZN(n4819)
         );
  OAI21D0BWP12T U993 ( .A1(n2103), .A2(n2104), .B(n2102), .ZN(n2106) );
  MOAI22D0BWP12T U994 ( .A1(n2773), .A2(n4896), .B1(n2773), .B2(n4896), .ZN(
        n362) );
  OAI22D1BWP12T U995 ( .A1(n2462), .A2(n362), .B1(n2464), .B2(n2463), .ZN(
        n2474) );
  MOAI22D0BWP12T U996 ( .A1(n5049), .A2(n26), .B1(n5049), .B2(n26), .ZN(n363)
         );
  OAI22D0BWP12T U997 ( .A1(n29), .A2(n2534), .B1(n2533), .B2(n363), .ZN(n2536)
         );
  IND2XD2BWP12T U998 ( .A1(n3588), .B1(n2825), .ZN(n3511) );
  IAO21D0BWP12T U999 ( .A1(n2250), .A2(n4568), .B(n2251), .ZN(n2253) );
  AOI222D0BWP12T U1000 ( .A1(n4301), .A2(n3790), .B1(n3948), .B2(n3827), .C1(
        n4178), .C2(n3789), .ZN(n364) );
  IND2D1BWP12T U1001 ( .A1(n3849), .B1(n364), .ZN(n5116) );
  CKND0BWP12T U1002 ( .I(n5196), .ZN(n365) );
  OAI221D0BWP12T U1003 ( .A1(n5196), .A2(n3574), .B1(n365), .B2(n3575), .C(
        n3905), .ZN(n2721) );
  INVD1BWP12T U1004 ( .I(n3362), .ZN(n366) );
  TPAOI21D1BWP12T U1005 ( .A1(n3241), .A2(n3246), .B(n366), .ZN(n3167) );
  OR4XD1BWP12T U1006 ( .A1(n5085), .A2(n5054), .A3(n3939), .A4(n5237), .Z(
        n2334) );
  IOA21D0BWP12T U1007 ( .A1(n3547), .A2(n3905), .B(n4657), .ZN(n4980) );
  CKND0BWP12T U1008 ( .I(n3948), .ZN(n367) );
  OAI221D0BWP12T U1009 ( .A1(n3948), .A2(n3846), .B1(n367), .B2(n3848), .C(
        n5214), .ZN(n4772) );
  CKND0BWP12T U1010 ( .I(n3937), .ZN(n368) );
  OAI221D0BWP12T U1011 ( .A1(n3937), .A2(n5295), .B1(n368), .B2(n5294), .C(
        n5254), .ZN(n2965) );
  OAI22D0BWP12T U1012 ( .A1(n4311), .A2(n4237), .B1(n4309), .B2(n4184), .ZN(
        n369) );
  OAI22D0BWP12T U1013 ( .A1(n4313), .A2(n4183), .B1(n4315), .B2(n4220), .ZN(
        n370) );
  OAI21D0BWP12T U1014 ( .A1(n369), .A2(n370), .B(n4208), .ZN(n371) );
  OAI211D0BWP12T U1015 ( .A1(n4294), .A2(n4815), .B(n4185), .C(n371), .ZN(n372) );
  AOI21D1BWP12T U1016 ( .A1(n4299), .A2(n4195), .B(n372), .ZN(n4956) );
  NR2D0BWP12T U1017 ( .A1(n5103), .A2(n5102), .ZN(n373) );
  AOI211D0BWP12T U1018 ( .A1(n5103), .A2(n5102), .B(n5104), .C(n373), .ZN(
        n5110) );
  NR2D0BWP12T U1019 ( .A1(n4683), .A2(n4682), .ZN(n374) );
  CKND2D0BWP12T U1020 ( .A1(n4685), .A2(n5297), .ZN(n375) );
  OAI211D1BWP12T U1021 ( .A1(n5312), .A2(n4684), .B(n374), .C(n375), .ZN(n376)
         );
  RCAOI21D1BWP12T U1022 ( .A1(n5313), .A2(n4670), .B(n376), .ZN(n377) );
  IOA21D1BWP12T U1023 ( .A1(n5303), .A2(n4686), .B(n377), .ZN(n378) );
  TPAOI21D1BWP12T U1024 ( .A1(n4687), .A2(n5308), .B(n378), .ZN(n4688) );
  OAI21D0BWP12T U1025 ( .A1(n3298), .A2(n3201), .B(n3210), .ZN(n379) );
  MOAI22D0BWP12T U1026 ( .A1(n3435), .A2(n379), .B1(n3435), .B2(n379), .ZN(
        n4665) );
  MAOI22D1BWP12T U1027 ( .A1(n5212), .A2(n3720), .B1(n3586), .B2(n5271), .ZN(
        n2671) );
  OAI22D0BWP12T U1028 ( .A1(n3589), .A2(n4790), .B1(n3588), .B2(n4578), .ZN(
        n380) );
  OAI22D0BWP12T U1029 ( .A1(n3587), .A2(n3890), .B1(n3591), .B2(n3889), .ZN(
        n381) );
  TPNR2D1BWP12T U1030 ( .A1(n380), .A2(n381), .ZN(n3558) );
  AOI222D0BWP12T U1031 ( .A1(n4501), .A2(n3569), .B1(n3570), .B2(n3595), .C1(
        n3596), .C2(n5192), .ZN(n382) );
  CKND0BWP12T U1032 ( .I(n3607), .ZN(n383) );
  CKND0BWP12T U1033 ( .I(n3707), .ZN(n384) );
  OAI22D1BWP12T U1034 ( .A1(n3573), .A2(n3609), .B1(n3568), .B2(n384), .ZN(
        n385) );
  AOI211D1BWP12T U1035 ( .A1(n3572), .A2(n383), .B(n3774), .C(n385), .ZN(n386)
         );
  OAI21D0BWP12T U1036 ( .A1(n3948), .A2(n382), .B(n386), .ZN(n5320) );
  AN2D0BWP12T U1037 ( .A1(n1550), .A2(n1549), .Z(n1548) );
  MOAI22D0BWP12T U1038 ( .A1(n4510), .A2(n4944), .B1(n4510), .B2(n4944), .ZN(
        n387) );
  OAI22D0BWP12T U1039 ( .A1(n2471), .A2(n2470), .B1(n2469), .B2(n387), .ZN(
        n2472) );
  MOAI22D0BWP12T U1040 ( .A1(n436), .A2(n5153), .B1(n436), .B2(n5153), .ZN(
        n388) );
  OAI22D0BWP12T U1041 ( .A1(n2523), .A2(n2522), .B1(n561), .B2(n388), .ZN(
        n2524) );
  CKND0BWP12T U1042 ( .I(n2129), .ZN(n2130) );
  IAO21D0BWP12T U1043 ( .A1(n3669), .A2(n2773), .B(n2254), .ZN(n3467) );
  IND4D0BWP12T U1044 ( .A1(n4529), .B1(n4635), .B2(n4916), .B3(n4572), .ZN(
        n4571) );
  IAO21D0BWP12T U1045 ( .A1(n3018), .A2(n3017), .B(n3019), .ZN(n4859) );
  IAO21D0BWP12T U1046 ( .A1(n2234), .A2(n4521), .B(n3361), .ZN(n3367) );
  CKND0BWP12T U1047 ( .I(n2849), .ZN(n389) );
  CKND0BWP12T U1048 ( .I(n3939), .ZN(n390) );
  OAI221D0BWP12T U1049 ( .A1(n3939), .A2(n5295), .B1(n390), .B2(n5294), .C(
        n5254), .ZN(n391) );
  OAI32D0BWP12T U1050 ( .A1(n390), .A2(n2848), .A3(n5255), .B1(n5254), .B2(
        n390), .ZN(n392) );
  AOI221D0BWP12T U1051 ( .A1(n5236), .A2(n389), .B1(n391), .B2(n2849), .C(n392), .ZN(n2850) );
  OAI21D0BWP12T U1052 ( .A1(n3421), .A2(n2959), .B(n2958), .ZN(n393) );
  CKND2D0BWP12T U1053 ( .A1(n2961), .A2(n2962), .ZN(n394) );
  MOAI22D0BWP12T U1054 ( .A1(n393), .A2(n394), .B1(n393), .B2(n394), .ZN(n3427) );
  IND2D0BWP12T U1055 ( .A1(n2184), .B1(n2351), .ZN(n4970) );
  TPND2D1BWP12T U1056 ( .A1(n822), .A2(n821), .ZN(n800) );
  TPND2D2BWP12T U1057 ( .A1(n1218), .A2(n1217), .ZN(n1219) );
  DCCKND4BWP12T U1058 ( .I(n750), .ZN(n894) );
  FA1D2BWP12T U1059 ( .A(n749), .B(n748), .CI(n747), .CO(n793), .S(n750) );
  XNR2D2BWP12T U1060 ( .A1(n4301), .A2(n4565), .ZN(n736) );
  INVD3BWP12T U1061 ( .I(n1268), .ZN(n395) );
  INVD4BWP12T U1062 ( .I(n395), .ZN(n396) );
  XNR2D2BWP12T U1063 ( .A1(n2123), .A2(n4770), .ZN(n757) );
  TPOAI22D2BWP12T U1064 ( .A1(n2518), .A2(n589), .B1(n2516), .B2(n588), .ZN(
        n634) );
  XNR2D2BWP12T U1065 ( .A1(n3899), .A2(n2014), .ZN(n2120) );
  XNR2D2BWP12T U1066 ( .A1(n2014), .A2(n3938), .ZN(n2015) );
  XNR2XD2BWP12T U1067 ( .A1(n48), .A2(n5196), .ZN(n1387) );
  OAI22D2BWP12T U1068 ( .A1(n2518), .A2(n865), .B1(n823), .B2(n2022), .ZN(n879) );
  INR2XD2BWP12T U1069 ( .A1(n3016), .B1(n2022), .ZN(n1335) );
  ND2D4BWP12T U1070 ( .A1(n2017), .A2(n2255), .ZN(n1912) );
  TPND2D1BWP12T U1071 ( .A1(n647), .A2(n781), .ZN(n648) );
  XOR2XD2BWP12T U1072 ( .A1(n1812), .A2(n4991), .Z(n1970) );
  TPND2D3BWP12T U1073 ( .A1(n1003), .A2(n1001), .ZN(n2627) );
  NR4D1BWP12T U1074 ( .A1(n3070), .A2(n4755), .A3(n3069), .A4(n5288), .ZN(
        n3071) );
  TPOAI21D1BWP12T U1075 ( .A1(n4381), .A2(n2278), .B(n2277), .ZN(n2279) );
  INVD4BWP12T U1076 ( .I(n2753), .ZN(n4491) );
  TPAOI21D2BWP12T U1077 ( .A1(n2635), .A2(n2280), .B(n2279), .ZN(n2753) );
  XOR3D2BWP12T U1078 ( .A1(n2485), .A2(n2484), .A3(n2483), .Z(n2490) );
  BUFFD8BWP12T U1079 ( .I(n2014), .Z(n4914) );
  ND2XD4BWP12T U1080 ( .A1(n469), .A2(n1869), .ZN(n397) );
  XOR3XD4BWP12T U1081 ( .A1(n1791), .A2(n1790), .A3(n1789), .Z(n398) );
  NR2XD1BWP12T U1082 ( .A1(n1887), .A2(n1886), .ZN(n1890) );
  CKND2D2BWP12T U1083 ( .A1(n1887), .A2(n1886), .ZN(n1888) );
  XOR3XD4BWP12T U1084 ( .A1(n1905), .A2(n1904), .A3(n1903), .Z(n1878) );
  ND2D1BWP12T U1085 ( .A1(n1905), .A2(n1903), .ZN(n400) );
  ND2D1BWP12T U1086 ( .A1(n1904), .A2(n1903), .ZN(n401) );
  ND3XD3BWP12T U1087 ( .A1(n399), .A2(n400), .A3(n401), .ZN(n1961) );
  TPNR2D2BWP12T U1088 ( .A1(n1962), .A2(n1961), .ZN(n1964) );
  TPND2D2BWP12T U1089 ( .A1(n1962), .A2(n1961), .ZN(n1963) );
  BUFFD2BWP12T U1090 ( .I(result[31]), .Z(n) );
  TPND2D1BWP12T U1091 ( .A1(n2084), .A2(n2083), .ZN(n2499) );
  OAI22D1BWP12T U1092 ( .A1(n2020), .A2(n1102), .B1(n14), .B2(n1143), .ZN(n459) );
  TPNR2D3BWP12T U1093 ( .A1(n1663), .A2(n1662), .ZN(n2991) );
  TPND2D3BWP12T U1094 ( .A1(n1594), .A2(n1593), .ZN(n3082) );
  TPND2D2BWP12T U1095 ( .A1(n1481), .A2(n1480), .ZN(n419) );
  CKND2D2BWP12T U1096 ( .A1(n1481), .A2(n1480), .ZN(n1519) );
  AN2XD2BWP12T U1097 ( .A1(n921), .A2(n922), .Z(n844) );
  CKND2D2BWP12T U1098 ( .A1(n4692), .A2(n5292), .ZN(n4724) );
  TPND2D2BWP12T U1099 ( .A1(n1002), .A2(n2627), .ZN(n1006) );
  DCCKND12BWP12T U1100 ( .I(n3838), .ZN(n3875) );
  NR2D2BWP12T U1101 ( .A1(n2331), .A2(n2330), .ZN(n2337) );
  NR3XD3BWP12T U1102 ( .A1(n2325), .A2(n2324), .A3(n2323), .ZN(n2338) );
  ND2D3BWP12T U1103 ( .A1(n1672), .A2(n1671), .ZN(n3131) );
  XNR2XD2BWP12T U1104 ( .A1(n2123), .A2(n5054), .ZN(n884) );
  XNR2XD2BWP12T U1105 ( .A1(n2123), .A2(b[22]), .ZN(n1871) );
  XNR2D2BWP12T U1106 ( .A1(n3948), .A2(n2123), .ZN(n1051) );
  TPND2D3BWP12T U1107 ( .A1(n1308), .A2(n1307), .ZN(n3051) );
  NR2XD3BWP12T U1108 ( .A1(n1308), .A2(n1307), .ZN(n3050) );
  INVD3BWP12T U1109 ( .I(n2314), .ZN(n402) );
  INVD2BWP12T U1110 ( .I(b[0]), .ZN(n2314) );
  CKND2D2BWP12T U1111 ( .A1(n1315), .A2(n5030), .ZN(n951) );
  XOR2XD2BWP12T U1112 ( .A1(n3930), .A2(n1812), .Z(n1021) );
  ND2XD4BWP12T U1113 ( .A1(n1838), .A2(n1837), .ZN(n3097) );
  TPNR2D3BWP12T U1114 ( .A1(n1207), .A2(n1208), .ZN(n1209) );
  INVD8BWP12T U1115 ( .I(a[13]), .ZN(n507) );
  INVD2BWP12T U1116 ( .I(a[9]), .ZN(n432) );
  XNR2D2BWP12T U1117 ( .A1(n3016), .A2(n4500), .ZN(n755) );
  XNR2D2BWP12T U1118 ( .A1(n3938), .A2(n4500), .ZN(n1786) );
  XNR2XD2BWP12T U1119 ( .A1(n3948), .A2(n4500), .ZN(n594) );
  OR2XD0BWP12T U1120 ( .A1(n1), .A2(n3667), .Z(n3280) );
  XNR2D2BWP12T U1121 ( .A1(n4503), .A2(n4609), .ZN(n413) );
  INVD2P3BWP12T U1122 ( .I(n4609), .ZN(n4607) );
  MUX2NXD1BWP12T U1123 ( .I0(n4608), .I1(n5299), .S(n4607), .ZN(n4613) );
  TPOAI22D1BWP12T U1124 ( .A1(n1689), .A2(n632), .B1(n2481), .B2(n614), .ZN(
        n640) );
  OAI21D1BWP12T U1125 ( .A1(n1783), .A2(n1782), .B(n1780), .ZN(n1781) );
  BUFFXD12BWP12T U1126 ( .I(n561), .Z(n2521) );
  CKND2D2BWP12T U1127 ( .A1(n847), .A2(n848), .ZN(n770) );
  INVD1BWP12T U1128 ( .I(n2773), .ZN(n405) );
  TPND2D2BWP12T U1129 ( .A1(n1628), .A2(n1627), .ZN(n1639) );
  FA1D2BWP12T U1130 ( .A(n1425), .B(n1424), .CI(n1423), .CO(n1581), .S(n1575)
         );
  FA1D2BWP12T U1131 ( .A(n1898), .B(n1897), .CI(n1896), .CO(n406) );
  INVD2BWP12T U1132 ( .I(n1173), .ZN(n1169) );
  TPND2D1BWP12T U1133 ( .A1(n1173), .A2(n1172), .ZN(n1174) );
  TPND2D3BWP12T U1134 ( .A1(n1347), .A2(n1346), .ZN(n1533) );
  NR2D0BWP12T U1135 ( .A1(n1), .A2(n5255), .ZN(n4611) );
  TPOAI22D2BWP12T U1136 ( .A1(n2518), .A2(n823), .B1(n726), .B2(n2516), .ZN(
        n805) );
  XNR2XD2BWP12T U1137 ( .A1(a[17]), .A2(n5033), .ZN(n726) );
  INVD3BWP12T U1138 ( .I(a[27]), .ZN(n2895) );
  BUFFD2BWP12T U1139 ( .I(n4993), .Z(n407) );
  DEL025D1BWP12T U1140 ( .I(n3134), .Z(n408) );
  INVD3BWP12T U1141 ( .I(n854), .ZN(n3134) );
  OAI22D2BWP12T U1142 ( .A1(n2532), .A2(n755), .B1(n754), .B2(n809), .ZN(n898)
         );
  TPOAI22D2BWP12T U1143 ( .A1(n2532), .A2(n3887), .B1(n727), .B2(n2530), .ZN(
        n903) );
  TPOAI22D1BWP12T U1144 ( .A1(n2529), .A2(n1711), .B1(n2), .B2(n1930), .ZN(
        n1849) );
  XOR2D2BWP12T U1145 ( .A1(n3003), .A2(n441), .Z(n4725) );
  INVD4BWP12T U1146 ( .I(n4503), .ZN(n3914) );
  XNR2XD2BWP12T U1147 ( .A1(n436), .A2(n4676), .ZN(n590) );
  ND2XD8BWP12T U1148 ( .A1(n4627), .A2(n4626), .ZN(result[28]) );
  TPOAI22D2BWP12T U1149 ( .A1(n560), .A2(n1969), .B1(n547), .B2(n3015), .ZN(
        n552) );
  XOR3XD4BWP12T U1150 ( .A1(n1844), .A2(n1845), .A3(n1843), .Z(n426) );
  TPND2D3BWP12T U1151 ( .A1(n649), .A2(n648), .ZN(n1845) );
  OR2D4BWP12T U1152 ( .A1(n1845), .A2(n1844), .Z(n1842) );
  XNR2XD4BWP12T U1153 ( .A1(n3068), .A2(n3067), .ZN(n5288) );
  XOR3D2BWP12T U1154 ( .A1(n1762), .A2(n1766), .A3(n1761), .Z(n409) );
  INVD2BWP12T U1155 ( .I(n939), .ZN(n942) );
  TPND2D2BWP12T U1156 ( .A1(n811), .A2(n810), .ZN(n813) );
  NR2XD1BWP12T U1157 ( .A1(n1639), .A2(n1640), .ZN(n1635) );
  TPND2D2BWP12T U1158 ( .A1(n833), .A2(n835), .ZN(n732) );
  CKND0BWP12T U1159 ( .I(n3684), .ZN(n410) );
  TPND2D2BWP12T U1160 ( .A1(n919), .A2(n918), .ZN(n1652) );
  CKND0BWP12T U1161 ( .I(n3075), .ZN(n411) );
  INVD1BWP12T U1162 ( .I(n411), .ZN(n412) );
  INVD2BWP12T U1163 ( .I(n2095), .ZN(n2098) );
  DCCKND4BWP12T U1164 ( .I(n719), .ZN(n574) );
  XNR2XD2BWP12T U1165 ( .A1(n5079), .A2(n5054), .ZN(n597) );
  AN2D1BWP12T U1166 ( .A1(n2131), .A2(n2130), .Z(n2133) );
  OR2XD1BWP12T U1167 ( .A1(n2131), .A2(n2130), .Z(n2132) );
  CKND2D2BWP12T U1168 ( .A1(n414), .A2(n415), .ZN(n417) );
  INVD2BWP12T U1169 ( .I(n1811), .ZN(n415) );
  TPNR2D1BWP12T U1170 ( .A1(n4668), .A2(n3073), .ZN(n3092) );
  TPND2D1BWP12T U1171 ( .A1(n3072), .A2(n3071), .ZN(n3073) );
  OR3D2BWP12T U1172 ( .A1(n3036), .A2(n3035), .A3(n3034), .Z(n3041) );
  XOR2XD2BWP12T U1173 ( .A1(n2875), .A2(n2874), .Z(n3036) );
  TPOAI21D1BWP12T U1174 ( .A1(n3011), .A2(n3008), .B(n3009), .ZN(n1002) );
  INVD18BWP12T U1175 ( .I(n1318), .ZN(n2005) );
  AN2XD2BWP12T U1176 ( .A1(n3152), .A2(n3154), .Z(n3142) );
  INVD1BWP12T U1177 ( .I(n822), .ZN(n798) );
  TPNR2D2BWP12T U1178 ( .A1(n1598), .A2(n1597), .ZN(n418) );
  TPNR2D2BWP12T U1179 ( .A1(n1598), .A2(n1597), .ZN(n3077) );
  TPND2D3BWP12T U1180 ( .A1(n487), .A2(n512), .ZN(n485) );
  XNR2XD2BWP12T U1181 ( .A1(n1812), .A2(n724), .ZN(n808) );
  BUFFXD8BWP12T U1182 ( .I(n2467), .Z(n420) );
  TPND2D1BWP12T U1183 ( .A1(n751), .A2(n752), .ZN(n567) );
  CKND2D2BWP12T U1184 ( .A1(n537), .A2(n536), .ZN(n539) );
  XNR2D2BWP12T U1185 ( .A1(n4788), .A2(n3016), .ZN(n1492) );
  NR2XD3BWP12T U1186 ( .A1(n1907), .A2(n1221), .ZN(n1284) );
  INVD2BWP12T U1187 ( .I(n1465), .ZN(n1460) );
  NR2D2BWP12T U1188 ( .A1(n1268), .A2(n1183), .ZN(n1184) );
  ND2D3BWP12T U1189 ( .A1(n5079), .A2(n2140), .ZN(n505) );
  TPOAI22D1BWP12T U1190 ( .A1(n2464), .A2(n2021), .B1(n2114), .B2(n2462), .ZN(
        n2064) );
  TPOAI22D2BWP12T U1191 ( .A1(n510), .A2(n2533), .B1(n554), .B2(n2535), .ZN(
        n607) );
  TPNR2D1BWP12T U1192 ( .A1(n2039), .A2(n2038), .ZN(n442) );
  CKND2D2BWP12T U1193 ( .A1(n4725), .A2(n5292), .ZN(n4754) );
  CKND0BWP12T U1194 ( .I(n3114), .ZN(n421) );
  INVD1BWP12T U1195 ( .I(n421), .ZN(n422) );
  TPOAI21D1BWP12T U1196 ( .A1(n3109), .A2(n3106), .B(n3110), .ZN(n3114) );
  INVD1BWP12T U1197 ( .I(n3085), .ZN(n3086) );
  TPOAI21D1BWP12T U1198 ( .A1(n1345), .A2(n1344), .B(n1343), .ZN(n423) );
  DCCKND4BWP12T U1199 ( .I(n1272), .ZN(n1345) );
  ND2D1BWP12T U1200 ( .A1(n1479), .A2(n1478), .ZN(n1480) );
  INVD2BWP12T U1201 ( .I(n1478), .ZN(n1474) );
  INR2D2BWP12T U1202 ( .A1(n3016), .B1(n2521), .ZN(n931) );
  TPND2D2BWP12T U1203 ( .A1(n1607), .A2(n1609), .ZN(n831) );
  TPND2D1BWP12T U1204 ( .A1(n910), .A2(n909), .ZN(n911) );
  TPND2D3BWP12T U1205 ( .A1(n843), .A2(n842), .ZN(n920) );
  XOR3D2BWP12T U1206 ( .A1(n746), .A2(n745), .A3(n744), .Z(n1649) );
  XNR2XD2BWP12T U1207 ( .A1(n2123), .A2(n5085), .ZN(n1450) );
  TPOAI22D2BWP12T U1208 ( .A1(n2467), .A2(n1447), .B1(n1446), .B2(n1799), .ZN(
        n1490) );
  DCCKND8BWP12T U1209 ( .I(a[5]), .ZN(n629) );
  INVD2P3BWP12T U1210 ( .I(n1767), .ZN(n1761) );
  XNR2XD2BWP12T U1211 ( .A1(n1906), .A2(n5237), .ZN(n1736) );
  XNR2XD2BWP12T U1212 ( .A1(n4511), .A2(n5237), .ZN(n828) );
  XNR2XD2BWP12T U1213 ( .A1(n5079), .A2(n5237), .ZN(n598) );
  XNR2XD2BWP12T U1214 ( .A1(a[17]), .A2(n5237), .ZN(n1925) );
  TPOAI21D1BWP12T U1215 ( .A1(n3084), .A2(n3083), .B(n438), .ZN(n3089) );
  XNR2XD2BWP12T U1216 ( .A1(n5079), .A2(n4826), .ZN(n1735) );
  TPND2D4BWP12T U1217 ( .A1(n4754), .A2(n4753), .ZN(result[18]) );
  INVD4BWP12T U1218 ( .I(n465), .ZN(n425) );
  INVD3BWP12T U1219 ( .I(n465), .ZN(n2146) );
  XOR3D2BWP12T U1220 ( .A1(n1844), .A2(n1845), .A3(n1843), .Z(n1677) );
  ND2XD8BWP12T U1221 ( .A1(n3875), .A2(n3882), .ZN(n3844) );
  XOR2XD2BWP12T U1222 ( .A1(n1812), .A2(n4676), .Z(n725) );
  AN2D4BWP12T U1223 ( .A1(n2600), .A2(n2599), .Z(n2601) );
  DCCKND4BWP12T U1224 ( .I(n2077), .ZN(n2025) );
  XOR3D2BWP12T U1225 ( .A1(n1748), .A2(n1747), .A3(n1745), .Z(n1844) );
  XNR2XD4BWP12T U1226 ( .A1(n1812), .A2(n1104), .ZN(n1120) );
  XOR2XD2BWP12T U1227 ( .A1(n3939), .A2(n1812), .Z(n1105) );
  TPOAI22D4BWP12T U1228 ( .A1(n866), .A2(n1969), .B1(n808), .B2(n3015), .ZN(
        n868) );
  BUFFXD8BWP12T U1229 ( .I(n1268), .Z(n2533) );
  INVD3BWP12T U1230 ( .I(n1430), .ZN(n1330) );
  BUFFXD16BWP12T U1231 ( .I(n2476), .Z(n1969) );
  XOR3XD4BWP12T U1232 ( .A1(n1433), .A2(n1469), .A3(n1468), .Z(n1565) );
  INVD3BWP12T U1233 ( .I(n1470), .ZN(n1433) );
  XOR3D2BWP12T U1234 ( .A1(n746), .A2(n745), .A3(n744), .Z(n427) );
  CKND2D2BWP12T U1235 ( .A1(n3147), .A2(n3146), .ZN(n3159) );
  BUFFD2BWP12T U1236 ( .I(n2140), .Z(n5234) );
  DCCKND4BWP12T U1237 ( .I(n2140), .ZN(n503) );
  CKND2D2BWP12T U1238 ( .A1(n3153), .A2(n3152), .ZN(n3155) );
  TPOAI21D1BWP12T U1239 ( .A1(n1986), .A2(n1985), .B(n1984), .ZN(n1988) );
  IND2D2BWP12T U1240 ( .A1(n1827), .B1(n1828), .ZN(n1832) );
  INR2D2BWP12T U1241 ( .A1(n1826), .B1(n1830), .ZN(n1827) );
  ND2D1BWP12T U1242 ( .A1(n1543), .A2(n69), .ZN(n1544) );
  BUFFD2BWP12T U1243 ( .I(n3150), .Z(n428) );
  CKND2D2BWP12T U1244 ( .A1(n1463), .A2(n1462), .ZN(n1467) );
  TPOAI22D1BWP12T U1245 ( .A1(n2518), .A2(n4790), .B1(n2022), .B2(n1429), .ZN(
        n429) );
  TPOAI22D1BWP12T U1246 ( .A1(n2518), .A2(n4790), .B1(n2516), .B2(n1429), .ZN(
        n1431) );
  HA1D2BWP12T U1247 ( .A(n1810), .B(n1809), .S(n430) );
  XNR2D2BWP12T U1248 ( .A1(a[17]), .A2(n3938), .ZN(n588) );
  IOA21D0BWP12T U1249 ( .A1(n1825), .A2(n1824), .B(n1823), .ZN(n1836) );
  TPOAI21D4BWP12T U1250 ( .A1(n1248), .A2(n1247), .B(n1246), .ZN(n1304) );
  TPND2D2BWP12T U1251 ( .A1(n1243), .A2(n1245), .ZN(n1246) );
  TPNR2D2BWP12T U1252 ( .A1(n1243), .A2(n1245), .ZN(n1248) );
  CKND2D2BWP12T U1253 ( .A1(a[10]), .A2(a[9]), .ZN(n433) );
  INVD2BWP12T U1254 ( .I(a[10]), .ZN(n431) );
  INVD3BWP12T U1255 ( .I(n2997), .ZN(n435) );
  ND2D4BWP12T U1256 ( .A1(n2996), .A2(n2995), .ZN(n2997) );
  RCOAI22D0BWP12T U1257 ( .A1(n1872), .A2(n1271), .B1(n2469), .B2(n1363), .ZN(
        n1367) );
  TPOAI22D1BWP12T U1258 ( .A1(n2469), .A2(n1271), .B1(n2020), .B2(n1234), .ZN(
        n1258) );
  INR2XD2BWP12T U1259 ( .A1(n3016), .B1(n2469), .ZN(n993) );
  NR2XD2BWP12T U1260 ( .A1(n2017), .A2(n2314), .ZN(n1904) );
  BUFFXD16BWP12T U1261 ( .I(a[3]), .Z(n436) );
  INVD3BWP12T U1262 ( .I(a[3]), .ZN(n512) );
  CKND0BWP12T U1263 ( .I(n71), .ZN(n437) );
  INVD1BWP12T U1264 ( .I(n3002), .ZN(n438) );
  XNR2XD2BWP12T U1265 ( .A1(a[1]), .A2(b[17]), .ZN(n439) );
  OAI21D1BWP12T U1266 ( .A1(n1439), .A2(n1440), .B(n1438), .ZN(n1442) );
  DEL100D1BWP12T U1267 ( .I(n4511), .Z(n2273) );
  INVD3BWP12T U1268 ( .I(n3140), .ZN(n3152) );
  TPNR2D3BWP12T U1269 ( .A1(n2041), .A2(n2040), .ZN(n3140) );
  INVD2BWP12T U1270 ( .I(b[28]), .ZN(n1811) );
  ND2XD4BWP12T U1271 ( .A1(n4936), .A2(n5292), .ZN(n4968) );
  NR2XD1BWP12T U1272 ( .A1(n3139), .A2(n3138), .ZN(n3166) );
  ND2XD8BWP12T U1273 ( .A1(n502), .A2(n501), .ZN(n2575) );
  XNR2XD2BWP12T U1274 ( .A1(n2067), .A2(n5264), .ZN(n1908) );
  TPNR2D2BWP12T U1275 ( .A1(n3124), .A2(n3125), .ZN(n2735) );
  BUFFXD8BWP12T U1276 ( .I(b[17]), .Z(n4794) );
  TPND2D3BWP12T U1277 ( .A1(n567), .A2(n566), .ZN(n745) );
  OR2D2BWP12T U1278 ( .A1(n1785), .A2(n51), .Z(n1738) );
  TPAOI21D1BWP12T U1279 ( .A1(n4896), .A2(n4895), .B(n4894), .ZN(n4897) );
  TPNR2D1BWP12T U1280 ( .A1(n3938), .A2(n4896), .ZN(n2317) );
  XNR2XD2BWP12T U1281 ( .A1(n2123), .A2(n4896), .ZN(n1187) );
  XNR2D2BWP12T U1282 ( .A1(n4511), .A2(n4896), .ZN(n1276) );
  XNR2D2BWP12T U1283 ( .A1(a[17]), .A2(n4896), .ZN(n589) );
  XNR2D2BWP12T U1284 ( .A1(n4896), .A2(n4500), .ZN(n1691) );
  XNR2D2BWP12T U1285 ( .A1(n5079), .A2(n4896), .ZN(n1382) );
  XNR2XD2BWP12T U1286 ( .A1(n48), .A2(n4896), .ZN(n861) );
  TPND2D3BWP12T U1287 ( .A1(n832), .A2(n831), .ZN(n1602) );
  OAI22D1BWP12T U1288 ( .A1(n1689), .A2(n796), .B1(n2115), .B2(n632), .ZN(n802) );
  TPOAI22D2BWP12T U1289 ( .A1(n2479), .A2(n1486), .B1(n1485), .B2(n2005), .ZN(
        n1508) );
  ND2XD0BWP12T U1290 ( .A1(n557), .A2(n568), .ZN(n559) );
  TPNR2D3BWP12T U1291 ( .A1(n1571), .A2(n1570), .ZN(n1643) );
  INVD2BWP12T U1292 ( .I(n1557), .ZN(n1513) );
  TPOAI22D1BWP12T U1293 ( .A1(n2471), .A2(n1051), .B1(n2469), .B2(n1102), .ZN(
        n1088) );
  TPOAI22D1BWP12T U1294 ( .A1(n2469), .A2(n1051), .B1(n2020), .B2(n1020), .ZN(
        n1053) );
  TPOAI22D2BWP12T U1295 ( .A1(n2471), .A2(n1143), .B1(n2469), .B2(n1187), .ZN(
        n1176) );
  TPND2D2BWP12T U1296 ( .A1(n769), .A2(n846), .ZN(n771) );
  INVD2BWP12T U1297 ( .I(n868), .ZN(n811) );
  RCOAI21D1BWP12T U1298 ( .A1(n840), .A2(n838), .B(n839), .ZN(n818) );
  XOR2XD2BWP12T U1299 ( .A1(b[1]), .A2(n3887), .Z(n754) );
  TPOAI22D2BWP12T U1300 ( .A1(n2519), .A2(n548), .B1(n2016), .B2(n4916), .ZN(
        n553) );
  XOR2XD4BWP12T U1301 ( .A1(n553), .A2(n552), .Z(n568) );
  TPNR2D2BWP12T U1302 ( .A1(n1428), .A2(n561), .ZN(n1378) );
  TPOAI21D1BWP12T U1303 ( .A1(n3006), .A2(n1422), .B(n1421), .ZN(n441) );
  TPOAI21D1BWP12T U1304 ( .A1(n3006), .A2(n1422), .B(n1421), .ZN(n3074) );
  IOA21D1BWP12T U1305 ( .A1(n572), .A2(n571), .B(n744), .ZN(n573) );
  XNR2XD2BWP12T U1306 ( .A1(n1812), .A2(n478), .ZN(n547) );
  XOR2XD2BWP12T U1307 ( .A1(n1812), .A2(b[25]), .Z(n690) );
  OR2XD1BWP12T U1308 ( .A1(n3098), .A2(n3097), .Z(n3099) );
  IOA21D2BWP12T U1309 ( .A1(n1783), .A2(n1782), .B(n1781), .ZN(n1883) );
  TPNR2D3BWP12T U1310 ( .A1(n3151), .A2(n2737), .ZN(n3144) );
  TPNR2D3BWP12T U1311 ( .A1(n3098), .A2(n3097), .ZN(n3151) );
  INVD2BWP12T U1312 ( .I(n1754), .ZN(n1709) );
  INVD2BWP12T U1313 ( .I(n2462), .ZN(n1680) );
  INVD1BWP12T U1314 ( .I(a[25]), .ZN(n691) );
  TPND2D1BWP12T U1315 ( .A1(n398), .A2(n1772), .ZN(n1773) );
  XOR2XD2BWP12T U1316 ( .A1(n1812), .A2(n5237), .Z(n1166) );
  XNR2XD2BWP12T U1317 ( .A1(n1812), .A2(n479), .ZN(n495) );
  XOR2XD2BWP12T U1318 ( .A1(n1812), .A2(n4700), .Z(n866) );
  XOR2XD8BWP12T U1319 ( .A1(n1812), .A2(b[27]), .Z(n1813) );
  TPNR2D3BWP12T U1320 ( .A1(n2039), .A2(n2038), .ZN(n2737) );
  INVD1BWP12T U1321 ( .I(n3157), .ZN(n3163) );
  TPOAI22D2BWP12T U1322 ( .A1(n1278), .A2(n1969), .B1(n1326), .B2(n3015), .ZN(
        n1332) );
  TPND2D2BWP12T U1323 ( .A1(n492), .A2(n491), .ZN(n585) );
  DEL025D1BWP12T U1324 ( .I(n1298), .Z(n443) );
  INVD3BWP12T U1325 ( .I(n1946), .ZN(n1942) );
  CKND2D2BWP12T U1326 ( .A1(n1876), .A2(n1875), .ZN(n1880) );
  OAI21D0BWP12T U1327 ( .A1(n1579), .A2(n1578), .B(n1577), .ZN(n1624) );
  XNR2XD0BWP12T U1328 ( .A1(n2944), .A2(n2943), .ZN(n3034) );
  AOI21D0BWP12T U1329 ( .A1(n2943), .A2(n2942), .B(n2870), .ZN(n2875) );
  TPNR2D1BWP12T U1330 ( .A1(n763), .A2(n766), .ZN(n643) );
  TPND2D2BWP12T U1331 ( .A1(n68), .A2(n1381), .ZN(n1491) );
  TPND2D2BWP12T U1332 ( .A1(n813), .A2(n867), .ZN(n815) );
  BUFFXD8BWP12T U1333 ( .I(b[19]), .Z(n4700) );
  IND2D4BWP12T U1334 ( .A1(n938), .B1(n937), .ZN(n2731) );
  INVD1BWP12T U1335 ( .I(n3013), .ZN(n938) );
  CKND2D2BWP12T U1336 ( .A1(n1468), .A2(n1435), .ZN(n1437) );
  XNR2XD4BWP12T U1337 ( .A1(n5030), .A2(n4794), .ZN(n756) );
  TPOAI22D1BWP12T U1338 ( .A1(n830), .A2(n2479), .B1(n2005), .B2(n756), .ZN(
        n897) );
  DCCKBD8BWP12T U1339 ( .I(n2141), .Z(n5118) );
  TPND2D3BWP12T U1340 ( .A1(n4565), .A2(n2141), .ZN(n452) );
  CKND4BWP12T U1341 ( .I(n2141), .ZN(n451) );
  BUFFXD3BWP12T U1342 ( .I(n2020), .Z(n2471) );
  TPND2D1BWP12T U1343 ( .A1(n1285), .A2(n1284), .ZN(n1286) );
  TPND2D2BWP12T U1344 ( .A1(n1079), .A2(n1073), .ZN(n446) );
  FA1D2BWP12T U1345 ( .A(n1898), .B(n1897), .CI(n1896), .CO(n1980), .S(n1937)
         );
  TPND2D2BWP12T U1346 ( .A1(n1399), .A2(n1398), .ZN(n1400) );
  INVD1BWP12T U1347 ( .I(n1593), .ZN(n1540) );
  INVD2BWP12T U1348 ( .I(n1561), .ZN(n1500) );
  INVD3BWP12T U1349 ( .I(n1420), .ZN(n1415) );
  TPND2D3BWP12T U1350 ( .A1(n3056), .A2(n3038), .ZN(n3044) );
  XOR3XD4BWP12T U1351 ( .A1(n699), .A2(n696), .A3(n698), .Z(n713) );
  ND2XD0BWP12T U1352 ( .A1(n2104), .A2(n2103), .ZN(n2105) );
  CKND0BWP12T U1353 ( .I(n4578), .ZN(n448) );
  INVD4BWP12T U1354 ( .I(n1409), .ZN(n2998) );
  RCOAI22D0BWP12T U1355 ( .A1(n405), .A2(n3591), .B1(n3587), .B2(n4607), .ZN(
        n2898) );
  OAI22D1BWP12T U1356 ( .A1(n29), .A2(n711), .B1(n2533), .B2(n1692), .ZN(n1684) );
  TPOAI22D1BWP12T U1357 ( .A1(n29), .A2(n1956), .B1(n2533), .B2(n2094), .ZN(
        n2058) );
  TPOAI22D1BWP12T U1358 ( .A1(n2535), .A2(n1229), .B1(n2533), .B2(n1228), .ZN(
        n1231) );
  TPOAI22D1BWP12T U1359 ( .A1(n2535), .A2(n862), .B1(n2533), .B2(n807), .ZN(
        n860) );
  XNR2XD8BWP12T U1360 ( .A1(n3495), .A2(n71), .ZN(n2481) );
  TPOAI21D1BWP12T U1361 ( .A1(n2467), .A2(n678), .B(n677), .ZN(n687) );
  INVD18BWP12T U1362 ( .I(n2904), .ZN(n4565) );
  INVD8BWP12T U1363 ( .I(a[19]), .ZN(n2904) );
  TPOAI22D2BWP12T U1364 ( .A1(n2535), .A2(n1269), .B1(n396), .B2(n1358), .ZN(
        n1369) );
  XNR2D2BWP12T U1365 ( .A1(n3948), .A2(n1858), .ZN(n1358) );
  INR2XD2BWP12T U1366 ( .A1(n3016), .B1(n1799), .ZN(n1098) );
  TPNR2D2BWP12T U1367 ( .A1(n984), .A2(n983), .ZN(n1011) );
  XNR2XD2BWP12T U1368 ( .A1(n4565), .A2(n3938), .ZN(n693) );
  INVD2BWP12T U1369 ( .I(n1479), .ZN(n1475) );
  INVD1BWP12T U1370 ( .I(n1590), .ZN(n449) );
  ND2XD8BWP12T U1371 ( .A1(n1152), .A2(n1151), .ZN(n3038) );
  XNR2XD2BWP12T U1372 ( .A1(n436), .A2(n3899), .ZN(n1108) );
  TPOAI22D1BWP12T U1373 ( .A1(n1908), .A2(n2575), .B1(n1907), .B2(n2007), .ZN(
        n2013) );
  OAI22D2BWP12T U1374 ( .A1(n2575), .A2(n3895), .B1(n1270), .B2(n1907), .ZN(
        n1368) );
  ND2D8BWP12T U1375 ( .A1(n450), .A2(n451), .ZN(n453) );
  ND2XD8BWP12T U1376 ( .A1(n452), .A2(n453), .ZN(n809) );
  BUFFXD12BWP12T U1377 ( .I(n809), .Z(n2530) );
  DCCKND4BWP12T U1378 ( .I(n809), .ZN(n709) );
  CKND0BWP12T U1379 ( .I(n4635), .ZN(n454) );
  TPNR2D1BWP12T U1380 ( .A1(n1938), .A2(n1937), .ZN(n1936) );
  XNR2D2BWP12T U1381 ( .A1(n436), .A2(b[22]), .ZN(n679) );
  XNR2XD2BWP12T U1382 ( .A1(n3911), .A2(b[22]), .ZN(n1687) );
  INVD3BWP12T U1383 ( .I(b[7]), .ZN(n473) );
  TPNR2D1BWP12T U1384 ( .A1(n1852), .A2(n1851), .ZN(n1854) );
  INVD6BWP12T U1385 ( .I(a[25]), .ZN(n3915) );
  XOR3XD4BWP12T U1386 ( .A1(n1722), .A2(n1721), .A3(n1720), .Z(n1825) );
  ND2D1BWP12T U1387 ( .A1(n1721), .A2(n1722), .ZN(n455) );
  CKND2D2BWP12T U1388 ( .A1(n1721), .A2(n1720), .ZN(n456) );
  TPOAI22D1BWP12T U1389 ( .A1(n1969), .A2(n690), .B1(n1739), .B2(n3015), .ZN(
        n1744) );
  XNR2D2BWP12T U1390 ( .A1(n1858), .A2(n3938), .ZN(n1503) );
  TPOAI21D1BWP12T U1391 ( .A1(n1817), .A2(n1818), .B(n1815), .ZN(n1816) );
  TPOAI22D1BWP12T U1392 ( .A1(n2523), .A2(n1683), .B1(n2521), .B2(n1814), .ZN(
        n1815) );
  XNR2XD2BWP12T U1393 ( .A1(n436), .A2(n2122), .ZN(n1814) );
  TPAOI21D2BWP12T U1394 ( .A1(n3057), .A2(n3038), .B(n1157), .ZN(n458) );
  TPOAI22D1BWP12T U1395 ( .A1(n2020), .A2(n1102), .B1(n14), .B2(n1143), .ZN(
        n1137) );
  XNR2XD2BWP12T U1396 ( .A1(n2123), .A2(n5033), .ZN(n1143) );
  TPND2D1BWP12T U1397 ( .A1(n1626), .A2(n1625), .ZN(n1627) );
  TPOAI22D2BWP12T U1398 ( .A1(n1872), .A2(n884), .B1(n2469), .B2(n824), .ZN(
        n878) );
  OAI22D1BWP12T U1399 ( .A1(n2532), .A2(n1857), .B1(n2004), .B2(n2530), .ZN(
        n1958) );
  ND2D8BWP12T U1400 ( .A1(n2384), .A2(n2383), .ZN(result[31]) );
  TPOAI22D2BWP12T U1401 ( .A1(n2031), .A2(n2030), .B1(n2029), .B2(n2028), .ZN(
        n2049) );
  RCOAI21D8BWP12T U1402 ( .A1(n4935), .A2(n5112), .B(n4934), .ZN(result[23])
         );
  XNR2D2BWP12T U1403 ( .A1(n5033), .A2(n1906), .ZN(n1502) );
  ND2D4BWP12T U1404 ( .A1(n2039), .A2(n2038), .ZN(n3150) );
  NR2D0BWP12T U1405 ( .A1(b[27]), .A2(n4944), .ZN(n2319) );
  INVD18BWP12T U1406 ( .I(n480), .ZN(n3015) );
  OR2XD1BWP12T U1407 ( .A1(n2250), .A2(n4568), .Z(n3268) );
  INVD4BWP12T U1408 ( .I(b[5]), .ZN(n2321) );
  INVD9BWP12T U1409 ( .I(n2321), .ZN(n5033) );
  BUFFXD4BWP12T U1410 ( .I(n2122), .Z(n4977) );
  INVD3BWP12T U1411 ( .I(n4977), .ZN(n2250) );
  BUFFXD3BWP12T U1412 ( .I(n1906), .Z(n2067) );
  OA21D1BWP12T U1413 ( .A1(n1087), .A2(n1086), .B(n1085), .Z(n460) );
  INVD8BWP12T U1414 ( .I(n950), .ZN(n5030) );
  BUFFD8BWP12T U1415 ( .I(a[0]), .Z(n480) );
  BUFFXD6BWP12T U1416 ( .I(n4502), .Z(n5049) );
  TPNR2D1BWP12T U1417 ( .A1(b[22]), .A2(n2825), .ZN(n4360) );
  BUFFD2BWP12T U1418 ( .I(n5033), .Z(n2190) );
  INVD2BWP12T U1419 ( .I(b[11]), .ZN(n1104) );
  INVD2BWP12T U1420 ( .I(n5085), .ZN(n2234) );
  INVD2BWP12T U1421 ( .I(n5085), .ZN(n2155) );
  NR2XD3BWP12T U1422 ( .A1(n4299), .A2(n4297), .ZN(n4208) );
  CKBD1BWP12T U1423 ( .I(n4501), .Z(n3684) );
  CKBD1BWP12T U1424 ( .I(n3948), .Z(n2269) );
  INVD1BWP12T U1425 ( .I(n4043), .ZN(n4044) );
  INVD2BWP12T U1426 ( .I(n4889), .ZN(n5321) );
  INVD1BWP12T U1427 ( .I(n2387), .ZN(n3217) );
  INVD1BWP12T U1428 ( .I(n2876), .ZN(n2962) );
  BUFFD2BWP12T U1429 ( .I(n4990), .Z(n2255) );
  BUFFD3BWP12T U1430 ( .I(n4896), .Z(n2271) );
  INVD2BWP12T U1431 ( .I(n2271), .ZN(n2227) );
  TPNR2D1BWP12T U1432 ( .A1(n4510), .A2(n2640), .ZN(n2661) );
  TPNR2D1BWP12T U1433 ( .A1(n2270), .A2(n2190), .ZN(n4417) );
  BUFFD2BWP12T U1434 ( .I(n4511), .Z(n2153) );
  INVD2BWP12T U1435 ( .I(n3237), .ZN(n3241) );
  INVD3BWP12T U1436 ( .I(n5104), .ZN(n5297) );
  TPND2D1BWP12T U1437 ( .A1(n2351), .A2(n2353), .ZN(n5104) );
  ND2D8BWP12T U1438 ( .A1(n4201), .A2(n2677), .ZN(n4309) );
  INVD6BWP12T U1439 ( .I(n4309), .ZN(n2839) );
  INVD1BWP12T U1440 ( .I(n5322), .ZN(n5271) );
  INR2D2BWP12T U1441 ( .A1(n2425), .B1(n2413), .ZN(n5322) );
  INVD1BWP12T U1442 ( .I(n4117), .ZN(n2203) );
  TPND2D2BWP12T U1443 ( .A1(n1165), .A2(n1164), .ZN(n1243) );
  NR2D2BWP12T U1444 ( .A1(n3507), .A2(n3506), .ZN(n5211) );
  DEL025D1BWP12T U1445 ( .I(n3939), .Z(n2195) );
  INVD4BWP12T U1446 ( .I(n3588), .ZN(n3498) );
  OR2D2BWP12T U1447 ( .A1(n1054), .A2(n1053), .Z(n462) );
  BUFFD6BWP12T U1448 ( .I(n4503), .Z(n2773) );
  OR2D2BWP12T U1449 ( .A1(n793), .A2(n794), .Z(n463) );
  INVD4BWP12T U1450 ( .I(a[14]), .ZN(n5260) );
  TPND2D2BWP12T U1451 ( .A1(n717), .A2(n716), .ZN(n1824) );
  INVD6BWP12T U1452 ( .I(n4635), .ZN(n2825) );
  BUFFXD4BWP12T U1453 ( .I(b[26]), .Z(n4944) );
  INVD2BWP12T U1454 ( .I(b[26]), .ZN(n689) );
  INVD8BWP12T U1455 ( .I(n70), .ZN(n5192) );
  INVD2BWP12T U1456 ( .I(b[14]), .ZN(n1222) );
  AN2XD2BWP12T U1457 ( .A1(n1788), .A2(n1787), .Z(n464) );
  INVD16BWP12T U1458 ( .I(n1106), .ZN(n5079) );
  ND2XD4BWP12T U1459 ( .A1(n488), .A2(n487), .ZN(n561) );
  BUFFXD4BWP12T U1460 ( .I(n629), .Z(n950) );
  TPOAI21D4BWP12T U1461 ( .A1(n3123), .A2(n3125), .B(n3126), .ZN(n2736) );
  BUFFXD3BWP12T U1462 ( .I(n1770), .Z(n1772) );
  TPND2D1BWP12T U1463 ( .A1(n3127), .A2(n3126), .ZN(n3128) );
  TPAOI21D4BWP12T U1464 ( .A1(n1185), .A2(n5049), .B(n1184), .ZN(n1213) );
  TPOAI22D2BWP12T U1465 ( .A1(n2467), .A2(n1167), .B1(n1799), .B2(n1235), .ZN(
        n1226) );
  XNR2XD2BWP12T U1466 ( .A1(n5079), .A2(n5196), .ZN(n1167) );
  CKND2D2BWP12T U1467 ( .A1(n1350), .A2(n1349), .ZN(n1351) );
  RCOAI21D1BWP12T U1468 ( .A1(n398), .A2(n1772), .B(n1771), .ZN(n1774) );
  ND2XD8BWP12T U1469 ( .A1(n469), .A2(n1869), .ZN(n2016) );
  ND2D3BWP12T U1470 ( .A1(a[1]), .A2(a[2]), .ZN(n487) );
  TPOAI22D4BWP12T U1471 ( .A1(n1689), .A2(n1186), .B1(n1225), .B2(n2115), .ZN(
        n1232) );
  FA1D2BWP12T U1472 ( .A(n2570), .B(n2569), .CI(n2568), .CO(n2580), .S(n2510)
         );
  IOA21D2BWP12T U1473 ( .A1(n2013), .A2(n2012), .B(n2011), .ZN(n2075) );
  OAI22D2BWP12T U1474 ( .A1(n2573), .A2(n1909), .B1(n2571), .B2(n1968), .ZN(
        n2012) );
  TPOAI21D1BWP12T U1475 ( .A1(n3151), .A2(n3150), .B(n3149), .ZN(n3153) );
  TPOAI22D2BWP12T U1476 ( .A1(n2523), .A2(n590), .B1(n679), .B2(n2521), .ZN(
        n549) );
  DCCKND4BWP12T U1477 ( .I(a[6]), .ZN(n465) );
  XNR2XD8BWP12T U1478 ( .A1(n513), .A2(n425), .ZN(n1384) );
  XNR2XD8BWP12T U1479 ( .A1(n2303), .A2(n2146), .ZN(n466) );
  ND2XD8BWP12T U1480 ( .A1(n1384), .A2(n466), .ZN(n2020) );
  XNR2XD2BWP12T U1481 ( .A1(n2123), .A2(n4794), .ZN(n600) );
  BUFFXD16BWP12T U1482 ( .I(n1384), .Z(n2469) );
  BUFFD8BWP12T U1483 ( .I(b[18]), .Z(n4732) );
  XNR2XD2BWP12T U1484 ( .A1(n2123), .A2(n4732), .ZN(n667) );
  OR2D4BWP12T U1485 ( .A1(n2469), .A2(n667), .Z(n467) );
  DCCKND4BWP12T U1486 ( .I(a[23]), .ZN(n468) );
  BUFFD6BWP12T U1487 ( .I(a[22]), .Z(n2142) );
  XOR2XD4BWP12T U1488 ( .A1(n2014), .A2(n2142), .Z(n469) );
  INVD3BWP12T U1489 ( .I(a[21]), .ZN(n2899) );
  INVD8BWP12T U1490 ( .I(n2899), .ZN(n4500) );
  XNR2XD8BWP12T U1491 ( .A1(n4500), .A2(n2142), .ZN(n1869) );
  INVD6BWP12T U1492 ( .I(b[2]), .ZN(n3906) );
  INVD18BWP12T U1493 ( .I(n3906), .ZN(n5196) );
  INVD1BWP12T U1494 ( .I(n5196), .ZN(n470) );
  CKND3BWP12T U1495 ( .I(n2014), .ZN(n4916) );
  XNR2XD4BWP12T U1496 ( .A1(n470), .A2(n4916), .ZN(n681) );
  XNR2XD4BWP12T U1497 ( .A1(n4500), .A2(n2142), .ZN(n2519) );
  TPOAI22D4BWP12T U1498 ( .A1(n397), .A2(n586), .B1(n681), .B2(n2519), .ZN(
        n620) );
  BUFFXD8BWP12T U1499 ( .I(a[16]), .Z(n4822) );
  XNR2XD8BWP12T U1500 ( .A1(n4822), .A2(n1906), .ZN(n472) );
  XOR2XD8BWP12T U1501 ( .A1(a[17]), .A2(n4822), .Z(n471) );
  ND2XD16BWP12T U1502 ( .A1(n472), .A2(n471), .ZN(n2518) );
  INVD6BWP12T U1503 ( .I(n474), .ZN(n3899) );
  XNR2D1BWP12T U1504 ( .A1(a[17]), .A2(n3899), .ZN(n494) );
  XNR2XD8BWP12T U1505 ( .A1(n4822), .A2(n1906), .ZN(n2516) );
  TPOAI22D1BWP12T U1506 ( .A1(n2518), .A2(n588), .B1(n494), .B2(n2022), .ZN(
        n617) );
  TPNR2D1BWP12T U1507 ( .A1(n620), .A2(n617), .ZN(n476) );
  CKND2D1BWP12T U1508 ( .A1(n620), .A2(n617), .ZN(n475) );
  BUFFXD16BWP12T U1509 ( .I(b[0]), .Z(n3016) );
  BUFFD6BWP12T U1510 ( .I(a[24]), .Z(n4649) );
  XNR2XD8BWP12T U1511 ( .A1(n4649), .A2(n2014), .ZN(n2527) );
  INR2XD2BWP12T U1512 ( .A1(n3016), .B1(n2527), .ZN(n551) );
  INVD1BWP12T U1513 ( .I(n551), .ZN(n483) );
  INVD18BWP12T U1514 ( .I(a[1]), .ZN(n1812) );
  CKND3BWP12T U1515 ( .I(b[23]), .ZN(n478) );
  CKND3BWP12T U1516 ( .I(b[24]), .ZN(n479) );
  TPNR2D3BWP12T U1517 ( .A1(n482), .A2(n481), .ZN(n550) );
  BUFFXD6BWP12T U1518 ( .I(b[21]), .Z(n4676) );
  TPND2D2BWP12T U1519 ( .A1(n489), .A2(n549), .ZN(n492) );
  TPND2D1BWP12T U1520 ( .A1(n490), .A2(n551), .ZN(n491) );
  INVD4BWP12T U1521 ( .I(b[9]), .ZN(n493) );
  INVD8BWP12T U1522 ( .I(n493), .ZN(n3930) );
  BUFFXD3BWP12T U1523 ( .I(b[25]), .Z(n2122) );
  TPOAI22D1BWP12T U1524 ( .A1(n690), .A2(n3015), .B1(n495), .B2(n1969), .ZN(
        n695) );
  OR2XD1BWP12T U1525 ( .A1(n584), .A2(n585), .Z(n496) );
  ND2D1BWP12T U1526 ( .A1(n583), .A2(n496), .ZN(n498) );
  ND2D1BWP12T U1527 ( .A1(n585), .A2(n584), .ZN(n497) );
  CKND2D2BWP12T U1528 ( .A1(n498), .A2(n497), .ZN(n1748) );
  CKND2D2BWP12T U1529 ( .A1(n3895), .A2(n1858), .ZN(n499) );
  ND2D4BWP12T U1530 ( .A1(n500), .A2(n5260), .ZN(n501) );
  XNR2XD8BWP12T U1531 ( .A1(a[14]), .A2(n1858), .ZN(n1907) );
  BUFFXD8BWP12T U1532 ( .I(b[11]), .Z(n5085) );
  TPOAI22D2BWP12T U1533 ( .A1(n2575), .A2(n546), .B1(n1907), .B2(n694), .ZN(
        n533) );
  BUFFXD4BWP12T U1534 ( .I(a[12]), .Z(n2140) );
  XOR2XD4BWP12T U1535 ( .A1(n1858), .A2(n2140), .Z(n506) );
  INVD8BWP12T U1536 ( .I(a[11]), .ZN(n1106) );
  ND2D8BWP12T U1537 ( .A1(n5081), .A2(n503), .ZN(n504) );
  ND2XD8BWP12T U1538 ( .A1(n505), .A2(n504), .ZN(n1268) );
  ND2XD8BWP12T U1539 ( .A1(n506), .A2(n1268), .ZN(n2535) );
  BUFFD6BWP12T U1540 ( .I(b[12]), .Z(n5237) );
  XNR2D1BWP12T U1541 ( .A1(n6), .A2(n5237), .ZN(n510) );
  INVD4BWP12T U1542 ( .I(n507), .ZN(n4502) );
  BUFFXD8BWP12T U1543 ( .I(b[13]), .Z(n5054) );
  XNR2D1BWP12T U1544 ( .A1(n4502), .A2(n5054), .ZN(n711) );
  XNR2XD8BWP12T U1545 ( .A1(a[17]), .A2(a[18]), .ZN(n2571) );
  ND2XD16BWP12T U1546 ( .A1(n2571), .A2(n508), .ZN(n2573) );
  INVD2BWP12T U1547 ( .I(b[6]), .ZN(n509) );
  INVD6BWP12T U1548 ( .I(n509), .ZN(n4896) );
  TPOAI22D2BWP12T U1549 ( .A1(n2573), .A2(n511), .B1(n2571), .B2(n693), .ZN(
        n534) );
  XOR3XD4BWP12T U1550 ( .A1(n533), .A2(n531), .A3(n534), .Z(n663) );
  XNR2D1BWP12T U1551 ( .A1(n1858), .A2(n5085), .ZN(n554) );
  XNR2D1BWP12T U1552 ( .A1(n4565), .A2(n5033), .ZN(n612) );
  TPOAI22D1BWP12T U1553 ( .A1(n2573), .A2(n612), .B1(n2571), .B2(n511), .ZN(
        n605) );
  XNR2D2BWP12T U1554 ( .A1(n3911), .A2(n4700), .ZN(n613) );
  INVD8BWP12T U1555 ( .I(a[4]), .ZN(n3912) );
  TPAOI21D8BWP12T U1556 ( .A1(n2185), .A2(n514), .B(n3912), .ZN(n517) );
  TPNR2D8BWP12T U1557 ( .A1(n517), .A2(n516), .ZN(n1315) );
  INVD12BWP12T U1558 ( .I(n1315), .ZN(n2479) );
  XOR2XD8BWP12T U1559 ( .A1(a[3]), .A2(a[4]), .Z(n1318) );
  XNR2D1BWP12T U1560 ( .A1(n3911), .A2(b[20]), .ZN(n665) );
  TPOAI22D2BWP12T U1561 ( .A1(n613), .A2(n2479), .B1(n2005), .B2(n665), .ZN(
        n608) );
  TPNR2D1BWP12T U1562 ( .A1(n605), .A2(n608), .ZN(n519) );
  ND2D1BWP12T U1563 ( .A1(n605), .A2(n608), .ZN(n518) );
  BUFFXD8BWP12T U1564 ( .I(a[8]), .Z(n3495) );
  DCCKND4BWP12T U1565 ( .I(a[7]), .ZN(n521) );
  XNR2XD4BWP12T U1566 ( .A1(n3495), .A2(n1007), .ZN(n523) );
  INVD15BWP12T U1567 ( .I(n2910), .ZN(n4511) );
  XOR2XD8BWP12T U1568 ( .A1(n56), .A2(n3495), .Z(n522) );
  ND2XD16BWP12T U1569 ( .A1(n523), .A2(n522), .ZN(n1689) );
  BUFFXD8BWP12T U1570 ( .I(b[15]), .Z(n4770) );
  XNR2D1BWP12T U1571 ( .A1(n4511), .A2(n4770), .ZN(n614) );
  BUFFD6BWP12T U1572 ( .I(b[16]), .Z(n4826) );
  OAI22D0BWP12T U1573 ( .A1(n1689), .A2(n614), .B1(n2481), .B2(n670), .ZN(n621) );
  XNR2XD4BWP12T U1574 ( .A1(n1106), .A2(a[10]), .ZN(n524) );
  ND2XD8BWP12T U1575 ( .A1(n524), .A2(n525), .ZN(n2467) );
  XNR2D1BWP12T U1576 ( .A1(n5079), .A2(n5264), .ZN(n678) );
  BUFFXD12BWP12T U1577 ( .I(n525), .Z(n1799) );
  TPOAI22D1BWP12T U1578 ( .A1(n2467), .A2(n597), .B1(n678), .B2(n1799), .ZN(
        n623) );
  INVD6BWP12T U1579 ( .I(b[4]), .ZN(n2311) );
  INVD12BWP12T U1580 ( .I(n2311), .ZN(n4301) );
  XNR2XD0BWP12T U1581 ( .A1(n4301), .A2(n4500), .ZN(n674) );
  INVD4BWP12T U1582 ( .I(b[3]), .ZN(n2362) );
  INVD12BWP12T U1583 ( .I(n2362), .ZN(n3948) );
  TPOAI22D2BWP12T U1584 ( .A1(n674), .A2(n2530), .B1(n2532), .B2(n594), .ZN(
        n622) );
  CKND2BWP12T U1585 ( .I(n622), .ZN(n526) );
  ND2D1BWP12T U1586 ( .A1(n623), .A2(n622), .ZN(n527) );
  IOA21D2BWP12T U1587 ( .A1(n621), .A2(n528), .B(n527), .ZN(n661) );
  ND2D2BWP12T U1588 ( .A1(n530), .A2(n529), .ZN(n1747) );
  IOA21D2BWP12T U1589 ( .A1(n534), .A2(n533), .B(n532), .ZN(n1750) );
  XNR2D2BWP12T U1590 ( .A1(n4301), .A2(n2014), .ZN(n1741) );
  TPOAI22D1BWP12T U1591 ( .A1(n2016), .A2(n680), .B1(n1741), .B2(n2519), .ZN(
        n1694) );
  INVD1BWP12T U1592 ( .I(n535), .ZN(n536) );
  XNR2D2BWP12T U1593 ( .A1(a[17]), .A2(n3939), .ZN(n1678) );
  OR2D2BWP12T U1594 ( .A1(n1678), .A2(n2516), .Z(n538) );
  TPND2D3BWP12T U1595 ( .A1(n539), .A2(n538), .ZN(n1697) );
  INVD6BWP12T U1596 ( .I(n2020), .ZN(n540) );
  INVD8BWP12T U1597 ( .I(n540), .ZN(n1872) );
  BUFFXD4BWP12T U1598 ( .I(b[20]), .Z(n5122) );
  XNR2XD2BWP12T U1599 ( .A1(n2123), .A2(n5122), .ZN(n1729) );
  TPOAI22D1BWP12T U1600 ( .A1(n1872), .A2(n666), .B1(n2469), .B2(n1729), .ZN(
        n1700) );
  XOR3XD4BWP12T U1601 ( .A1(n1694), .A2(n1697), .A3(n1700), .Z(n1751) );
  XNR2XD4BWP12T U1602 ( .A1(n5079), .A2(n4770), .ZN(n675) );
  INVD1P75BWP12T U1603 ( .I(n1735), .ZN(n541) );
  CKND3BWP12T U1604 ( .I(n1799), .ZN(n1110) );
  TPND2D2BWP12T U1605 ( .A1(n541), .A2(n1110), .ZN(n542) );
  TPOAI21D2BWP12T U1606 ( .A1(n2467), .A2(n675), .B(n542), .ZN(n1702) );
  TPOAI22D1BWP12T U1607 ( .A1(n1689), .A2(n671), .B1(n2481), .B2(n1688), .ZN(
        n1701) );
  XOR2XD4BWP12T U1608 ( .A1(n4568), .A2(n4649), .Z(n543) );
  XNR2D2BWP12T U1609 ( .A1(b[1]), .A2(n4568), .ZN(n668) );
  XNR2D1BWP12T U1610 ( .A1(n5196), .A2(n4568), .ZN(n1690) );
  TPOAI22D2BWP12T U1611 ( .A1(n2529), .A2(n668), .B1(n1690), .B2(n23), .ZN(
        n1703) );
  INVD1P75BWP12T U1612 ( .I(n1703), .ZN(n544) );
  XNR3XD4BWP12T U1613 ( .A1(n1702), .A2(n1701), .A3(n544), .ZN(n1749) );
  CKND3BWP12T U1614 ( .I(n1749), .ZN(n545) );
  XNR3XD4BWP12T U1615 ( .A1(n1750), .A2(n1751), .A3(n545), .ZN(n1745) );
  TPOAI22D1BWP12T U1616 ( .A1(n51), .A2(n546), .B1(n2575), .B2(n555), .ZN(n579) );
  XOR2D2BWP12T U1617 ( .A1(b[22]), .A2(n1812), .Z(n560) );
  IND2D1BWP12T U1618 ( .A1(b[0]), .B1(n4914), .ZN(n548) );
  AN2XD2BWP12T U1619 ( .A1(n553), .A2(n552), .Z(n578) );
  XNR3XD4BWP12T U1620 ( .A1(n551), .A2(n550), .A3(n549), .ZN(n577) );
  XOR3XD4BWP12T U1621 ( .A1(n579), .A2(n578), .A3(n577), .Z(n719) );
  XNR2XD0BWP12T U1622 ( .A1(n1858), .A2(b[10]), .ZN(n737) );
  TPOAI22D1BWP12T U1623 ( .A1(n2535), .A2(n737), .B1(n2533), .B2(n554), .ZN(
        n569) );
  XNR2XD2BWP12T U1624 ( .A1(n48), .A2(n3899), .ZN(n735) );
  TPOAI22D2BWP12T U1625 ( .A1(n2575), .A2(n735), .B1(n1907), .B2(n555), .ZN(
        n570) );
  IND2D2BWP12T U1626 ( .A1(n569), .B1(n556), .ZN(n557) );
  INVD1BWP12T U1627 ( .I(n720), .ZN(n575) );
  NR2XD2BWP12T U1628 ( .A1(n2519), .A2(n3233), .ZN(n723) );
  TPOAI22D2BWP12T U1629 ( .A1(n560), .A2(n3015), .B1(n725), .B2(n1969), .ZN(
        n722) );
  XNR2XD2BWP12T U1630 ( .A1(n436), .A2(n4700), .ZN(n729) );
  XNR2D1BWP12T U1631 ( .A1(n436), .A2(b[20]), .ZN(n591) );
  OAI22D1BWP12T U1632 ( .A1(n2523), .A2(n729), .B1(n2521), .B2(n591), .ZN(n721) );
  OAI21D1BWP12T U1633 ( .A1(n723), .A2(n722), .B(n721), .ZN(n563) );
  ND2D2BWP12T U1634 ( .A1(n563), .A2(n562), .ZN(n746) );
  XNR2XD2BWP12T U1635 ( .A1(n2123), .A2(n4826), .ZN(n601) );
  ND2D3BWP12T U1636 ( .A1(n565), .A2(n564), .ZN(n751) );
  TPOAI22D2BWP12T U1637 ( .A1(n2518), .A2(n726), .B1(n589), .B2(n2516), .ZN(
        n752) );
  XNR2D1BWP12T U1638 ( .A1(n1104), .A2(n1106), .ZN(n728) );
  TPOAI22D2BWP12T U1639 ( .A1(n2467), .A2(n728), .B1(n598), .B2(n1799), .ZN(
        n753) );
  TPOAI21D2BWP12T U1640 ( .A1(n751), .A2(n752), .B(n753), .ZN(n566) );
  CKND2BWP12T U1641 ( .I(n745), .ZN(n571) );
  XOR3XD4BWP12T U1642 ( .A1(n570), .A2(n569), .A3(n568), .Z(n744) );
  IOA21D2BWP12T U1643 ( .A1(n574), .A2(n575), .B(n718), .ZN(n576) );
  IOA21D2BWP12T U1644 ( .A1(n719), .A2(n720), .B(n576), .ZN(n781) );
  INVD2BWP12T U1645 ( .I(n577), .ZN(n582) );
  TPNR2D1BWP12T U1646 ( .A1(n578), .A2(n579), .ZN(n581) );
  ND2D1BWP12T U1647 ( .A1(n579), .A2(n578), .ZN(n580) );
  TPOAI21D2BWP12T U1648 ( .A1(n582), .A2(n581), .B(n580), .ZN(n778) );
  XOR3XD4BWP12T U1649 ( .A1(n585), .A2(n584), .A3(n583), .Z(n777) );
  XNR2D2BWP12T U1650 ( .A1(n3016), .A2(n2014), .ZN(n587) );
  ND2D1BWP12T U1651 ( .A1(n633), .A2(n634), .ZN(n592) );
  TPND2D1BWP12T U1652 ( .A1(n593), .A2(n592), .ZN(n625) );
  XOR2D2BWP12T U1653 ( .A1(n3887), .A2(n5196), .Z(n631) );
  TPNR2D2BWP12T U1654 ( .A1(n2532), .A2(n631), .ZN(n596) );
  NR2D1BWP12T U1655 ( .A1(n594), .A2(n809), .ZN(n595) );
  NR2D2BWP12T U1656 ( .A1(n596), .A2(n595), .ZN(n739) );
  TPOAI22D2BWP12T U1657 ( .A1(n2467), .A2(n598), .B1(n597), .B2(n1799), .ZN(
        n740) );
  TPND2D1BWP12T U1658 ( .A1(n739), .A2(n599), .ZN(n602) );
  IND2D2BWP12T U1659 ( .A1(n739), .B1(n740), .ZN(n603) );
  CKND2D2BWP12T U1660 ( .A1(n604), .A2(n603), .ZN(n628) );
  INVD1BWP12T U1661 ( .I(n605), .ZN(n606) );
  XNR3XD4BWP12T U1662 ( .A1(n608), .A2(n607), .A3(n606), .ZN(n627) );
  OA21XD2BWP12T U1663 ( .A1(n611), .A2(n610), .B(n609), .Z(n776) );
  TPOAI22D1BWP12T U1664 ( .A1(n2573), .A2(n736), .B1(n2571), .B2(n612), .ZN(
        n637) );
  XNR2D1BWP12T U1665 ( .A1(n3911), .A2(n4732), .ZN(n630) );
  OAI22D2BWP12T U1666 ( .A1(n2479), .A2(n630), .B1(n2005), .B2(n613), .ZN(n636) );
  XNR2D1BWP12T U1667 ( .A1(n4511), .A2(n5264), .ZN(n632) );
  OAI21D1BWP12T U1668 ( .A1(n637), .A2(n636), .B(n640), .ZN(n616) );
  ND2D1BWP12T U1669 ( .A1(n637), .A2(n636), .ZN(n615) );
  CKND2D2BWP12T U1670 ( .A1(n616), .A2(n615), .ZN(n656) );
  CKND2BWP12T U1671 ( .I(n617), .ZN(n619) );
  XOR3XD4BWP12T U1672 ( .A1(n620), .A2(n619), .A3(n618), .Z(n655) );
  INVD1BWP12T U1673 ( .I(n653), .ZN(n624) );
  XOR3D2BWP12T U1674 ( .A1(n656), .A2(n655), .A3(n624), .Z(n789) );
  INVD1P75BWP12T U1675 ( .I(n789), .ZN(n646) );
  INVD1BWP12T U1676 ( .I(n625), .ZN(n626) );
  XNR3XD4BWP12T U1677 ( .A1(n628), .A2(n627), .A3(n626), .ZN(n790) );
  XNR2D2BWP12T U1678 ( .A1(n4511), .A2(n5054), .ZN(n796) );
  XNR2D2BWP12T U1679 ( .A1(n3495), .A2(n1007), .ZN(n2115) );
  XOR3XD4BWP12T U1680 ( .A1(n635), .A2(n634), .A3(n633), .Z(n766) );
  CKND3BWP12T U1681 ( .I(n636), .ZN(n639) );
  INVD1P25BWP12T U1682 ( .I(n637), .ZN(n638) );
  XOR3XD4BWP12T U1683 ( .A1(n640), .A2(n639), .A3(n638), .Z(n765) );
  INVD1BWP12T U1684 ( .I(n765), .ZN(n642) );
  TPOAI21D1BWP12T U1685 ( .A1(n643), .A2(n642), .B(n641), .ZN(n791) );
  ND2D1BWP12T U1686 ( .A1(n790), .A2(n791), .ZN(n644) );
  TPOAI21D2BWP12T U1687 ( .A1(n646), .A2(n645), .B(n644), .ZN(n779) );
  TPNR2D1BWP12T U1688 ( .A1(n777), .A2(n778), .ZN(n651) );
  ND2D1BWP12T U1689 ( .A1(n777), .A2(n778), .ZN(n650) );
  TPOAI21D1BWP12T U1690 ( .A1(n776), .A2(n651), .B(n650), .ZN(n1829) );
  CKND2BWP12T U1691 ( .I(n656), .ZN(n652) );
  TPND2D2BWP12T U1692 ( .A1(n655), .A2(n652), .ZN(n654) );
  TPND2D2BWP12T U1693 ( .A1(n654), .A2(n653), .ZN(n659) );
  TPND2D2BWP12T U1694 ( .A1(n657), .A2(n656), .ZN(n658) );
  TPND2D4BWP12T U1695 ( .A1(n659), .A2(n658), .ZN(n775) );
  CKND3BWP12T U1696 ( .I(n660), .ZN(n664) );
  INVD1P75BWP12T U1697 ( .I(n661), .ZN(n662) );
  XOR3XD4BWP12T U1698 ( .A1(n664), .A2(n663), .A3(n662), .Z(n772) );
  TPOAI22D2BWP12T U1699 ( .A1(n2479), .A2(n665), .B1(n2005), .B2(n706), .ZN(
        n699) );
  XNR2D1BWP12T U1700 ( .A1(n3016), .A2(n4568), .ZN(n669) );
  TPOAI22D2BWP12T U1701 ( .A1(n2529), .A2(n669), .B1(n2), .B2(n668), .ZN(n698)
         );
  INVD1BWP12T U1702 ( .I(n4568), .ZN(n4975) );
  IND2D1BWP12T U1703 ( .A1(b[0]), .B1(n4568), .ZN(n672) );
  TPOAI22D2BWP12T U1704 ( .A1(n2529), .A2(n4975), .B1(n2527), .B2(n672), .ZN(
        n702) );
  XOR3XD4BWP12T U1705 ( .A1(n700), .A2(n702), .A3(n704), .Z(n712) );
  INVD1P75BWP12T U1706 ( .I(n676), .ZN(n677) );
  BUFFXD4BWP12T U1707 ( .I(b[23]), .Z(n4920) );
  XNR2D1BWP12T U1708 ( .A1(n436), .A2(n4920), .ZN(n692) );
  TPOAI22D1BWP12T U1709 ( .A1(n2523), .A2(n679), .B1(n692), .B2(n2521), .ZN(
        n685) );
  INVD1BWP12T U1710 ( .I(n688), .ZN(n682) );
  XNR3XD4BWP12T U1711 ( .A1(n687), .A2(n685), .A3(n682), .ZN(n715) );
  XNR3XD4BWP12T U1712 ( .A1(n713), .A2(n712), .A3(n715), .ZN(n774) );
  RCOAI21D2BWP12T U1713 ( .A1(n775), .A2(n772), .B(n774), .ZN(n684) );
  ND2D3BWP12T U1714 ( .A1(n772), .A2(n775), .ZN(n683) );
  TPND2D3BWP12T U1715 ( .A1(n684), .A2(n683), .ZN(n1830) );
  OAI21D1BWP12T U1716 ( .A1(n688), .A2(n687), .B(n685), .ZN(n686) );
  BUFFD8BWP12T U1717 ( .I(a[26]), .Z(n4943) );
  ND2XD4BWP12T U1718 ( .A1(n1679), .A2(n1731), .ZN(n2462) );
  XNR2D1BWP12T U1719 ( .A1(n436), .A2(n4655), .ZN(n1683) );
  XNR2D1BWP12T U1720 ( .A1(n4565), .A2(n3899), .ZN(n1693) );
  TPOAI22D1BWP12T U1721 ( .A1(n2575), .A2(n694), .B1(n1907), .B2(n1736), .ZN(
        n1727) );
  TPOAI21D1BWP12T U1722 ( .A1(n699), .A2(n698), .B(n58), .ZN(n697) );
  TPNR2D1BWP12T U1723 ( .A1(n702), .A2(n701), .ZN(n705) );
  INVD1BWP12T U1724 ( .I(n702), .ZN(n703) );
  XNR2D1BWP12T U1725 ( .A1(n4502), .A2(n5264), .ZN(n1692) );
  INVD1BWP12T U1726 ( .I(n712), .ZN(n714) );
  RCOAI21D1BWP12T U1727 ( .A1(n715), .A2(n714), .B(n713), .ZN(n717) );
  ND2D1BWP12T U1728 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR3XD4BWP12T U1729 ( .A1(n1825), .A2(n1822), .A3(n1824), .Z(n1828) );
  XOR3XD4BWP12T U1730 ( .A1(n1829), .A2(n1830), .A3(n1828), .Z(n1843) );
  XOR3D2BWP12T U1731 ( .A1(n723), .A2(n722), .A3(n721), .Z(n833) );
  INVD2BWP12T U1732 ( .I(b[20]), .ZN(n724) );
  TPOAI22D1BWP12T U1733 ( .A1(n808), .A2(n1969), .B1(n725), .B2(n3015), .ZN(
        n806) );
  XNR2D2BWP12T U1734 ( .A1(a[17]), .A2(n4301), .ZN(n823) );
  TPNR2D1BWP12T U1735 ( .A1(n833), .A2(n835), .ZN(n734) );
  OR2XD1BWP12T U1736 ( .A1(b[0]), .A2(n3887), .Z(n727) );
  ND2D1BWP12T U1737 ( .A1(n903), .A2(n904), .ZN(n731) );
  XNR2D2BWP12T U1738 ( .A1(n436), .A2(n4732), .ZN(n812) );
  TPOAI22D1BWP12T U1739 ( .A1(n2523), .A2(n812), .B1(n2521), .B2(n729), .ZN(
        n901) );
  INVD0BWP12T U1740 ( .I(n834), .ZN(n733) );
  TPOAI21D2BWP12T U1741 ( .A1(n734), .A2(n733), .B(n732), .ZN(n792) );
  TPOAI22D1BWP12T U1742 ( .A1(n2575), .A2(n795), .B1(n1907), .B2(n735), .ZN(
        n749) );
  XNR2D1BWP12T U1743 ( .A1(n3948), .A2(n4565), .ZN(n797) );
  TPOAI22D2BWP12T U1744 ( .A1(n2573), .A2(n797), .B1(n2571), .B2(n736), .ZN(
        n748) );
  XNR2D1BWP12T U1745 ( .A1(n4502), .A2(n3930), .ZN(n807) );
  OAI22D1BWP12T U1746 ( .A1(n2535), .A2(n807), .B1(n2533), .B2(n737), .ZN(n747) );
  XNR3XD4BWP12T U1747 ( .A1(n740), .A2(n739), .A3(n738), .ZN(n794) );
  TPND2D2BWP12T U1748 ( .A1(n792), .A2(n463), .ZN(n742) );
  CKND2D2BWP12T U1749 ( .A1(n793), .A2(n794), .ZN(n741) );
  TPND2D2BWP12T U1750 ( .A1(n742), .A2(n741), .ZN(n848) );
  CKND2BWP12T U1751 ( .I(n848), .ZN(n743) );
  XOR3XD4BWP12T U1752 ( .A1(n753), .A2(n752), .A3(n751), .Z(n895) );
  XNR2D1BWP12T U1753 ( .A1(n3911), .A2(n4826), .ZN(n830) );
  ND2D1BWP12T U1754 ( .A1(n898), .A2(n897), .ZN(n760) );
  XNR2XD2BWP12T U1755 ( .A1(n2123), .A2(n5264), .ZN(n824) );
  TPND2D1BWP12T U1756 ( .A1(n899), .A2(n897), .ZN(n759) );
  ND3XD3BWP12T U1757 ( .A1(n760), .A2(n758), .A3(n759), .ZN(n896) );
  TPNR2D2BWP12T U1758 ( .A1(n895), .A2(n896), .ZN(n762) );
  TPOAI21D4BWP12T U1759 ( .A1(n894), .A2(n762), .B(n761), .ZN(n1650) );
  CKND3BWP12T U1760 ( .I(n763), .ZN(n764) );
  ND2D1BWP12T U1761 ( .A1(n1650), .A2(n427), .ZN(n767) );
  TPND2D3BWP12T U1762 ( .A1(n771), .A2(n770), .ZN(n787) );
  CKND3BWP12T U1763 ( .I(n772), .ZN(n773) );
  XOR3XD4BWP12T U1764 ( .A1(n775), .A2(n774), .A3(n773), .Z(n788) );
  INVD3BWP12T U1765 ( .I(n788), .ZN(n783) );
  OR2XD1BWP12T U1766 ( .A1(n787), .A2(n783), .Z(n782) );
  XNR3XD4BWP12T U1767 ( .A1(n778), .A2(n777), .A3(n776), .ZN(n780) );
  XOR3XD4BWP12T U1768 ( .A1(n781), .A2(n780), .A3(n779), .Z(n786) );
  CKND2D2BWP12T U1769 ( .A1(n782), .A2(n440), .ZN(n785) );
  ND2D1BWP12T U1770 ( .A1(n787), .A2(n783), .ZN(n784) );
  TPND2D3BWP12T U1771 ( .A1(n785), .A2(n784), .ZN(n1676) );
  NR2XD3BWP12T U1772 ( .A1(n426), .A2(n1676), .ZN(n3125) );
  XNR3XD4BWP12T U1773 ( .A1(n788), .A2(n787), .A3(n786), .ZN(n1674) );
  XOR3D2BWP12T U1774 ( .A1(n791), .A2(n790), .A3(n789), .Z(n857) );
  INVD1BWP12T U1775 ( .I(n857), .ZN(n851) );
  XOR3XD4BWP12T U1776 ( .A1(n794), .A2(n793), .A3(n792), .Z(n921) );
  TPOAI22D2BWP12T U1777 ( .A1(n861), .A2(n2575), .B1(n795), .B2(n1907), .ZN(
        n821) );
  TPOAI22D2BWP12T U1778 ( .A1(n1689), .A2(n828), .B1(n2115), .B2(n796), .ZN(
        n822) );
  XNR2D1BWP12T U1779 ( .A1(n5196), .A2(n4565), .ZN(n829) );
  TPOAI22D1BWP12T U1780 ( .A1(n2573), .A2(n829), .B1(n2571), .B2(n797), .ZN(
        n820) );
  IOA21D2BWP12T U1781 ( .A1(n799), .A2(n798), .B(n820), .ZN(n801) );
  TPND2D2BWP12T U1782 ( .A1(n801), .A2(n800), .ZN(n840) );
  FA1D2BWP12T U1783 ( .A(n804), .B(n803), .CI(n802), .CO(n763), .S(n838) );
  HA1D2BWP12T U1784 ( .A(n806), .B(n805), .CO(n835), .S(n858) );
  XNR2D2BWP12T U1785 ( .A1(n1858), .A2(n3899), .ZN(n862) );
  NR2XD1BWP12T U1786 ( .A1(n809), .A2(n2314), .ZN(n869) );
  INVD1BWP12T U1787 ( .I(n869), .ZN(n810) );
  XNR2D2BWP12T U1788 ( .A1(n436), .A2(n4794), .ZN(n872) );
  TPND2D2BWP12T U1789 ( .A1(n815), .A2(n814), .ZN(n859) );
  TPOAI21D1BWP12T U1790 ( .A1(n858), .A2(n860), .B(n859), .ZN(n816) );
  IOA21D2BWP12T U1791 ( .A1(n858), .A2(n860), .B(n816), .ZN(n839) );
  ND2D1BWP12T U1792 ( .A1(n838), .A2(n840), .ZN(n817) );
  TPND2D2BWP12T U1793 ( .A1(n818), .A2(n817), .ZN(n922) );
  TPNR2D1BWP12T U1794 ( .A1(n921), .A2(n922), .ZN(n819) );
  INVD1BWP12T U1795 ( .I(n819), .ZN(n845) );
  XOR3XD4BWP12T U1796 ( .A1(n822), .A2(n821), .A3(n820), .Z(n1607) );
  XNR2XD4BWP12T U1797 ( .A1(n4822), .A2(n1906), .ZN(n2022) );
  XNR2D1BWP12T U1798 ( .A1(n5079), .A2(n3930), .ZN(n870) );
  OR2D2BWP12T U1799 ( .A1(n879), .A2(n880), .Z(n825) );
  ND2D3BWP12T U1800 ( .A1(n825), .A2(n878), .ZN(n827) );
  ND2D4BWP12T U1801 ( .A1(n827), .A2(n826), .ZN(n1609) );
  XNR2D1BWP12T U1802 ( .A1(n4511), .A2(n5085), .ZN(n1505) );
  TPOAI22D1BWP12T U1803 ( .A1(n1689), .A2(n1505), .B1(n2481), .B2(n828), .ZN(
        n887) );
  TPOAI22D2BWP12T U1804 ( .A1(n2573), .A2(n882), .B1(n2571), .B2(n829), .ZN(
        n886) );
  XNR2D2BWP12T U1805 ( .A1(n5030), .A2(n32), .ZN(n871) );
  DEL025D1BWP12T U1806 ( .I(n2005), .Z(n2477) );
  TPOAI22D1BWP12T U1807 ( .A1(n52), .A2(n871), .B1(n2477), .B2(n830), .ZN(n885) );
  RCOAI21D2BWP12T U1808 ( .A1(n1607), .A2(n1609), .B(n1608), .ZN(n832) );
  XOR3XD4BWP12T U1809 ( .A1(n835), .A2(n834), .A3(n833), .Z(n1603) );
  INVD1BWP12T U1810 ( .I(n1603), .ZN(n836) );
  XOR3XD4BWP12T U1811 ( .A1(n840), .A2(n839), .A3(n838), .Z(n1601) );
  ND2D2BWP12T U1812 ( .A1(n841), .A2(n1601), .ZN(n843) );
  ND2D1BWP12T U1813 ( .A1(n1602), .A2(n1603), .ZN(n842) );
  TPAOI21D2BWP12T U1814 ( .A1(n845), .A2(n920), .B(n844), .ZN(n856) );
  TPND2D1BWP12T U1815 ( .A1(n851), .A2(n856), .ZN(n849) );
  XOR3XD4BWP12T U1816 ( .A1(n848), .A2(n847), .A3(n846), .Z(n855) );
  TPND2D2BWP12T U1817 ( .A1(n849), .A2(n855), .ZN(n853) );
  IND2D2BWP12T U1818 ( .A1(n851), .B1(n850), .ZN(n852) );
  TPNR2D3BWP12T U1819 ( .A1(n1674), .A2(n1673), .ZN(n854) );
  XNR3XD4BWP12T U1820 ( .A1(n857), .A2(n856), .A3(n855), .ZN(n1672) );
  INVD2BWP12T U1821 ( .I(n1672), .ZN(n927) );
  XOR3D2BWP12T U1822 ( .A1(n1650), .A2(n427), .A3(n1648), .Z(n925) );
  XOR3D2BWP12T U1823 ( .A1(n860), .A2(n859), .A3(n858), .Z(n1631) );
  TPOAI22D2BWP12T U1824 ( .A1(n2575), .A2(n1502), .B1(n861), .B2(n1907), .ZN(
        n909) );
  DCCKND4BWP12T U1825 ( .I(n2535), .ZN(n1185) );
  CKND3BWP12T U1826 ( .I(n1503), .ZN(n864) );
  NR2D2BWP12T U1827 ( .A1(n862), .A2(n1268), .ZN(n863) );
  RCAOI21D4BWP12T U1828 ( .A1(n1185), .A2(n864), .B(n863), .ZN(n908) );
  TPOAI22D2BWP12T U1829 ( .A1(n866), .A2(n3015), .B1(n1426), .B2(n1969), .ZN(
        n1443) );
  CKND2D2BWP12T U1830 ( .A1(n1444), .A2(n1443), .ZN(n905) );
  XOR3XD4BWP12T U1831 ( .A1(n869), .A2(n868), .A3(n867), .Z(n1574) );
  BUFFD4BWP12T U1832 ( .I(n1574), .Z(n875) );
  XNR2D1BWP12T U1833 ( .A1(n5079), .A2(n3899), .ZN(n1446) );
  TPOAI22D1BWP12T U1834 ( .A1(n2467), .A2(n1446), .B1(n870), .B2(n1799), .ZN(
        n1511) );
  OAI22D1BWP12T U1835 ( .A1(n871), .A2(n2005), .B1(n2479), .B2(n1485), .ZN(
        n1510) );
  XNR2D1BWP12T U1836 ( .A1(n436), .A2(n4826), .ZN(n1427) );
  OAI21D1BWP12T U1837 ( .A1(n1511), .A2(n1510), .B(n1512), .ZN(n874) );
  ND2D1BWP12T U1838 ( .A1(n1511), .A2(n1510), .ZN(n873) );
  ND2D1BWP12T U1839 ( .A1(n874), .A2(n873), .ZN(n1573) );
  ND2D3BWP12T U1840 ( .A1(n1572), .A2(n875), .ZN(n876) );
  TPND2D2BWP12T U1841 ( .A1(n877), .A2(n876), .ZN(n1630) );
  XNR3XD4BWP12T U1842 ( .A1(n880), .A2(n879), .A3(n878), .ZN(n1582) );
  INVD1BWP12T U1843 ( .I(n4565), .ZN(n3890) );
  IND2D1BWP12T U1844 ( .A1(b[0]), .B1(n4565), .ZN(n881) );
  XNR2D1BWP12T U1845 ( .A1(n3016), .A2(n4565), .ZN(n883) );
  TPOAI22D2BWP12T U1846 ( .A1(n2573), .A2(n883), .B1(n2571), .B2(n882), .ZN(
        n1424) );
  XNR2XD2BWP12T U1847 ( .A1(n2123), .A2(n5237), .ZN(n1449) );
  TPOAI22D1BWP12T U1848 ( .A1(n2471), .A2(n1449), .B1(n2469), .B2(n884), .ZN(
        n1423) );
  FA1D2BWP12T U1849 ( .A(n887), .B(n886), .CI(n885), .CO(n1608), .S(n888) );
  INVD1P75BWP12T U1850 ( .I(n888), .ZN(n1580) );
  ND2D1BWP12T U1851 ( .A1(n889), .A2(n1581), .ZN(n890) );
  OAI21D1BWP12T U1852 ( .A1(n891), .A2(n1580), .B(n890), .ZN(n1629) );
  OAI21D1BWP12T U1853 ( .A1(n1631), .A2(n1630), .B(n1629), .ZN(n893) );
  ND2D1BWP12T U1854 ( .A1(n1631), .A2(n1630), .ZN(n892) );
  TPND2D2BWP12T U1855 ( .A1(n893), .A2(n892), .ZN(n1621) );
  XNR3XD4BWP12T U1856 ( .A1(n896), .A2(n895), .A3(n894), .ZN(n1622) );
  XNR2D2BWP12T U1857 ( .A1(n897), .A2(n898), .ZN(n900) );
  XNR2XD4BWP12T U1858 ( .A1(n900), .A2(n899), .ZN(n1604) );
  INVD1BWP12T U1859 ( .I(n1604), .ZN(n915) );
  INVD1P75BWP12T U1860 ( .I(n901), .ZN(n902) );
  XNR3XD4BWP12T U1861 ( .A1(n904), .A2(n903), .A3(n902), .ZN(n1605) );
  CKND3BWP12T U1862 ( .I(n905), .ZN(n907) );
  IND2D2BWP12T U1863 ( .A1(n909), .B1(n908), .ZN(n906) );
  CKND2D2BWP12T U1864 ( .A1(n907), .A2(n906), .ZN(n912) );
  TPND2D2BWP12T U1865 ( .A1(n912), .A2(n911), .ZN(n1606) );
  TPNR2D1BWP12T U1866 ( .A1(n1605), .A2(n1606), .ZN(n914) );
  ND2D1BWP12T U1867 ( .A1(n1606), .A2(n1605), .ZN(n913) );
  TPOAI21D2BWP12T U1868 ( .A1(n915), .A2(n914), .B(n913), .ZN(n1623) );
  IND2D2BWP12T U1869 ( .A1(n1622), .B1(n916), .ZN(n917) );
  ND2D1BWP12T U1870 ( .A1(n1622), .A2(n1623), .ZN(n918) );
  XOR3XD4BWP12T U1871 ( .A1(n922), .A2(n921), .A3(n920), .Z(n1651) );
  ND2D1BWP12T U1872 ( .A1(n1651), .A2(n923), .ZN(n924) );
  IOA21D2BWP12T U1873 ( .A1(n925), .A2(n1652), .B(n924), .ZN(n1671) );
  INVD1P75BWP12T U1874 ( .I(n1671), .ZN(n926) );
  TPND2D2BWP12T U1875 ( .A1(n927), .A2(n926), .ZN(n3130) );
  BUFFXD8BWP12T U1876 ( .I(a[1]), .Z(n4501) );
  XNR2XD2BWP12T U1877 ( .A1(n4501), .A2(n5196), .ZN(n930) );
  XNR2XD4BWP12T U1878 ( .A1(n4501), .A2(n3948), .ZN(n944) );
  TPOAI22D2BWP12T U1879 ( .A1(n930), .A2(n1969), .B1(n3015), .B2(n944), .ZN(
        n947) );
  XNR2XD2BWP12T U1880 ( .A1(b[1]), .A2(n3570), .ZN(n945) );
  TPOAI22D2BWP12T U1881 ( .A1(n2523), .A2(n928), .B1(n2521), .B2(n945), .ZN(
        n946) );
  BUFFD2BWP12T U1882 ( .I(a[3]), .Z(n3570) );
  IND2D1BWP12T U1883 ( .A1(b[0]), .B1(n436), .ZN(n929) );
  OAI22D1BWP12T U1884 ( .A1(n2523), .A2(n512), .B1(n2521), .B2(n929), .ZN(n940) );
  OR2XD4BWP12T U1885 ( .A1(n939), .A2(n940), .Z(n2729) );
  TPND2D1BWP12T U1886 ( .A1(n932), .A2(n931), .ZN(n3013) );
  TPNR2D2BWP12T U1887 ( .A1(n932), .A2(n931), .ZN(n3014) );
  INVD1BWP12T U1888 ( .I(n3014), .ZN(n936) );
  TPOAI22D1BWP12T U1889 ( .A1(n1969), .A2(n3016), .B1(n933), .B2(n3015), .ZN(
        n3018) );
  INVD1P75BWP12T U1890 ( .I(n3018), .ZN(n935) );
  INVD1BWP12T U1891 ( .I(n3017), .ZN(n934) );
  TPNR2D2BWP12T U1892 ( .A1(n935), .A2(n934), .ZN(n3019) );
  INVD1P75BWP12T U1893 ( .I(n940), .ZN(n941) );
  TPAOI21D2BWP12T U1894 ( .A1(n2729), .A2(n2731), .B(n2730), .ZN(n3027) );
  INVD1BWP12T U1895 ( .I(n3016), .ZN(n943) );
  XNR2XD4BWP12T U1896 ( .A1(n4301), .A2(a[1]), .ZN(n953) );
  TPOAI22D2BWP12T U1897 ( .A1(n944), .A2(n1969), .B1(n953), .B2(n3015), .ZN(
        n956) );
  TPOAI22D1BWP12T U1898 ( .A1(n2523), .A2(n945), .B1(n2521), .B2(n949), .ZN(
        n954) );
  XOR3XD4BWP12T U1899 ( .A1(n955), .A2(n956), .A3(n954), .Z(n961) );
  HA1D2BWP12T U1900 ( .A(n947), .B(n946), .CO(n960), .S(n939) );
  ND2D3BWP12T U1901 ( .A1(n961), .A2(n960), .ZN(n3025) );
  TPND2D2BWP12T U1902 ( .A1(n3027), .A2(n3025), .ZN(n966) );
  XNR2D2BWP12T U1903 ( .A1(n3911), .A2(b[1]), .ZN(n971) );
  TPOAI22D2BWP12T U1904 ( .A1(n948), .A2(n2479), .B1(n2005), .B2(n971), .ZN(
        n979) );
  XNR2D1BWP12T U1905 ( .A1(n3948), .A2(n3570), .ZN(n967) );
  TPOAI22D2BWP12T U1906 ( .A1(n2523), .A2(n949), .B1(n2521), .B2(n967), .ZN(
        n978) );
  IND2D1BWP12T U1907 ( .A1(b[0]), .B1(n3911), .ZN(n952) );
  TPOAI21D2BWP12T U1908 ( .A1(n2005), .A2(n952), .B(n951), .ZN(n969) );
  XNR2D2BWP12T U1909 ( .A1(n5033), .A2(a[1]), .ZN(n968) );
  TPOAI22D2BWP12T U1910 ( .A1(n968), .A2(n3015), .B1(n953), .B2(n2476), .ZN(
        n970) );
  XOR3XD4BWP12T U1911 ( .A1(n979), .A2(n978), .A3(n974), .Z(n963) );
  CKND3BWP12T U1912 ( .I(n954), .ZN(n959) );
  TPNR2D2BWP12T U1913 ( .A1(n956), .A2(n955), .ZN(n958) );
  ND2D2BWP12T U1914 ( .A1(n956), .A2(n955), .ZN(n957) );
  TPOAI21D2BWP12T U1915 ( .A1(n959), .A2(n958), .B(n957), .ZN(n962) );
  TPNR2D3BWP12T U1916 ( .A1(n963), .A2(n962), .ZN(n3023) );
  DCCKND4BWP12T U1917 ( .I(n3023), .ZN(n965) );
  OR2XD4BWP12T U1918 ( .A1(n961), .A2(n960), .Z(n3024) );
  XNR2D1BWP12T U1919 ( .A1(n4301), .A2(n436), .ZN(n989) );
  OAI22D1BWP12T U1920 ( .A1(n967), .A2(n2523), .B1(n989), .B2(n2521), .ZN(n992) );
  TPOAI22D2BWP12T U1921 ( .A1(n982), .A2(n3015), .B1(n968), .B2(n1969), .ZN(
        n994) );
  XNR2XD4BWP12T U1922 ( .A1(n994), .A2(n993), .ZN(n973) );
  CKAN2D2BWP12T U1923 ( .A1(n969), .A2(n970), .Z(n998) );
  XNR2D2BWP12T U1924 ( .A1(n3911), .A2(n5196), .ZN(n985) );
  OAI22D1BWP12T U1925 ( .A1(n2479), .A2(n971), .B1(n2005), .B2(n985), .ZN(n997) );
  XNR2D2BWP12T U1926 ( .A1(n998), .A2(n997), .ZN(n972) );
  XOR3XD4BWP12T U1927 ( .A1(n992), .A2(n973), .A3(n972), .Z(n981) );
  CKND3BWP12T U1928 ( .I(n978), .ZN(n976) );
  CKND3BWP12T U1929 ( .I(n979), .ZN(n975) );
  IOA21D2BWP12T U1930 ( .A1(n979), .A2(n978), .B(n977), .ZN(n980) );
  TPND2D2BWP12T U1931 ( .A1(n981), .A2(n980), .ZN(n3009) );
  TPOAI22D2BWP12T U1932 ( .A1(n2479), .A2(n985), .B1(n2005), .B2(n1009), .ZN(
        n1010) );
  XNR2XD4BWP12T U1933 ( .A1(n1011), .A2(n1010), .ZN(n1043) );
  OAI21D1BWP12T U1934 ( .A1(n993), .A2(n994), .B(n992), .ZN(n987) );
  ND2D1BWP12T U1935 ( .A1(n994), .A2(n993), .ZN(n986) );
  TPND2D2BWP12T U1936 ( .A1(n987), .A2(n986), .ZN(n1044) );
  IND2D1BWP12T U1937 ( .A1(b[0]), .B1(n2123), .ZN(n988) );
  TPOAI22D1BWP12T U1938 ( .A1(n2469), .A2(n988), .B1(n2020), .B2(n437), .ZN(
        n1030) );
  XNR2D1BWP12T U1939 ( .A1(n436), .A2(n5033), .ZN(n1026) );
  TPOAI22D1BWP12T U1940 ( .A1(n2523), .A2(n989), .B1(n2521), .B2(n1026), .ZN(
        n1029) );
  BUFFD2BWP12T U1941 ( .I(n1007), .Z(n4510) );
  XNR2XD4BWP12T U1942 ( .A1(n4510), .A2(b[1]), .ZN(n1008) );
  TPOAI22D1BWP12T U1943 ( .A1(n2020), .A2(n990), .B1(n2469), .B2(n1008), .ZN(
        n1031) );
  INVD1BWP12T U1944 ( .I(n1031), .ZN(n991) );
  XOR3XD4BWP12T U1945 ( .A1(n1030), .A2(n1029), .A3(n991), .Z(n1046) );
  XOR3D2BWP12T U1946 ( .A1(n994), .A2(n993), .A3(n992), .Z(n996) );
  OR2D2BWP12T U1947 ( .A1(n998), .A2(n997), .Z(n995) );
  TPND2D1BWP12T U1948 ( .A1(n996), .A2(n995), .ZN(n1000) );
  ND2D1BWP12T U1949 ( .A1(n998), .A2(n997), .ZN(n999) );
  TPND2D2BWP12T U1950 ( .A1(n1000), .A2(n999), .ZN(n1004) );
  INVD1P75BWP12T U1951 ( .I(n1004), .ZN(n1001) );
  CKND3BWP12T U1952 ( .I(n1003), .ZN(n1005) );
  ND2XD3BWP12T U1953 ( .A1(n1005), .A2(n1004), .ZN(n2626) );
  XNR2D1BWP12T U1954 ( .A1(n5196), .A2(n71), .ZN(n1020) );
  TPOAI22D1BWP12T U1955 ( .A1(n2020), .A2(n1008), .B1(n14), .B2(n1020), .ZN(
        n1038) );
  TPOAI22D1BWP12T U1956 ( .A1(n2479), .A2(n1009), .B1(n1022), .B2(n2005), .ZN(
        n1039) );
  CKND2BWP12T U1957 ( .I(n1010), .ZN(n1012) );
  NR2XD0BWP12T U1958 ( .A1(n1012), .A2(n1011), .ZN(n1037) );
  CKND2BWP12T U1959 ( .I(n1038), .ZN(n1014) );
  CKND2BWP12T U1960 ( .I(n1039), .ZN(n1013) );
  TPND2D1BWP12T U1961 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  TPND2D1BWP12T U1962 ( .A1(n1037), .A2(n1015), .ZN(n1016) );
  IOA21D2BWP12T U1963 ( .A1(n1038), .A2(n1039), .B(n1016), .ZN(n1070) );
  INVD1BWP12T U1964 ( .I(n4511), .ZN(n3898) );
  IND2D1BWP12T U1965 ( .A1(b[0]), .B1(n4511), .ZN(n1017) );
  XNR2D2BWP12T U1966 ( .A1(n436), .A2(n4896), .ZN(n1025) );
  XNR2D1BWP12T U1967 ( .A1(n436), .A2(n3938), .ZN(n1059) );
  OAI22D1BWP12T U1968 ( .A1(n2523), .A2(n1025), .B1(n2521), .B2(n1059), .ZN(
        n1061) );
  XNR2D1BWP12T U1969 ( .A1(n3016), .A2(n4511), .ZN(n1018) );
  XNR2XD2BWP12T U1970 ( .A1(b[1]), .A2(n4511), .ZN(n1050) );
  XNR3XD4BWP12T U1971 ( .A1(n1063), .A2(n1061), .A3(n1019), .ZN(n1069) );
  XOR2XD2BWP12T U1972 ( .A1(n3899), .A2(n1812), .Z(n1023) );
  TPOAI22D2BWP12T U1973 ( .A1(n1023), .A2(n1969), .B1(n1021), .B2(n3015), .ZN(
        n1058) );
  XNR2D2BWP12T U1974 ( .A1(n3911), .A2(n5033), .ZN(n1049) );
  NR2XD2BWP12T U1975 ( .A1(n3334), .A2(n2481), .ZN(n1036) );
  TPOAI22D1BWP12T U1976 ( .A1(n2523), .A2(n1026), .B1(n2521), .B2(n1025), .ZN(
        n1034) );
  OAI21D1BWP12T U1977 ( .A1(n1036), .A2(n1035), .B(n1034), .ZN(n1028) );
  CKND2D2BWP12T U1978 ( .A1(n1028), .A2(n1027), .ZN(n1052) );
  XOR3XD4BWP12T U1979 ( .A1(n1053), .A2(n1054), .A3(n1052), .Z(n1067) );
  XOR3XD4BWP12T U1980 ( .A1(n1070), .A2(n1069), .A3(n1067), .Z(n1078) );
  OAI21D1BWP12T U1981 ( .A1(n1030), .A2(n1031), .B(n1029), .ZN(n1033) );
  ND2D1BWP12T U1982 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  ND2D1BWP12T U1983 ( .A1(n1033), .A2(n1032), .ZN(n1042) );
  XOR3XD4BWP12T U1984 ( .A1(n1036), .A2(n1035), .A3(n1034), .Z(n1041) );
  XOR3D2BWP12T U1985 ( .A1(n1039), .A2(n1038), .A3(n1037), .Z(n1040) );
  TPNR2D4BWP12T U1986 ( .A1(n1078), .A2(n1077), .ZN(n2871) );
  FA1D4BWP12T U1987 ( .A(n1042), .B(n1041), .CI(n1040), .CO(n1077), .S(n1076)
         );
  NR2D0BWP12T U1988 ( .A1(n1044), .A2(n1043), .ZN(n1047) );
  ND2D1BWP12T U1989 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  TPOAI21D2BWP12T U1990 ( .A1(n1047), .A2(n1046), .B(n1045), .ZN(n1075) );
  NR2D4BWP12T U1991 ( .A1(n1076), .A2(n1075), .ZN(n2869) );
  CKND2BWP12T U1992 ( .I(n2801), .ZN(n1074) );
  XNR2D1BWP12T U1993 ( .A1(n5030), .A2(n4896), .ZN(n1113) );
  OAI22D1BWP12T U1994 ( .A1(n1049), .A2(n2479), .B1(n1113), .B2(n2005), .ZN(
        n1090) );
  XNR2D1BWP12T U1995 ( .A1(n5196), .A2(n4511), .ZN(n1103) );
  TPOAI22D1BWP12T U1996 ( .A1(n1689), .A2(n1050), .B1(n2481), .B2(n1103), .ZN(
        n1089) );
  CKND2D2BWP12T U1997 ( .A1(n1052), .A2(n462), .ZN(n1056) );
  CKND2D2BWP12T U1998 ( .A1(n1056), .A2(n1055), .ZN(n1083) );
  HA1D2BWP12T U1999 ( .A(n1058), .B(n1057), .CO(n1092), .S(n1054) );
  TPOAI22D2BWP12T U2000 ( .A1(n1105), .A2(n3015), .B1(n3930), .B2(n1969), .ZN(
        n1099) );
  TPOAI22D2BWP12T U2001 ( .A1(n2521), .A2(n1108), .B1(n1059), .B2(n2523), .ZN(
        n1097) );
  CKND3BWP12T U2002 ( .I(n1097), .ZN(n1060) );
  XNR3XD4BWP12T U2003 ( .A1(n1098), .A2(n1099), .A3(n1060), .ZN(n1091) );
  TPOAI21D0BWP12T U2004 ( .A1(n1063), .A2(n1062), .B(n1061), .ZN(n1065) );
  CKND2D0BWP12T U2005 ( .A1(n1063), .A2(n1062), .ZN(n1064) );
  CKAN2D2BWP12T U2006 ( .A1(n1065), .A2(n1064), .Z(n1095) );
  XOR3XD4BWP12T U2007 ( .A1(n1092), .A2(n1091), .A3(n1095), .Z(n1087) );
  XOR3XD4BWP12T U2008 ( .A1(n1084), .A2(n1083), .A3(n1087), .Z(n1079) );
  INVD1BWP12T U2009 ( .I(n1069), .ZN(n1066) );
  IND2XD1BWP12T U2010 ( .A1(n1070), .B1(n1066), .ZN(n1068) );
  ND2D1BWP12T U2011 ( .A1(n1068), .A2(n1067), .ZN(n1072) );
  ND2D1BWP12T U2012 ( .A1(n1070), .A2(n1069), .ZN(n1071) );
  CKND2D2BWP12T U2013 ( .A1(n1072), .A2(n1071), .ZN(n1080) );
  INVD1BWP12T U2014 ( .I(n1080), .ZN(n1073) );
  TPND2D2BWP12T U2015 ( .A1(n1074), .A2(n447), .ZN(n1082) );
  TPND2D3BWP12T U2016 ( .A1(n1076), .A2(n1075), .ZN(n2941) );
  CKND2D2BWP12T U2017 ( .A1(n1078), .A2(n1077), .ZN(n2872) );
  TPOAI21D1BWP12T U2018 ( .A1(n2871), .A2(n2941), .B(n2872), .ZN(n2800) );
  INR2D4BWP12T U2019 ( .A1(n1080), .B1(n1079), .ZN(n2804) );
  TPAOI21D2BWP12T U2020 ( .A1(n2800), .A2(n446), .B(n2804), .ZN(n1081) );
  ND2XD3BWP12T U2021 ( .A1(n1082), .A2(n1081), .ZN(n3058) );
  DCCKND4BWP12T U2022 ( .I(n3058), .ZN(n3045) );
  NR2D1BWP12T U2023 ( .A1(n1084), .A2(n1083), .ZN(n1086) );
  ND2D1BWP12T U2024 ( .A1(n1084), .A2(n1083), .ZN(n1085) );
  FA1D2BWP12T U2025 ( .A(n1090), .B(n1089), .CI(n1088), .CO(n1147), .S(n1084)
         );
  TPNR2D1BWP12T U2026 ( .A1(n1091), .A2(n1092), .ZN(n1096) );
  INVD1BWP12T U2027 ( .I(n1091), .ZN(n1094) );
  INVD1BWP12T U2028 ( .I(n1092), .ZN(n1093) );
  TPOAI22D1BWP12T U2029 ( .A1(n1096), .A2(n1095), .B1(n1094), .B2(n1093), .ZN(
        n1148) );
  OAI21D1BWP12T U2030 ( .A1(n1098), .A2(n1099), .B(n1097), .ZN(n1101) );
  ND2D1BWP12T U2031 ( .A1(n1099), .A2(n1098), .ZN(n1100) );
  CKND2D2BWP12T U2032 ( .A1(n1101), .A2(n1100), .ZN(n1124) );
  XNR2D1BWP12T U2033 ( .A1(n3948), .A2(n4511), .ZN(n1117) );
  TPOAI22D2BWP12T U2034 ( .A1(n1689), .A2(n1103), .B1(n1117), .B2(n2481), .ZN(
        n1138) );
  TPOAI22D2BWP12T U2035 ( .A1(n1105), .A2(n1969), .B1(n1120), .B2(n3015), .ZN(
        n1119) );
  TPOAI22D2BWP12T U2036 ( .A1(n2467), .A2(n5081), .B1(n1799), .B2(n1107), .ZN(
        n1118) );
  XOR3XD4BWP12T U2037 ( .A1(n1137), .A2(n1138), .A3(n1136), .Z(n1123) );
  XNR2D2BWP12T U2038 ( .A1(n436), .A2(n3930), .ZN(n1121) );
  TPOAI22D1BWP12T U2039 ( .A1(n2523), .A2(n1108), .B1(n2521), .B2(n1121), .ZN(
        n1128) );
  XNR2D1BWP12T U2040 ( .A1(n5079), .A2(n3016), .ZN(n1112) );
  INVD1BWP12T U2041 ( .I(n1142), .ZN(n1109) );
  TPND2D2BWP12T U2042 ( .A1(n1110), .A2(n1109), .ZN(n1111) );
  XNR2D1BWP12T U2043 ( .A1(n3911), .A2(n3938), .ZN(n1141) );
  INVD1BWP12T U2044 ( .I(n1130), .ZN(n1114) );
  XNR3XD4BWP12T U2045 ( .A1(n1128), .A2(n1129), .A3(n1114), .ZN(n1125) );
  CKND3BWP12T U2046 ( .I(n1125), .ZN(n1115) );
  XNR3XD4BWP12T U2047 ( .A1(n1124), .A2(n1123), .A3(n1115), .ZN(n1144) );
  XOR3XD4BWP12T U2048 ( .A1(n1147), .A2(n1148), .A3(n1144), .Z(n1153) );
  INR2D2BWP12T U2049 ( .A1(n460), .B1(n1153), .ZN(n1116) );
  INVD1P75BWP12T U2050 ( .I(n1116), .ZN(n3056) );
  XNR2D2BWP12T U2051 ( .A1(n4301), .A2(n4511), .ZN(n1186) );
  TPOAI22D1BWP12T U2052 ( .A1(n1689), .A2(n1117), .B1(n2481), .B2(n1186), .ZN(
        n1190) );
  INVD1BWP12T U2053 ( .I(n1190), .ZN(n1122) );
  HA1D2BWP12T U2054 ( .A(n1119), .B(n1118), .CO(n1191), .S(n1136) );
  TPOAI22D4BWP12T U2055 ( .A1(n1120), .A2(n1969), .B1(n1166), .B2(n3015), .ZN(
        n1173) );
  INR2D2BWP12T U2056 ( .A1(n3016), .B1(n1268), .ZN(n1172) );
  XNR2D2BWP12T U2057 ( .A1(n436), .A2(n3939), .ZN(n1182) );
  TPOAI22D2BWP12T U2058 ( .A1(n2523), .A2(n1121), .B1(n2521), .B2(n1182), .ZN(
        n1170) );
  XOR3XD4BWP12T U2059 ( .A1(n1172), .A2(n1173), .A3(n1170), .Z(n1189) );
  XOR3XD4BWP12T U2060 ( .A1(n1122), .A2(n1191), .A3(n1189), .Z(n1195) );
  TPND2D2BWP12T U2061 ( .A1(n1127), .A2(n1126), .ZN(n1194) );
  TPOAI21D1BWP12T U2062 ( .A1(n1130), .A2(n1129), .B(n1128), .ZN(n1132) );
  ND2D1BWP12T U2063 ( .A1(n1130), .A2(n1129), .ZN(n1131) );
  ND2D2BWP12T U2064 ( .A1(n1132), .A2(n1131), .ZN(n1162) );
  CKND2BWP12T U2065 ( .I(n1138), .ZN(n1134) );
  INVD2BWP12T U2066 ( .I(n459), .ZN(n1133) );
  TPND2D2BWP12T U2067 ( .A1(n1134), .A2(n1133), .ZN(n1135) );
  TPND2D2BWP12T U2068 ( .A1(n1136), .A2(n1135), .ZN(n1140) );
  ND2D1BWP12T U2069 ( .A1(n1138), .A2(n459), .ZN(n1139) );
  TPND2D2BWP12T U2070 ( .A1(n1140), .A2(n1139), .ZN(n1163) );
  XNR2D2BWP12T U2071 ( .A1(n3911), .A2(n3899), .ZN(n1181) );
  TPOAI22D1BWP12T U2072 ( .A1(n2479), .A2(n1141), .B1(n1181), .B2(n2005), .ZN(
        n1177) );
  OAI22D1BWP12T U2073 ( .A1(n2467), .A2(n1142), .B1(n1167), .B2(n1799), .ZN(
        n1178) );
  XOR3XD4BWP12T U2074 ( .A1(n1177), .A2(n1178), .A3(n1176), .Z(n1160) );
  XOR3XD4BWP12T U2075 ( .A1(n1162), .A2(n1163), .A3(n1160), .Z(n1193) );
  XNR3XD4BWP12T U2076 ( .A1(n1195), .A2(n1194), .A3(n1193), .ZN(n1156) );
  DCCKND4BWP12T U2077 ( .I(n1156), .ZN(n1152) );
  INVD1BWP12T U2078 ( .I(n1148), .ZN(n1146) );
  INVD1BWP12T U2079 ( .I(n1147), .ZN(n1145) );
  IOA21D2BWP12T U2080 ( .A1(n1146), .A2(n1145), .B(n1144), .ZN(n1150) );
  ND2D1BWP12T U2081 ( .A1(n1148), .A2(n1147), .ZN(n1149) );
  ND2XD3BWP12T U2082 ( .A1(n1150), .A2(n1149), .ZN(n1155) );
  CKND2BWP12T U2083 ( .I(n1155), .ZN(n1151) );
  TPNR2D3BWP12T U2084 ( .A1(n1154), .A2(n460), .ZN(n3057) );
  ND2D3BWP12T U2085 ( .A1(n1156), .A2(n1155), .ZN(n3037) );
  INVD1P75BWP12T U2086 ( .I(n3037), .ZN(n1157) );
  TPAOI21D2BWP12T U2087 ( .A1(n3057), .A2(n3038), .B(n1157), .ZN(n3043) );
  TPOAI21D2BWP12T U2088 ( .A1(n3045), .A2(n3044), .B(n3043), .ZN(n1312) );
  INVD1P75BWP12T U2089 ( .I(n1163), .ZN(n1159) );
  TPND2D2BWP12T U2090 ( .A1(n1159), .A2(n1158), .ZN(n1161) );
  TPND2D2BWP12T U2091 ( .A1(n1161), .A2(n1160), .ZN(n1165) );
  ND2D1BWP12T U2092 ( .A1(n1163), .A2(n1162), .ZN(n1164) );
  XOR2XD2BWP12T U2093 ( .A1(n1812), .A2(n5054), .Z(n1223) );
  TPOAI22D1BWP12T U2094 ( .A1(n1166), .A2(n1969), .B1(n1223), .B2(n3015), .ZN(
        n1227) );
  INVD1BWP12T U2095 ( .I(n1172), .ZN(n1168) );
  CKND2D1BWP12T U2096 ( .A1(n1169), .A2(n1168), .ZN(n1171) );
  CKND2D2BWP12T U2097 ( .A1(n1171), .A2(n1170), .ZN(n1175) );
  TPND2D2BWP12T U2098 ( .A1(n1175), .A2(n1174), .ZN(n1239) );
  OAI21D1BWP12T U2099 ( .A1(n1178), .A2(n1177), .B(n1176), .ZN(n1180) );
  TPND2D2BWP12T U2100 ( .A1(n1180), .A2(n1179), .ZN(n1237) );
  XNR3XD2BWP12T U2101 ( .A1(n1238), .A2(n1239), .A3(n1237), .ZN(n1244) );
  XNR2D2BWP12T U2102 ( .A1(n3911), .A2(b[9]), .ZN(n1233) );
  TPOAI22D4BWP12T U2103 ( .A1(n2479), .A2(n1181), .B1(n2005), .B2(n1233), .ZN(
        n1216) );
  XNR2XD2BWP12T U2104 ( .A1(n2185), .A2(n5085), .ZN(n1224) );
  TPOAI22D2BWP12T U2105 ( .A1(n2523), .A2(n1182), .B1(n2521), .B2(n1224), .ZN(
        n1214) );
  IND2D1BWP12T U2106 ( .A1(b[0]), .B1(n4502), .ZN(n1183) );
  XOR3XD4BWP12T U2107 ( .A1(n1216), .A2(n1214), .A3(n1218), .Z(n1208) );
  XNR2XD8BWP12T U2108 ( .A1(n4511), .A2(n5033), .ZN(n1225) );
  XNR2D2BWP12T U2109 ( .A1(n3016), .A2(n1858), .ZN(n1229) );
  XNR2XD4BWP12T U2110 ( .A1(b[1]), .A2(n1858), .ZN(n1228) );
  TPOAI22D2BWP12T U2111 ( .A1(n2535), .A2(n1229), .B1(n2533), .B2(n1228), .ZN(
        n1188) );
  XNR2XD2BWP12T U2112 ( .A1(n2123), .A2(n3938), .ZN(n1234) );
  INVD4BWP12T U2113 ( .I(n1189), .ZN(n1203) );
  NR2D1BWP12T U2114 ( .A1(n1191), .A2(n1190), .ZN(n1202) );
  ND2D1BWP12T U2115 ( .A1(n1191), .A2(n1190), .ZN(n1204) );
  OAI21D1BWP12T U2116 ( .A1(n1203), .A2(n1202), .B(n1204), .ZN(n1192) );
  XNR3XD4BWP12T U2117 ( .A1(n1207), .A2(n1208), .A3(n1192), .ZN(n1247) );
  XNR3XD4BWP12T U2118 ( .A1(n1243), .A2(n1244), .A3(n1247), .ZN(n1302) );
  INVD1BWP12T U2119 ( .I(n1193), .ZN(n1200) );
  DEL025D1BWP12T U2120 ( .I(n1194), .Z(n1197) );
  INR2D1BWP12T U2121 ( .A1(n1195), .B1(n1197), .ZN(n1199) );
  INVD1BWP12T U2122 ( .I(n1195), .ZN(n1196) );
  ND2D1BWP12T U2123 ( .A1(n1197), .A2(n1196), .ZN(n1198) );
  TPOAI21D1BWP12T U2124 ( .A1(n1200), .A2(n1199), .B(n1198), .ZN(n1303) );
  INVD1BWP12T U2125 ( .I(n1303), .ZN(n1201) );
  TPND2D2BWP12T U2126 ( .A1(n1302), .A2(n1201), .ZN(n3062) );
  TPNR2D3BWP12T U2127 ( .A1(n1203), .A2(n1202), .ZN(n1206) );
  INVD1BWP12T U2128 ( .I(n1204), .ZN(n1205) );
  RCAOI21D4BWP12T U2129 ( .A1(n1211), .A2(n1210), .B(n1209), .ZN(n1298) );
  DEL025D1BWP12T U2130 ( .I(n1216), .Z(n1217) );
  INVD2BWP12T U2131 ( .I(n3016), .ZN(n1221) );
  XNR2D2BWP12T U2132 ( .A1(n1812), .A2(n1222), .ZN(n1278) );
  TPOAI22D2BWP12T U2133 ( .A1(n1223), .A2(n1969), .B1(n1278), .B2(n3015), .ZN(
        n1285) );
  XNR2D1BWP12T U2134 ( .A1(n436), .A2(n5237), .ZN(n1275) );
  TPOAI22D1BWP12T U2135 ( .A1(n2523), .A2(n1224), .B1(n2521), .B2(n1275), .ZN(
        n1283) );
  XOR3XD4BWP12T U2136 ( .A1(n1284), .A2(n1285), .A3(n1283), .Z(n1293) );
  TPOAI22D4BWP12T U2137 ( .A1(n1689), .A2(n1225), .B1(n1276), .B2(n2481), .ZN(
        n1263) );
  XNR2XD8BWP12T U2138 ( .A1(n6), .A2(n5196), .ZN(n1269) );
  TPOAI22D2BWP12T U2139 ( .A1(n2535), .A2(n1228), .B1(n1269), .B2(n396), .ZN(
        n1264) );
  HA1D1BWP12T U2140 ( .A(n1227), .B(n1226), .CO(n1266), .S(n1238) );
  XOR3D2BWP12T U2141 ( .A1(n1263), .A2(n1264), .A3(n1266), .Z(n1291) );
  XOR3XD4BWP12T U2142 ( .A1(n1292), .A2(n1293), .A3(n1291), .Z(n1299) );
  IOA21D2BWP12T U2143 ( .A1(n1232), .A2(n1231), .B(n1230), .ZN(n1254) );
  INVD1P75BWP12T U2144 ( .I(n1254), .ZN(n1252) );
  XNR2D2BWP12T U2145 ( .A1(n3911), .A2(n3939), .ZN(n1274) );
  TPOAI22D2BWP12T U2146 ( .A1(n1233), .A2(n2479), .B1(n1274), .B2(n2005), .ZN(
        n1260) );
  XNR2XD2BWP12T U2147 ( .A1(n2123), .A2(n3899), .ZN(n1271) );
  XNR2XD2BWP12T U2148 ( .A1(n5079), .A2(n4301), .ZN(n1279) );
  TPOAI22D1BWP12T U2149 ( .A1(n2467), .A2(n1235), .B1(n1799), .B2(n1279), .ZN(
        n1259) );
  INVD1BWP12T U2150 ( .I(n1259), .ZN(n1236) );
  XOR3XD4BWP12T U2151 ( .A1(n1260), .A2(n1258), .A3(n1236), .Z(n1253) );
  INVD2P3BWP12T U2152 ( .I(n1237), .ZN(n1242) );
  ND2D1BWP12T U2153 ( .A1(n1239), .A2(n1238), .ZN(n1240) );
  TPOAI21D4BWP12T U2154 ( .A1(n1242), .A2(n1241), .B(n1240), .ZN(n1251) );
  XOR3XD4BWP12T U2155 ( .A1(n1252), .A2(n1253), .A3(n1251), .Z(n1297) );
  XOR3XD4BWP12T U2156 ( .A1(n1298), .A2(n1299), .A3(n1297), .Z(n1305) );
  CKND3BWP12T U2157 ( .I(n1305), .ZN(n1250) );
  INVD2BWP12T U2158 ( .I(n1244), .ZN(n1245) );
  ND2D1BWP12T U2159 ( .A1(n1255), .A2(n1254), .ZN(n1256) );
  TPND2D2BWP12T U2160 ( .A1(n1257), .A2(n1256), .ZN(n1410) );
  ND2D1BWP12T U2161 ( .A1(n1259), .A2(n1260), .ZN(n1262) );
  OAI21D1BWP12T U2162 ( .A1(n1259), .A2(n1260), .B(n1258), .ZN(n1261) );
  CKND2D2BWP12T U2163 ( .A1(n1262), .A2(n1261), .ZN(n1341) );
  AN2XD2BWP12T U2164 ( .A1(n1264), .A2(n1263), .Z(n1265) );
  AO21D4BWP12T U2165 ( .A1(n1267), .A2(n1266), .B(n1265), .Z(n1342) );
  IND2D1BWP12T U2166 ( .A1(b[0]), .B1(n4508), .ZN(n1270) );
  XNR2XD2BWP12T U2167 ( .A1(n2123), .A2(n3930), .ZN(n1363) );
  XNR3XD4BWP12T U2168 ( .A1(n1341), .A2(n1342), .A3(n1345), .ZN(n1411) );
  XNR2D2BWP12T U2169 ( .A1(n3016), .A2(n2067), .ZN(n1273) );
  TPOAI22D2BWP12T U2170 ( .A1(n1273), .A2(n2575), .B1(n1907), .B2(n1355), .ZN(
        n1337) );
  XNR2XD2BWP12T U2171 ( .A1(n3911), .A2(n5085), .ZN(n1316) );
  TPOAI22D1BWP12T U2172 ( .A1(n2479), .A2(n1274), .B1(n2005), .B2(n1316), .ZN(
        n1336) );
  XNR2D1BWP12T U2173 ( .A1(n436), .A2(n5054), .ZN(n1327) );
  OAI22D1BWP12T U2174 ( .A1(n1275), .A2(n2523), .B1(n1327), .B2(n2521), .ZN(
        n1338) );
  XOR3XD4BWP12T U2175 ( .A1(n1337), .A2(n1336), .A3(n1338), .Z(n1398) );
  CKND4BWP12T U2176 ( .I(n1398), .ZN(n1296) );
  XNR2D1BWP12T U2177 ( .A1(n4511), .A2(n3938), .ZN(n1354) );
  TPOAI22D1BWP12T U2178 ( .A1(n1689), .A2(n1276), .B1(n2115), .B2(n1354), .ZN(
        n1394) );
  INVD1BWP12T U2179 ( .I(b[15]), .ZN(n1277) );
  XNR2XD4BWP12T U2180 ( .A1(n5033), .A2(n5079), .ZN(n1314) );
  TPOAI22D2BWP12T U2181 ( .A1(n1279), .A2(n2467), .B1(n1799), .B2(n1314), .ZN(
        n1331) );
  INVD2BWP12T U2182 ( .I(n1285), .ZN(n1281) );
  INVD3BWP12T U2183 ( .I(n1284), .ZN(n1280) );
  XOR3XD4BWP12T U2184 ( .A1(n1394), .A2(n1395), .A3(n1393), .Z(n1399) );
  INVD1BWP12T U2185 ( .I(n1292), .ZN(n1288) );
  TPND2D1BWP12T U2186 ( .A1(n1289), .A2(n1288), .ZN(n1290) );
  ND2D1BWP12T U2187 ( .A1(n1291), .A2(n1290), .ZN(n1295) );
  ND2D1BWP12T U2188 ( .A1(n1293), .A2(n1292), .ZN(n1294) );
  TPND2D2BWP12T U2189 ( .A1(n1295), .A2(n1294), .ZN(n1396) );
  XOR3XD4BWP12T U2190 ( .A1(n1296), .A2(n1399), .A3(n1396), .Z(n1413) );
  XNR3XD4BWP12T U2191 ( .A1(n1410), .A2(n1411), .A3(n1413), .ZN(n1308) );
  OAI21D1BWP12T U2192 ( .A1(n1299), .A2(n443), .B(n1297), .ZN(n1301) );
  ND2D1BWP12T U2193 ( .A1(n1299), .A2(n443), .ZN(n1300) );
  CKND2D2BWP12T U2194 ( .A1(n1301), .A2(n1300), .ZN(n1307) );
  TPNR2D1BWP12T U2195 ( .A1(n3046), .A2(n3050), .ZN(n1311) );
  INR2D4BWP12T U2196 ( .A1(n1303), .B1(n1302), .ZN(n3061) );
  TPND2D3BWP12T U2197 ( .A1(n1305), .A2(n1304), .ZN(n1306) );
  INVD3BWP12T U2198 ( .I(n1306), .ZN(n3065) );
  RCAOI21D2BWP12T U2199 ( .A1(n3061), .A2(n3064), .B(n3065), .ZN(n1309) );
  TPAOI21D2BWP12T U2200 ( .A1(n1312), .A2(n1311), .B(n1310), .ZN(n3006) );
  XNR2XD2BWP12T U2201 ( .A1(n2123), .A2(n3939), .ZN(n1385) );
  ND2D1BWP12T U2202 ( .A1(n1872), .A2(n1362), .ZN(n1322) );
  ND2D1BWP12T U2203 ( .A1(n1362), .A2(n1363), .ZN(n1321) );
  TPOAI22D2BWP12T U2204 ( .A1(n1314), .A2(n2467), .B1(n1382), .B2(n1799), .ZN(
        n1366) );
  ND3D1BWP12T U2205 ( .A1(n1322), .A2(n1321), .A3(n1366), .ZN(n1325) );
  IND2D1BWP12T U2206 ( .A1(n1316), .B1(n1315), .ZN(n1320) );
  XNR2XD2BWP12T U2207 ( .A1(n3911), .A2(n5237), .ZN(n1386) );
  CKND2BWP12T U2208 ( .I(n1386), .ZN(n1317) );
  ND2D2BWP12T U2209 ( .A1(n63), .A2(n1317), .ZN(n1319) );
  ND3D1BWP12T U2210 ( .A1(n1322), .A2(n1321), .A3(n1365), .ZN(n1324) );
  ND3D2BWP12T U2211 ( .A1(n1325), .A2(n1324), .A3(n1323), .ZN(n1479) );
  XNR2XD4BWP12T U2212 ( .A1(n436), .A2(n5264), .ZN(n1377) );
  OAI21D1BWP12T U2213 ( .A1(n1335), .A2(n55), .B(n1333), .ZN(n1328) );
  XNR2D1BWP12T U2214 ( .A1(n4511), .A2(n3930), .ZN(n1487) );
  XNR2D1BWP12T U2215 ( .A1(n1858), .A2(n5033), .ZN(n1432) );
  XNR2D1BWP12T U2216 ( .A1(n4301), .A2(n1858), .ZN(n1356) );
  TPOAI22D2BWP12T U2217 ( .A1(n2533), .A2(n1432), .B1(n2535), .B2(n1356), .ZN(
        n1465) );
  INVD1BWP12T U2218 ( .I(a[17]), .ZN(n4790) );
  BUFFXD4BWP12T U2219 ( .I(a[17]), .Z(n4788) );
  IND2D1BWP12T U2220 ( .A1(b[0]), .B1(n4788), .ZN(n1429) );
  TPOAI22D2BWP12T U2221 ( .A1(n1329), .A2(n1969), .B1(n439), .B2(n3015), .ZN(
        n1430) );
  XNR2XD4BWP12T U2222 ( .A1(n1431), .A2(n1330), .ZN(n1463) );
  XOR3XD4BWP12T U2223 ( .A1(n1464), .A2(n1465), .A3(n1463), .Z(n1476) );
  XOR3D2BWP12T U2224 ( .A1(n1479), .A2(n1478), .A3(n1476), .Z(n1538) );
  HA1D2BWP12T U2225 ( .A(n1332), .B(n1331), .CO(n1349), .S(n1395) );
  OAI21D1BWP12T U2226 ( .A1(n1338), .A2(n1337), .B(n1336), .ZN(n1340) );
  TPND2D1BWP12T U2227 ( .A1(n1338), .A2(n1337), .ZN(n1339) );
  TPND2D2BWP12T U2228 ( .A1(n1340), .A2(n1339), .ZN(n1348) );
  XOR3XD4BWP12T U2229 ( .A1(n1349), .A2(n1350), .A3(n1348), .Z(n1391) );
  ND2D1BWP12T U2230 ( .A1(n1391), .A2(n1392), .ZN(n1347) );
  NR2XD2BWP12T U2231 ( .A1(n1342), .A2(n1341), .ZN(n1344) );
  ND2D3BWP12T U2232 ( .A1(n1342), .A2(n1341), .ZN(n1343) );
  TPOAI21D2BWP12T U2233 ( .A1(n1392), .A2(n1391), .B(n1389), .ZN(n1346) );
  INVD3BWP12T U2234 ( .I(n1348), .ZN(n1353) );
  TPOAI21D4BWP12T U2235 ( .A1(n1353), .A2(n1352), .B(n1351), .ZN(n1521) );
  TPOAI22D2BWP12T U2236 ( .A1(n2575), .A2(n1355), .B1(n1387), .B2(n1907), .ZN(
        n1373) );
  TPNR2D1BWP12T U2237 ( .A1(n2533), .A2(n1356), .ZN(n1357) );
  CKND2BWP12T U2238 ( .I(n1357), .ZN(n1361) );
  TPNR2D2BWP12T U2239 ( .A1(n2535), .A2(n1358), .ZN(n1359) );
  INVD1P75BWP12T U2240 ( .I(n1359), .ZN(n1360) );
  ND2D4BWP12T U2241 ( .A1(n1361), .A2(n1360), .ZN(n1374) );
  XOR3XD4BWP12T U2242 ( .A1(n1372), .A2(n1373), .A3(n1374), .Z(n1402) );
  OAI21D1BWP12T U2243 ( .A1(n1872), .A2(n1363), .B(n1362), .ZN(n1364) );
  XOR3XD4BWP12T U2244 ( .A1(n1366), .A2(n1365), .A3(n1364), .Z(n1403) );
  FA1D2BWP12T U2245 ( .A(n1368), .B(n1369), .CI(n1367), .CO(n1404), .S(n1272)
         );
  RCOAI21D2BWP12T U2246 ( .A1(n1402), .A2(n1403), .B(n1404), .ZN(n1371) );
  ND2D3BWP12T U2247 ( .A1(n1403), .A2(n1402), .ZN(n1370) );
  TPND2D3BWP12T U2248 ( .A1(n1371), .A2(n1370), .ZN(n1520) );
  TPOAI21D1BWP12T U2249 ( .A1(n1374), .A2(n1373), .B(n1372), .ZN(n1376) );
  ND2D1BWP12T U2250 ( .A1(n1376), .A2(n1375), .ZN(n1471) );
  INVD3BWP12T U2251 ( .I(n2523), .ZN(n1380) );
  XNR2XD8BWP12T U2252 ( .A1(n436), .A2(n4770), .ZN(n1428) );
  RCAOI21D4BWP12T U2253 ( .A1(n1380), .A2(n1379), .B(n1378), .ZN(n1494) );
  XNR2D2BWP12T U2254 ( .A1(a[17]), .A2(b[1]), .ZN(n1445) );
  INVD1P75BWP12T U2255 ( .I(n1445), .ZN(n1381) );
  XNR2D2BWP12T U2256 ( .A1(n5079), .A2(n3938), .ZN(n1447) );
  TPOAI22D1BWP12T U2257 ( .A1(n1382), .A2(n2467), .B1(n1447), .B2(n1799), .ZN(
        n1496) );
  INVD1BWP12T U2258 ( .I(n1496), .ZN(n1383) );
  TPOAI22D1BWP12T U2259 ( .A1(n2020), .A2(n1385), .B1(n14), .B2(n1450), .ZN(
        n1455) );
  XNR2XD2BWP12T U2260 ( .A1(n3911), .A2(n5054), .ZN(n1486) );
  OAI22D1BWP12T U2261 ( .A1(n1484), .A2(n1907), .B1(n2575), .B2(n1387), .ZN(
        n1457) );
  XNR3XD4BWP12T U2262 ( .A1(n1471), .A2(n1472), .A3(n1473), .ZN(n1524) );
  XOR3XD4BWP12T U2263 ( .A1(n1388), .A2(n1520), .A3(n1524), .Z(n1534) );
  XOR3XD4BWP12T U2264 ( .A1(n1538), .A2(n1533), .A3(n1534), .Z(n2996) );
  INVD1P75BWP12T U2265 ( .I(n423), .ZN(n1390) );
  XNR3XD4BWP12T U2266 ( .A1(n1392), .A2(n1391), .A3(n1390), .ZN(n1417) );
  FA1D2BWP12T U2267 ( .A(n1394), .B(n1395), .CI(n1393), .CO(n1392), .S(n1397)
         );
  XOR3XD4BWP12T U2268 ( .A1(n1404), .A2(n1403), .A3(n1402), .Z(n1419) );
  NR2XD2BWP12T U2269 ( .A1(n1418), .A2(n1419), .ZN(n1405) );
  INVD1P75BWP12T U2270 ( .I(n1405), .ZN(n1406) );
  CKND2D2BWP12T U2271 ( .A1(n1417), .A2(n1406), .ZN(n1408) );
  ND2XD3BWP12T U2272 ( .A1(n1408), .A2(n1407), .ZN(n2995) );
  NR2XD2BWP12T U2273 ( .A1(n2996), .A2(n2995), .ZN(n1409) );
  XOR3D2BWP12T U2274 ( .A1(n1419), .A2(n1418), .A3(n1417), .Z(n1416) );
  TPNR2D1BWP12T U2275 ( .A1(n1411), .A2(n1410), .ZN(n1414) );
  ND2D1BWP12T U2276 ( .A1(n1411), .A2(n1410), .ZN(n1412) );
  OA21D1BWP12T U2277 ( .A1(n1414), .A2(n1413), .B(n1412), .Z(n1420) );
  TPNR2D2BWP12T U2278 ( .A1(n1416), .A2(n1415), .ZN(n2994) );
  INVD2BWP12T U2279 ( .I(n2994), .ZN(n3005) );
  TPND2D2BWP12T U2280 ( .A1(n2998), .A2(n3005), .ZN(n1422) );
  TPAOI21D2BWP12T U2281 ( .A1(n2998), .A2(n2993), .B(n435), .ZN(n1421) );
  INR2XD2BWP12T U2282 ( .A1(n3016), .B1(n2571), .ZN(n1440) );
  TPOAI22D2BWP12T U2283 ( .A1(n2523), .A2(n1428), .B1(n1427), .B2(n2521), .ZN(
        n1438) );
  XOR3XD4BWP12T U2284 ( .A1(n1439), .A2(n1440), .A3(n1438), .Z(n1468) );
  AN2XD2BWP12T U2285 ( .A1(n429), .A2(n1430), .Z(n1469) );
  XNR2D2BWP12T U2286 ( .A1(n4502), .A2(n4896), .ZN(n1504) );
  ND2D1BWP12T U2287 ( .A1(n1469), .A2(n1470), .ZN(n1436) );
  TPND2D2BWP12T U2288 ( .A1(n1437), .A2(n1436), .ZN(n1576) );
  TPND2D2BWP12T U2289 ( .A1(n1442), .A2(n1441), .ZN(n1549) );
  XOR2XD4BWP12T U2290 ( .A1(n1444), .A2(n1443), .Z(n1550) );
  INVD1BWP12T U2291 ( .I(n1490), .ZN(n1448) );
  IND2XD2BWP12T U2292 ( .A1(n1489), .B1(n1448), .ZN(n1451) );
  TPOAI22D1BWP12T U2293 ( .A1(n1872), .A2(n1450), .B1(n2469), .B2(n1449), .ZN(
        n1488) );
  ND2D2BWP12T U2294 ( .A1(n1451), .A2(n1488), .ZN(n1453) );
  ND2D1BWP12T U2295 ( .A1(n1489), .A2(n1490), .ZN(n1452) );
  TPND2D2BWP12T U2296 ( .A1(n1453), .A2(n1452), .ZN(n1547) );
  XOR3XD4BWP12T U2297 ( .A1(n1549), .A2(n1454), .A3(n1547), .Z(n1579) );
  XOR3XD4BWP12T U2298 ( .A1(n1575), .A2(n1576), .A3(n1579), .Z(n1588) );
  OAI21D1BWP12T U2299 ( .A1(n1457), .A2(n1456), .B(n1455), .ZN(n1459) );
  CKND2D2BWP12T U2300 ( .A1(n1459), .A2(n1458), .ZN(n1482) );
  INVD1BWP12T U2301 ( .I(n1464), .ZN(n1461) );
  ND2D1BWP12T U2302 ( .A1(n1465), .A2(n1464), .ZN(n1466) );
  TPND2D2BWP12T U2303 ( .A1(n1475), .A2(n1474), .ZN(n1477) );
  ND2D3BWP12T U2304 ( .A1(n1477), .A2(n1476), .ZN(n1481) );
  CKND2D2BWP12T U2305 ( .A1(n1518), .A2(n419), .ZN(n1583) );
  TPNR2D1BWP12T U2306 ( .A1(n1483), .A2(n1482), .ZN(n1564) );
  TPND2D1BWP12T U2307 ( .A1(n1483), .A2(n1482), .ZN(n1563) );
  TPOAI21D2BWP12T U2308 ( .A1(n1565), .A2(n1564), .B(n1563), .ZN(n1515) );
  XNR2D1BWP12T U2309 ( .A1(n4511), .A2(n3939), .ZN(n1506) );
  XOR3XD4BWP12T U2310 ( .A1(n1490), .A2(n1489), .A3(n1488), .Z(n1525) );
  TPOAI21D1BWP12T U2311 ( .A1(n2518), .A2(n1492), .B(n1491), .ZN(n1495) );
  TPNR2D1BWP12T U2312 ( .A1(n1495), .A2(n1496), .ZN(n1493) );
  TPNR2D1BWP12T U2313 ( .A1(n1494), .A2(n1493), .ZN(n1498) );
  AN2XD2BWP12T U2314 ( .A1(n1496), .A2(n1495), .Z(n1497) );
  TPNR2D2BWP12T U2315 ( .A1(n1498), .A2(n1497), .ZN(n1526) );
  INVD2BWP12T U2316 ( .I(n1526), .ZN(n1499) );
  AN2D4BWP12T U2317 ( .A1(n1501), .A2(n1500), .Z(n1514) );
  TPOAI22D2BWP12T U2318 ( .A1(n1504), .A2(n2535), .B1(n2533), .B2(n1503), .ZN(
        n1543) );
  OA22D2BWP12T U2319 ( .A1(n1689), .A2(n1506), .B1(n2481), .B2(n1505), .Z(
        n1546) );
  XOR3XD4BWP12T U2320 ( .A1(n1542), .A2(n1543), .A3(n1546), .Z(n1553) );
  FA1D2BWP12T U2321 ( .A(n1509), .B(n1508), .CI(n1507), .CO(n1556), .S(n1559)
         );
  XOR3D2BWP12T U2322 ( .A1(n1512), .A2(n1511), .A3(n1510), .Z(n1557) );
  XOR3XD4BWP12T U2323 ( .A1(n1553), .A2(n1556), .A3(n1513), .Z(n1558) );
  XOR3XD4BWP12T U2324 ( .A1(n1515), .A2(n1514), .A3(n1558), .Z(n1586) );
  XOR3XD4BWP12T U2325 ( .A1(n1588), .A2(n1516), .A3(n1586), .Z(n1596) );
  XNR3XD4BWP12T U2326 ( .A1(n1519), .A2(n1518), .A3(n1517), .ZN(n1530) );
  TPND2D1BWP12T U2327 ( .A1(n1521), .A2(n1520), .ZN(n1522) );
  TPOAI21D2BWP12T U2328 ( .A1(n1524), .A2(n1523), .B(n1522), .ZN(n1531) );
  XNR3XD4BWP12T U2329 ( .A1(n1526), .A2(n1525), .A3(n1559), .ZN(n1529) );
  TPNR2D1BWP12T U2330 ( .A1(n1531), .A2(n1529), .ZN(n1528) );
  ND2D1BWP12T U2331 ( .A1(n1531), .A2(n1529), .ZN(n1527) );
  OA21D2BWP12T U2332 ( .A1(n1528), .A2(n1530), .B(n1527), .Z(n1595) );
  TPND2D3BWP12T U2333 ( .A1(n1596), .A2(n1595), .ZN(n3087) );
  INVD2BWP12T U2334 ( .I(n1529), .ZN(n1532) );
  XOR3XD4BWP12T U2335 ( .A1(n1532), .A2(n1531), .A3(n1530), .Z(n1594) );
  INVD2BWP12T U2336 ( .I(n1594), .ZN(n1541) );
  INVD2BWP12T U2337 ( .I(n1533), .ZN(n1535) );
  INVD1BWP12T U2338 ( .I(n1535), .ZN(n1539) );
  CKND0BWP12T U2339 ( .I(n1538), .ZN(n1536) );
  IOA21D1BWP12T U2340 ( .A1(n1535), .A2(n1536), .B(n1534), .ZN(n1537) );
  IOA21D2BWP12T U2341 ( .A1(n1539), .A2(n1538), .B(n1537), .ZN(n1593) );
  TPND2D2BWP12T U2342 ( .A1(n1541), .A2(n1540), .ZN(n3001) );
  CKND2D2BWP12T U2343 ( .A1(n3001), .A2(n3087), .ZN(n3076) );
  NR2D1BWP12T U2344 ( .A1(n69), .A2(n1543), .ZN(n1545) );
  TPNR2D1BWP12T U2345 ( .A1(n1548), .A2(n1547), .ZN(n1552) );
  TPNR2D1BWP12T U2346 ( .A1(n1549), .A2(n1550), .ZN(n1551) );
  TPNR2D2BWP12T U2347 ( .A1(n1552), .A2(n1551), .ZN(n1613) );
  INVD1BWP12T U2348 ( .I(n1553), .ZN(n1554) );
  TPOAI21D1BWP12T U2349 ( .A1(n1557), .A2(n1556), .B(n1554), .ZN(n1555) );
  IOA21D2BWP12T U2350 ( .A1(n1557), .A2(n1556), .B(n1555), .ZN(n1611) );
  XOR3D2BWP12T U2351 ( .A1(n1612), .A2(n1613), .A3(n1611), .Z(n1644) );
  CKND3BWP12T U2352 ( .I(n1558), .ZN(n1567) );
  CKND0BWP12T U2353 ( .I(n1559), .ZN(n1562) );
  XOR3XD4BWP12T U2354 ( .A1(n1574), .A2(n1573), .A3(n1572), .Z(n1625) );
  ND2D1BWP12T U2355 ( .A1(n1576), .A2(n1575), .ZN(n1577) );
  XOR3XD4BWP12T U2356 ( .A1(n1625), .A2(n444), .A3(n1626), .Z(n1641) );
  XNR3XD4BWP12T U2357 ( .A1(n1644), .A2(n1643), .A3(n1641), .ZN(n1598) );
  TPND2D1BWP12T U2358 ( .A1(n1584), .A2(n1583), .ZN(n1589) );
  INVD1BWP12T U2359 ( .I(n1589), .ZN(n1585) );
  CKND2D1BWP12T U2360 ( .A1(n1585), .A2(n449), .ZN(n1587) );
  ND2D1BWP12T U2361 ( .A1(n1587), .A2(n1586), .ZN(n1592) );
  INVD1BWP12T U2362 ( .I(n1588), .ZN(n1590) );
  ND2D1BWP12T U2363 ( .A1(n1590), .A2(n1589), .ZN(n1591) );
  TPND2D2BWP12T U2364 ( .A1(n1592), .A2(n1591), .ZN(n1597) );
  TPNR2D2BWP12T U2365 ( .A1(n1596), .A2(n1595), .ZN(n3085) );
  TPAOI21D2BWP12T U2366 ( .A1(n3002), .A2(n3087), .B(n3085), .ZN(n3075) );
  ND2D3BWP12T U2367 ( .A1(n1598), .A2(n1597), .ZN(n3078) );
  TPOAI21D1BWP12T U2368 ( .A1(n3075), .A2(n3077), .B(n3078), .ZN(n1599) );
  TPAOI21D2BWP12T U2369 ( .A1(n3074), .A2(n1600), .B(n1599), .ZN(n2990) );
  XOR3XD4BWP12T U2370 ( .A1(n1603), .A2(n1602), .A3(n1601), .Z(n1658) );
  XOR3XD4BWP12T U2371 ( .A1(n1606), .A2(n1605), .A3(n1604), .Z(n1634) );
  NR2D1BWP12T U2372 ( .A1(n1613), .A2(n1612), .ZN(n1616) );
  INVD1BWP12T U2373 ( .I(n1611), .ZN(n1615) );
  ND2D1BWP12T U2374 ( .A1(n1613), .A2(n1612), .ZN(n1614) );
  TPOAI21D2BWP12T U2375 ( .A1(n1616), .A2(n1615), .B(n1614), .ZN(n1632) );
  ND2D2BWP12T U2376 ( .A1(n1617), .A2(n1632), .ZN(n1620) );
  TPND2D2BWP12T U2377 ( .A1(n1620), .A2(n1619), .ZN(n1657) );
  XNR3XD4BWP12T U2378 ( .A1(n1623), .A2(n1622), .A3(n1621), .ZN(n1654) );
  XNR3XD4BWP12T U2379 ( .A1(n1658), .A2(n1657), .A3(n1654), .ZN(n1665) );
  TPOAI21D1BWP12T U2380 ( .A1(n1625), .A2(n1626), .B(n1624), .ZN(n1628) );
  XOR3D2BWP12T U2381 ( .A1(n1631), .A2(n1630), .A3(n1629), .Z(n1640) );
  XNR3XD4BWP12T U2382 ( .A1(n1634), .A2(n1633), .A3(n1632), .ZN(n1638) );
  IND2D2BWP12T U2383 ( .A1(n1635), .B1(n1638), .ZN(n1637) );
  ND2D1BWP12T U2384 ( .A1(n1639), .A2(n1640), .ZN(n1636) );
  TPND2D2BWP12T U2385 ( .A1(n1637), .A2(n1636), .ZN(n1664) );
  NR2XD2BWP12T U2386 ( .A1(n1665), .A2(n1664), .ZN(n3109) );
  XOR3XD4BWP12T U2387 ( .A1(n1640), .A2(n1639), .A3(n1638), .Z(n1663) );
  IND2D1BWP12T U2388 ( .A1(n1644), .B1(n1643), .ZN(n1642) );
  INVD1BWP12T U2389 ( .I(n1643), .ZN(n1645) );
  ND2D1BWP12T U2390 ( .A1(n1645), .A2(n1644), .ZN(n1646) );
  TPND2D2BWP12T U2391 ( .A1(n1647), .A2(n1646), .ZN(n1662) );
  XOR3XD4BWP12T U2392 ( .A1(n1650), .A2(n1649), .A3(n1648), .Z(n1653) );
  XOR3XD4BWP12T U2393 ( .A1(n1653), .A2(n1652), .A3(n1651), .Z(n1667) );
  OR2D2BWP12T U2394 ( .A1(n1658), .A2(n1657), .Z(n1656) );
  INVD2BWP12T U2395 ( .I(n1654), .ZN(n1655) );
  TPND2D2BWP12T U2396 ( .A1(n1656), .A2(n1655), .ZN(n1660) );
  ND2D1BWP12T U2397 ( .A1(n1658), .A2(n1657), .ZN(n1659) );
  NR2XD2BWP12T U2398 ( .A1(n1667), .A2(n1666), .ZN(n1661) );
  INVD3BWP12T U2399 ( .I(n1661), .ZN(n3118) );
  CKND2D2BWP12T U2400 ( .A1(n3115), .A2(n3118), .ZN(n1670) );
  INVD1P75BWP12T U2401 ( .I(n3117), .ZN(n1668) );
  TPAOI21D1BWP12T U2402 ( .A1(n3114), .A2(n3118), .B(n1668), .ZN(n1669) );
  TPOAI21D1BWP12T U2403 ( .A1(n2990), .A2(n1670), .B(n1669), .ZN(n3104) );
  ND2D3BWP12T U2404 ( .A1(n1677), .A2(n1676), .ZN(n3126) );
  AOI21D0BWP12T U2405 ( .A1(n2735), .A2(n3104), .B(n2736), .ZN(n2048) );
  XNR2D1BWP12T U2406 ( .A1(a[17]), .A2(n5085), .ZN(n1713) );
  TPOAI22D2BWP12T U2407 ( .A1(n2518), .A2(n1678), .B1(n1713), .B2(n2516), .ZN(
        n1818) );
  INVD8BWP12T U2408 ( .I(n2895), .ZN(n4503) );
  XNR2D1BWP12T U2409 ( .A1(n3016), .A2(n2773), .ZN(n1682) );
  IND2D2BWP12T U2410 ( .A1(n1794), .B1(n1680), .ZN(n1681) );
  FA1D4BWP12T U2411 ( .A(n1686), .B(n1685), .CI(n1684), .CO(n1759), .S(n1723)
         );
  XNR2D1BWP12T U2412 ( .A1(n3911), .A2(b[23]), .ZN(n1710) );
  XNR2D1BWP12T U2413 ( .A1(n4511), .A2(n4700), .ZN(n1801) );
  XNR2XD0BWP12T U2414 ( .A1(n1858), .A2(b[15]), .ZN(n1712) );
  TPOAI22D1BWP12T U2415 ( .A1(n2535), .A2(n1692), .B1(n2533), .B2(n1712), .ZN(
        n1715) );
  XNR2D1BWP12T U2416 ( .A1(n4565), .A2(n3930), .ZN(n1784) );
  OAI22D1BWP12T U2417 ( .A1(n2573), .A2(n1693), .B1(n2571), .B2(n1784), .ZN(
        n1718) );
  XOR3XD4BWP12T U2418 ( .A1(n1717), .A2(n1715), .A3(n1718), .Z(n1754) );
  INVD2BWP12T U2419 ( .I(n1694), .ZN(n1696) );
  TPND2D2BWP12T U2420 ( .A1(n1696), .A2(n1695), .ZN(n1699) );
  INR2D4BWP12T U2421 ( .A1(n1697), .B1(n1696), .ZN(n1698) );
  INVD1P75BWP12T U2422 ( .I(n1755), .ZN(n1706) );
  TPND2D2BWP12T U2423 ( .A1(n1705), .A2(n1704), .ZN(n1756) );
  INVD1BWP12T U2424 ( .I(n1756), .ZN(n1707) );
  XNR2D1BWP12T U2425 ( .A1(n3911), .A2(n4655), .ZN(n1856) );
  OAI22D1BWP12T U2426 ( .A1(n2479), .A2(n1710), .B1(n1856), .B2(n2005), .ZN(
        n1850) );
  XNR2XD2BWP12T U2427 ( .A1(n4301), .A2(n4568), .ZN(n1930) );
  XNR2XD0BWP12T U2428 ( .A1(n4502), .A2(n4826), .ZN(n1859) );
  OAI22D0BWP12T U2429 ( .A1(n2535), .A2(n1712), .B1(n2533), .B2(n1859), .ZN(
        n1848) );
  OAI22D1BWP12T U2430 ( .A1(n2518), .A2(n1713), .B1(n1925), .B2(n2022), .ZN(
        n1914) );
  TPOAI22D2BWP12T U2431 ( .A1(n397), .A2(n1740), .B1(n2519), .B2(n1870), .ZN(
        n1916) );
  XNR2XD2BWP12T U2432 ( .A1(n2123), .A2(n4676), .ZN(n1730) );
  TPOAI22D1BWP12T U2433 ( .A1(n1872), .A2(n1730), .B1(n2469), .B2(n1871), .ZN(
        n1915) );
  CKND2BWP12T U2434 ( .I(n1915), .ZN(n1714) );
  XNR3XD4BWP12T U2435 ( .A1(n1914), .A2(n1916), .A3(n1714), .ZN(n1902) );
  IOA21D2BWP12T U2436 ( .A1(n1718), .A2(n1717), .B(n1716), .ZN(n1901) );
  INVD1BWP12T U2437 ( .I(n1901), .ZN(n1719) );
  XNR3XD4BWP12T U2438 ( .A1(n1899), .A2(n1902), .A3(n1719), .ZN(n1896) );
  FA1D2BWP12T U2439 ( .A(n1725), .B(n1724), .CI(n1723), .CO(n1771), .S(n1822)
         );
  FA1D2BWP12T U2440 ( .A(n1728), .B(n1727), .CI(n1726), .CO(n1791), .S(n1720)
         );
  TPOAI22D1BWP12T U2441 ( .A1(n2469), .A2(n1730), .B1(n2020), .B2(n1729), .ZN(
        n1775) );
  ND2D3BWP12T U2442 ( .A1(n3914), .A2(n1731), .ZN(n1732) );
  TPND2D2BWP12T U2443 ( .A1(n1733), .A2(n1732), .ZN(n1868) );
  OR2D2BWP12T U2444 ( .A1(n1799), .A2(n1800), .Z(n1734) );
  OAI21D1BWP12T U2445 ( .A1(n2467), .A2(n1735), .B(n1734), .ZN(n1777) );
  XOR3D2BWP12T U2446 ( .A1(n1775), .A2(n1776), .A3(n1777), .Z(n1790) );
  XNR2D1BWP12T U2447 ( .A1(n2067), .A2(n5054), .ZN(n1785) );
  TPOAI22D1BWP12T U2448 ( .A1(n1739), .A2(n1969), .B1(n1813), .B2(n3015), .ZN(
        n1810) );
  FA1D2BWP12T U2449 ( .A(n1744), .B(n1743), .CI(n1742), .CO(n1804), .S(n1721)
         );
  XOR3XD4BWP12T U2450 ( .A1(n1805), .A2(n1806), .A3(n1804), .Z(n1789) );
  XOR3XD4BWP12T U2451 ( .A1(n1770), .A2(n1771), .A3(n398), .Z(n1820) );
  IOA21D2BWP12T U2452 ( .A1(n1748), .A2(n1747), .B(n1746), .ZN(n1821) );
  XNR3XD4BWP12T U2453 ( .A1(n1756), .A2(n1755), .A3(n1754), .ZN(n1766) );
  CKND3BWP12T U2454 ( .I(n1757), .ZN(n1758) );
  XNR3XD4BWP12T U2455 ( .A1(n1760), .A2(n1759), .A3(n1758), .ZN(n1767) );
  XOR3XD4BWP12T U2456 ( .A1(n1762), .A2(n1766), .A3(n1761), .Z(n1819) );
  TPOAI21D1BWP12T U2457 ( .A1(n1820), .A2(n1821), .B(n1819), .ZN(n1764) );
  TPND2D1BWP12T U2458 ( .A1(n1820), .A2(n1821), .ZN(n1763) );
  TPND2D2BWP12T U2459 ( .A1(n1764), .A2(n1763), .ZN(n1938) );
  ND2D3BWP12T U2460 ( .A1(n1767), .A2(n1766), .ZN(n1768) );
  TPND2D2BWP12T U2461 ( .A1(n1774), .A2(n1773), .ZN(n1887) );
  ND2D1BWP12T U2462 ( .A1(n1777), .A2(n1776), .ZN(n1778) );
  XNR2D1BWP12T U2463 ( .A1(n4565), .A2(n3939), .ZN(n1909) );
  TPOAI22D1BWP12T U2464 ( .A1(n2573), .A2(n1784), .B1(n2571), .B2(n1909), .ZN(
        n1923) );
  OAI22D1BWP12T U2465 ( .A1(n2575), .A2(n1785), .B1(n1908), .B2(n1907), .ZN(
        n1921) );
  XNR2D1BWP12T U2466 ( .A1(n3887), .A2(n3653), .ZN(n1857) );
  TPOAI22D1BWP12T U2467 ( .A1(n2532), .A2(n1786), .B1(n1857), .B2(n2530), .ZN(
        n1924) );
  XOR3D2BWP12T U2468 ( .A1(n1923), .A2(n1921), .A3(n1924), .Z(n1881) );
  XOR3XD4BWP12T U2469 ( .A1(n1882), .A2(n1883), .A3(n1881), .Z(n1891) );
  CKND2BWP12T U2470 ( .I(n1791), .ZN(n1788) );
  CKND3BWP12T U2471 ( .I(n1789), .ZN(n1793) );
  ND2D1BWP12T U2472 ( .A1(n1791), .A2(n1790), .ZN(n1792) );
  TPOAI21D2BWP12T U2473 ( .A1(n464), .A2(n1793), .B(n1792), .ZN(n1892) );
  INVD1P75BWP12T U2474 ( .I(n2464), .ZN(n1796) );
  TPND2D2BWP12T U2475 ( .A1(n1796), .A2(n1795), .ZN(n1798) );
  OR2D2BWP12T U2476 ( .A1(n2462), .A2(n1867), .Z(n1797) );
  XNR2XD2BWP12T U2477 ( .A1(n5079), .A2(n4732), .ZN(n1932) );
  TPOAI22D1BWP12T U2478 ( .A1(n420), .A2(n1800), .B1(n2465), .B2(n1932), .ZN(
        n1852) );
  XNR2D1BWP12T U2479 ( .A1(n4511), .A2(n5122), .ZN(n1931) );
  OA22D2BWP12T U2480 ( .A1(n1689), .A2(n1801), .B1(n2115), .B2(n1931), .Z(
        n1855) );
  TPNR2D2BWP12T U2481 ( .A1(n430), .A2(n1805), .ZN(n1802) );
  INVD1P75BWP12T U2482 ( .I(n1802), .ZN(n1803) );
  ND2D2BWP12T U2483 ( .A1(n1804), .A2(n1803), .ZN(n1808) );
  TPND2D2BWP12T U2484 ( .A1(n1808), .A2(n1807), .ZN(n1861) );
  BUFFD6BWP12T U2485 ( .I(a[28]), .Z(n4609) );
  XNR2XD8BWP12T U2486 ( .A1(n4503), .A2(n4609), .ZN(n2017) );
  TPOAI22D1BWP12T U2487 ( .A1(n2523), .A2(n1814), .B1(n2521), .B2(n1928), .ZN(
        n1903) );
  IOA21D2BWP12T U2488 ( .A1(n1818), .A2(n1817), .B(n1816), .ZN(n1875) );
  XOR3XD4BWP12T U2489 ( .A1(n1877), .A2(n1878), .A3(n1875), .Z(n1860) );
  XNR3XD4BWP12T U2490 ( .A1(n1862), .A2(n1861), .A3(n1860), .ZN(n1894) );
  XOR3XD4BWP12T U2491 ( .A1(n1891), .A2(n1892), .A3(n1894), .Z(n1889) );
  XNR3XD4BWP12T U2492 ( .A1(n1886), .A2(n1887), .A3(n1889), .ZN(n1935) );
  XOR3XD4BWP12T U2493 ( .A1(n1937), .A2(n1938), .A3(n1935), .Z(n3098) );
  XNR3XD4BWP12T U2494 ( .A1(n1821), .A2(n1820), .A3(n409), .ZN(n1839) );
  INVD2BWP12T U2495 ( .I(n1839), .ZN(n1835) );
  OAI21D1BWP12T U2496 ( .A1(n1825), .A2(n1824), .B(n1822), .ZN(n1823) );
  INVD1P75BWP12T U2497 ( .I(n1836), .ZN(n1841) );
  CKND1BWP12T U2498 ( .I(n1829), .ZN(n1826) );
  ND2D1BWP12T U2499 ( .A1(n1830), .A2(n1829), .ZN(n1831) );
  TPND2D2BWP12T U2500 ( .A1(n1832), .A2(n1831), .ZN(n1840) );
  INR2D2BWP12T U2501 ( .A1(n1841), .B1(n1840), .ZN(n1833) );
  INVD1P75BWP12T U2502 ( .I(n1833), .ZN(n1834) );
  TPND2D2BWP12T U2503 ( .A1(n1835), .A2(n1834), .ZN(n1838) );
  XOR3XD4BWP12T U2504 ( .A1(n1841), .A2(n1840), .A3(n1839), .Z(n2039) );
  CKND2D2BWP12T U2505 ( .A1(n1843), .A2(n1842), .ZN(n1847) );
  TPND2D1BWP12T U2506 ( .A1(n1845), .A2(n1844), .ZN(n1846) );
  TPND2D3BWP12T U2507 ( .A1(n1847), .A2(n1846), .ZN(n2038) );
  FA1D2BWP12T U2508 ( .A(n1849), .B(n1850), .CI(n1848), .CO(n1975), .S(n1899)
         );
  TPOAI21D2BWP12T U2509 ( .A1(n1855), .A2(n1854), .B(n1853), .ZN(n1974) );
  XNR2D1BWP12T U2510 ( .A1(n2122), .A2(n3911), .ZN(n2006) );
  XOR2D1BWP12T U2511 ( .A1(n3887), .A2(n3930), .Z(n2004) );
  XNR2XD1BWP12T U2512 ( .A1(n4502), .A2(n4794), .ZN(n1956) );
  OAI22D0BWP12T U2513 ( .A1(n29), .A2(n1859), .B1(n2533), .B2(n1956), .ZN(
        n1957) );
  INVD1BWP12T U2514 ( .I(n1860), .ZN(n1866) );
  NR2D1BWP12T U2515 ( .A1(n1861), .A2(n1862), .ZN(n1865) );
  INVD1BWP12T U2516 ( .I(n1861), .ZN(n1864) );
  INVD1BWP12T U2517 ( .I(n1862), .ZN(n1863) );
  TPOAI22D2BWP12T U2518 ( .A1(n1866), .A2(n1865), .B1(n1864), .B2(n1863), .ZN(
        n2027) );
  TPOAI22D2BWP12T U2519 ( .A1(n1868), .A2(n1867), .B1(n2462), .B2(n2021), .ZN(
        n2000) );
  OAI22D1BWP12T U2520 ( .A1(n2016), .A2(n1870), .B1(n2015), .B2(n1869), .ZN(
        n2001) );
  XNR2XD2BWP12T U2521 ( .A1(n2123), .A2(n4920), .ZN(n2019) );
  TPOAI22D1BWP12T U2522 ( .A1(n1872), .A2(n1871), .B1(n2469), .B2(n2019), .ZN(
        n1999) );
  XOR3XD4BWP12T U2523 ( .A1(n1999), .A2(n2001), .A3(n2000), .Z(n1945) );
  CKND3BWP12T U2524 ( .I(n1878), .ZN(n1874) );
  INVD1BWP12T U2525 ( .I(n1877), .ZN(n1873) );
  TPND2D2BWP12T U2526 ( .A1(n1874), .A2(n1873), .ZN(n1876) );
  ND2D1BWP12T U2527 ( .A1(n1878), .A2(n1877), .ZN(n1879) );
  CKND2D4BWP12T U2528 ( .A1(n1880), .A2(n1879), .ZN(n1946) );
  XNR3XD4BWP12T U2529 ( .A1(n1945), .A2(n1946), .A3(n1943), .ZN(n2030) );
  INVD3BWP12T U2530 ( .I(n2030), .ZN(n1885) );
  XNR3XD4BWP12T U2531 ( .A1(n2028), .A2(n2027), .A3(n1885), .ZN(n2032) );
  OA21XD4BWP12T U2532 ( .A1(n1889), .A2(n1890), .B(n1888), .Z(n2034) );
  ND2D1BWP12T U2533 ( .A1(n1892), .A2(n1891), .ZN(n1893) );
  TPOAI21D2BWP12T U2534 ( .A1(n1894), .A2(n1895), .B(n1893), .ZN(n1979) );
  OAI21D1BWP12T U2535 ( .A1(n1902), .A2(n1901), .B(n1899), .ZN(n1900) );
  IOA21D2BWP12T U2536 ( .A1(n1902), .A2(n1901), .B(n1900), .ZN(n1985) );
  XNR2D1BWP12T U2537 ( .A1(n4565), .A2(n5085), .ZN(n1968) );
  BUFFD6BWP12T U2538 ( .I(b[29]), .Z(n4991) );
  TPOAI22D1BWP12T U2539 ( .A1(n1910), .A2(n1969), .B1(n1970), .B2(n3015), .ZN(
        n1967) );
  DCCKND4BWP12T U2540 ( .I(a[29]), .ZN(n4993) );
  INVD9BWP12T U2541 ( .I(n4993), .ZN(n4990) );
  XOR2XD4BWP12T U2542 ( .A1(n4990), .A2(n4609), .Z(n1926) );
  CKND3BWP12T U2543 ( .I(n1926), .ZN(n1913) );
  TPOAI22D2BWP12T U2544 ( .A1(n1913), .A2(n1912), .B1(n1911), .B2(n2017), .ZN(
        n1966) );
  XOR3XD4BWP12T U2545 ( .A1(n2013), .A2(n2012), .A3(n2008), .Z(n1960) );
  BUFFD2BWP12T U2546 ( .I(n1914), .Z(n1917) );
  TPOAI21D2BWP12T U2547 ( .A1(n1917), .A2(n1916), .B(n1915), .ZN(n1919) );
  ND2D3BWP12T U2548 ( .A1(n1917), .A2(n1916), .ZN(n1918) );
  TPND2D3BWP12T U2549 ( .A1(n1919), .A2(n1918), .ZN(n1962) );
  INVD1BWP12T U2550 ( .I(n1962), .ZN(n1920) );
  XNR3XD4BWP12T U2551 ( .A1(n1961), .A2(n1960), .A3(n1920), .ZN(n1986) );
  OAI21D1BWP12T U2552 ( .A1(n1924), .A2(n1923), .B(n1921), .ZN(n1922) );
  IOA21D2BWP12T U2553 ( .A1(n1924), .A2(n1923), .B(n1922), .ZN(n1989) );
  XNR2D1BWP12T U2554 ( .A1(a[17]), .A2(n5054), .ZN(n2023) );
  XNR2D1BWP12T U2555 ( .A1(n3016), .A2(n4990), .ZN(n1927) );
  XNR2D2BWP12T U2556 ( .A1(n4990), .A2(b[1]), .ZN(n2018) );
  TPOAI22D2BWP12T U2557 ( .A1(n2545), .A2(n1927), .B1(n413), .B2(n2018), .ZN(
        n1995) );
  XNR2D1BWP12T U2558 ( .A1(n436), .A2(b[27]), .ZN(n1972) );
  OAI22D1BWP12T U2559 ( .A1(n2523), .A2(n1928), .B1(n2521), .B2(n1972), .ZN(
        n1929) );
  INVD1BWP12T U2560 ( .I(n1929), .ZN(n1997) );
  XNR3XD4BWP12T U2561 ( .A1(n1994), .A2(n1995), .A3(n1997), .ZN(n1990) );
  XNR2D1BWP12T U2562 ( .A1(n4568), .A2(n5033), .ZN(n1954) );
  XNR2XD0BWP12T U2563 ( .A1(n4511), .A2(n4676), .ZN(n2024) );
  XNR2XD0BWP12T U2564 ( .A1(n5079), .A2(n4700), .ZN(n1955) );
  TPOAI22D1BWP12T U2565 ( .A1(n420), .A2(n1932), .B1(n1955), .B2(n2465), .ZN(
        n1951) );
  XNR3XD4BWP12T U2566 ( .A1(n1950), .A2(n1949), .A3(n1951), .ZN(n1993) );
  XNR3XD4BWP12T U2567 ( .A1(n1989), .A2(n1990), .A3(n1993), .ZN(n1984) );
  INVD1BWP12T U2568 ( .I(n1984), .ZN(n1933) );
  XNR3XD4BWP12T U2569 ( .A1(n1985), .A2(n1986), .A3(n1933), .ZN(n1981) );
  XOR3XD4BWP12T U2570 ( .A1(n1979), .A2(n1980), .A3(n1934), .Z(n2036) );
  XOR3XD4BWP12T U2571 ( .A1(n2032), .A2(n2034), .A3(n2036), .Z(n2041) );
  IND2XD2BWP12T U2572 ( .A1(n1936), .B1(n1935), .ZN(n1940) );
  ND2D1BWP12T U2573 ( .A1(n1938), .A2(n1937), .ZN(n1939) );
  TPND2D2BWP12T U2574 ( .A1(n1942), .A2(n1941), .ZN(n1944) );
  TPND2D2BWP12T U2575 ( .A1(n1944), .A2(n1943), .ZN(n1948) );
  ND2D1BWP12T U2576 ( .A1(n1946), .A2(n1945), .ZN(n1947) );
  CKND2D2BWP12T U2577 ( .A1(n1948), .A2(n1947), .ZN(n2127) );
  CKND2D1BWP12T U2578 ( .A1(n1951), .A2(n1950), .ZN(n1953) );
  OAI21D1BWP12T U2579 ( .A1(n1951), .A2(n1950), .B(n1949), .ZN(n1952) );
  ND2D1BWP12T U2580 ( .A1(n1953), .A2(n1952), .ZN(n2081) );
  XNR2D1BWP12T U2581 ( .A1(n4568), .A2(n4896), .ZN(n2092) );
  TPOAI22D2BWP12T U2582 ( .A1(n2529), .A2(n1954), .B1(n2), .B2(n2092), .ZN(
        n2060) );
  XNR2D1BWP12T U2583 ( .A1(n5079), .A2(n5122), .ZN(n2113) );
  TPOAI22D1BWP12T U2584 ( .A1(n2113), .A2(n2465), .B1(n1955), .B2(n2467), .ZN(
        n2061) );
  XNR2D1BWP12T U2585 ( .A1(n4502), .A2(n25), .ZN(n2094) );
  XOR3XD4BWP12T U2586 ( .A1(n2060), .A2(n2061), .A3(n2058), .Z(n2080) );
  FA1D2BWP12T U2587 ( .A(n1959), .B(n1958), .CI(n1957), .CO(n2082), .S(n1973)
         );
  XOR3D2BWP12T U2588 ( .A1(n2081), .A2(n2080), .A3(n2082), .Z(n2126) );
  RCOAI21D2BWP12T U2589 ( .A1(n1965), .A2(n1964), .B(n1963), .ZN(n2057) );
  HA1D2BWP12T U2590 ( .A(n1967), .B(n1966), .CO(n2119), .S(n2008) );
  XNR2XD0BWP12T U2591 ( .A1(n4565), .A2(n5237), .ZN(n2065) );
  TPOAI22D1BWP12T U2592 ( .A1(n2573), .A2(n1968), .B1(n2571), .B2(n2065), .ZN(
        n2118) );
  XOR2XD2BWP12T U2593 ( .A1(n1812), .A2(b[30]), .Z(n2100) );
  TPNR2D2BWP12T U2594 ( .A1(n2100), .A2(n3015), .ZN(n1971) );
  BUFFD6BWP12T U2595 ( .I(a[30]), .Z(n5146) );
  XNR2D2BWP12T U2596 ( .A1(n4990), .A2(a[30]), .ZN(n2547) );
  TPNR2D1BWP12T U2597 ( .A1(n2547), .A2(n3233), .ZN(n2099) );
  BUFFXD6BWP12T U2598 ( .I(b[28]), .Z(n4610) );
  XNR2D1BWP12T U2599 ( .A1(n436), .A2(n4610), .ZN(n2088) );
  OAI22D1BWP12T U2600 ( .A1(n2523), .A2(n1972), .B1(n2521), .B2(n2088), .ZN(
        n2096) );
  XNR3XD4BWP12T U2601 ( .A1(n2095), .A2(n2099), .A3(n2096), .ZN(n2117) );
  NR2D1BWP12T U2602 ( .A1(n1975), .A2(n1974), .ZN(n1977) );
  CKND2D1BWP12T U2603 ( .A1(n1975), .A2(n1974), .ZN(n1976) );
  OAI21D1BWP12T U2604 ( .A1(n1978), .A2(n1977), .B(n1976), .ZN(n2055) );
  TPOAI21D1BWP12T U2605 ( .A1(n1981), .A2(n406), .B(n1979), .ZN(n1983) );
  TPND2D1BWP12T U2606 ( .A1(n1981), .A2(n406), .ZN(n1982) );
  TPND2D2BWP12T U2607 ( .A1(n1983), .A2(n1982), .ZN(n2128) );
  ND2D2BWP12T U2608 ( .A1(n1988), .A2(n1987), .ZN(n2053) );
  CKND2BWP12T U2609 ( .I(n2053), .ZN(n2050) );
  TPNR2D2BWP12T U2610 ( .A1(n1990), .A2(n1989), .ZN(n1992) );
  TPOAI21D2BWP12T U2611 ( .A1(n1993), .A2(n1992), .B(n1991), .ZN(n2070) );
  TPNR2D1BWP12T U2612 ( .A1(n1994), .A2(n1995), .ZN(n1998) );
  ND2D1BWP12T U2613 ( .A1(n1995), .A2(n1994), .ZN(n1996) );
  TPOAI21D2BWP12T U2614 ( .A1(n1998), .A2(n1997), .B(n1996), .ZN(n2108) );
  TPOAI21D1BWP12T U2615 ( .A1(n2001), .A2(n2000), .B(n1999), .ZN(n2003) );
  TPND2D2BWP12T U2616 ( .A1(n2003), .A2(n2002), .ZN(n2109) );
  XNR2D1BWP12T U2617 ( .A1(n3887), .A2(n3652), .ZN(n2066) );
  TPOAI22D1BWP12T U2618 ( .A1(n2532), .A2(n2004), .B1(n2066), .B2(n2530), .ZN(
        n2091) );
  XNR2D1BWP12T U2619 ( .A1(n5030), .A2(n4944), .ZN(n2093) );
  XNR2XD0BWP12T U2620 ( .A1(n4508), .A2(n4826), .ZN(n2068) );
  OAI22D1BWP12T U2621 ( .A1(n2575), .A2(n2007), .B1(n2068), .B2(n51), .ZN(
        n2089) );
  XOR3XD4BWP12T U2622 ( .A1(n2108), .A2(n2109), .A3(n2107), .Z(n2069) );
  INVD1BWP12T U2623 ( .I(n2013), .ZN(n2009) );
  XNR2D1BWP12T U2624 ( .A1(n5196), .A2(n4990), .ZN(n2085) );
  XNR2XD0BWP12T U2625 ( .A1(n2123), .A2(n4655), .ZN(n2124) );
  OAI22D0BWP12T U2626 ( .A1(n2124), .A2(n2469), .B1(n2019), .B2(n2020), .ZN(
        n2102) );
  XOR3D2BWP12T U2627 ( .A1(n2104), .A2(n2103), .A3(n2102), .Z(n2076) );
  XNR2D1BWP12T U2628 ( .A1(n4301), .A2(n4503), .ZN(n2114) );
  XNR2D1BWP12T U2629 ( .A1(a[17]), .A2(n5264), .ZN(n2121) );
  OAI22D1BWP12T U2630 ( .A1(n2518), .A2(n2023), .B1(n2121), .B2(n2516), .ZN(
        n2063) );
  XNR2XD0BWP12T U2631 ( .A1(n4511), .A2(b[22]), .ZN(n2116) );
  OAI22D0BWP12T U2632 ( .A1(n1689), .A2(n2024), .B1(n2481), .B2(n2116), .ZN(
        n2062) );
  XNR3XD4BWP12T U2633 ( .A1(n2075), .A2(n2076), .A3(n2025), .ZN(n2071) );
  XNR3XD4BWP12T U2634 ( .A1(n2070), .A2(n2069), .A3(n2071), .ZN(n2051) );
  INVD1BWP12T U2635 ( .I(n2028), .ZN(n2026) );
  TPNR2D1BWP12T U2636 ( .A1(n2026), .A2(n2027), .ZN(n2031) );
  INVD1BWP12T U2637 ( .I(n2027), .ZN(n2029) );
  XNR3XD4BWP12T U2638 ( .A1(n2050), .A2(n2051), .A3(n2049), .ZN(n2131) );
  INVD2BWP12T U2639 ( .I(n2032), .ZN(n2035) );
  TPND2D1BWP12T U2640 ( .A1(n2034), .A2(n2035), .ZN(n2033) );
  INVD1P75BWP12T U2641 ( .I(n2033), .ZN(n2037) );
  OAI22D2BWP12T U2642 ( .A1(n2037), .A2(n2036), .B1(n2035), .B2(n2034), .ZN(
        n2042) );
  NR2D2BWP12T U2643 ( .A1(n3140), .A2(n3145), .ZN(n2044) );
  TPND2D1BWP12T U2644 ( .A1(n2044), .A2(n3144), .ZN(n2047) );
  TPOAI21D1BWP12T U2645 ( .A1(n3151), .A2(n3150), .B(n3149), .ZN(n2045) );
  TPOAI21D1BWP12T U2646 ( .A1(n3145), .A2(n3141), .B(n3146), .ZN(n2043) );
  TPAOI21D1BWP12T U2647 ( .A1(n2045), .A2(n2044), .B(n2043), .ZN(n2046) );
  TPOAI21D1BWP12T U2648 ( .A1(n2048), .A2(n2047), .B(n2046), .ZN(n2461) );
  INVD1BWP12T U2649 ( .I(n2051), .ZN(n2054) );
  IOA21D1BWP12T U2650 ( .A1(n2051), .A2(n2050), .B(n2049), .ZN(n2052) );
  IOA21D1BWP12T U2651 ( .A1(n2053), .A2(n2054), .B(n2052), .ZN(n2595) );
  FA1D2BWP12T U2652 ( .A(n2056), .B(n2057), .CI(n2055), .CO(n2587), .S(n2125)
         );
  FA1D2BWP12T U2653 ( .A(n2064), .B(n2063), .CI(n2062), .CO(n2508), .S(n2077)
         );
  XNR2XD0BWP12T U2654 ( .A1(n4565), .A2(n5054), .ZN(n2572) );
  OAI22D0BWP12T U2655 ( .A1(n2573), .A2(n2065), .B1(n2571), .B2(n2572), .ZN(
        n2515) );
  XNR2D1BWP12T U2656 ( .A1(n3887), .A2(n2234), .ZN(n2531) );
  OAI22D1BWP12T U2657 ( .A1(n2532), .A2(n2066), .B1(n2531), .B2(n2530), .ZN(
        n2514) );
  XNR2XD0BWP12T U2658 ( .A1(n4508), .A2(n4794), .ZN(n2574) );
  OAI22D0BWP12T U2659 ( .A1(n2575), .A2(n2068), .B1(n2574), .B2(n51), .ZN(
        n2513) );
  TPND2D0BWP12T U2660 ( .A1(n2069), .A2(n2070), .ZN(n2074) );
  ND2D1BWP12T U2661 ( .A1(n2069), .A2(n2071), .ZN(n2073) );
  ND2D1BWP12T U2662 ( .A1(n2071), .A2(n2070), .ZN(n2072) );
  ND3D1BWP12T U2663 ( .A1(n2074), .A2(n2073), .A3(n2072), .ZN(n2585) );
  ND2D1BWP12T U2664 ( .A1(n2077), .A2(n2076), .ZN(n2079) );
  OAI21D1BWP12T U2665 ( .A1(n2077), .A2(n2076), .B(n2075), .ZN(n2078) );
  ND2D1BWP12T U2666 ( .A1(n2079), .A2(n2078), .ZN(n2500) );
  OAI21D0BWP12T U2667 ( .A1(n2082), .A2(n2081), .B(n2080), .ZN(n2084) );
  CKND2D1BWP12T U2668 ( .A1(n2082), .A2(n2081), .ZN(n2083) );
  XNR2D1BWP12T U2669 ( .A1(n3948), .A2(n4990), .ZN(n2546) );
  INVD3BWP12T U2670 ( .I(a[31]), .ZN(n3564) );
  INVD9BWP12T U2671 ( .I(n3564), .ZN(n5108) );
  XOR2D1BWP12T U2672 ( .A1(n5108), .A2(n5146), .Z(n2086) );
  TPND2D1BWP12T U2673 ( .A1(n2086), .A2(n2547), .ZN(n2549) );
  XNR2D1BWP12T U2674 ( .A1(n3016), .A2(n5108), .ZN(n2087) );
  XNR2XD0BWP12T U2675 ( .A1(n5108), .A2(b[1]), .ZN(n2548) );
  TPOAI22D1BWP12T U2676 ( .A1(n2549), .A2(n2087), .B1(n2548), .B2(n2547), .ZN(
        n2553) );
  XNR2D1BWP12T U2677 ( .A1(n436), .A2(n31), .ZN(n2522) );
  OAI22D0BWP12T U2678 ( .A1(n2523), .A2(n2088), .B1(n2521), .B2(n2522), .ZN(
        n2550) );
  FA1D2BWP12T U2679 ( .A(n2091), .B(n2090), .CI(n2089), .CO(n2511), .S(n2107)
         );
  XNR2XD0BWP12T U2680 ( .A1(n4568), .A2(n3938), .ZN(n2528) );
  OAI22D0BWP12T U2681 ( .A1(n2529), .A2(n2092), .B1(n23), .B2(n2528), .ZN(
        n2570) );
  XNR2D1BWP12T U2682 ( .A1(n3911), .A2(n21), .ZN(n2478) );
  XNR2XD0BWP12T U2683 ( .A1(n5049), .A2(n4700), .ZN(n2534) );
  OAI22D0BWP12T U2684 ( .A1(n29), .A2(n2094), .B1(n2533), .B2(n2534), .ZN(
        n2568) );
  OAI21D1BWP12T U2685 ( .A1(n2099), .A2(n2098), .B(n2096), .ZN(n2097) );
  IOA21D1BWP12T U2686 ( .A1(n2099), .A2(n2098), .B(n2097), .ZN(n2488) );
  BUFFD6BWP12T U2687 ( .I(b[31]), .Z(n3936) );
  XOR2XD0BWP12T U2688 ( .A1(n1812), .A2(n3936), .Z(n2475) );
  OAI22D1BWP12T U2689 ( .A1(n2476), .A2(n2100), .B1(n2475), .B2(n3015), .ZN(
        n2577) );
  INVD1BWP12T U2690 ( .I(n5108), .ZN(n2612) );
  IND2D1BWP12T U2691 ( .A1(n3016), .B1(n5108), .ZN(n2101) );
  OAI22D1BWP12T U2692 ( .A1(n2549), .A2(n2612), .B1(n2101), .B2(n2547), .ZN(
        n2576) );
  TPND2D1BWP12T U2693 ( .A1(n2106), .A2(n2105), .ZN(n2486) );
  INVD1BWP12T U2694 ( .I(n2107), .ZN(n2112) );
  TPNR2D1BWP12T U2695 ( .A1(n2109), .A2(n2108), .ZN(n2111) );
  CKND2D0BWP12T U2696 ( .A1(n2109), .A2(n2108), .ZN(n2110) );
  OAI21D1BWP12T U2697 ( .A1(n2112), .A2(n2111), .B(n2110), .ZN(n2497) );
  XNR2XD0BWP12T U2698 ( .A1(n5079), .A2(n4676), .ZN(n2468) );
  OAI22D1BWP12T U2699 ( .A1(n2113), .A2(n2467), .B1(n2468), .B2(n2465), .ZN(
        n2556) );
  XNR2D1BWP12T U2700 ( .A1(n4503), .A2(n5033), .ZN(n2463) );
  XNR2XD0BWP12T U2701 ( .A1(n4511), .A2(n4920), .ZN(n2482) );
  OAI22D0BWP12T U2702 ( .A1(n1689), .A2(n2116), .B1(n2115), .B2(n2482), .ZN(
        n2554) );
  FA1D2BWP12T U2703 ( .A(n2119), .B(n2118), .CI(n2117), .CO(n2560), .S(n2056)
         );
  XNR2XD0BWP12T U2704 ( .A1(n4914), .A2(n3930), .ZN(n2520) );
  OAI22D1BWP12T U2705 ( .A1(n397), .A2(n2120), .B1(n2520), .B2(n2519), .ZN(
        n2567) );
  XNR2D1BWP12T U2706 ( .A1(n4788), .A2(n32), .ZN(n2517) );
  OAI22D1BWP12T U2707 ( .A1(n2518), .A2(n2121), .B1(n2517), .B2(n2022), .ZN(
        n2566) );
  XNR2XD0BWP12T U2708 ( .A1(n2123), .A2(n4977), .ZN(n2470) );
  OAI22D0BWP12T U2709 ( .A1(n2471), .A2(n2124), .B1(n2469), .B2(n2470), .ZN(
        n2565) );
  XOR3XD4BWP12T U2710 ( .A1(n2496), .A2(n2497), .A3(n2492), .Z(n2505) );
  FA1D2BWP12T U2711 ( .A(n2127), .B(n2126), .CI(n2125), .CO(n2504), .S(n2129)
         );
  INVD1BWP12T U2712 ( .I(n2128), .ZN(n2134) );
  OAI21D2BWP12T U2713 ( .A1(n2134), .A2(n2133), .B(n2132), .ZN(n2136) );
  TPNR2D2BWP12T U2714 ( .A1(n2137), .A2(n2136), .ZN(n2135) );
  CKND2D2BWP12T U2715 ( .A1(n2137), .A2(n2136), .ZN(n2458) );
  TPND2D2BWP12T U2716 ( .A1(n2460), .A2(n2458), .ZN(n2138) );
  XNR2XD4BWP12T U2717 ( .A1(n2461), .A2(n2138), .ZN(n5100) );
  INVD1P75BWP12T U2718 ( .I(op[0]), .ZN(n2183) );
  INR2D4BWP12T U2719 ( .A1(op[3]), .B1(n2183), .ZN(n2351) );
  INR2D2BWP12T U2720 ( .A1(op[2]), .B1(op[1]), .ZN(n2139) );
  CKBD1BWP12T U2721 ( .I(n5079), .Z(n4521) );
  OR2D2BWP12T U2722 ( .A1(n2155), .A2(n4521), .Z(n3242) );
  INVD3BWP12T U2723 ( .I(n5237), .ZN(n3650) );
  OR2D2BWP12T U2724 ( .A1(n3650), .A2(n5234), .Z(n3246) );
  ND2D1BWP12T U2725 ( .A1(n3242), .A2(n3246), .ZN(n3168) );
  INVD3BWP12T U2726 ( .I(n5054), .ZN(n3651) );
  OR2D2BWP12T U2727 ( .A1(n3651), .A2(n5049), .Z(n3176) );
  NR2D1BWP12T U2728 ( .A1(n1222), .A2(a[14]), .ZN(n2235) );
  INVD1BWP12T U2729 ( .I(n2235), .ZN(n3181) );
  ND2D1BWP12T U2730 ( .A1(n3176), .A2(n3181), .ZN(n2158) );
  NR2D1BWP12T U2731 ( .A1(n3168), .A2(n2158), .ZN(n3302) );
  INVD2BWP12T U2732 ( .I(n3930), .ZN(n3658) );
  OR2D2BWP12T U2733 ( .A1(n3658), .A2(n2153), .Z(n2878) );
  BUFFD2BWP12T U2734 ( .I(a[10]), .Z(n2848) );
  OR2D2BWP12T U2735 ( .A1(n2232), .A2(n2848), .Z(n2811) );
  ND2D1BWP12T U2736 ( .A1(n2878), .A2(n2811), .ZN(n2154) );
  BUFFD2BWP12T U2737 ( .I(n3899), .Z(n3937) );
  NR2D1BWP12T U2738 ( .A1(n3653), .A2(n3495), .ZN(n2876) );
  NR2D1BWP12T U2739 ( .A1(n2154), .A2(n2876), .ZN(n3240) );
  ND2D1BWP12T U2740 ( .A1(n3302), .A2(n3240), .ZN(n3250) );
  INVD2BWP12T U2741 ( .I(n4794), .ZN(n3648) );
  NR2D1BWP12T U2742 ( .A1(n3648), .A2(n4788), .ZN(n3384) );
  INVD1BWP12T U2743 ( .I(n3384), .ZN(n3379) );
  NR2D1BWP12T U2744 ( .A1(n3641), .A2(a[18]), .ZN(n2243) );
  INVD1BWP12T U2745 ( .I(n2243), .ZN(n3192) );
  ND2D1BWP12T U2746 ( .A1(n3379), .A2(n3192), .ZN(n2164) );
  INVD2BWP12T U2747 ( .I(n32), .ZN(n3649) );
  OR2D2BWP12T U2748 ( .A1(n3649), .A2(n4508), .Z(n3448) );
  INVD2BWP12T U2749 ( .I(n4826), .ZN(n3643) );
  NR2D1BWP12T U2750 ( .A1(n3643), .A2(n4822), .ZN(n2242) );
  ND2D1BWP12T U2751 ( .A1(n3448), .A2(n3308), .ZN(n3310) );
  TPNR2D1BWP12T U2752 ( .A1(n2164), .A2(n3310), .ZN(n3194) );
  INVD3BWP12T U2753 ( .I(n16), .ZN(n3642) );
  BUFFD2BWP12T U2754 ( .I(n4565), .Z(n4696) );
  NR2D2BWP12T U2755 ( .A1(n3642), .A2(n4696), .ZN(n3393) );
  INVD1BWP12T U2756 ( .I(n3393), .ZN(n3390) );
  INVD3BWP12T U2757 ( .I(n26), .ZN(n3639) );
  OR2D2BWP12T U2758 ( .A1(n3639), .A2(n5118), .Z(n3188) );
  ND2D1BWP12T U2759 ( .A1(n3390), .A2(n3188), .ZN(n3259) );
  INVD3BWP12T U2760 ( .I(n17), .ZN(n3640) );
  OR2D2BWP12T U2761 ( .A1(n3640), .A2(n4672), .Z(n3263) );
  INVD3BWP12T U2762 ( .I(n2142), .ZN(n4635) );
  OR2XD1BWP12T U2763 ( .A1(n3637), .A2(n2825), .Z(n3265) );
  ND2D1BWP12T U2764 ( .A1(n3263), .A2(n3265), .ZN(n2169) );
  NR2D1BWP12T U2765 ( .A1(n3259), .A2(n2169), .ZN(n2171) );
  ND2D1BWP12T U2766 ( .A1(n3194), .A2(n2171), .ZN(n2173) );
  NR2D1BWP12T U2767 ( .A1(n3250), .A2(n2173), .ZN(n2175) );
  TPNR2D1BWP12T U2768 ( .A1(n3334), .A2(n480), .ZN(n5290) );
  INVD3BWP12T U2769 ( .I(n4849), .ZN(n2834) );
  NR2D1BWP12T U2770 ( .A1(n2834), .A2(n4501), .ZN(n2219) );
  ND2D1BWP12T U2771 ( .A1(n2834), .A2(n4501), .ZN(n3231) );
  OAI21D1BWP12T U2772 ( .A1(n5290), .A2(n2219), .B(n3231), .ZN(n2692) );
  INVD1BWP12T U2773 ( .I(n3948), .ZN(n2143) );
  BUFFXD4BWP12T U2774 ( .I(n3570), .Z(n3661) );
  NR2D1BWP12T U2775 ( .A1(n2143), .A2(n3661), .ZN(n2693) );
  INVD3BWP12T U2776 ( .I(n5196), .ZN(n3539) );
  NR2D1BWP12T U2777 ( .A1(n3539), .A2(n5192), .ZN(n3227) );
  NR2D1BWP12T U2778 ( .A1(n2693), .A2(n3227), .ZN(n2145) );
  ND2D1BWP12T U2779 ( .A1(n3539), .A2(n5192), .ZN(n3228) );
  ND2D1BWP12T U2780 ( .A1(n2143), .A2(n3661), .ZN(n2694) );
  OAI21D1BWP12T U2781 ( .A1(n2693), .A2(n3228), .B(n2694), .ZN(n2144) );
  AOI21D1BWP12T U2782 ( .A1(n2692), .A2(n2145), .B(n2144), .ZN(n2386) );
  INVD1BWP12T U2783 ( .I(n4301), .ZN(n2147) );
  INVD4BWP12T U2784 ( .I(n3912), .ZN(n4541) );
  NR2D1BWP12T U2785 ( .A1(n2147), .A2(n4541), .ZN(n2387) );
  INVD1BWP12T U2786 ( .I(n5033), .ZN(n3660) );
  BUFFXD0BWP12T U2787 ( .I(n5030), .Z(n2148) );
  TPNR2D2BWP12T U2788 ( .A1(n3660), .A2(n2148), .ZN(n3346) );
  NR2XD0BWP12T U2789 ( .A1(n2387), .A2(n3346), .ZN(n3221) );
  INVD2BWP12T U2790 ( .I(n3938), .ZN(n3659) );
  BUFFD2BWP12T U2791 ( .I(n4510), .Z(n3679) );
  TPNR2D1BWP12T U2792 ( .A1(n3659), .A2(n3679), .ZN(n2631) );
  BUFFD3BWP12T U2793 ( .I(n2146), .Z(n4891) );
  TPNR2D2BWP12T U2794 ( .A1(n2227), .A2(n4891), .ZN(n3223) );
  NR2XD0BWP12T U2795 ( .A1(n2631), .A2(n3223), .ZN(n2150) );
  ND2D1BWP12T U2796 ( .A1(n3221), .A2(n2150), .ZN(n2152) );
  ND2D1BWP12T U2797 ( .A1(n2147), .A2(n4541), .ZN(n3215) );
  ND2D1BWP12T U2798 ( .A1(n3660), .A2(n2148), .ZN(n3345) );
  OAI21D1BWP12T U2799 ( .A1(n3215), .A2(n3346), .B(n3345), .ZN(n3220) );
  ND2D1BWP12T U2800 ( .A1(n2227), .A2(n4891), .ZN(n3224) );
  ND2D1BWP12T U2801 ( .A1(n3659), .A2(n3679), .ZN(n2632) );
  OAI21D1BWP12T U2802 ( .A1(n2631), .A2(n3224), .B(n2632), .ZN(n2149) );
  AOI21D1BWP12T U2803 ( .A1(n3220), .A2(n2150), .B(n2149), .ZN(n2151) );
  TPOAI21D1BWP12T U2804 ( .A1(n2386), .A2(n2152), .B(n2151), .ZN(n2807) );
  INVD2BWP12T U2805 ( .I(n3495), .ZN(n3900) );
  INVD2BWP12T U2806 ( .I(n3900), .ZN(n4509) );
  ND2D1BWP12T U2807 ( .A1(n3658), .A2(n2153), .ZN(n2877) );
  BUFFD2BWP12T U2808 ( .I(n2848), .Z(n2849) );
  ND2D1BWP12T U2809 ( .A1(n2232), .A2(n2849), .ZN(n2819) );
  ND2D1BWP12T U2810 ( .A1(n2155), .A2(n4521), .ZN(n3237) );
  ND2D1BWP12T U2811 ( .A1(n3650), .A2(n5234), .ZN(n3362) );
  ND2D1BWP12T U2812 ( .A1(n3651), .A2(n5049), .ZN(n3171) );
  INVD1BWP12T U2813 ( .I(n3171), .ZN(n3175) );
  ND2D1BWP12T U2814 ( .A1(n1222), .A2(a[14]), .ZN(n3180) );
  INVD1BWP12T U2815 ( .I(n3180), .ZN(n2156) );
  AOI21D1BWP12T U2816 ( .A1(n3181), .A2(n3175), .B(n2156), .ZN(n2157) );
  OAI21D1BWP12T U2817 ( .A1(n3167), .A2(n2158), .B(n2157), .ZN(n2159) );
  AOI21D1BWP12T U2818 ( .A1(n3243), .A2(n3302), .B(n2159), .ZN(n3249) );
  INVD2BWP12T U2819 ( .I(n3447), .ZN(n3376) );
  ND2D1BWP12T U2820 ( .A1(n3643), .A2(n4822), .ZN(n3307) );
  INVD1BWP12T U2821 ( .I(n3307), .ZN(n2160) );
  AOI21D1BWP12T U2822 ( .A1(n3308), .A2(n3376), .B(n2160), .ZN(n3312) );
  ND2D1BWP12T U2823 ( .A1(n3648), .A2(n4788), .ZN(n3383) );
  INVD0BWP12T U2824 ( .I(n3383), .ZN(n2162) );
  ND2D1BWP12T U2825 ( .A1(n3641), .A2(a[18]), .ZN(n3191) );
  INVD1BWP12T U2826 ( .I(n3191), .ZN(n2161) );
  AOI21D1BWP12T U2827 ( .A1(n3192), .A2(n2162), .B(n2161), .ZN(n2163) );
  OAI21D1BWP12T U2828 ( .A1(n3312), .A2(n2164), .B(n2163), .ZN(n3193) );
  ND2D1BWP12T U2829 ( .A1(n3642), .A2(n4696), .ZN(n3198) );
  CKND0BWP12T U2830 ( .I(n3198), .ZN(n2166) );
  ND2D1BWP12T U2831 ( .A1(n3639), .A2(n5118), .ZN(n3187) );
  INVD1BWP12T U2832 ( .I(n3187), .ZN(n2165) );
  AOI21D1BWP12T U2833 ( .A1(n3188), .A2(n2166), .B(n2165), .ZN(n3261) );
  ND2D1BWP12T U2834 ( .A1(n3640), .A2(n4672), .ZN(n3410) );
  INVD1BWP12T U2835 ( .I(n3410), .ZN(n3262) );
  ND2D1BWP12T U2836 ( .A1(n3637), .A2(n2825), .ZN(n3414) );
  INVD0BWP12T U2837 ( .I(n3414), .ZN(n2167) );
  AOI21D1BWP12T U2838 ( .A1(n3265), .A2(n3262), .B(n2167), .ZN(n2168) );
  OAI21D1BWP12T U2839 ( .A1(n3261), .A2(n2169), .B(n2168), .ZN(n2170) );
  AOI21D1BWP12T U2840 ( .A1(n3193), .A2(n2171), .B(n2170), .ZN(n2172) );
  OAI21D1BWP12T U2841 ( .A1(n3249), .A2(n2173), .B(n2172), .ZN(n2174) );
  TPAOI21D2BWP12T U2842 ( .A1(n2175), .A2(n2807), .B(n2174), .ZN(n3298) );
  INVD2BWP12T U2843 ( .I(n21), .ZN(n3669) );
  OR2D2BWP12T U2844 ( .A1(n3669), .A2(n2773), .Z(n3453) );
  INVD2BWP12T U2845 ( .I(n22), .ZN(n3667) );
  ND2D1BWP12T U2846 ( .A1(n3453), .A2(n3280), .ZN(n3284) );
  INVD3BWP12T U2847 ( .I(n31), .ZN(n3668) );
  INVD2BWP12T U2848 ( .I(n5153), .ZN(n3666) );
  OR2XD1BWP12T U2849 ( .A1(n3666), .A2(n5146), .Z(n3300) );
  CKND2D1BWP12T U2850 ( .A1(n3294), .A2(n3300), .ZN(n2177) );
  OR2XD1BWP12T U2851 ( .A1(n3284), .A2(n2177), .Z(n2178) );
  INVD3BWP12T U2852 ( .I(n4920), .ZN(n3638) );
  NR2D1BWP12T U2853 ( .A1(n3638), .A2(n4914), .ZN(n3201) );
  INVD3BWP12T U2854 ( .I(n4655), .ZN(n3670) );
  NR2D1BWP12T U2855 ( .A1(n3670), .A2(n4649), .ZN(n3202) );
  NR2D1BWP12T U2856 ( .A1(n3201), .A2(n3202), .ZN(n3266) );
  OR2D2BWP12T U2857 ( .A1(n689), .A2(n4943), .Z(n3273) );
  AN2XD1BWP12T U2858 ( .A1(n3268), .A2(n3273), .Z(n2176) );
  ND2D1BWP12T U2859 ( .A1(n3266), .A2(n2176), .ZN(n3282) );
  NR2D1BWP12T U2860 ( .A1(n2178), .A2(n3282), .ZN(n2603) );
  INVD1BWP12T U2861 ( .I(n2603), .ZN(n2180) );
  ND2D1BWP12T U2862 ( .A1(n3638), .A2(n4914), .ZN(n3210) );
  ND2D1BWP12T U2863 ( .A1(n3670), .A2(n4649), .ZN(n3203) );
  OAI21D1BWP12T U2864 ( .A1(n3202), .A2(n3210), .B(n3203), .ZN(n3269) );
  ND2D1BWP12T U2865 ( .A1(n2250), .A2(n4568), .ZN(n3207) );
  INVD1BWP12T U2866 ( .I(n3207), .ZN(n3267) );
  ND2D1BWP12T U2867 ( .A1(n689), .A2(n4943), .ZN(n3272) );
  CKND2D2BWP12T U2868 ( .A1(n3669), .A2(n2773), .ZN(n2744) );
  INVD2BWP12T U2869 ( .I(n2744), .ZN(n3452) );
  ND2D1BWP12T U2870 ( .A1(n3667), .A2(n1), .ZN(n3279) );
  ND2D1BWP12T U2871 ( .A1(n4990), .A2(n3668), .ZN(n3288) );
  INVD1BWP12T U2872 ( .I(n3288), .ZN(n3293) );
  ND2D1BWP12T U2873 ( .A1(n3666), .A2(n5146), .ZN(n3299) );
  INVD1BWP12T U2874 ( .I(n2606), .ZN(n2179) );
  OAI21D1BWP12T U2875 ( .A1(n3298), .A2(n2180), .B(n2179), .ZN(n2182) );
  OR2XD1BWP12T U2876 ( .A1(n2612), .A2(n3936), .Z(n2605) );
  ND2D1BWP12T U2877 ( .A1(n2612), .A2(n3936), .ZN(n2604) );
  ND2D1BWP12T U2878 ( .A1(n2605), .A2(n2604), .ZN(n2181) );
  XNR2D1BWP12T U2879 ( .A1(n2182), .A2(n2181), .ZN(n3315) );
  IND2XD1BWP12T U2880 ( .A1(op[2]), .B1(op[1]), .ZN(n2184) );
  INR2D2BWP12T U2881 ( .A1(n2183), .B1(n2184), .ZN(n2344) );
  CKND2D2BWP12T U2882 ( .A1(n2344), .A2(op[3]), .ZN(n5203) );
  INVD6BWP12T U2883 ( .I(n5203), .ZN(n5305) );
  CKND2D1BWP12T U2884 ( .A1(n480), .A2(n3016), .ZN(n4059) );
  NR2D1BWP12T U2885 ( .A1(n4849), .A2(n4501), .ZN(n4058) );
  ND2D1BWP12T U2886 ( .A1(n4849), .A2(n4501), .ZN(n4433) );
  OAI21D1BWP12T U2887 ( .A1(n4059), .A2(n4058), .B(n4433), .ZN(n2701) );
  DEL025D1BWP12T U2888 ( .I(n3948), .Z(n2186) );
  NR2D1BWP12T U2889 ( .A1(n2186), .A2(n2185), .ZN(n2702) );
  TPNR2D2BWP12T U2890 ( .A1(n5196), .A2(n5192), .ZN(n4056) );
  NR2D1BWP12T U2891 ( .A1(n2702), .A2(n4056), .ZN(n2188) );
  ND2D1BWP12T U2892 ( .A1(n5196), .A2(n5192), .ZN(n4429) );
  ND2D1BWP12T U2893 ( .A1(n2186), .A2(n2185), .ZN(n2703) );
  OAI21D1BWP12T U2894 ( .A1(n2702), .A2(n4429), .B(n2703), .ZN(n2187) );
  AOI21D1BWP12T U2895 ( .A1(n2701), .A2(n2188), .B(n2187), .ZN(n2442) );
  CKBD1BWP12T U2896 ( .I(n4301), .Z(n2189) );
  NR2D1BWP12T U2897 ( .A1(n2189), .A2(n4541), .ZN(n2443) );
  NR2D1BWP12T U2898 ( .A1(n2443), .A2(n4046), .ZN(n4049) );
  BUFFD2BWP12T U2899 ( .I(n3938), .Z(n2640) );
  NR2D1BWP12T U2900 ( .A1(n2271), .A2(n4891), .ZN(n4051) );
  NR2D1BWP12T U2901 ( .A1(n2661), .A2(n4051), .ZN(n2192) );
  ND2D1BWP12T U2902 ( .A1(n4049), .A2(n2192), .ZN(n2194) );
  ND2D1BWP12T U2903 ( .A1(n2189), .A2(n4541), .ZN(n4043) );
  CKND2D1BWP12T U2904 ( .A1(n2271), .A2(n4891), .ZN(n4422) );
  ND2D1BWP12T U2905 ( .A1(n4510), .A2(n2640), .ZN(n2945) );
  OAI21D1BWP12T U2906 ( .A1(n2661), .A2(n4422), .B(n2945), .ZN(n2191) );
  AOI21D1BWP12T U2907 ( .A1(n4048), .A2(n2192), .B(n2191), .ZN(n2193) );
  TPOAI21D1BWP12T U2908 ( .A1(n2442), .A2(n2194), .B(n2193), .ZN(n2865) );
  BUFFD2BWP12T U2909 ( .I(n3930), .Z(n2909) );
  TPNR2D2BWP12T U2910 ( .A1(n2273), .A2(n2909), .ZN(n2859) );
  NR2D1BWP12T U2911 ( .A1(n3937), .A2(n4509), .ZN(n2930) );
  NR2D1BWP12T U2912 ( .A1(n2859), .A2(n2930), .ZN(n4084) );
  NR2D1BWP12T U2913 ( .A1(n4521), .A2(n5085), .ZN(n4091) );
  TPNR2D2BWP12T U2914 ( .A1(n2195), .A2(n2849), .ZN(n2863) );
  NR2D1BWP12T U2915 ( .A1(n4091), .A2(n2863), .ZN(n2196) );
  ND2D1BWP12T U2916 ( .A1(n4084), .A2(n2196), .ZN(n4095) );
  NR2D1BWP12T U2917 ( .A1(n5049), .A2(n5054), .ZN(n4406) );
  TPNR2D1BWP12T U2918 ( .A1(n5237), .A2(n5234), .ZN(n4387) );
  TPNR2D1BWP12T U2919 ( .A1(n4406), .A2(n4387), .ZN(n4023) );
  NR2D1BWP12T U2920 ( .A1(n4508), .A2(n32), .ZN(n4029) );
  NR2D1BWP12T U2921 ( .A1(n5264), .A2(a[14]), .ZN(n4027) );
  NR2D1BWP12T U2922 ( .A1(n4029), .A2(n4027), .ZN(n2197) );
  ND2D1BWP12T U2923 ( .A1(n4023), .A2(n2197), .ZN(n2199) );
  TPNR2D1BWP12T U2924 ( .A1(n4095), .A2(n2199), .ZN(n2201) );
  CKND2D1BWP12T U2925 ( .A1(n3937), .A2(n4509), .ZN(n2948) );
  ND2D1BWP12T U2926 ( .A1(n2153), .A2(n2909), .ZN(n2931) );
  OAI21D1BWP12T U2927 ( .A1(n2859), .A2(n2948), .B(n2931), .ZN(n4088) );
  CKND2D2BWP12T U2928 ( .A1(n2195), .A2(n2849), .ZN(n4085) );
  ND2D1BWP12T U2929 ( .A1(n4521), .A2(n5085), .ZN(n4382) );
  ND2D1BWP12T U2930 ( .A1(n5237), .A2(n5234), .ZN(n4388) );
  ND2D1BWP12T U2931 ( .A1(n5049), .A2(n5054), .ZN(n4405) );
  OAI21D1BWP12T U2932 ( .A1(n4406), .A2(n4388), .B(n4405), .ZN(n4025) );
  ND2D1BWP12T U2933 ( .A1(n5264), .A2(a[14]), .ZN(n4026) );
  ND2D1BWP12T U2934 ( .A1(n4508), .A2(n32), .ZN(n4393) );
  TPOAI21D1BWP12T U2935 ( .A1(n4094), .A2(n2199), .B(n2198), .ZN(n2200) );
  TPAOI21D4BWP12T U2936 ( .A1(n2865), .A2(n2201), .B(n2200), .ZN(n4116) );
  OR2D2BWP12T U2937 ( .A1(n4914), .A2(n4920), .Z(n4366) );
  NR2D1BWP12T U2938 ( .A1(b[22]), .A2(n2825), .ZN(n4075) );
  INVD1BWP12T U2939 ( .I(n4075), .ZN(n4072) );
  ND2D1BWP12T U2940 ( .A1(n4366), .A2(n4072), .ZN(n4100) );
  OR2XD1BWP12T U2941 ( .A1(n4568), .A2(n4977), .Z(n4118) );
  OR2XD1BWP12T U2942 ( .A1(n4655), .A2(n4649), .Z(n4106) );
  ND2D1BWP12T U2943 ( .A1(n4118), .A2(n4106), .ZN(n2205) );
  NR2D1BWP12T U2944 ( .A1(n4100), .A2(n2205), .ZN(n2207) );
  NR2D1BWP12T U2945 ( .A1(n4672), .A2(n17), .ZN(n4356) );
  NR2D1BWP12T U2946 ( .A1(n26), .A2(n5118), .ZN(n4008) );
  NR2D1BWP12T U2947 ( .A1(n4356), .A2(n4008), .ZN(n4069) );
  ND2D1BWP12T U2948 ( .A1(n2207), .A2(n4069), .ZN(n2209) );
  NR2D1BWP12T U2949 ( .A1(n4788), .A2(n4794), .ZN(n4030) );
  NR2D1BWP12T U2950 ( .A1(n4826), .A2(n448), .ZN(n4061) );
  NR2D1BWP12T U2951 ( .A1(n4030), .A2(n4061), .ZN(n3998) );
  NR2D1BWP12T U2952 ( .A1(n4696), .A2(n16), .ZN(n4005) );
  NR2D1BWP12T U2953 ( .A1(n25), .A2(a[18]), .ZN(n3996) );
  NR2D1BWP12T U2954 ( .A1(n4005), .A2(n3996), .ZN(n2202) );
  ND2D1BWP12T U2955 ( .A1(n3998), .A2(n2202), .ZN(n4010) );
  TPNR2D1BWP12T U2956 ( .A1(n2209), .A2(n4010), .ZN(n3985) );
  OR2D2BWP12T U2957 ( .A1(n2773), .A2(n21), .Z(n4461) );
  NR2D1BWP12T U2958 ( .A1(n4944), .A2(n4943), .ZN(n2287) );
  INVD1BWP12T U2959 ( .I(n2287), .ZN(n3983) );
  ND2D1BWP12T U2960 ( .A1(n4461), .A2(n3983), .ZN(n3972) );
  OR2D2BWP12T U2961 ( .A1(n2255), .A2(n31), .Z(n3980) );
  NR2D1BWP12T U2962 ( .A1(n22), .A2(n1), .ZN(n3974) );
  INVD1BWP12T U2963 ( .I(n3974), .ZN(n3970) );
  CKND2D1BWP12T U2964 ( .A1(n3980), .A2(n3970), .ZN(n2210) );
  NR2D1BWP12T U2965 ( .A1(n3972), .A2(n2210), .ZN(n3987) );
  NR2D1BWP12T U2966 ( .A1(n5153), .A2(n5146), .ZN(n2290) );
  INVD1BWP12T U2967 ( .I(n2290), .ZN(n3992) );
  CKND2D1BWP12T U2968 ( .A1(n3987), .A2(n3992), .ZN(n2616) );
  INVD1BWP12T U2969 ( .I(n2616), .ZN(n2213) );
  TPND2D0BWP12T U2970 ( .A1(n3985), .A2(n2213), .ZN(n2215) );
  CKND2D0BWP12T U2971 ( .A1(n4826), .A2(n4822), .ZN(n4062) );
  ND2D1BWP12T U2972 ( .A1(n4788), .A2(n4794), .ZN(n4031) );
  OAI21D1BWP12T U2973 ( .A1(n4030), .A2(n4062), .B(n4031), .ZN(n4002) );
  ND2D1BWP12T U2974 ( .A1(n25), .A2(a[18]), .ZN(n3999) );
  ND2D1BWP12T U2975 ( .A1(n4696), .A2(n16), .ZN(n4342) );
  ND2D1BWP12T U2976 ( .A1(n26), .A2(n5118), .ZN(n4012) );
  ND2D1BWP12T U2977 ( .A1(n4672), .A2(n17), .ZN(n4355) );
  OAI21D1BWP12T U2978 ( .A1(n4356), .A2(n4012), .B(n4355), .ZN(n4068) );
  ND2D1BWP12T U2979 ( .A1(b[22]), .A2(n2825), .ZN(n4361) );
  ND2D1BWP12T U2980 ( .A1(n4914), .A2(n4920), .ZN(n4080) );
  ND2D1BWP12T U2981 ( .A1(n4655), .A2(n4649), .ZN(n4374) );
  INVD1BWP12T U2982 ( .I(n4374), .ZN(n4105) );
  ND2D1BWP12T U2983 ( .A1(n4568), .A2(n4977), .ZN(n4117) );
  AOI21D1BWP12T U2984 ( .A1(n4118), .A2(n4105), .B(n2203), .ZN(n2204) );
  OAI21D1BWP12T U2985 ( .A1(n4104), .A2(n2205), .B(n2204), .ZN(n2206) );
  AOI21D1BWP12T U2986 ( .A1(n2207), .A2(n4068), .B(n2206), .ZN(n2208) );
  TPOAI21D1BWP12T U2987 ( .A1(n2209), .A2(n4011), .B(n2208), .ZN(n3988) );
  ND2D1BWP12T U2988 ( .A1(n4944), .A2(n4943), .ZN(n3982) );
  INVD1BWP12T U2989 ( .I(n3982), .ZN(n2747) );
  ND2D1BWP12T U2990 ( .A1(n2773), .A2(n21), .ZN(n2750) );
  INVD1BWP12T U2991 ( .I(n2750), .ZN(n4460) );
  AOI21D1BWP12T U2992 ( .A1(n4461), .A2(n2747), .B(n4460), .ZN(n3975) );
  ND2D1BWP12T U2993 ( .A1(n22), .A2(n1), .ZN(n3973) );
  ND2D1BWP12T U2994 ( .A1(n2255), .A2(n31), .ZN(n4480) );
  ND2D1BWP12T U2995 ( .A1(n5153), .A2(n5146), .ZN(n3991) );
  INVD1BWP12T U2996 ( .I(n3991), .ZN(n2211) );
  AOI21D1BWP12T U2997 ( .A1(n3986), .A2(n3992), .B(n2211), .ZN(n2619) );
  INVD1BWP12T U2998 ( .I(n2619), .ZN(n2212) );
  AOI21D1BWP12T U2999 ( .A1(n3988), .A2(n2213), .B(n2212), .ZN(n2214) );
  OAI21D1BWP12T U3000 ( .A1(n4116), .A2(n2215), .B(n2214), .ZN(n2218) );
  NR2D1BWP12T U3001 ( .A1(n2612), .A2(n2355), .ZN(n2618) );
  INVD1BWP12T U3002 ( .I(n2618), .ZN(n2216) );
  ND2D1BWP12T U3003 ( .A1(n2612), .A2(n2355), .ZN(n2617) );
  ND2D1BWP12T U3004 ( .A1(n2216), .A2(n2617), .ZN(n2217) );
  XNR2D1BWP12T U3005 ( .A1(n2218), .A2(n2217), .ZN(n4036) );
  CKND0BWP12T U3006 ( .I(n2219), .ZN(n3336) );
  NR2D1BWP12T U3007 ( .A1(n480), .A2(c_in), .ZN(n3332) );
  CKND2D1BWP12T U3008 ( .A1(n480), .A2(c_in), .ZN(n3333) );
  OAI21D1BWP12T U3009 ( .A1(b[0]), .A2(n3332), .B(n3333), .ZN(n3325) );
  ND2D1BWP12T U3010 ( .A1(n3336), .A2(n3325), .ZN(n2221) );
  INVD1BWP12T U3011 ( .I(n5196), .ZN(n2835) );
  TPNR2D1BWP12T U3012 ( .A1(n2835), .A2(n5192), .ZN(n2222) );
  TPNR2D1BWP12T U3013 ( .A1(n2221), .A2(n2222), .ZN(n2224) );
  CKND2D0BWP12T U3014 ( .A1(n2834), .A2(n4501), .ZN(n3671) );
  ND2D1BWP12T U3015 ( .A1(n2835), .A2(n5192), .ZN(n3328) );
  TPOAI21D1BWP12T U3016 ( .A1(n2222), .A2(n3671), .B(n3328), .ZN(n2223) );
  TPNR2D2BWP12T U3017 ( .A1(n2224), .A2(n2223), .ZN(n2716) );
  INVD1BWP12T U3018 ( .I(n3948), .ZN(n2225) );
  NR2D1BWP12T U3019 ( .A1(n2225), .A2(n3661), .ZN(n2436) );
  INVD1BWP12T U3020 ( .I(n4301), .ZN(n2226) );
  TPNR2D1BWP12T U3021 ( .A1(n2226), .A2(n4541), .ZN(n2438) );
  NR2D1BWP12T U3022 ( .A1(n2436), .A2(n2438), .ZN(n3342) );
  NR2D1BWP12T U3023 ( .A1(n3223), .A2(n3346), .ZN(n2229) );
  ND2D1BWP12T U3024 ( .A1(n3342), .A2(n2229), .ZN(n2231) );
  ND2D1BWP12T U3025 ( .A1(n2225), .A2(n3661), .ZN(n2713) );
  ND2D1BWP12T U3026 ( .A1(n2226), .A2(n4541), .ZN(n2439) );
  OAI21D1BWP12T U3027 ( .A1(n2438), .A2(n2713), .B(n2439), .ZN(n3344) );
  ND2D1BWP12T U3028 ( .A1(n2227), .A2(n4891), .ZN(n3351) );
  OAI21D1BWP12T U3029 ( .A1(n3223), .A2(n3345), .B(n3351), .ZN(n2228) );
  AOI21D1BWP12T U3030 ( .A1(n3344), .A2(n2229), .B(n2228), .ZN(n2230) );
  TPOAI21D1BWP12T U3031 ( .A1(n2716), .A2(n2231), .B(n2230), .ZN(n2630) );
  NR2D1BWP12T U3032 ( .A1(n3659), .A2(n3679), .ZN(n2959) );
  NR2D1BWP12T U3033 ( .A1(n3653), .A2(n4509), .ZN(n2960) );
  NR2D1BWP12T U3034 ( .A1(n2959), .A2(n2960), .ZN(n2881) );
  NR2D1BWP12T U3035 ( .A1(n2232), .A2(n2849), .ZN(n2818) );
  NR2D1BWP12T U3036 ( .A1(n3658), .A2(n2153), .ZN(n2814) );
  NR2D1BWP12T U3037 ( .A1(n2818), .A2(n2814), .ZN(n2233) );
  ND2D1BWP12T U3038 ( .A1(n2881), .A2(n2233), .ZN(n3420) );
  NR2D1BWP12T U3039 ( .A1(n3650), .A2(n5234), .ZN(n3361) );
  NR2D1BWP12T U3040 ( .A1(n3651), .A2(n5049), .ZN(n3371) );
  NR2D1BWP12T U3041 ( .A1(n2235), .A2(n3371), .ZN(n2237) );
  ND2D1BWP12T U3042 ( .A1(n3367), .A2(n2237), .ZN(n2239) );
  NR2D1BWP12T U3043 ( .A1(n3420), .A2(n2239), .ZN(n2241) );
  ND2D1BWP12T U3044 ( .A1(n3659), .A2(n3679), .ZN(n2958) );
  OAI21D1BWP12T U3045 ( .A1(n2960), .A2(n2958), .B(n2961), .ZN(n2882) );
  ND2D1BWP12T U3046 ( .A1(n3658), .A2(n2153), .ZN(n2885) );
  ND2D1BWP12T U3047 ( .A1(n2234), .A2(n4521), .ZN(n3422) );
  OAI21D1BWP12T U3048 ( .A1(n3361), .A2(n3422), .B(n3362), .ZN(n3366) );
  ND2D1BWP12T U3049 ( .A1(n3651), .A2(n5049), .ZN(n3372) );
  OAI21D1BWP12T U3050 ( .A1(n2235), .A2(n3372), .B(n3180), .ZN(n2236) );
  AOI21D1BWP12T U3051 ( .A1(n2237), .A2(n3366), .B(n2236), .ZN(n2238) );
  OAI21D1BWP12T U3052 ( .A1(n3419), .A2(n2239), .B(n2238), .ZN(n2240) );
  TPAOI21D1BWP12T U3053 ( .A1(n2630), .A2(n2241), .B(n2240), .ZN(n2741) );
  NR2D1BWP12T U3054 ( .A1(n3639), .A2(n5118), .ZN(n3397) );
  NR2D1BWP12T U3055 ( .A1(n3397), .A2(n3393), .ZN(n3403) );
  NR2D1BWP12T U3056 ( .A1(n3637), .A2(n2825), .ZN(n3413) );
  NR2D1BWP12T U3057 ( .A1(n3640), .A2(n4672), .ZN(n3411) );
  NR2D1BWP12T U3058 ( .A1(n3413), .A2(n3411), .ZN(n2247) );
  ND2D1BWP12T U3059 ( .A1(n3403), .A2(n2247), .ZN(n2249) );
  NR2D1BWP12T U3060 ( .A1(n2243), .A2(n3384), .ZN(n2245) );
  ND2D1BWP12T U3061 ( .A1(n3380), .A2(n2245), .ZN(n3391) );
  TPNR2D1BWP12T U3062 ( .A1(n2249), .A2(n3391), .ZN(n3433) );
  NR2D1BWP12T U3063 ( .A1(n3638), .A2(n4914), .ZN(n3434) );
  NR2D1BWP12T U3064 ( .A1(n3202), .A2(n3434), .ZN(n3442) );
  NR2D1BWP12T U3065 ( .A1(n689), .A2(n4943), .ZN(n2251) );
  ND2D1BWP12T U3066 ( .A1(n3442), .A2(n2253), .ZN(n3450) );
  NR2D1BWP12T U3067 ( .A1(n3667), .A2(n1), .ZN(n2254) );
  NR2D1BWP12T U3068 ( .A1(n3666), .A2(n5146), .ZN(n2256) );
  NR2D1BWP12T U3069 ( .A1(n3668), .A2(n2255), .ZN(n3473) );
  NR2D1BWP12T U3070 ( .A1(n2256), .A2(n3473), .ZN(n2258) );
  CKND2D1BWP12T U3071 ( .A1(n3467), .A2(n2258), .ZN(n2260) );
  NR2D1BWP12T U3072 ( .A1(n3450), .A2(n2260), .ZN(n2262) );
  TPND2D0BWP12T U3073 ( .A1(n3433), .A2(n2262), .ZN(n2264) );
  OAI21D1BWP12T U3074 ( .A1(n2242), .A2(n3447), .B(n3307), .ZN(n3382) );
  OAI21D1BWP12T U3075 ( .A1(n2243), .A2(n3383), .B(n3191), .ZN(n2244) );
  AOI21D1BWP12T U3076 ( .A1(n2245), .A2(n3382), .B(n2244), .ZN(n3394) );
  ND2D1BWP12T U3077 ( .A1(n3642), .A2(n4696), .ZN(n3392) );
  ND2D1BWP12T U3078 ( .A1(n3639), .A2(n5118), .ZN(n3398) );
  OAI21D1BWP12T U3079 ( .A1(n3397), .A2(n3392), .B(n3398), .ZN(n3402) );
  TPOAI21D0BWP12T U3080 ( .A1(n3413), .A2(n3410), .B(n3414), .ZN(n2246) );
  AOI21D1BWP12T U3081 ( .A1(n2247), .A2(n3402), .B(n2246), .ZN(n2248) );
  OAI21D1BWP12T U3082 ( .A1(n3394), .A2(n2249), .B(n2248), .ZN(n3415) );
  ND2D1BWP12T U3083 ( .A1(n3638), .A2(n4914), .ZN(n3432) );
  OAI21D1BWP12T U3084 ( .A1(n3202), .A2(n3432), .B(n3203), .ZN(n3444) );
  ND2D1BWP12T U3085 ( .A1(n2250), .A2(n4568), .ZN(n3443) );
  TPOAI21D0BWP12T U3086 ( .A1(n2251), .A2(n3443), .B(n3272), .ZN(n2252) );
  AOI21D1BWP12T U3087 ( .A1(n2253), .A2(n3444), .B(n2252), .ZN(n3451) );
  OAI21D1BWP12T U3088 ( .A1(n2254), .A2(n2744), .B(n3279), .ZN(n3471) );
  ND2D1BWP12T U3089 ( .A1(n3668), .A2(n2255), .ZN(n3472) );
  OAI21D0BWP12T U3090 ( .A1(n2256), .A2(n3472), .B(n3299), .ZN(n2257) );
  TPAOI21D0BWP12T U3091 ( .A1(n2258), .A2(n3471), .B(n2257), .ZN(n2259) );
  TPOAI21D0BWP12T U3092 ( .A1(n3451), .A2(n2260), .B(n2259), .ZN(n2261) );
  TPAOI21D0BWP12T U3093 ( .A1(n3415), .A2(n2262), .B(n2261), .ZN(n2263) );
  TPOAI21D0BWP12T U3094 ( .A1(n2741), .A2(n2264), .B(n2263), .ZN(n2609) );
  OR2XD1BWP12T U3095 ( .A1(n3936), .A2(n2612), .Z(n2608) );
  ND2D1BWP12T U3096 ( .A1(n3936), .A2(n2612), .ZN(n2607) );
  ND2D1BWP12T U3097 ( .A1(n2608), .A2(n2607), .ZN(n2265) );
  XNR2D1BWP12T U3098 ( .A1(n2609), .A2(n2265), .ZN(n3324) );
  INR2D2BWP12T U3099 ( .A1(op[2]), .B1(op[3]), .ZN(n2412) );
  INR2D1BWP12T U3100 ( .A1(op[1]), .B1(op[0]), .ZN(n2348) );
  INVD6BWP12T U3101 ( .I(n5105), .ZN(n5308) );
  INR2XD0BWP12T U3102 ( .A1(op[0]), .B1(op[1]), .ZN(n2266) );
  INVD4BWP12T U3103 ( .I(n4965), .ZN(n5313) );
  TPNR2D1BWP12T U3104 ( .A1(n3908), .A2(n4501), .ZN(n4428) );
  NR2D1BWP12T U3105 ( .A1(n4056), .A2(n4428), .ZN(n2268) );
  CKND2D1BWP12T U3106 ( .A1(n480), .A2(c_in), .ZN(n4436) );
  OAI21D1BWP12T U3107 ( .A1(n3233), .A2(n3332), .B(n4436), .ZN(n4427) );
  OA21D1BWP12T U3108 ( .A1(n4056), .A2(n4433), .B(n4429), .Z(n2267) );
  IOA21D2BWP12T U3109 ( .A1(n2268), .A2(n4427), .B(n2267), .ZN(n4421) );
  NR2D1BWP12T U3110 ( .A1(n2269), .A2(n3661), .ZN(n2416) );
  CKBD1BWP12T U3111 ( .I(n4301), .Z(n2272) );
  NR2D1BWP12T U3112 ( .A1(n2272), .A2(n4541), .ZN(n2418) );
  NR2D1BWP12T U3113 ( .A1(n2416), .A2(n2418), .ZN(n4413) );
  BUFFXD0BWP12T U3114 ( .I(n5030), .Z(n2270) );
  BUFFD1BWP12T U3115 ( .I(n2271), .Z(n4892) );
  NR2D1BWP12T U3116 ( .A1(n3679), .A2(n2640), .ZN(n2946) );
  NR2D1BWP12T U3117 ( .A1(n3937), .A2(n3495), .ZN(n2947) );
  NR2D1BWP12T U3118 ( .A1(n2946), .A2(n2947), .ZN(n2923) );
  NR2D1BWP12T U3119 ( .A1(n2859), .A2(n2863), .ZN(n2274) );
  ND2D1BWP12T U3120 ( .A1(n2923), .A2(n2274), .ZN(n4380) );
  NR2D1BWP12T U3121 ( .A1(n4521), .A2(n5085), .ZN(n4377) );
  NR2D1BWP12T U3122 ( .A1(n4377), .A2(n4387), .ZN(n4402) );
  NR2D1BWP12T U3123 ( .A1(n4406), .A2(n4027), .ZN(n2276) );
  ND2D1BWP12T U3124 ( .A1(n4402), .A2(n2276), .ZN(n2278) );
  NR2D1BWP12T U3125 ( .A1(n4380), .A2(n2278), .ZN(n2280) );
  OAI21D1BWP12T U3126 ( .A1(n2947), .A2(n2945), .B(n2948), .ZN(n2924) );
  ND2D1BWP12T U3127 ( .A1(n2273), .A2(n2909), .ZN(n2927) );
  OAI21D1BWP12T U3128 ( .A1(n4387), .A2(n4382), .B(n4388), .ZN(n4404) );
  OAI21D1BWP12T U3129 ( .A1(n4027), .A2(n4405), .B(n4026), .ZN(n2275) );
  AOI21D1BWP12T U3130 ( .A1(n2276), .A2(n4404), .B(n2275), .ZN(n2277) );
  NR2D1BWP12T U3131 ( .A1(n4788), .A2(n4794), .ZN(n4334) );
  NR2D1BWP12T U3132 ( .A1(n4334), .A2(n3996), .ZN(n2281) );
  NR2D1BWP12T U3133 ( .A1(n4029), .A2(n4061), .ZN(n4330) );
  ND2D1BWP12T U3134 ( .A1(n2281), .A2(n4330), .ZN(n4341) );
  NR2D1BWP12T U3135 ( .A1(n4696), .A2(n16), .ZN(n4343) );
  NR2D1BWP12T U3136 ( .A1(n26), .A2(n5118), .ZN(n2282) );
  NR2D1BWP12T U3137 ( .A1(n4343), .A2(n2282), .ZN(n4351) );
  NR2D1BWP12T U3138 ( .A1(n4356), .A2(n4360), .ZN(n2284) );
  ND2D1BWP12T U3139 ( .A1(n4351), .A2(n2284), .ZN(n2286) );
  NR2D1BWP12T U3140 ( .A1(n4341), .A2(n2286), .ZN(n4365) );
  NR2D1BWP12T U3141 ( .A1(n4914), .A2(n4920), .ZN(n4370) );
  NR2D1BWP12T U3142 ( .A1(n4655), .A2(n4649), .ZN(n4373) );
  NR2D1BWP12T U3143 ( .A1(n4370), .A2(n4373), .ZN(n4453) );
  NR2D1BWP12T U3144 ( .A1(n4568), .A2(n4977), .ZN(n4452) );
  NR2D1BWP12T U3145 ( .A1(n4452), .A2(n2287), .ZN(n2289) );
  ND2D1BWP12T U3146 ( .A1(n4453), .A2(n2289), .ZN(n4458) );
  NR2D1BWP12T U3147 ( .A1(n2255), .A2(n31), .ZN(n4481) );
  NR2D1BWP12T U3148 ( .A1(n4481), .A2(n2290), .ZN(n2292) );
  ND2D1BWP12T U3149 ( .A1(n4475), .A2(n2292), .ZN(n2294) );
  NR2D1BWP12T U3150 ( .A1(n4458), .A2(n2294), .ZN(n2296) );
  TPND2D0BWP12T U3151 ( .A1(n4365), .A2(n2296), .ZN(n2298) );
  OAI21D1BWP12T U3152 ( .A1(n4061), .A2(n4393), .B(n4062), .ZN(n4332) );
  ND2D1BWP12T U3153 ( .A1(n4788), .A2(n4794), .ZN(n4333) );
  TPOAI21D0BWP12T U3154 ( .A1(n2282), .A2(n4342), .B(n4012), .ZN(n4350) );
  OAI21D1BWP12T U3155 ( .A1(n4360), .A2(n4355), .B(n4361), .ZN(n2283) );
  AOI21D1BWP12T U3156 ( .A1(n2284), .A2(n4350), .B(n2283), .ZN(n2285) );
  OAI21D1BWP12T U3157 ( .A1(n4344), .A2(n2286), .B(n2285), .ZN(n4364) );
  ND2D1BWP12T U3158 ( .A1(n4914), .A2(n4920), .ZN(n4369) );
  OAI21D1BWP12T U3159 ( .A1(n4373), .A2(n4369), .B(n4374), .ZN(n4456) );
  ND2D1BWP12T U3160 ( .A1(n4568), .A2(n4977), .ZN(n4454) );
  OAI21D0BWP12T U3161 ( .A1(n2287), .A2(n4454), .B(n3982), .ZN(n2288) );
  AOI21D1BWP12T U3162 ( .A1(n2289), .A2(n4456), .B(n2288), .ZN(n4459) );
  ND2D1BWP12T U3163 ( .A1(n2773), .A2(n21), .ZN(n2756) );
  OAI21D0BWP12T U3164 ( .A1(n3974), .A2(n2756), .B(n3973), .ZN(n4479) );
  OAI21D0BWP12T U3165 ( .A1(n2290), .A2(n4480), .B(n3991), .ZN(n2291) );
  TPAOI21D0BWP12T U3166 ( .A1(n2292), .A2(n4479), .B(n2291), .ZN(n2293) );
  TPOAI21D0BWP12T U3167 ( .A1(n4459), .A2(n2294), .B(n2293), .ZN(n2295) );
  TPAOI21D0BWP12T U3168 ( .A1(n4364), .A2(n2296), .B(n2295), .ZN(n2297) );
  OAI21D1BWP12T U3169 ( .A1(n2753), .A2(n2298), .B(n2297), .ZN(n2622) );
  OR2XD1BWP12T U3170 ( .A1(n5108), .A2(n3936), .Z(n2621) );
  ND2D1BWP12T U3171 ( .A1(n5108), .A2(n3936), .ZN(n2620) );
  ND2D1BWP12T U3172 ( .A1(n2621), .A2(n2620), .ZN(n2299) );
  XNR2XD1BWP12T U3173 ( .A1(n2622), .A2(n2299), .ZN(n4450) );
  INVD1P75BWP12T U3174 ( .I(n4822), .ZN(n4578) );
  ND2D1BWP12T U3175 ( .A1(n4790), .A2(n4578), .ZN(n4580) );
  INVD2BWP12T U3176 ( .I(a[18]), .ZN(n3889) );
  INVD1P75BWP12T U3177 ( .I(n5118), .ZN(n3888) );
  ND2D1BWP12T U3178 ( .A1(n3887), .A2(n3888), .ZN(n4529) );
  CKND2BWP12T U3179 ( .I(n4649), .ZN(n4651) );
  ND2D1BWP12T U3180 ( .A1(n4975), .A2(n4651), .ZN(n4570) );
  ND2D1BWP12T U3181 ( .A1(n3898), .A2(n3900), .ZN(n4519) );
  INVD1P25BWP12T U3182 ( .I(n2848), .ZN(n3897) );
  INVD1BWP12T U3183 ( .I(n4502), .ZN(n3896) );
  INVD1P75BWP12T U3184 ( .I(n5234), .ZN(n5235) );
  ND2D1BWP12T U3185 ( .A1(n3896), .A2(n5235), .ZN(n4575) );
  INVD1BWP12T U3186 ( .I(n4508), .ZN(n2300) );
  CKND2D1BWP12T U3187 ( .A1(n2300), .A2(n5260), .ZN(n2301) );
  NR2D1BWP12T U3188 ( .A1(n4575), .A2(n2301), .ZN(n2302) );
  ND2D1BWP12T U3189 ( .A1(n4574), .A2(n2302), .ZN(n2306) );
  ND2D1BWP12T U3190 ( .A1(n3015), .A2(n1812), .ZN(n2706) );
  NR3D2BWP12T U3191 ( .A1(n5192), .A2(n3661), .A3(n2706), .ZN(n2634) );
  ND2D1BWP12T U3192 ( .A1(n5032), .A2(n3912), .ZN(n4542) );
  INVD1BWP12T U3193 ( .I(n4891), .ZN(n3910) );
  ND2D1BWP12T U3194 ( .A1(n2303), .A2(n3910), .ZN(n2304) );
  NR2D1BWP12T U3195 ( .A1(n4542), .A2(n2304), .ZN(n2305) );
  ND2D1BWP12T U3196 ( .A1(n2634), .A2(n2305), .ZN(n2822) );
  NR2D3BWP12T U3197 ( .A1(n2306), .A2(n2822), .ZN(n4582) );
  INVD1BWP12T U3198 ( .I(n2612), .ZN(n2615) );
  NR2XD0BWP12T U3199 ( .A1(op[2]), .A2(op[1]), .ZN(n2353) );
  ND2XD4BWP12T U3200 ( .A1(n4849), .A2(n5196), .ZN(n3869) );
  MUX2XD0BWP12T U3201 ( .I0(n5030), .I1(n4541), .S(b[0]), .Z(n4134) );
  IND2XD16BWP12T U3202 ( .A1(n5196), .B1(n3908), .ZN(n3871) );
  TPOAI22D0BWP12T U3203 ( .A1(n4133), .A2(n3869), .B1(n4134), .B2(n3871), .ZN(
        n2308) );
  MUX2XD0BWP12T U3204 ( .I0(n4510), .I1(n4891), .S(b[0]), .Z(n2890) );
  TPND2D3BWP12T U3205 ( .A1(n2834), .A2(n4175), .ZN(n3872) );
  MUX2XD0BWP12T U3206 ( .I0(n3570), .I1(n5192), .S(b[0]), .Z(n4132) );
  IND2XD2BWP12T U3207 ( .A1(n3908), .B1(n5196), .ZN(n3870) );
  TPOAI22D0BWP12T U3208 ( .A1(n2890), .A2(n3872), .B1(n4132), .B2(n3870), .ZN(
        n2307) );
  NR2D1BWP12T U3209 ( .A1(n2308), .A2(n2307), .ZN(n3848) );
  CKND2D2BWP12T U3210 ( .A1(n3948), .A2(n4301), .ZN(n3858) );
  MUX2XD0BWP12T U3211 ( .I0(n4502), .I1(n5234), .S(b[0]), .Z(n4140) );
  MUX2XD0BWP12T U3212 ( .I0(n4508), .I1(a[14]), .S(b[0]), .Z(n4131) );
  OAI22D0BWP12T U3213 ( .A1(n4140), .A2(n3871), .B1(n4131), .B2(n3872), .ZN(
        n2310) );
  MUX2XD0BWP12T U3214 ( .I0(n4511), .I1(n3495), .S(b[0]), .Z(n2889) );
  MUX2D1BWP12T U3215 ( .I0(n5079), .I1(n2848), .S(b[0]), .Z(n4152) );
  OAI22D0BWP12T U3216 ( .A1(n2889), .A2(n3869), .B1(n4152), .B2(n3870), .ZN(
        n2309) );
  NR2D1BWP12T U3217 ( .A1(n2310), .A2(n2309), .ZN(n3846) );
  BUFFD3BWP12T U3218 ( .I(n2311), .Z(n3882) );
  NR2D1BWP12T U3219 ( .A1(n3882), .A2(n3948), .ZN(n4262) );
  INVD1BWP12T U3220 ( .I(n4262), .ZN(n3859) );
  OAI22D0BWP12T U3221 ( .A1(n3848), .A2(n3858), .B1(n3846), .B2(n3859), .ZN(
        n2342) );
  INVD4BWP12T U3222 ( .I(n3872), .ZN(n3855) );
  MUX2ND0BWP12T U3223 ( .I0(n4914), .I1(n2825), .S(b[0]), .ZN(n4164) );
  MUX2ND0BWP12T U3224 ( .I0(n4672), .I1(n5118), .S(b[0]), .ZN(n4166) );
  INVD2BWP12T U3225 ( .I(n3871), .ZN(n3854) );
  AOI22D0BWP12T U3226 ( .A1(n3855), .A2(n4164), .B1(n4166), .B2(n3854), .ZN(
        n2313) );
  INVD2BWP12T U3227 ( .I(n3869), .ZN(n3853) );
  MUX2ND0BWP12T U3228 ( .I0(n4788), .I1(n4822), .S(b[0]), .ZN(n3757) );
  MUX2ND0BWP12T U3229 ( .I0(n4565), .I1(a[18]), .S(b[0]), .ZN(n4163) );
  INVD1P75BWP12T U3230 ( .I(n3870), .ZN(n3852) );
  AOI22D0BWP12T U3231 ( .A1(n3853), .A2(n3757), .B1(n4163), .B2(n3852), .ZN(
        n2312) );
  ND2D1BWP12T U3232 ( .A1(n2313), .A2(n2312), .ZN(n3845) );
  IND2D1BWP12T U3233 ( .A1(n4301), .B1(n3948), .ZN(n3861) );
  INR2D0BWP12T U3234 ( .A1(n3845), .B1(n3861), .ZN(n2341) );
  OR2XD8BWP12T U3235 ( .A1(n4849), .A2(b[0]), .Z(n3588) );
  INR2XD2BWP12T U3236 ( .A1(n3906), .B1(n3588), .ZN(n2363) );
  INVD4BWP12T U3237 ( .I(n2363), .ZN(n3594) );
  OR2D2BWP12T U3238 ( .A1(n3948), .A2(n4301), .Z(n4953) );
  NR2D1BWP12T U3239 ( .A1(n3594), .A2(n4953), .ZN(n4170) );
  INVD1BWP12T U3240 ( .I(n4170), .ZN(n4185) );
  MUX2ND0BWP12T U3241 ( .I0(n4568), .I1(n4649), .S(b[0]), .ZN(n4165) );
  INVD1BWP12T U3242 ( .I(n4165), .ZN(n4241) );
  MUX2ND0BWP12T U3243 ( .I0(n4990), .I1(n1), .S(n402), .ZN(n3794) );
  INVD0BWP12T U3244 ( .I(n3794), .ZN(n4247) );
  OAI22D0BWP12T U3245 ( .A1(n4241), .A2(n3869), .B1(n4247), .B2(n3871), .ZN(
        n2316) );
  MUX2ND4BWP12T U3246 ( .I0(n2773), .I1(n4943), .S(n402), .ZN(n3793) );
  INVD1BWP12T U3247 ( .I(n3793), .ZN(n4246) );
  OAI22D1BWP12T U3248 ( .A1(n4246), .A2(n3870), .B1(n3806), .B2(n5146), .ZN(
        n2315) );
  INVD1BWP12T U3249 ( .I(n4953), .ZN(n4178) );
  OAI21D0BWP12T U3250 ( .A1(n2316), .A2(n2315), .B(n4178), .ZN(n2339) );
  NR2D1BWP12T U3251 ( .A1(n3930), .A2(n3937), .ZN(n2318) );
  CKND2D1BWP12T U3252 ( .A1(n2318), .A2(n2317), .ZN(n2325) );
  TPNR2D1BWP12T U3253 ( .A1(n31), .A2(n22), .ZN(n2320) );
  TPNR2D1BWP12T U3254 ( .A1(n3936), .A2(n5153), .ZN(n2322) );
  TPND2D1BWP12T U3255 ( .A1(n2322), .A2(n2321), .ZN(n2323) );
  TPNR2D1BWP12T U3256 ( .A1(n4977), .A2(n4655), .ZN(n2327) );
  ND2D1BWP12T U3257 ( .A1(n2327), .A2(n2326), .ZN(n2331) );
  TPNR2D1BWP12T U3258 ( .A1(n17), .A2(n26), .ZN(n2329) );
  TPNR2D1BWP12T U3259 ( .A1(n16), .A2(n25), .ZN(n2328) );
  ND2D1BWP12T U3260 ( .A1(n2329), .A2(n2328), .ZN(n2330) );
  NR2D1BWP12T U3261 ( .A1(n4794), .A2(n4826), .ZN(n2333) );
  NR2D1BWP12T U3262 ( .A1(n5264), .A2(n32), .ZN(n2332) );
  ND2D1BWP12T U3263 ( .A1(n2333), .A2(n2332), .ZN(n2335) );
  TPNR2D2BWP12T U3264 ( .A1(n2335), .A2(n2334), .ZN(n2336) );
  ND3XD8BWP12T U3265 ( .A1(n2338), .A2(n2337), .A3(n2336), .ZN(n3838) );
  OAI211D0BWP12T U3266 ( .A1(n5108), .A2(n4185), .B(n2339), .C(n3875), .ZN(
        n2340) );
  NR3D1BWP12T U3267 ( .A1(n2342), .A2(n2341), .A3(n2340), .ZN(n3805) );
  CKND0BWP12T U3268 ( .I(op[3]), .ZN(n2343) );
  TPND2D2BWP12T U3269 ( .A1(n2344), .A2(n2343), .ZN(n5232) );
  INVD2BWP12T U3270 ( .I(n5232), .ZN(n5252) );
  CKND2D1BWP12T U3271 ( .A1(op[0]), .A2(op[1]), .ZN(n2346) );
  INVD1BWP12T U3272 ( .I(n2346), .ZN(n2345) );
  INVD4BWP12T U3273 ( .I(n5312), .ZN(n5281) );
  IND2XD2BWP12T U3274 ( .A1(n4301), .B1(n5281), .ZN(n4889) );
  NR3D1BWP12T U3275 ( .A1(n2346), .A2(op[3]), .A3(op[2]), .ZN(n5212) );
  INR2D2BWP12T U3276 ( .A1(n5212), .B1(n3844), .ZN(n4974) );
  INR2D2BWP12T U3277 ( .A1(n4889), .B1(n4974), .ZN(n4924) );
  INVD1BWP12T U3278 ( .I(n4924), .ZN(n5126) );
  IND2D1BWP12T U3279 ( .A1(n3948), .B1(n5108), .ZN(n2347) );
  NR2D1BWP12T U3280 ( .A1(n3594), .A2(n2347), .ZN(n3726) );
  ND2D0BWP12T U3281 ( .A1(op[3]), .A2(op[2]), .ZN(n2354) );
  INR2D4BWP12T U3282 ( .A1(n2348), .B1(n2354), .ZN(n3925) );
  CKND0BWP12T U3283 ( .I(n3925), .ZN(n2350) );
  NR2D1BWP12T U3284 ( .A1(op[0]), .A2(op[1]), .ZN(n2425) );
  OAI21D1BWP12T U3285 ( .A1(n3936), .A2(op[2]), .B(n2425), .ZN(n2349) );
  OAI21D1BWP12T U3286 ( .A1(n3936), .A2(n2350), .B(n2349), .ZN(n2352) );
  MUX2ND0BWP12T U3287 ( .I0(n2352), .I1(n5236), .S(n3564), .ZN(n2358) );
  XOR2D1BWP12T U3288 ( .A1(n3936), .A2(n5108), .Z(n5106) );
  INVD1BWP12T U3289 ( .I(n2423), .ZN(n5289) );
  INR2D2BWP12T U3290 ( .A1(n2425), .B1(n2354), .ZN(n5296) );
  INVD4BWP12T U3291 ( .I(n5296), .ZN(n5254) );
  NR2XD0BWP12T U3292 ( .A1(n2355), .A2(n5254), .ZN(n2356) );
  AOI21D1BWP12T U3293 ( .A1(n5106), .A2(n5289), .B(n2356), .ZN(n2357) );
  CKND2D1BWP12T U3294 ( .A1(n2358), .A2(n2357), .ZN(n2359) );
  AOI21D1BWP12T U3295 ( .A1(n5126), .A2(n3726), .B(n2359), .ZN(n2360) );
  IOA21D1BWP12T U3296 ( .A1(n3805), .A2(n5252), .B(n2360), .ZN(n2361) );
  AOI21D1BWP12T U3297 ( .A1(n5102), .A2(n5297), .B(n2361), .ZN(n2377) );
  BUFFD3BWP12T U3298 ( .I(n2362), .Z(n3905) );
  XNR2XD4BWP12T U3299 ( .A1(n2363), .A2(n2269), .ZN(n4297) );
  INVD2BWP12T U3300 ( .I(n4297), .ZN(n4277) );
  INVD3BWP12T U3301 ( .I(n3858), .ZN(n4260) );
  TPAOI21D4BWP12T U3302 ( .A1(n3594), .A2(n4301), .B(n4260), .ZN(n4299) );
  NR2D2BWP12T U3303 ( .A1(n4277), .A2(n4299), .ZN(n4267) );
  INVD2BWP12T U3304 ( .I(n4267), .ZN(n4815) );
  INVD2BWP12T U3305 ( .I(n5196), .ZN(n4175) );
  TPNR2D2BWP12T U3306 ( .A1(n3498), .A2(n4175), .ZN(n2364) );
  INVD1P75BWP12T U3307 ( .I(n2364), .ZN(n2678) );
  ND2D3BWP12T U3308 ( .A1(n2678), .A2(n3594), .ZN(n4201) );
  INVD2BWP12T U3309 ( .I(n4201), .ZN(n2976) );
  ND2XD8BWP12T U3310 ( .A1(n3908), .A2(b[0]), .ZN(n3587) );
  ND2D3BWP12T U3311 ( .A1(n3588), .A2(n3587), .ZN(n2677) );
  TPND2D3BWP12T U3312 ( .A1(n2976), .A2(n2677), .ZN(n4311) );
  TPND2D0BWP12T U3313 ( .A1(n4242), .A2(n4163), .ZN(n2367) );
  INVD1P75BWP12T U3314 ( .I(n2677), .ZN(n2974) );
  TPND2D2BWP12T U3315 ( .A1(n2974), .A2(n2364), .ZN(n4313) );
  INVD1BWP12T U3316 ( .I(n4313), .ZN(n4245) );
  IND2D2BWP12T U3317 ( .A1(n2364), .B1(n2974), .ZN(n4315) );
  INVD1P75BWP12T U3318 ( .I(n4315), .ZN(n4244) );
  AOI22D0BWP12T U3319 ( .A1(n4245), .A2(n4166), .B1(n4244), .B2(n3757), .ZN(
        n2366) );
  CKND2D1BWP12T U3320 ( .A1(n2839), .A2(n4164), .ZN(n2365) );
  ND3D1BWP12T U3321 ( .A1(n2367), .A2(n2366), .A3(n2365), .ZN(n4192) );
  INVD1P75BWP12T U3322 ( .I(n4299), .ZN(n4281) );
  NR2D1BWP12T U3323 ( .A1(n4281), .A2(n4170), .ZN(n2368) );
  ND2D1BWP12T U3324 ( .A1(n2368), .A2(n4277), .ZN(n4817) );
  INVD1BWP12T U3325 ( .I(n4131), .ZN(n4150) );
  TPNR2D0BWP12T U3326 ( .A1(n4309), .A2(n4150), .ZN(n2371) );
  INVD1BWP12T U3327 ( .I(n4152), .ZN(n4138) );
  NR2D1BWP12T U3328 ( .A1(n4311), .A2(n4138), .ZN(n2370) );
  INVD1BWP12T U3329 ( .I(n2889), .ZN(n4137) );
  INVD1BWP12T U3330 ( .I(n4140), .ZN(n4151) );
  OAI22D1BWP12T U3331 ( .A1(n4315), .A2(n4137), .B1(n4313), .B2(n4151), .ZN(
        n2369) );
  NR3D1BWP12T U3332 ( .A1(n2371), .A2(n2370), .A3(n2369), .ZN(n4266) );
  INVD3BWP12T U3333 ( .I(n4208), .ZN(n5183) );
  TPNR2D0BWP12T U3334 ( .A1(n4311), .A2(n3793), .ZN(n2373) );
  OAI22D0BWP12T U3335 ( .A1(n4315), .A2(n4165), .B1(n4313), .B2(n3794), .ZN(
        n2372) );
  RCAOI211D0BWP12T U3336 ( .A1(n2839), .A2(n5146), .B(n2373), .C(n2372), .ZN(
        n2374) );
  OAI222D1BWP12T U3337 ( .A1(n4815), .A2(n4192), .B1(n4817), .B2(n4266), .C1(
        n5183), .C2(n2374), .ZN(n4324) );
  INVD1BWP12T U3338 ( .I(n2890), .ZN(n4139) );
  INVD1BWP12T U3339 ( .I(n4132), .ZN(n3762) );
  INVD1BWP12T U3340 ( .I(n4133), .ZN(n3760) );
  INVD1BWP12T U3341 ( .I(n4134), .ZN(n3761) );
  ND2D1BWP12T U3342 ( .A1(n4297), .A2(n4299), .ZN(n5162) );
  NR2D1BWP12T U3343 ( .A1(n4203), .A2(n5162), .ZN(n2375) );
  OAI21D1BWP12T U3344 ( .A1(n4324), .A2(n2375), .B(n5281), .ZN(n2376) );
  ND2D1BWP12T U3345 ( .A1(n2377), .A2(n2376), .ZN(n2378) );
  AOI21D1BWP12T U3346 ( .A1(n5313), .A2(n4450), .B(n2378), .ZN(n2379) );
  IOA21D1BWP12T U3347 ( .A1(n3324), .A2(n5308), .B(n2379), .ZN(n2380) );
  AOI21D1BWP12T U3348 ( .A1(n5303), .A2(n4036), .B(n2380), .ZN(n2381) );
  IOA21D2BWP12T U3349 ( .A1(n3315), .A2(n5305), .B(n2381), .ZN(n2382) );
  INVD3BWP12T U3350 ( .I(n2382), .ZN(n2383) );
  ND2D3BWP12T U3351 ( .A1(n3024), .A2(n3025), .ZN(n2385) );
  XOR2D2BWP12T U3352 ( .A1(n2385), .A2(n3027), .Z(n3031) );
  INVD1BWP12T U3353 ( .I(n3031), .ZN(n2457) );
  INVD1BWP12T U3354 ( .I(n2386), .ZN(n3222) );
  INVD1BWP12T U3355 ( .I(n3213), .ZN(n2435) );
  IND2XD8BWP12T U3356 ( .A1(b[1]), .B1(b[0]), .ZN(n3589) );
  OA22D1BWP12T U3357 ( .A1(n3588), .A2(n4651), .B1(n3589), .B2(n4975), .Z(
        n2389) );
  MUX2XD2BWP12T U3358 ( .I0(n4943), .I1(n4503), .S(b[0]), .Z(n2831) );
  ND2D1BWP12T U3359 ( .A1(n2831), .A2(n3908), .ZN(n2388) );
  ND2D1BWP12T U3360 ( .A1(n2389), .A2(n2388), .ZN(n3536) );
  INVD1BWP12T U3361 ( .I(n5196), .ZN(n3553) );
  OR2D2BWP12T U3362 ( .A1(n3536), .A2(n3553), .Z(n2391) );
  IND2XD8BWP12T U3363 ( .A1(b[0]), .B1(n4849), .ZN(n3591) );
  TPND2D1BWP12T U3364 ( .A1(n3535), .A2(n3553), .ZN(n2390) );
  NR2D2BWP12T U3365 ( .A1(n3905), .A2(n5196), .ZN(n3707) );
  INVD3BWP12T U3366 ( .I(n3707), .ZN(n3618) );
  OAI22D1BWP12T U3367 ( .A1(n3588), .A2(n4607), .B1(n3564), .B2(n3587), .ZN(
        n2393) );
  INVD1BWP12T U3368 ( .I(n5146), .ZN(n5148) );
  OAI22D1BWP12T U3369 ( .A1(n3591), .A2(n5148), .B1(n3589), .B2(n407), .ZN(
        n2392) );
  TPNR2D1BWP12T U3370 ( .A1(n2393), .A2(n2392), .ZN(n3731) );
  INVD1P75BWP12T U3371 ( .I(n3731), .ZN(n4602) );
  INVD2BWP12T U3372 ( .I(n4602), .ZN(n2394) );
  ND2D1BWP12T U3373 ( .A1(n3948), .A2(n5108), .ZN(n3524) );
  OAI21D0BWP12T U3374 ( .A1(n3524), .A2(n3906), .B(n4301), .ZN(n2395) );
  TPNR2D1BWP12T U3375 ( .A1(n5127), .A2(n2395), .ZN(n2411) );
  INVD2P3BWP12T U3376 ( .I(n3587), .ZN(n3497) );
  AOI22D0BWP12T U3377 ( .A1(n3498), .A2(n3900), .B1(n3497), .B2(n5081), .ZN(
        n2399) );
  NR2D0BWP12T U3378 ( .A1(n3591), .A2(n2848), .ZN(n2397) );
  NR2D1BWP12T U3379 ( .A1(n3589), .A2(n4511), .ZN(n2396) );
  NR2D1BWP12T U3380 ( .A1(n2397), .A2(n2396), .ZN(n2398) );
  CKND2D1BWP12T U3381 ( .A1(n2399), .A2(n2398), .ZN(n3568) );
  IND2XD2BWP12T U3382 ( .A1(n3948), .B1(n5196), .ZN(n3607) );
  TPOAI21D0BWP12T U3383 ( .A1(n3568), .A2(n3607), .B(n3882), .ZN(n2401) );
  ND2D1BWP12T U3384 ( .A1(n3948), .A2(n5196), .ZN(n3609) );
  NR2D1BWP12T U3385 ( .A1(n3558), .A2(n3609), .ZN(n2400) );
  TPNR2D1BWP12T U3386 ( .A1(n2401), .A2(n2400), .ZN(n2409) );
  INVD1P75BWP12T U3387 ( .I(n3591), .ZN(n3496) );
  INVD2BWP12T U3388 ( .I(n3589), .ZN(n3494) );
  AOI22D0BWP12T U3389 ( .A1(n3496), .A2(n4891), .B1(n3494), .B2(n5030), .ZN(
        n2403) );
  AOI22D0BWP12T U3390 ( .A1(n3498), .A2(n4541), .B1(n3497), .B2(n4510), .ZN(
        n2402) );
  CKND2D1BWP12T U3391 ( .A1(n2403), .A2(n2402), .ZN(n3572) );
  OR2D4BWP12T U3392 ( .A1(n3948), .A2(n5196), .Z(n3730) );
  INVD2BWP12T U3393 ( .I(n3730), .ZN(n4601) );
  AOI22D1BWP12T U3394 ( .A1(n3498), .A2(n5234), .B1(n3497), .B2(n4508), .ZN(
        n2407) );
  NR2D1BWP12T U3395 ( .A1(n3591), .A2(n5260), .ZN(n2405) );
  NR2D1BWP12T U3396 ( .A1(n3589), .A2(n3896), .ZN(n2404) );
  NR2D1BWP12T U3397 ( .A1(n2405), .A2(n2404), .ZN(n2406) );
  TPND2D1BWP12T U3398 ( .A1(n2407), .A2(n2406), .ZN(n3559) );
  AOI22D1BWP12T U3399 ( .A1(n3572), .A2(n4601), .B1(n3707), .B2(n3559), .ZN(
        n2408) );
  TPND2D1BWP12T U3400 ( .A1(n2409), .A2(n2408), .ZN(n2446) );
  CKND2D1BWP12T U3401 ( .A1(n2446), .A2(n3875), .ZN(n2410) );
  ND2D4BWP12T U3402 ( .A1(n3838), .A2(n5108), .ZN(n3565) );
  OAI21D1BWP12T U3403 ( .A1(n2411), .A2(n2410), .B(n3565), .ZN(n3566) );
  INVD1P75BWP12T U3404 ( .I(n2412), .ZN(n2413) );
  CKND2D1BWP12T U3405 ( .A1(n3566), .A2(n5322), .ZN(n2434) );
  MUX2ND0BWP12T U3406 ( .I0(n5192), .I1(n4501), .S(b[0]), .ZN(n4198) );
  INR2D2BWP12T U3407 ( .A1(n480), .B1(n3588), .ZN(n2964) );
  INVD1BWP12T U3408 ( .I(n2964), .ZN(n3571) );
  AOI22D0BWP12T U3409 ( .A1(n3854), .A2(n4198), .B1(n3571), .B2(n5196), .ZN(
        n2415) );
  MUX2XD0BWP12T U3410 ( .I0(n3912), .I1(n512), .S(b[0]), .Z(n4199) );
  CKND2D1BWP12T U3411 ( .A1(n4199), .A2(n3855), .ZN(n2414) );
  TPND2D1BWP12T U3412 ( .A1(n2415), .A2(n2414), .ZN(n3790) );
  INVD1BWP12T U3413 ( .I(n3790), .ZN(n3828) );
  INR2D1BWP12T U3414 ( .A1(n5252), .B1(n3948), .ZN(n2664) );
  ND2XD0BWP12T U3415 ( .A1(n3828), .A2(n2664), .ZN(n2422) );
  INVD1BWP12T U3416 ( .I(n2416), .ZN(n2691) );
  INVD1BWP12T U3417 ( .I(n2703), .ZN(n2417) );
  TPAOI21D1BWP12T U3418 ( .A1(n4421), .A2(n2691), .B(n2417), .ZN(n2420) );
  NR2D1BWP12T U3419 ( .A1(n4044), .A2(n2418), .ZN(n2419) );
  XNR2D2BWP12T U3420 ( .A1(n2420), .A2(n2419), .ZN(n4412) );
  CKND2D1BWP12T U3421 ( .A1(n4412), .A2(n5313), .ZN(n2421) );
  OAI21D1BWP12T U3422 ( .A1(n3844), .A2(n2422), .B(n2421), .ZN(n2432) );
  INVD1BWP12T U3423 ( .I(n2446), .ZN(n4288) );
  INVD2BWP12T U3424 ( .I(n5289), .ZN(n5255) );
  OAI21D0BWP12T U3425 ( .A1(n4541), .A2(n5255), .B(n5254), .ZN(n2429) );
  INR2XD2BWP12T U3426 ( .A1(n2423), .B1(n3925), .ZN(n5295) );
  INVD2BWP12T U3427 ( .I(n5295), .ZN(n5258) );
  CKND0BWP12T U3428 ( .I(op[2]), .ZN(n2424) );
  ND2D1BWP12T U3429 ( .A1(n2425), .A2(n2424), .ZN(n5294) );
  INVD1P75BWP12T U3430 ( .I(n5294), .ZN(n5257) );
  MUX2D1BWP12T U3431 ( .I0(n5258), .I1(n5257), .S(n4301), .Z(n2426) );
  NR2D0BWP12T U3432 ( .A1(n2426), .A2(n5296), .ZN(n2427) );
  INVD2BWP12T U3433 ( .I(n5236), .ZN(n5299) );
  MUX2NXD0BWP12T U3434 ( .I0(n2427), .I1(n5299), .S(n3912), .ZN(n2428) );
  AOI21D1BWP12T U3435 ( .A1(n4301), .A2(n2429), .B(n2428), .ZN(n2430) );
  OAI21D1BWP12T U3436 ( .A1(n4288), .A2(n4889), .B(n2430), .ZN(n2431) );
  TPNR2D1BWP12T U3437 ( .A1(n2432), .A2(n2431), .ZN(n2433) );
  OAI211D1BWP12T U3438 ( .A1(n5203), .A2(n2435), .B(n2434), .C(n2433), .ZN(
        n2455) );
  INVD1BWP12T U3439 ( .I(n2436), .ZN(n2714) );
  CKND2BWP12T U3440 ( .I(n2716), .ZN(n3350) );
  INVD1BWP12T U3441 ( .I(n2713), .ZN(n2437) );
  RCAOI21D1BWP12T U3442 ( .A1(n2714), .A2(n3350), .B(n2437), .ZN(n2441) );
  CKND2D1BWP12T U3443 ( .A1(n3217), .A2(n2439), .ZN(n2440) );
  XOR2XD1BWP12T U3444 ( .A1(n2441), .A2(n2440), .Z(n3339) );
  INVD1BWP12T U3445 ( .I(n3339), .ZN(n2445) );
  INVD1BWP12T U3446 ( .I(n2442), .ZN(n4050) );
  INVD1BWP12T U3447 ( .I(n2443), .ZN(n4045) );
  XNR2XD1BWP12T U3448 ( .A1(n2634), .A2(n4541), .ZN(n4539) );
  AOI22D1BWP12T U3449 ( .A1(n4055), .A2(n5303), .B1(n5297), .B2(n4539), .ZN(
        n2444) );
  TPOAI21D0BWP12T U3450 ( .A1(n2445), .A2(n5105), .B(n2444), .ZN(n2454) );
  NR2D1BWP12T U3451 ( .A1(n3737), .A2(n5327), .ZN(n2453) );
  ND2D1BWP12T U3452 ( .A1(n5127), .A2(n2446), .ZN(n2451) );
  INVD1BWP12T U3453 ( .I(n4198), .ZN(n2975) );
  INR2D1BWP12T U3454 ( .A1(n2975), .B1(n4313), .ZN(n2449) );
  INVD1BWP12T U3455 ( .I(n4199), .ZN(n3781) );
  INR2D1BWP12T U3456 ( .A1(n3781), .B1(n4309), .ZN(n2448) );
  INR2D1BWP12T U3457 ( .A1(n3594), .B1(n3571), .ZN(n2447) );
  TPNR3D1BWP12T U3458 ( .A1(n2449), .A2(n2448), .A3(n2447), .ZN(n4319) );
  TPNR2D1BWP12T U3459 ( .A1(n4319), .A2(n5183), .ZN(n2450) );
  INR2D1BWP12T U3460 ( .A1(n2451), .B1(n2450), .ZN(n4273) );
  TPNR2D1BWP12T U3461 ( .A1(n4273), .A2(n5312), .ZN(n2452) );
  NR4D0BWP12T U3462 ( .A1(n2455), .A2(n2454), .A3(n2453), .A4(n2452), .ZN(
        n2456) );
  RCOAI21D2BWP12T U3463 ( .A1(n2457), .A2(n5112), .B(n2456), .ZN(result[4]) );
  TPAOI21D1BWP12T U3464 ( .A1(n2461), .A2(n2460), .B(n2459), .ZN(n2602) );
  XNR2XD0BWP12T U3465 ( .A1(n5079), .A2(b[22]), .ZN(n2466) );
  OAI22D0BWP12T U3466 ( .A1(n2468), .A2(n420), .B1(n2466), .B2(n2465), .ZN(
        n2473) );
  XOR3D1BWP12T U3467 ( .A1(n2474), .A2(n2473), .A3(n2472), .Z(n2491) );
  AO21D0BWP12T U3468 ( .A1(n2476), .A2(n3015), .B(n2475), .Z(n2485) );
  XNR2XD0BWP12T U3469 ( .A1(n4511), .A2(n4655), .ZN(n2480) );
  OAI22D0BWP12T U3470 ( .A1(n1689), .A2(n2482), .B1(n2481), .B2(n2480), .ZN(
        n2483) );
  FA1D2BWP12T U3471 ( .A(n2488), .B(n2487), .CI(n2486), .CO(n2489), .S(n2496)
         );
  XOR3D1BWP12T U3472 ( .A1(n2491), .A2(n2490), .A3(n2489), .Z(n2503) );
  CKND2BWP12T U3473 ( .I(n2496), .ZN(n2494) );
  CKND1BWP12T U3474 ( .I(n2497), .ZN(n2493) );
  IOA21D2BWP12T U3475 ( .A1(n2494), .A2(n2493), .B(n2492), .ZN(n2495) );
  IOA21D2BWP12T U3476 ( .A1(n2497), .A2(n2496), .B(n2495), .ZN(n2502) );
  FA1D2BWP12T U3477 ( .A(n2500), .B(n2499), .CI(n2498), .CO(n2501), .S(n2506)
         );
  FA1D2BWP12T U3478 ( .A(n2506), .B(n2505), .CI(n2504), .CO(n2592), .S(n2593)
         );
  FA1D2BWP12T U3479 ( .A(n2509), .B(n2508), .CI(n2507), .CO(n2544), .S(n2586)
         );
  FA1D2BWP12T U3480 ( .A(n2512), .B(n2511), .CI(n2510), .CO(n2543), .S(n2498)
         );
  FA1D0BWP12T U3481 ( .A(n2515), .B(n2514), .CI(n2513), .CO(n2541), .S(n2507)
         );
  XOR3D1BWP12T U3482 ( .A1(n2526), .A2(n2525), .A3(n2524), .Z(n2540) );
  XOR3D1BWP12T U3483 ( .A1(n2538), .A2(n2537), .A3(n2536), .Z(n2539) );
  XOR3D2BWP12T U3484 ( .A1(n2541), .A2(n2540), .A3(n2539), .Z(n2542) );
  XOR3D2BWP12T U3485 ( .A1(n2544), .A2(n2543), .A3(n2542), .Z(n2590) );
  OAI21D1BWP12T U3486 ( .A1(n2553), .A2(n2552), .B(n2550), .ZN(n2551) );
  IOA21D1BWP12T U3487 ( .A1(n2553), .A2(n2552), .B(n2551), .ZN(n2558) );
  FA1D2BWP12T U3488 ( .A(n2556), .B(n2555), .CI(n2554), .CO(n2557), .S(n2561)
         );
  XOR3D1BWP12T U3489 ( .A1(n2559), .A2(n2558), .A3(n2557), .Z(n2584) );
  OAI21D1BWP12T U3490 ( .A1(n2562), .A2(n2561), .B(n2560), .ZN(n2564) );
  ND2D1BWP12T U3491 ( .A1(n2564), .A2(n2563), .ZN(n2583) );
  FA1D2BWP12T U3492 ( .A(n2567), .B(n2566), .CI(n2565), .CO(n2581), .S(n2562)
         );
  HA1D1BWP12T U3493 ( .A(n2577), .B(n2576), .CO(n2578), .S(n2487) );
  XOR3D1BWP12T U3494 ( .A1(n2581), .A2(n2580), .A3(n2579), .Z(n2582) );
  XOR3D2BWP12T U3495 ( .A1(n2584), .A2(n2583), .A3(n2582), .Z(n2589) );
  FA1D2BWP12T U3496 ( .A(n2587), .B(n2586), .CI(n2585), .CO(n2588), .S(n2594)
         );
  XOR3D2BWP12T U3497 ( .A1(n2590), .A2(n2589), .A3(n2588), .Z(n2591) );
  FA1D2BWP12T U3498 ( .A(n2595), .B(n2594), .CI(n2593), .CO(n2597), .S(n2137)
         );
  INVD1P75BWP12T U3499 ( .I(n2597), .ZN(n2596) );
  IND2D2BWP12T U3500 ( .A1(n2598), .B1(n2596), .ZN(n2600) );
  ND2D1BWP12T U3501 ( .A1(n2598), .A2(n2597), .ZN(n2599) );
  XNR2XD4BWP12T U3502 ( .A1(n2602), .A2(n2601), .ZN(n5101) );
  NR2D0BWP12T U3503 ( .A1(n5148), .A2(n2615), .ZN(n2610) );
  MUX2ND0BWP12T U3504 ( .I0(n2610), .I1(n2612), .S(n4557), .ZN(n2611) );
  MUX2NXD0BWP12T U3505 ( .I0(n2615), .I1(n2611), .S(n4559), .ZN(n2613) );
  MUX2ND0BWP12T U3506 ( .I0(n2613), .I1(n2612), .S(n4571), .ZN(n2614) );
  MUX2ND0BWP12T U3507 ( .I0(n2615), .I1(n2614), .S(n4582), .ZN(n5103) );
  TPND2D0BWP12T U3508 ( .A1(n5103), .A2(n5297), .ZN(n2624) );
  ND3D1BWP12T U3509 ( .A1(n5107), .A2(n2624), .A3(n2623), .ZN(n2625) );
  AO21D2BWP12T U3510 ( .A1(n5101), .A2(n5292), .B(n2625), .Z(c_out) );
  ND2D1BWP12T U3511 ( .A1(n2627), .A2(n2626), .ZN(n2629) );
  XNR2D2BWP12T U3512 ( .A1(n2629), .A2(n2628), .ZN(n3032) );
  CKND2D2BWP12T U3513 ( .A1(n3032), .A2(n5292), .ZN(n2676) );
  INVD1P75BWP12T U3514 ( .I(n2630), .ZN(n3421) );
  ND2D1BWP12T U3515 ( .A1(n3355), .A2(n5308), .ZN(n2674) );
  CKND0BWP12T U3516 ( .I(n2631), .ZN(n2633) );
  INVD1BWP12T U3517 ( .I(n2634), .ZN(n4543) );
  AOI22D1BWP12T U3518 ( .A1(n5305), .A2(n3212), .B1(n4535), .B2(n5297), .ZN(
        n2673) );
  INVD0BWP12T U3519 ( .I(n2946), .ZN(n2636) );
  ND2D1BWP12T U3520 ( .A1(n4208), .A2(n5281), .ZN(n5017) );
  OAI21D0BWP12T U3521 ( .A1(n71), .A2(n5255), .B(n5254), .ZN(n2639) );
  CKND0BWP12T U3522 ( .I(n3679), .ZN(n3909) );
  MUX2ND0BWP12T U3523 ( .I0(n2637), .I1(n5299), .S(n3909), .ZN(n2638) );
  RCAOI21D0BWP12T U3524 ( .A1(n2640), .A2(n2639), .B(n2638), .ZN(n2641) );
  OAI21D1BWP12T U3525 ( .A1(n4203), .A2(n5017), .B(n2641), .ZN(n2667) );
  OAI22D1BWP12T U3526 ( .A1(n3588), .A2(n4916), .B1(n3587), .B2(n7), .ZN(n2643) );
  OAI22D0BWP12T U3527 ( .A1(n3591), .A2(n3915), .B1(n3589), .B2(n4651), .ZN(
        n2642) );
  OAI22D0BWP12T U3528 ( .A1(n3588), .A2(n2895), .B1(n3587), .B2(n5148), .ZN(
        n2645) );
  OAI22D1BWP12T U3529 ( .A1(n3591), .A2(n407), .B1(n3589), .B2(n4607), .ZN(
        n2644) );
  TPNR2D1BWP12T U3530 ( .A1(n2645), .A2(n2644), .ZN(n2779) );
  MUX2XD2BWP12T U3531 ( .I0(n3575), .I1(n2779), .S(n5196), .Z(n3605) );
  NR2D1BWP12T U3532 ( .A1(n3605), .A2(n3948), .ZN(n3548) );
  NR2D0BWP12T U3533 ( .A1(n3594), .A2(n3524), .ZN(n2646) );
  NR2D1BWP12T U3534 ( .A1(n3548), .A2(n2646), .ZN(n4925) );
  OAI22D0BWP12T U3535 ( .A1(n3588), .A2(n3895), .B1(n3587), .B2(n3889), .ZN(
        n2648) );
  OAI22D0BWP12T U3536 ( .A1(n3591), .A2(n4790), .B1(n3589), .B2(n4578), .ZN(
        n2647) );
  NR2D1BWP12T U3537 ( .A1(n2648), .A2(n2647), .ZN(n3577) );
  OAI22D0BWP12T U3538 ( .A1(n3588), .A2(n2904), .B1(n3587), .B2(n4635), .ZN(
        n2650) );
  OAI22D1BWP12T U3539 ( .A1(n3887), .A2(n3591), .B1(n3589), .B2(n3888), .ZN(
        n2649) );
  TPNR2D1BWP12T U3540 ( .A1(n2650), .A2(n2649), .ZN(n3574) );
  MUX2XD2BWP12T U3541 ( .I0(n3577), .I1(n3574), .S(n5196), .Z(n3606) );
  AOI22D0BWP12T U3542 ( .A1(n3496), .A2(n4511), .B1(n3494), .B2(n3495), .ZN(
        n2652) );
  AOI22D0BWP12T U3543 ( .A1(n3498), .A2(n3679), .B1(n3497), .B2(n2848), .ZN(
        n2651) );
  CKND2D1BWP12T U3544 ( .A1(n2652), .A2(n2651), .ZN(n2679) );
  OAI22D0BWP12T U3545 ( .A1(n3588), .A2(n5081), .B1(n3587), .B2(n5260), .ZN(
        n2654) );
  OAI22D0BWP12T U3546 ( .A1(n3591), .A2(n3896), .B1(n3589), .B2(n5235), .ZN(
        n2653) );
  NR2D1BWP12T U3547 ( .A1(n2654), .A2(n2653), .ZN(n3576) );
  NR2D1BWP12T U3548 ( .A1(n3576), .A2(n3607), .ZN(n2655) );
  AOI211D1BWP12T U3549 ( .A1(n2679), .A2(n4601), .B(n2655), .C(n4301), .ZN(
        n2656) );
  OAI21D1BWP12T U3550 ( .A1(n3606), .A2(n3905), .B(n2656), .ZN(n4285) );
  CKND0BWP12T U3551 ( .I(n4049), .ZN(n2657) );
  TPNR2D0BWP12T U3552 ( .A1(n2657), .A2(n4051), .ZN(n2660) );
  CKND1BWP12T U3553 ( .I(n4048), .ZN(n2658) );
  TPOAI21D0BWP12T U3554 ( .A1(n2658), .A2(n4051), .B(n4422), .ZN(n2659) );
  AOI21D1BWP12T U3555 ( .A1(n4050), .A2(n2660), .B(n2659), .ZN(n2663) );
  CKND2D0BWP12T U3556 ( .A1(n2636), .A2(n2945), .ZN(n2662) );
  XOR2XD1BWP12T U3557 ( .A1(n2663), .A2(n2662), .Z(n4054) );
  CKND2D1BWP12T U3558 ( .A1(n4054), .A2(n5303), .ZN(n2665) );
  INR2XD2BWP12T U3559 ( .A1(n2664), .B1(n3844), .ZN(n5181) );
  INVD4BWP12T U3560 ( .I(n3844), .ZN(n5214) );
  CKND0BWP12T U3561 ( .I(n3605), .ZN(n2668) );
  NR2XD0BWP12T U3562 ( .A1(n2668), .A2(n3882), .ZN(n2669) );
  TPOAI21D0BWP12T U3563 ( .A1(n2669), .A2(n4260), .B(n3524), .ZN(n2670) );
  INVD4BWP12T U3564 ( .I(n3565), .ZN(n5323) );
  AOI31D1BWP12T U3565 ( .A1(n2670), .A2(n3875), .A3(n4285), .B(n5323), .ZN(
        n3586) );
  AN4D2BWP12T U3566 ( .A1(n2674), .A2(n2673), .A3(n2672), .A4(n2671), .Z(n2675) );
  ND2D4BWP12T U3567 ( .A1(n2676), .A2(n2675), .ZN(result[7]) );
  AOI22D1BWP12T U3568 ( .A1(n3854), .A2(n4133), .B1(n4132), .B2(n3855), .ZN(
        n3778) );
  NR2D1BWP12T U3569 ( .A1(n2976), .A2(n2677), .ZN(n2888) );
  AOI22D1BWP12T U3570 ( .A1(n4133), .A2(n2888), .B1(n2839), .B2(n4132), .ZN(
        n4202) );
  OAI21D1BWP12T U3571 ( .A1(n2772), .A2(n3905), .B(n2721), .ZN(n4710) );
  INVD1BWP12T U3572 ( .I(n2679), .ZN(n2680) );
  TPOAI21D0BWP12T U3573 ( .A1(n2680), .A2(n3607), .B(n3882), .ZN(n2685) );
  INVD1BWP12T U3574 ( .I(n3806), .ZN(n3569) );
  INR2XD0BWP12T U3575 ( .A1(n3661), .B1(n3594), .ZN(n2681) );
  AOI21D1BWP12T U3576 ( .A1(n3569), .A2(n4541), .B(n2681), .ZN(n2683) );
  INR2D1BWP12T U3577 ( .A1(b[0]), .B1(n3871), .ZN(n3595) );
  NR2D1BWP12T U3578 ( .A1(n3871), .A2(b[0]), .ZN(n3596) );
  AOI22D0BWP12T U3579 ( .A1(n4891), .A2(n3595), .B1(n3596), .B2(n5030), .ZN(
        n2682) );
  AOI21D1BWP12T U3580 ( .A1(n2683), .A2(n2682), .B(n3948), .ZN(n2684) );
  NR2D1BWP12T U3581 ( .A1(n2685), .A2(n2684), .ZN(n2689) );
  INVD1BWP12T U3582 ( .I(n3609), .ZN(n3703) );
  CKND0BWP12T U3583 ( .I(n3577), .ZN(n2687) );
  INVD1BWP12T U3584 ( .I(n3576), .ZN(n2686) );
  AOI22D1BWP12T U3585 ( .A1(n3703), .A2(n2687), .B1(n2686), .B2(n3707), .ZN(
        n2688) );
  ND2D1BWP12T U3586 ( .A1(n2689), .A2(n2688), .ZN(n2722) );
  INVD1BWP12T U3587 ( .I(n2722), .ZN(n2690) );
  AOI21D1BWP12T U3588 ( .A1(n4710), .A2(n4301), .B(n2690), .ZN(n3725) );
  ND2D1BWP12T U3589 ( .A1(n3875), .A2(n5212), .ZN(n5275) );
  ND2D1BWP12T U3590 ( .A1(n5275), .A2(n5312), .ZN(n5072) );
  TPND2D1BWP12T U3591 ( .A1(n3725), .A2(n5072), .ZN(n2727) );
  CKND2D1BWP12T U3592 ( .A1(n4426), .A2(n5313), .ZN(n2719) );
  INVD1BWP12T U3593 ( .I(n2692), .ZN(n3230) );
  OAI21D1BWP12T U3594 ( .A1(n3230), .A2(n3227), .B(n3228), .ZN(n2696) );
  CKND2D0BWP12T U3595 ( .A1(n2714), .A2(n2694), .ZN(n2695) );
  XNR2D1BWP12T U3596 ( .A1(n2696), .A2(n2695), .ZN(n3234) );
  TPND2D0BWP12T U3597 ( .A1(n3234), .A2(n5305), .ZN(n2712) );
  OAI21D0BWP12T U3598 ( .A1(n3661), .A2(n5255), .B(n5254), .ZN(n2700) );
  MUX2D1BWP12T U3599 ( .I0(n5295), .I1(n5294), .S(n3948), .Z(n2697) );
  CKND2D0BWP12T U3600 ( .A1(n2697), .A2(n5254), .ZN(n2698) );
  MUX2XD0BWP12T U3601 ( .I0(n5236), .I1(n2698), .S(n436), .Z(n2699) );
  AOI21D1BWP12T U3602 ( .A1(n3948), .A2(n2700), .B(n2699), .ZN(n2711) );
  CKND1BWP12T U3603 ( .I(n2701), .ZN(n4057) );
  OAI21D1BWP12T U3604 ( .A1(n4057), .A2(n4056), .B(n4429), .ZN(n2705) );
  CKND2D0BWP12T U3605 ( .A1(n2691), .A2(n2703), .ZN(n2704) );
  XNR2D1BWP12T U3606 ( .A1(n2705), .A2(n2704), .ZN(n4064) );
  CKND2D1BWP12T U3607 ( .A1(n4064), .A2(n5303), .ZN(n2710) );
  CKND1BWP12T U3608 ( .I(n2706), .ZN(n4536) );
  CKND0BWP12T U3609 ( .I(n5192), .ZN(n2707) );
  ND2D1BWP12T U3610 ( .A1(n4536), .A2(n2707), .ZN(n2708) );
  XOR2XD1BWP12T U3611 ( .A1(n2708), .A2(n3661), .Z(n4537) );
  CKND2D0BWP12T U3612 ( .A1(n4537), .A2(n5297), .ZN(n2709) );
  ND4D1BWP12T U3613 ( .A1(n2712), .A2(n2711), .A3(n2710), .A4(n2709), .ZN(
        n2718) );
  CKAN2D2BWP12T U3614 ( .A1(n2714), .A2(n2713), .Z(n2715) );
  XNR2XD2BWP12T U3615 ( .A1(n2716), .A2(n2715), .ZN(n3340) );
  AN2XD1BWP12T U3616 ( .A1(n3340), .A2(n5308), .Z(n2717) );
  AOI22D0BWP12T U3617 ( .A1(n2779), .A2(n3707), .B1(n3703), .B2(n3564), .ZN(
        n2720) );
  TPND2D1BWP12T U3618 ( .A1(n2721), .A2(n2720), .ZN(n4703) );
  TPOAI21D1BWP12T U3619 ( .A1(n4703), .A2(n3838), .B(n3844), .ZN(n2723) );
  AOI21D1BWP12T U3620 ( .A1(n2723), .A2(n2722), .B(n5323), .ZN(n3604) );
  NR2D1BWP12T U3621 ( .A1(n3604), .A2(n5271), .ZN(n2724) );
  ND2D2BWP12T U3622 ( .A1(n2727), .A2(n2726), .ZN(n2728) );
  INR2D4BWP12T U3623 ( .A1(n461), .B1(n2728), .ZN(n2734) );
  IND2D2BWP12T U3624 ( .A1(n2730), .B1(n2729), .ZN(n2732) );
  XNR2XD4BWP12T U3625 ( .A1(n2732), .A2(n2731), .ZN(n3021) );
  CKND2D8BWP12T U3626 ( .A1(n2734), .A2(n2733), .ZN(result[3]) );
  TPND2D1BWP12T U3627 ( .A1(n3104), .A2(n2735), .ZN(n3094) );
  INVD2BWP12T U3628 ( .I(n2736), .ZN(n3093) );
  TPND2D2BWP12T U3629 ( .A1(n3094), .A2(n3093), .ZN(n3157) );
  INVD2BWP12T U3630 ( .I(n442), .ZN(n3095) );
  ND2D1BWP12T U3631 ( .A1(n3095), .A2(n3150), .ZN(n2738) );
  OAI21D1BWP12T U3632 ( .A1(n3298), .A2(n3282), .B(n3285), .ZN(n2740) );
  CKND2D1BWP12T U3633 ( .A1(n3453), .A2(n2744), .ZN(n2739) );
  XNR2D1BWP12T U3634 ( .A1(n2740), .A2(n2739), .ZN(n3291) );
  INVD3BWP12T U3635 ( .I(n2741), .ZN(n3483) );
  INVD1BWP12T U3636 ( .I(n3433), .ZN(n3470) );
  NR2D0BWP12T U3637 ( .A1(n3470), .A2(n3450), .ZN(n2743) );
  INVD1BWP12T U3638 ( .I(n3415), .ZN(n3480) );
  TPOAI21D0BWP12T U3639 ( .A1(n3480), .A2(n3450), .B(n3451), .ZN(n2742) );
  TPAOI21D0BWP12T U3640 ( .A1(n3483), .A2(n2743), .B(n2742), .ZN(n2746) );
  ND2D1BWP12T U3641 ( .A1(n3453), .A2(n2744), .ZN(n2745) );
  XOR2XD1BWP12T U3642 ( .A1(n2746), .A2(n2745), .Z(n3446) );
  TPND2D0BWP12T U3643 ( .A1(n3985), .A2(n3983), .ZN(n2749) );
  AOI21D1BWP12T U3644 ( .A1(n3988), .A2(n3983), .B(n2747), .ZN(n2748) );
  OAI21D1BWP12T U3645 ( .A1(n4116), .A2(n2749), .B(n2748), .ZN(n2752) );
  ND2D1BWP12T U3646 ( .A1(n4461), .A2(n2750), .ZN(n2751) );
  XNR2D1BWP12T U3647 ( .A1(n2752), .A2(n2751), .ZN(n3984) );
  INR2D1BWP12T U3648 ( .A1(n3984), .B1(n4970), .ZN(n2797) );
  INVD1BWP12T U3649 ( .I(n4365), .ZN(n4478) );
  NR2D0BWP12T U3650 ( .A1(n4478), .A2(n4458), .ZN(n2755) );
  INVD1BWP12T U3651 ( .I(n4364), .ZN(n4488) );
  TPOAI21D0BWP12T U3652 ( .A1(n4488), .A2(n4458), .B(n4459), .ZN(n2754) );
  TPAOI21D0BWP12T U3653 ( .A1(n4491), .A2(n2755), .B(n2754), .ZN(n2758) );
  CKND2D1BWP12T U3654 ( .A1(n4461), .A2(n2756), .ZN(n2757) );
  XOR2XD1BWP12T U3655 ( .A1(n2758), .A2(n2757), .Z(n4468) );
  INVD1BWP12T U3656 ( .I(n4468), .ZN(n2795) );
  CKND0BWP12T U3657 ( .I(n4570), .ZN(n2759) );
  TPND2D0BWP12T U3658 ( .A1(n2759), .A2(n7), .ZN(n2760) );
  TPNR2D0BWP12T U3659 ( .A1(n4571), .A2(n2760), .ZN(n2761) );
  TPND2D0BWP12T U3660 ( .A1(n2761), .A2(n4582), .ZN(n2762) );
  XOR2XD1BWP12T U3661 ( .A1(n2762), .A2(n2773), .Z(n4563) );
  OAI22D0BWP12T U3662 ( .A1(n2889), .A2(n3871), .B1(n4152), .B2(n3872), .ZN(
        n2764) );
  OAI22D0BWP12T U3663 ( .A1(n4134), .A2(n3869), .B1(n2890), .B2(n3870), .ZN(
        n2763) );
  NR2D1BWP12T U3664 ( .A1(n2764), .A2(n2763), .ZN(n3749) );
  INVD0BWP12T U3665 ( .I(n3778), .ZN(n3748) );
  MUX2ND0BWP12T U3666 ( .I0(n3749), .I1(n3748), .S(n3948), .ZN(n5087) );
  CKND0BWP12T U3667 ( .I(n5087), .ZN(n2771) );
  INVD1BWP12T U3668 ( .I(n3861), .ZN(n3880) );
  AOI22D0BWP12T U3669 ( .A1(n3855), .A2(n4163), .B1(n3757), .B2(n3854), .ZN(
        n2766) );
  AOI22D0BWP12T U3670 ( .A1(n3853), .A2(n4151), .B1(n4150), .B2(n3852), .ZN(
        n2765) );
  CKND2D1BWP12T U3671 ( .A1(n2766), .A2(n2765), .ZN(n3750) );
  AOI22D0BWP12T U3672 ( .A1(n3855), .A2(n3793), .B1(n4165), .B2(n3854), .ZN(
        n2768) );
  AOI22D0BWP12T U3673 ( .A1(n3853), .A2(n4166), .B1(n4164), .B2(n3852), .ZN(
        n2767) );
  AOI21D0BWP12T U3674 ( .A1(n2768), .A2(n2767), .B(n4953), .ZN(n2769) );
  AOI211D0BWP12T U3675 ( .A1(n3880), .A2(n3750), .B(n2769), .C(n3838), .ZN(
        n2770) );
  TPOAI21D0BWP12T U3676 ( .A1(n2771), .A2(n3882), .B(n2770), .ZN(n3884) );
  NR2XD0BWP12T U3677 ( .A1(n3884), .A2(n5232), .ZN(n2784) );
  CKND2D1BWP12T U3678 ( .A1(n2772), .A2(n3905), .ZN(n3724) );
  OAI21D1BWP12T U3679 ( .A1(n2773), .A2(n5255), .B(n5254), .ZN(n2777) );
  MUX2D0BWP12T U3680 ( .I0(n5295), .I1(n5294), .S(n21), .Z(n2774) );
  CKND2D0BWP12T U3681 ( .A1(n2774), .A2(n5254), .ZN(n2775) );
  MUX2D1BWP12T U3682 ( .I0(n5236), .I1(n2775), .S(n4503), .Z(n2776) );
  RCAOI21D0BWP12T U3683 ( .A1(n21), .A2(n2777), .B(n2776), .ZN(n2781) );
  NR2D1BWP12T U3684 ( .A1(n3882), .A2(n5108), .ZN(n2778) );
  TPNR2D1BWP12T U3685 ( .A1(n3838), .A2(n2778), .ZN(n4633) );
  INVD1P75BWP12T U3686 ( .I(n3607), .ZN(n3617) );
  INVD1BWP12T U3687 ( .I(n3524), .ZN(n3625) );
  CKND2D0BWP12T U3688 ( .A1(n4633), .A2(n3578), .ZN(n3581) );
  NR2D0BWP12T U3689 ( .A1(n3581), .A2(n5271), .ZN(n2780) );
  ND2D2BWP12T U3690 ( .A1(n3844), .A2(n5108), .ZN(n3580) );
  INR2D2BWP12T U3691 ( .A1(n5322), .B1(n3580), .ZN(n5151) );
  INR3D0BWP12T U3692 ( .A1(n2781), .B1(n2780), .B2(n5151), .ZN(n2782) );
  TPOAI21D0BWP12T U3693 ( .A1(n4924), .A2(n3724), .B(n2782), .ZN(n2783) );
  AOI211XD0BWP12T U3694 ( .A1(n4563), .A2(n5297), .B(n2784), .C(n2783), .ZN(
        n2794) );
  MUX2D1BWP12T U3695 ( .I0(n4202), .I1(n4189), .S(n4277), .Z(n5071) );
  INVD1BWP12T U3696 ( .I(n4163), .ZN(n4130) );
  TPNR2D0BWP12T U3697 ( .A1(n4309), .A2(n4130), .ZN(n2787) );
  TPNR2D0BWP12T U3698 ( .A1(n4311), .A2(n4131), .ZN(n2786) );
  INVD1BWP12T U3699 ( .I(n3757), .ZN(n4153) );
  OAI22D1BWP12T U3700 ( .A1(n4315), .A2(n4140), .B1(n4313), .B2(n4153), .ZN(
        n2785) );
  NR3D1BWP12T U3701 ( .A1(n2787), .A2(n2786), .A3(n2785), .ZN(n4187) );
  INVD0BWP12T U3702 ( .I(n4166), .ZN(n4129) );
  TPOAI22D0BWP12T U3703 ( .A1(n4315), .A2(n4129), .B1(n4313), .B2(n4241), .ZN(
        n2790) );
  INVD0BWP12T U3704 ( .I(n4164), .ZN(n4243) );
  TPNR2D0BWP12T U3705 ( .A1(n4311), .A2(n4243), .ZN(n2789) );
  TPNR2D0BWP12T U3706 ( .A1(n4309), .A2(n4246), .ZN(n2788) );
  TPOAI31D0BWP12T U3707 ( .A1(n2790), .A2(n2789), .A3(n2788), .B(n4208), .ZN(
        n2791) );
  OAI211D1BWP12T U3708 ( .A1(n4187), .A2(n4815), .B(n2791), .C(n4185), .ZN(
        n2792) );
  AOI21D1BWP12T U3709 ( .A1(n5071), .A2(n4299), .B(n2792), .ZN(n4186) );
  CKND2D1BWP12T U3710 ( .A1(n4186), .A2(n5281), .ZN(n2793) );
  OAI211D1BWP12T U3711 ( .A1(n4965), .A2(n2795), .B(n2794), .C(n2793), .ZN(
        n2796) );
  AOI211XD1BWP12T U3712 ( .A1(n3446), .A2(n5308), .B(n2797), .C(n2796), .ZN(
        n2798) );
  IOA21D2BWP12T U3713 ( .A1(n3291), .A2(n5305), .B(n2798), .ZN(n2799) );
  INR2D1BWP12T U3714 ( .A1(n2801), .B1(n2800), .ZN(n2806) );
  INVD1BWP12T U3715 ( .I(n2802), .ZN(n2803) );
  TPNR2D1BWP12T U3716 ( .A1(n2804), .A2(n2803), .ZN(n2805) );
  XNR2D2BWP12T U3717 ( .A1(n2806), .A2(n2805), .ZN(n3042) );
  INVD3BWP12T U3718 ( .I(n2807), .ZN(n3314) );
  CKND2D0BWP12T U3719 ( .A1(n2878), .A2(n2962), .ZN(n2810) );
  CKND0BWP12T U3720 ( .I(n2961), .ZN(n2808) );
  TPAOI21D0BWP12T U3721 ( .A1(n2878), .A2(n2808), .B(n2815), .ZN(n2809) );
  OAI21D1BWP12T U3722 ( .A1(n3314), .A2(n2810), .B(n2809), .ZN(n2813) );
  CKND2D1BWP12T U3723 ( .A1(n2811), .A2(n2819), .ZN(n2812) );
  XNR2D1BWP12T U3724 ( .A1(n2813), .A2(n2812), .ZN(n3253) );
  CKND2D0BWP12T U3725 ( .A1(n2881), .A2(n2878), .ZN(n2817) );
  INVD0BWP12T U3726 ( .I(n2885), .ZN(n2815) );
  TPAOI21D0BWP12T U3727 ( .A1(n2882), .A2(n2878), .B(n2815), .ZN(n2816) );
  OAI21D1BWP12T U3728 ( .A1(n3421), .A2(n2817), .B(n2816), .ZN(n2821) );
  TPND2D0BWP12T U3729 ( .A1(n2811), .A2(n2819), .ZN(n2820) );
  XNR2XD1BWP12T U3730 ( .A1(n2821), .A2(n2820), .ZN(n3425) );
  INVD1P75BWP12T U3731 ( .I(n2822), .ZN(n4577) );
  CKND0BWP12T U3732 ( .I(n4519), .ZN(n2823) );
  CKND2D1BWP12T U3733 ( .A1(n4577), .A2(n2823), .ZN(n2824) );
  INVD1BWP12T U3734 ( .I(n3897), .ZN(n4518) );
  XOR2D1BWP12T U3735 ( .A1(n2824), .A2(n4518), .Z(n4523) );
  INVD1BWP12T U3736 ( .I(n4523), .ZN(n2837) );
  ND2D1BWP12T U3737 ( .A1(n3496), .A2(n4649), .ZN(n3510) );
  AOI22D1BWP12T U3738 ( .A1(n3494), .A2(n4914), .B1(n3497), .B2(n4568), .ZN(
        n3512) );
  CKND2D1BWP12T U3739 ( .A1(n3510), .A2(n3512), .ZN(n3491) );
  ND2D1BWP12T U3740 ( .A1(n3511), .A2(n5196), .ZN(n2826) );
  NR2D1BWP12T U3741 ( .A1(n3491), .A2(n2826), .ZN(n2828) );
  OAI22D1BWP12T U3742 ( .A1(n3591), .A2(n3888), .B1(n3589), .B2(n2904), .ZN(
        n3517) );
  INR3D0BWP12T U3743 ( .A1(n3539), .B1(n3517), .B2(n3518), .ZN(n2827) );
  NR2D1BWP12T U3744 ( .A1(n2828), .A2(n2827), .ZN(n4261) );
  AOI21D0BWP12T U3745 ( .A1(n3515), .A2(n4601), .B(n4301), .ZN(n2829) );
  OAI21D0BWP12T U3746 ( .A1(n3513), .A2(n3607), .B(n2829), .ZN(n2830) );
  AOI21D1BWP12T U3747 ( .A1(n3948), .A2(n4261), .B(n2830), .ZN(n4270) );
  AOI22D1BWP12T U3748 ( .A1(n3498), .A2(n5146), .B1(n3494), .B2(n5108), .ZN(
        n3727) );
  INVD1BWP12T U3749 ( .I(n2831), .ZN(n2833) );
  OAI22D1BWP12T U3750 ( .A1(n3591), .A2(n4609), .B1(n3587), .B2(n4990), .ZN(
        n2832) );
  TPAOI21D2BWP12T U3751 ( .A1(n2834), .A2(n2833), .B(n2832), .ZN(n3527) );
  INVD1BWP12T U3752 ( .I(n3527), .ZN(n2856) );
  MUX2XD2BWP12T U3753 ( .I0(n3727), .I1(n2856), .S(n2835), .Z(n4954) );
  INR2D2BWP12T U3754 ( .A1(n3905), .B1(n4954), .ZN(n4945) );
  AOI21D0BWP12T U3755 ( .A1(n4945), .A2(n5281), .B(n5321), .ZN(n2836) );
  OAI22D0BWP12T U3756 ( .A1(n2837), .A2(n5104), .B1(n4270), .B2(n2836), .ZN(
        n2854) );
  INR2D1BWP12T U3757 ( .A1(n5281), .B1(n4299), .ZN(n5074) );
  MUX2ND0BWP12T U3758 ( .I0(n4891), .I1(n5030), .S(b[0]), .ZN(n4216) );
  MUX2ND0BWP12T U3759 ( .I0(n3495), .I1(n4510), .S(b[0]), .ZN(n4228) );
  MUX2XD0BWP12T U3760 ( .I0(n3897), .I1(n2910), .S(b[0]), .Z(n4226) );
  CKND2D1BWP12T U3761 ( .A1(n4296), .A2(n4277), .ZN(n2841) );
  INR2D1BWP12T U3762 ( .A1(n480), .B1(n3591), .ZN(n3779) );
  INVD1BWP12T U3763 ( .I(n3779), .ZN(n4200) );
  NR2D1BWP12T U3764 ( .A1(n2976), .A2(n4200), .ZN(n2838) );
  TPOAI21D1BWP12T U3765 ( .A1(n2839), .A2(n2838), .B(n2845), .ZN(n5182) );
  INVD1P75BWP12T U3766 ( .I(n4277), .ZN(n4274) );
  CKND2D1BWP12T U3767 ( .A1(n5182), .A2(n4274), .ZN(n2840) );
  ND2D1BWP12T U3768 ( .A1(n2841), .A2(n2840), .ZN(n4195) );
  INR2D1BWP12T U3769 ( .A1(n5074), .B1(n4195), .ZN(n2853) );
  INVD1BWP12T U3770 ( .I(n4945), .ZN(n2842) );
  INR2D1BWP12T U3771 ( .A1(n3875), .B1(n2842), .ZN(n2844) );
  INVD1BWP12T U3772 ( .I(n4270), .ZN(n2843) );
  OAI21D1BWP12T U3773 ( .A1(n2844), .A2(n5214), .B(n2843), .ZN(n3714) );
  NR2D1BWP12T U3774 ( .A1(n3714), .A2(n5327), .ZN(n2852) );
  AOI22D1BWP12T U3775 ( .A1(n3854), .A2(n4228), .B1(n4226), .B2(n3855), .ZN(
        n2847) );
  AOI22D1BWP12T U3776 ( .A1(n3852), .A2(n4216), .B1(n4199), .B2(n3853), .ZN(
        n2846) );
  ND2D1BWP12T U3777 ( .A1(n2847), .A2(n2846), .ZN(n3837) );
  MUX2D1BWP12T U3778 ( .I0(n3821), .I1(n3837), .S(n3905), .Z(n3867) );
  ND2D1BWP12T U3779 ( .A1(n5214), .A2(n5252), .ZN(n5317) );
  OAI21D1BWP12T U3780 ( .A1(n3867), .A2(n5317), .B(n2850), .ZN(n2851) );
  NR4D0BWP12T U3781 ( .A1(n2854), .A2(n2853), .A3(n2852), .A4(n2851), .ZN(
        n2855) );
  IOA21D1BWP12T U3782 ( .A1(n3425), .A2(n5308), .B(n2855), .ZN(n2868) );
  INVD1BWP12T U3783 ( .I(n3509), .ZN(n3492) );
  MUX2XD0BWP12T U3784 ( .I0(n3492), .I1(n2856), .S(n3539), .Z(n2857) );
  OAI21D1BWP12T U3785 ( .A1(n2857), .A2(n3948), .B(n3524), .ZN(n4942) );
  AOI21D0BWP12T U3786 ( .A1(n4942), .A2(n3875), .B(n5214), .ZN(n2858) );
  TPOAI21D0BWP12T U3787 ( .A1(n2858), .A2(n4270), .B(n3565), .ZN(n3545) );
  INVD2BWP12T U3788 ( .I(n2859), .ZN(n2932) );
  CKND2D0BWP12T U3789 ( .A1(n2923), .A2(n2932), .ZN(n2862) );
  INVD0BWP12T U3790 ( .I(n2927), .ZN(n2860) );
  TPAOI21D0BWP12T U3791 ( .A1(n2924), .A2(n2932), .B(n2860), .ZN(n2861) );
  OAI21D1BWP12T U3792 ( .A1(n4408), .A2(n2862), .B(n2861), .ZN(n2864) );
  INVD1BWP12T U3793 ( .I(n2863), .ZN(n4087) );
  ND2D1BWP12T U3794 ( .A1(n4087), .A2(n4085), .ZN(n2866) );
  XNR2XD1BWP12T U3795 ( .A1(n2864), .A2(n2866), .ZN(n4391) );
  INVD1P75BWP12T U3796 ( .I(n2865), .ZN(n4096) );
  AOI22D1BWP12T U3797 ( .A1(n5313), .A2(n4391), .B1(n4098), .B2(n5303), .ZN(
        n2867) );
  INVD1BWP12T U3798 ( .I(n2869), .ZN(n2942) );
  INVD1BWP12T U3799 ( .I(n2941), .ZN(n2870) );
  INVD1BWP12T U3800 ( .I(n2871), .ZN(n2873) );
  ND2D1BWP12T U3801 ( .A1(n2873), .A2(n2872), .ZN(n2874) );
  INVD1BWP12T U3802 ( .I(n3036), .ZN(n2940) );
  OAI21D1BWP12T U3803 ( .A1(n3314), .A2(n2876), .B(n2961), .ZN(n2880) );
  ND2D1BWP12T U3804 ( .A1(n2878), .A2(n2877), .ZN(n2879) );
  XNR2D1BWP12T U3805 ( .A1(n2880), .A2(n2879), .ZN(n3235) );
  CKND0BWP12T U3806 ( .I(n2881), .ZN(n2884) );
  INVD1BWP12T U3807 ( .I(n2882), .ZN(n2883) );
  OAI21D1BWP12T U3808 ( .A1(n3421), .A2(n2884), .B(n2883), .ZN(n2887) );
  CKND2D1BWP12T U3809 ( .A1(n2878), .A2(n2885), .ZN(n2886) );
  XNR2XD1BWP12T U3810 ( .A1(n2887), .A2(n2886), .ZN(n3426) );
  CKND1BWP12T U3811 ( .I(n2888), .ZN(n2973) );
  OAI22D1BWP12T U3812 ( .A1(n2890), .A2(n2973), .B1(n4309), .B2(n2889), .ZN(
        n2892) );
  OAI22D0BWP12T U3813 ( .A1(n4311), .A2(n4134), .B1(n4132), .B2(n4315), .ZN(
        n2891) );
  NR2D1BWP12T U3814 ( .A1(n2892), .A2(n2891), .ZN(n4158) );
  INVD1BWP12T U3815 ( .I(n4158), .ZN(n2894) );
  TPNR2D1BWP12T U3816 ( .A1(n4309), .A2(n3760), .ZN(n4207) );
  CKND2D1BWP12T U3817 ( .A1(n4274), .A2(n4207), .ZN(n2893) );
  TPOAI21D1BWP12T U3818 ( .A1(n2894), .A2(n4274), .B(n2893), .ZN(n4174) );
  AOI22D1BWP12T U3819 ( .A1(n3498), .A2(n4990), .B1(n3494), .B2(n5146), .ZN(
        n3537) );
  NR2D0BWP12T U3820 ( .A1(n3588), .A2(n3915), .ZN(n2897) );
  NR2D1BWP12T U3821 ( .A1(n3589), .A2(n7), .ZN(n2896) );
  NR3D1BWP12T U3822 ( .A1(n2898), .A2(n2897), .A3(n2896), .ZN(n4176) );
  INVD1BWP12T U3823 ( .I(n4176), .ZN(n3615) );
  AOI22D1BWP12T U3824 ( .A1(n3617), .A2(n4995), .B1(n3615), .B2(n4601), .ZN(
        n4978) );
  OAI22D0BWP12T U3825 ( .A1(n3588), .A2(n445), .B1(n3587), .B2(n4651), .ZN(
        n2901) );
  OAI22D0BWP12T U3826 ( .A1(n3591), .A2(n4916), .B1(n3589), .B2(n4635), .ZN(
        n2900) );
  NR2D1BWP12T U3827 ( .A1(n2901), .A2(n2900), .ZN(n3619) );
  OAI22D0BWP12T U3828 ( .A1(n3588), .A2(n3896), .B1(n3587), .B2(n4578), .ZN(
        n2903) );
  OAI22D0BWP12T U3829 ( .A1(n3591), .A2(n3895), .B1(n3589), .B2(n5260), .ZN(
        n2902) );
  OAI22D0BWP12T U3830 ( .A1(n3588), .A2(n4790), .B1(n3589), .B2(n3889), .ZN(
        n2906) );
  OAI22D0BWP12T U3831 ( .A1(n3591), .A2(n2904), .B1(n3587), .B2(n3888), .ZN(
        n2905) );
  TPNR2D1BWP12T U3832 ( .A1(n2906), .A2(n2905), .ZN(n3614) );
  OAI22D0BWP12T U3833 ( .A1(n3588), .A2(n2910), .B1(n3587), .B2(n5235), .ZN(
        n2908) );
  OAI22D1BWP12T U3834 ( .A1(n3591), .A2(n5081), .B1(n3589), .B2(n3897), .ZN(
        n2907) );
  NR2D1BWP12T U3835 ( .A1(n2908), .A2(n2907), .ZN(n3608) );
  TPNR2D1BWP12T U3836 ( .A1(n4323), .A2(n5312), .ZN(n2918) );
  ND2D1BWP12T U3837 ( .A1(n4133), .A2(n3855), .ZN(n3777) );
  MUX2D1BWP12T U3838 ( .I0(n3777), .I1(n3768), .S(n3905), .Z(n3775) );
  OAI21D1BWP12T U3839 ( .A1(n3775), .A2(n5317), .B(n2911), .ZN(n2916) );
  CKND2D1BWP12T U3840 ( .A1(n4524), .A2(n5297), .ZN(n2915) );
  CKND0BWP12T U3841 ( .I(n2920), .ZN(n2913) );
  OAI21D0BWP12T U3842 ( .A1(n4978), .A2(n3838), .B(n3844), .ZN(n2912) );
  ND2D1BWP12T U3843 ( .A1(n2913), .A2(n2912), .ZN(n3718) );
  OR2XD1BWP12T U3844 ( .A1(n3718), .A2(n5327), .Z(n2914) );
  IND3D1BWP12T U3845 ( .A1(n2916), .B1(n2915), .B2(n2914), .ZN(n2917) );
  TPNR2D1BWP12T U3846 ( .A1(n2918), .A2(n2917), .ZN(n2919) );
  IOA21D1BWP12T U3847 ( .A1(n3426), .A2(n5308), .B(n2919), .ZN(n2938) );
  NR2D1BWP12T U3848 ( .A1(n3838), .A2(n4260), .ZN(n3817) );
  OAI21D0BWP12T U3849 ( .A1(n3547), .A2(n3882), .B(n3817), .ZN(n2921) );
  TPAOI21D0BWP12T U3850 ( .A1(n2921), .A2(n3524), .B(n2920), .ZN(n2922) );
  INR2D1BWP12T U3851 ( .A1(n3565), .B1(n2922), .ZN(n3551) );
  INVD1BWP12T U3852 ( .I(n3551), .ZN(n2936) );
  INVD0BWP12T U3853 ( .I(n2923), .ZN(n2926) );
  INVD1BWP12T U3854 ( .I(n2924), .ZN(n2925) );
  OAI21D1BWP12T U3855 ( .A1(n4408), .A2(n2926), .B(n2925), .ZN(n2929) );
  CKND2D1BWP12T U3856 ( .A1(n2932), .A2(n2927), .ZN(n2928) );
  XNR2XD1BWP12T U3857 ( .A1(n2929), .A2(n2928), .ZN(n4392) );
  OAI21D1BWP12T U3858 ( .A1(n4096), .A2(n2930), .B(n2948), .ZN(n2934) );
  ND2D1BWP12T U3859 ( .A1(n2932), .A2(n2931), .ZN(n2933) );
  XNR2XD1BWP12T U3860 ( .A1(n2934), .A2(n2933), .ZN(n4099) );
  AOI22D1BWP12T U3861 ( .A1(n5313), .A2(n4392), .B1(n4099), .B2(n5303), .ZN(
        n2935) );
  IOA21D1BWP12T U3862 ( .A1(n5322), .A2(n2936), .B(n2935), .ZN(n2937) );
  TPOAI21D1BWP12T U3863 ( .A1(n2940), .A2(n5112), .B(n2939), .ZN(result[9]) );
  ND2D1BWP12T U3864 ( .A1(n2942), .A2(n2941), .ZN(n2944) );
  TPOAI21D0BWP12T U3865 ( .A1(n4408), .A2(n2946), .B(n2945), .ZN(n2949) );
  XNR2XD1BWP12T U3866 ( .A1(n2949), .A2(n2953), .ZN(n4451) );
  AOI22D1BWP12T U3867 ( .A1(n3617), .A2(n4602), .B1(n3536), .B2(n4601), .ZN(
        n3583) );
  INVD1BWP12T U3868 ( .I(n3583), .ZN(n4660) );
  OAI22D1BWP12T U3869 ( .A1(n3568), .A2(n3730), .B1(n3535), .B2(n3609), .ZN(
        n2952) );
  INVD1BWP12T U3870 ( .I(n3559), .ZN(n3573) );
  TPOAI21D0BWP12T U3871 ( .A1(n3573), .A2(n3607), .B(n3882), .ZN(n2951) );
  TPNR2D0BWP12T U3872 ( .A1(n3558), .A2(n3618), .ZN(n2950) );
  NR3D1BWP12T U3873 ( .A1(n2952), .A2(n2951), .A3(n2950), .ZN(n2981) );
  XOR2XD1BWP12T U3874 ( .A1(n4096), .A2(n2953), .Z(n4063) );
  CKND2D1BWP12T U3875 ( .A1(n4063), .A2(n5303), .ZN(n2954) );
  IOA21D1BWP12T U3876 ( .A1(n5212), .A2(n3713), .B(n2954), .ZN(n2957) );
  TPOAI21D0BWP12T U3877 ( .A1(n2981), .A2(n3524), .B(n3565), .ZN(n2955) );
  NR2D1BWP12T U3878 ( .A1(n3713), .A2(n2955), .ZN(n3629) );
  NR2D1BWP12T U3879 ( .A1(n3629), .A2(n5271), .ZN(n2956) );
  AOI211D1BWP12T U3880 ( .A1(n4451), .A2(n5313), .B(n2957), .C(n2956), .ZN(
        n2987) );
  CKND2D1BWP12T U3881 ( .A1(n3427), .A2(n5308), .ZN(n2972) );
  ND2XD0BWP12T U3882 ( .A1(n2962), .A2(n2961), .ZN(n2963) );
  XOR2XD1BWP12T U3883 ( .A1(n3314), .A2(n2963), .Z(n3214) );
  CKND2D1BWP12T U3884 ( .A1(n3214), .A2(n5305), .ZN(n2970) );
  ND2D1BWP12T U3885 ( .A1(n2964), .A2(n3539), .ZN(n4816) );
  INVD1BWP12T U3886 ( .I(n4816), .ZN(n4144) );
  INVD1BWP12T U3887 ( .I(n4216), .ZN(n3780) );
  INVD1BWP12T U3888 ( .I(n4228), .ZN(n4215) );
  OAI21D0BWP12T U3889 ( .A1(n3495), .A2(n5255), .B(n5254), .ZN(n2967) );
  MUX2D0BWP12T U3890 ( .I0(n5236), .I1(n2965), .S(n3495), .Z(n2966) );
  RCAOI21D0BWP12T U3891 ( .A1(n3937), .A2(n2967), .B(n2966), .ZN(n2968) );
  OAI21D1BWP12T U3892 ( .A1(n3842), .A2(n5232), .B(n2968), .ZN(n2969) );
  INR2D1BWP12T U3893 ( .A1(n2970), .B1(n2969), .ZN(n2971) );
  ND2D1BWP12T U3894 ( .A1(n2972), .A2(n2971), .ZN(n2986) );
  XNR2D1BWP12T U3895 ( .A1(n4577), .A2(n4509), .ZN(n4540) );
  INVD1BWP12T U3896 ( .I(n4540), .ZN(n2984) );
  OAI22D1BWP12T U3897 ( .A1(n2973), .A2(n4216), .B1(n4311), .B2(n4199), .ZN(
        n2979) );
  ND3D0BWP12T U3898 ( .A1(n2976), .A2(n2975), .A3(n2974), .ZN(n2977) );
  OAI21D0BWP12T U3899 ( .A1(n4309), .A2(n4228), .B(n2977), .ZN(n2978) );
  NR2D1BWP12T U3900 ( .A1(n2979), .A2(n2978), .ZN(n4814) );
  OAI22D1BWP12T U3901 ( .A1(n4814), .A2(n5183), .B1(n4816), .B2(n4815), .ZN(
        n2983) );
  NR2XD0BWP12T U3902 ( .A1(n4660), .A2(n3882), .ZN(n2980) );
  NR2D1BWP12T U3903 ( .A1(n2981), .A2(n2980), .ZN(n2982) );
  NR2D1BWP12T U3904 ( .A1(n2983), .A2(n2982), .ZN(n4159) );
  OAI22D1BWP12T U3905 ( .A1(n2984), .A2(n5104), .B1(n4159), .B2(n5312), .ZN(
        n2985) );
  INR3D2BWP12T U3906 ( .A1(n2987), .B1(n2986), .B2(n2985), .ZN(n2988) );
  TPND2D3BWP12T U3907 ( .A1(n2989), .A2(n2988), .ZN(result[8]) );
  INVD2BWP12T U3908 ( .I(n2990), .ZN(n3116) );
  INVD2BWP12T U3909 ( .I(n2991), .ZN(n3108) );
  ND2D1BWP12T U3910 ( .A1(n3108), .A2(n3106), .ZN(n2992) );
  XNR2XD4BWP12T U3911 ( .A1(n3116), .A2(n2992), .ZN(n4668) );
  INVD1BWP12T U3912 ( .I(n2993), .ZN(n3004) );
  OA21D2BWP12T U3913 ( .A1(n3006), .A2(n2994), .B(n3004), .Z(n3000) );
  AN2XD2BWP12T U3914 ( .A1(n2997), .A2(n2998), .Z(n2999) );
  XNR2XD4BWP12T U3915 ( .A1(n3000), .A2(n2999), .ZN(n4785) );
  INVD1P75BWP12T U3916 ( .I(n3001), .ZN(n3083) );
  NR2XD0BWP12T U3917 ( .A1(n3083), .A2(n3002), .ZN(n3003) );
  ND2D1BWP12T U3918 ( .A1(n3005), .A2(n3004), .ZN(n3007) );
  XOR2D1BWP12T U3919 ( .A1(n3007), .A2(n3006), .Z(n4811) );
  NR3D0BWP12T U3920 ( .A1(n4785), .A2(n4725), .A3(n4811), .ZN(n3072) );
  INVD2BWP12T U3921 ( .I(n3008), .ZN(n3010) );
  ND2D1BWP12T U3922 ( .A1(n3010), .A2(n3009), .ZN(n3012) );
  XOR2D2BWP12T U3923 ( .A1(n3012), .A2(n53), .Z(n4876) );
  INR2D1BWP12T U3924 ( .A1(n3016), .B1(n3015), .ZN(n5293) );
  OR3D0BWP12T U3925 ( .A1(n5293), .A2(n5112), .A3(n4859), .Z(n3020) );
  INVD1BWP12T U3926 ( .I(n3022), .ZN(n3030) );
  INVD2BWP12T U3927 ( .I(n3024), .ZN(n3026) );
  OAI21D1BWP12T U3928 ( .A1(n3026), .A2(n3027), .B(n3025), .ZN(n3028) );
  XNR2D2BWP12T U3929 ( .A1(n3029), .A2(n3028), .ZN(n5039) );
  OR3XD4BWP12T U3930 ( .A1(n3031), .A2(n3030), .A3(n5039), .Z(n3033) );
  OR3XD4BWP12T U3931 ( .A1(n4876), .A2(n3033), .A3(n3032), .Z(n3035) );
  TPAOI21D1BWP12T U3932 ( .A1(n3058), .A2(n3056), .B(n3057), .ZN(n3040) );
  ND2D1BWP12T U3933 ( .A1(n3038), .A2(n3037), .ZN(n3039) );
  TPOAI21D2BWP12T U3934 ( .A1(n3045), .A2(n3044), .B(n458), .ZN(n3063) );
  INVD1BWP12T U3935 ( .I(n3046), .ZN(n3047) );
  AOI21D0BWP12T U3936 ( .A1(n3061), .A2(n3064), .B(n3065), .ZN(n3048) );
  TPND2D1BWP12T U3937 ( .A1(n3049), .A2(n3048), .ZN(n3054) );
  INVD1BWP12T U3938 ( .I(n3050), .ZN(n3052) );
  ND2D1BWP12T U3939 ( .A1(n3052), .A2(n3051), .ZN(n3053) );
  XNR2XD4BWP12T U3940 ( .A1(n3054), .A2(n3053), .ZN(n4755) );
  IND2D2BWP12T U3941 ( .A1(n3057), .B1(n3056), .ZN(n3059) );
  XNR2D2BWP12T U3942 ( .A1(n3059), .A2(n3058), .ZN(n5099) );
  CKND0BWP12T U3943 ( .I(n5099), .ZN(n3060) );
  TPAOI21D1BWP12T U3944 ( .A1(n3063), .A2(n3062), .B(n3061), .ZN(n3068) );
  IND2XD0BWP12T U3945 ( .A1(n3065), .B1(n3064), .ZN(n3066) );
  INVD1BWP12T U3946 ( .I(n3066), .ZN(n3067) );
  INVD1BWP12T U3947 ( .I(n441), .ZN(n3084) );
  INVD1BWP12T U3948 ( .I(n418), .ZN(n3079) );
  AN2XD2BWP12T U3949 ( .A1(n3079), .A2(n3078), .Z(n3080) );
  XNR2XD4BWP12T U3950 ( .A1(n3081), .A2(n3080), .ZN(n5144) );
  INVD2BWP12T U3951 ( .I(n5144), .ZN(n3090) );
  ND2D1BWP12T U3952 ( .A1(n3086), .A2(n3087), .ZN(n3088) );
  XNR2XD4BWP12T U3953 ( .A1(n3089), .A2(n3088), .ZN(n4692) );
  NR2XD0BWP12T U3954 ( .A1(n3090), .A2(n4692), .ZN(n3091) );
  TPND2D1BWP12T U3955 ( .A1(n3092), .A2(n3091), .ZN(n3102) );
  TPND3D1BWP12T U3956 ( .A1(n3094), .A2(n3093), .A3(n428), .ZN(n3096) );
  TPND2D2BWP12T U3957 ( .A1(n3096), .A2(n3095), .ZN(n3101) );
  AN2XD2BWP12T U3958 ( .A1(n3149), .A2(n3099), .Z(n3100) );
  XNR2XD4BWP12T U3959 ( .A1(n3101), .A2(n3100), .ZN(n4597) );
  INVD1BWP12T U3960 ( .I(n3103), .ZN(n3122) );
  INVD1P75BWP12T U3961 ( .I(n3104), .ZN(n3133) );
  ND2D1BWP12T U3962 ( .A1(n3130), .A2(n3131), .ZN(n3105) );
  XOR2XD4BWP12T U3963 ( .A1(n3133), .A2(n3105), .Z(n4644) );
  INVD1BWP12T U3964 ( .I(n3106), .ZN(n3107) );
  TPAOI21D1BWP12T U3965 ( .A1(n3116), .A2(n3108), .B(n3107), .ZN(n3113) );
  INVD1BWP12T U3966 ( .I(n3109), .ZN(n3111) );
  AN2XD2BWP12T U3967 ( .A1(n3111), .A2(n3110), .Z(n3112) );
  XNR2XD4BWP12T U3968 ( .A1(n3113), .A2(n3112), .ZN(n4628) );
  TPAOI21D1BWP12T U3969 ( .A1(n3116), .A2(n50), .B(n422), .ZN(n3120) );
  AN2XD2BWP12T U3970 ( .A1(n3118), .A2(n3117), .Z(n3119) );
  XNR2XD4BWP12T U3971 ( .A1(n3120), .A2(n3119), .ZN(n4909) );
  TPNR3D1BWP12T U3972 ( .A1(n4644), .A2(n4628), .A3(n4909), .ZN(n3121) );
  TPND2D1BWP12T U3973 ( .A1(n3122), .A2(n3121), .ZN(n3139) );
  TPOAI21D1BWP12T U3974 ( .A1(n3133), .A2(n3124), .B(n72), .ZN(n3129) );
  INVD1BWP12T U3975 ( .I(n3125), .ZN(n3127) );
  XNR2XD4BWP12T U3976 ( .A1(n3129), .A2(n3128), .ZN(n4936) );
  INVD1BWP12T U3977 ( .I(n3130), .ZN(n3132) );
  TPOAI21D1BWP12T U3978 ( .A1(n3133), .A2(n3132), .B(n3131), .ZN(n3136) );
  CKND2D2BWP12T U3979 ( .A1(n408), .A2(n404), .ZN(n3135) );
  XNR2XD4BWP12T U3980 ( .A1(n3136), .A2(n3135), .ZN(n4969) );
  CKND3BWP12T U3981 ( .I(n4969), .ZN(n3137) );
  IND2D2BWP12T U3982 ( .A1(n4936), .B1(n3137), .ZN(n3138) );
  TPAOI21D1BWP12T U3983 ( .A1(n3157), .A2(n3144), .B(n2045), .ZN(n3143) );
  INVD1P75BWP12T U3984 ( .I(n54), .ZN(n3154) );
  XNR2XD4BWP12T U3985 ( .A1(n3143), .A2(n3142), .ZN(n4988) );
  INVD1BWP12T U3986 ( .I(n3145), .ZN(n3147) );
  INVD1P75BWP12T U3987 ( .I(n3148), .ZN(n3156) );
  TPND2D2BWP12T U3988 ( .A1(n3155), .A2(n3154), .ZN(n3160) );
  AOI22D1BWP12T U3989 ( .A1(n3156), .A2(n3157), .B1(n3160), .B2(n3159), .ZN(
        n3165) );
  INVD1BWP12T U3990 ( .I(n3158), .ZN(n3162) );
  TPOAI21D1BWP12T U3991 ( .A1(n3163), .A2(n3162), .B(n3161), .ZN(n3164) );
  INVD1BWP12T U3992 ( .I(n3240), .ZN(n3304) );
  NR2D1BWP12T U3993 ( .A1(n3304), .A2(n3168), .ZN(n3174) );
  INVD0BWP12T U3994 ( .I(n3174), .ZN(n3170) );
  INVD1BWP12T U3995 ( .I(n3243), .ZN(n3236) );
  OAI21D1BWP12T U3996 ( .A1(n3236), .A2(n3168), .B(n3167), .ZN(n3177) );
  INVD1BWP12T U3997 ( .I(n3177), .ZN(n3169) );
  OAI21D1BWP12T U3998 ( .A1(n3314), .A2(n3170), .B(n3169), .ZN(n3173) );
  CKND2D1BWP12T U3999 ( .A1(n3176), .A2(n3171), .ZN(n3172) );
  XNR2D1BWP12T U4000 ( .A1(n3173), .A2(n3172), .ZN(n5061) );
  CKND2D1BWP12T U4001 ( .A1(n3174), .A2(n3176), .ZN(n3179) );
  AOI21D1BWP12T U4002 ( .A1(n3177), .A2(n3176), .B(n3175), .ZN(n3178) );
  OAI21D1BWP12T U4003 ( .A1(n3314), .A2(n3179), .B(n3178), .ZN(n3182) );
  CKND2D1BWP12T U4004 ( .A1(n3181), .A2(n3180), .ZN(n3322) );
  XNR2D1BWP12T U4005 ( .A1(n3182), .A2(n3322), .ZN(n5251) );
  INVD1BWP12T U4006 ( .I(n3194), .ZN(n3260) );
  NR2D1BWP12T U4007 ( .A1(n3260), .A2(n3393), .ZN(n3184) );
  INVD1BWP12T U4008 ( .I(n3250), .ZN(n3311) );
  CKND2D1BWP12T U4009 ( .A1(n3184), .A2(n3311), .ZN(n3186) );
  INVD1BWP12T U4010 ( .I(n3249), .ZN(n3313) );
  INVD1BWP12T U4011 ( .I(n3193), .ZN(n3264) );
  OAI21D1BWP12T U4012 ( .A1(n3264), .A2(n3393), .B(n3198), .ZN(n3183) );
  AOI21D1BWP12T U4013 ( .A1(n3313), .A2(n3184), .B(n3183), .ZN(n3185) );
  OAI21D1BWP12T U4014 ( .A1(n3314), .A2(n3186), .B(n3185), .ZN(n3190) );
  ND2D1BWP12T U4015 ( .A1(n3188), .A2(n3187), .ZN(n3189) );
  XNR2D1BWP12T U4016 ( .A1(n3190), .A2(n3189), .ZN(n5141) );
  CKND2D1BWP12T U4017 ( .A1(n3192), .A2(n3191), .ZN(n3388) );
  AOI21D0BWP12T U4018 ( .A1(n3313), .A2(n3194), .B(n3193), .ZN(n3197) );
  INR3XD0BWP12T U4019 ( .A1(n3194), .B1(n3314), .B2(n3250), .ZN(n3195) );
  INVD1BWP12T U4020 ( .I(n3195), .ZN(n3196) );
  ND2D1BWP12T U4021 ( .A1(n3197), .A2(n3196), .ZN(n3200) );
  CKND2D1BWP12T U4022 ( .A1(n3390), .A2(n3198), .ZN(n3199) );
  XNR2D1BWP12T U4023 ( .A1(n3200), .A2(n3199), .ZN(n4693) );
  INVD0BWP12T U4024 ( .I(n3202), .ZN(n3204) );
  ND2D1BWP12T U4025 ( .A1(n3204), .A2(n3203), .ZN(n3435) );
  INVD0BWP12T U4026 ( .I(n3266), .ZN(n3206) );
  INVD1BWP12T U4027 ( .I(n3269), .ZN(n3205) );
  OAI21D1BWP12T U4028 ( .A1(n3298), .A2(n3206), .B(n3205), .ZN(n3209) );
  ND2D1BWP12T U4029 ( .A1(n3268), .A2(n3207), .ZN(n3208) );
  XNR2D1BWP12T U4030 ( .A1(n3209), .A2(n3208), .ZN(n4984) );
  INVD0BWP12T U4031 ( .I(n3434), .ZN(n3416) );
  CKND2D1BWP12T U4032 ( .A1(n3416), .A2(n3210), .ZN(n3211) );
  XOR2XD1BWP12T U4033 ( .A1(n3298), .A2(n3211), .Z(n4910) );
  INVD0BWP12T U4034 ( .I(n3215), .ZN(n3216) );
  AOI21D1BWP12T U4035 ( .A1(n3222), .A2(n3217), .B(n3216), .ZN(n3219) );
  CKND0BWP12T U4036 ( .I(n3346), .ZN(n3218) );
  CKND2D1BWP12T U4037 ( .A1(n3218), .A2(n3345), .ZN(n3341) );
  XOR2XD1BWP12T U4038 ( .A1(n3219), .A2(n3341), .Z(n5021) );
  AOI21D1BWP12T U4039 ( .A1(n3222), .A2(n3221), .B(n3220), .ZN(n3226) );
  CKND0BWP12T U4040 ( .I(n3223), .ZN(n3352) );
  CKND2D1BWP12T U4041 ( .A1(n3352), .A2(n3224), .ZN(n3225) );
  XOR2XD1BWP12T U4042 ( .A1(n3226), .A2(n3225), .Z(n4884) );
  INVD1BWP12T U4043 ( .I(n3227), .ZN(n3329) );
  CKND2D1BWP12T U4044 ( .A1(n3329), .A2(n3228), .ZN(n3229) );
  XNR2D2BWP12T U4045 ( .A1(n3230), .A2(n3229), .ZN(n5204) );
  ND2XD0BWP12T U4046 ( .A1(n3336), .A2(n3231), .ZN(n3232) );
  XOR2XD1BWP12T U4047 ( .A1(n3232), .A2(n5290), .Z(n4853) );
  INVD1BWP12T U4048 ( .I(b[0]), .ZN(n3233) );
  XNR2D1BWP12T U4049 ( .A1(n3233), .A2(n480), .ZN(n5306) );
  OAI21D1BWP12T U4050 ( .A1(n3314), .A2(n3304), .B(n3236), .ZN(n3239) );
  ND2D1BWP12T U4051 ( .A1(n3242), .A2(n3237), .ZN(n3238) );
  XNR2D1BWP12T U4052 ( .A1(n3239), .A2(n3238), .ZN(n5097) );
  TPND2D0BWP12T U4053 ( .A1(n3240), .A2(n3242), .ZN(n3245) );
  TPAOI21D0BWP12T U4054 ( .A1(n3243), .A2(n3242), .B(n3241), .ZN(n3244) );
  OAI21D1BWP12T U4055 ( .A1(n3314), .A2(n3245), .B(n3244), .ZN(n3248) );
  ND2D1BWP12T U4056 ( .A1(n3246), .A2(n3362), .ZN(n3247) );
  XNR2D1BWP12T U4057 ( .A1(n3248), .A2(n3247), .ZN(n5226) );
  OAI21D0BWP12T U4058 ( .A1(n3314), .A2(n3250), .B(n3249), .ZN(n3252) );
  CKND2D1BWP12T U4059 ( .A1(n3448), .A2(n3447), .ZN(n3251) );
  XNR2XD1BWP12T U4060 ( .A1(n3252), .A2(n3251), .ZN(n4779) );
  NR2D1BWP12T U4061 ( .A1(n3260), .A2(n3259), .ZN(n3255) );
  CKND2D1BWP12T U4062 ( .A1(n3255), .A2(n3311), .ZN(n3257) );
  OAI21D1BWP12T U4063 ( .A1(n3264), .A2(n3259), .B(n3261), .ZN(n3254) );
  AOI21D1BWP12T U4064 ( .A1(n3313), .A2(n3255), .B(n3254), .ZN(n3256) );
  OAI21D1BWP12T U4065 ( .A1(n3314), .A2(n3257), .B(n3256), .ZN(n3258) );
  ND2D1BWP12T U4066 ( .A1(n3263), .A2(n3410), .ZN(n3407) );
  XNR2D1BWP12T U4067 ( .A1(n3258), .A2(n3407), .ZN(n4669) );
  ND2D0BWP12T U4068 ( .A1(n3266), .A2(n3268), .ZN(n3271) );
  TPAOI21D0BWP12T U4069 ( .A1(n3269), .A2(n3268), .B(n3267), .ZN(n3270) );
  OAI21D1BWP12T U4070 ( .A1(n3298), .A2(n3271), .B(n3270), .ZN(n3274) );
  ND2D1BWP12T U4071 ( .A1(n3273), .A2(n3272), .ZN(n3445) );
  XNR2D1BWP12T U4072 ( .A1(n3274), .A2(n3445), .ZN(n4938) );
  CKND0BWP12T U4073 ( .I(n3282), .ZN(n3275) );
  CKND2D1BWP12T U4074 ( .A1(n3275), .A2(n3453), .ZN(n3278) );
  CKND0BWP12T U4075 ( .I(n3285), .ZN(n3276) );
  TPAOI21D0BWP12T U4076 ( .A1(n3276), .A2(n3453), .B(n3452), .ZN(n3277) );
  OAI21D1BWP12T U4077 ( .A1(n3298), .A2(n3278), .B(n3277), .ZN(n3281) );
  ND2D1BWP12T U4078 ( .A1(n3280), .A2(n3279), .ZN(n3458) );
  XNR2D1BWP12T U4079 ( .A1(n3281), .A2(n3458), .ZN(n4624) );
  NR2D1BWP12T U4080 ( .A1(n3282), .A2(n3284), .ZN(n3292) );
  INVD1BWP12T U4081 ( .I(n3292), .ZN(n3287) );
  OAI21D1BWP12T U4082 ( .A1(n3285), .A2(n3284), .B(n3283), .ZN(n3295) );
  INVD1BWP12T U4083 ( .I(n3295), .ZN(n3286) );
  OAI21D1BWP12T U4084 ( .A1(n3298), .A2(n3287), .B(n3286), .ZN(n3290) );
  ND2D1BWP12T U4085 ( .A1(n3294), .A2(n3288), .ZN(n3289) );
  XNR2D2BWP12T U4086 ( .A1(n3290), .A2(n3289), .ZN(n5002) );
  CKND2D1BWP12T U4087 ( .A1(n3292), .A2(n3294), .ZN(n3297) );
  AOI21D1BWP12T U4088 ( .A1(n3295), .A2(n3294), .B(n3293), .ZN(n3296) );
  OAI21D1BWP12T U4089 ( .A1(n3298), .A2(n3297), .B(n3296), .ZN(n3301) );
  ND2D1BWP12T U4090 ( .A1(n3300), .A2(n3299), .ZN(n3484) );
  XNR2D2BWP12T U4091 ( .A1(n3301), .A2(n3484), .ZN(n5175) );
  AOI21D1BWP12T U4092 ( .A1(n3313), .A2(n3448), .B(n3376), .ZN(n3306) );
  INR2XD0BWP12T U4093 ( .A1(n3448), .B1(n3314), .ZN(n3303) );
  IND3D1BWP12T U4094 ( .A1(n3304), .B1(n3303), .B2(n3302), .ZN(n3305) );
  ND2D1BWP12T U4095 ( .A1(n3306), .A2(n3305), .ZN(n3309) );
  TPND2D0BWP12T U4096 ( .A1(n3308), .A2(n3307), .ZN(n3377) );
  XNR2D1BWP12T U4097 ( .A1(n3309), .A2(n3377), .ZN(n4839) );
  CKND0BWP12T U4098 ( .I(n3367), .ZN(n3316) );
  NR2D0BWP12T U4099 ( .A1(n3316), .A2(n3371), .ZN(n3319) );
  INVD1BWP12T U4100 ( .I(n3420), .ZN(n3365) );
  ND2D0BWP12T U4101 ( .A1(n3319), .A2(n3365), .ZN(n3321) );
  INVD1BWP12T U4102 ( .I(n3419), .ZN(n3368) );
  CKND0BWP12T U4103 ( .I(n3366), .ZN(n3317) );
  OAI21D0BWP12T U4104 ( .A1(n3317), .A2(n3371), .B(n3372), .ZN(n3318) );
  AOI21D1BWP12T U4105 ( .A1(n3368), .A2(n3319), .B(n3318), .ZN(n3320) );
  OAI21D1BWP12T U4106 ( .A1(n3421), .A2(n3321), .B(n3320), .ZN(n3323) );
  XNR2D1BWP12T U4107 ( .A1(n3323), .A2(n3322), .ZN(n5283) );
  CKND0BWP12T U4108 ( .I(n3324), .ZN(n3358) );
  INVD1BWP12T U4109 ( .I(n3325), .ZN(n3337) );
  INVD1BWP12T U4110 ( .I(n3908), .ZN(n3326) );
  TPNR2D1BWP12T U4111 ( .A1(n3326), .A2(n3684), .ZN(n3327) );
  OAI21D1BWP12T U4112 ( .A1(n3337), .A2(n3327), .B(n3671), .ZN(n3331) );
  ND2XD0BWP12T U4113 ( .A1(n3329), .A2(n3328), .ZN(n3330) );
  XNR2D1BWP12T U4114 ( .A1(n3331), .A2(n3330), .ZN(n5205) );
  INVD1BWP12T U4115 ( .I(n3332), .ZN(n4437) );
  ND2D1BWP12T U4116 ( .A1(n4437), .A2(n3333), .ZN(n3335) );
  INVD1BWP12T U4117 ( .I(b[0]), .ZN(n3334) );
  XNR2D1BWP12T U4118 ( .A1(n3335), .A2(n3334), .ZN(n5307) );
  OR3D0BWP12T U4119 ( .A1(n5307), .A2(n5105), .A3(n4854), .Z(n3338) );
  NR4D0BWP12T U4120 ( .A1(n3340), .A2(n3339), .A3(n5205), .A4(n3338), .ZN(
        n3357) );
  CKND0BWP12T U4121 ( .I(n3342), .ZN(n3343) );
  NR2XD0BWP12T U4122 ( .A1(n3343), .A2(n3346), .ZN(n3349) );
  CKND0BWP12T U4123 ( .I(n3344), .ZN(n3347) );
  OAI21D0BWP12T U4124 ( .A1(n3347), .A2(n3346), .B(n3345), .ZN(n3348) );
  AOI21D1BWP12T U4125 ( .A1(n3350), .A2(n3349), .B(n3348), .ZN(n3354) );
  ND2XD0BWP12T U4126 ( .A1(n3352), .A2(n3351), .ZN(n3353) );
  XOR2XD1BWP12T U4127 ( .A1(n3354), .A2(n3353), .Z(n4879) );
  NR3D0BWP12T U4128 ( .A1(n3355), .A2(n5014), .A3(n4879), .ZN(n3356) );
  IND4D1BWP12T U4129 ( .A1(n5283), .B1(n3358), .B2(n3357), .B3(n3356), .ZN(
        n3375) );
  CKND2D1BWP12T U4130 ( .A1(n3365), .A2(n3242), .ZN(n3360) );
  AOI21D1BWP12T U4131 ( .A1(n3368), .A2(n3242), .B(n3241), .ZN(n3359) );
  OAI21D1BWP12T U4132 ( .A1(n3421), .A2(n3360), .B(n3359), .ZN(n3364) );
  CKND2D1BWP12T U4133 ( .A1(n3246), .A2(n3362), .ZN(n3363) );
  XNR2D1BWP12T U4134 ( .A1(n3364), .A2(n3363), .ZN(n5225) );
  TPND2D0BWP12T U4135 ( .A1(n3365), .A2(n3367), .ZN(n3370) );
  AOI21D1BWP12T U4136 ( .A1(n3368), .A2(n3367), .B(n3366), .ZN(n3369) );
  OAI21D1BWP12T U4137 ( .A1(n3421), .A2(n3370), .B(n3369), .ZN(n3374) );
  ND2D1BWP12T U4138 ( .A1(n3176), .A2(n3372), .ZN(n3373) );
  XNR2D1BWP12T U4139 ( .A1(n3374), .A2(n3373), .ZN(n5065) );
  NR3XD0BWP12T U4140 ( .A1(n3375), .A2(n5225), .A3(n5065), .ZN(n3431) );
  AOI21D1BWP12T U4141 ( .A1(n3483), .A2(n3448), .B(n3376), .ZN(n3378) );
  XOR2XD1BWP12T U4142 ( .A1(n3378), .A2(n3377), .Z(n4837) );
  CKND0BWP12T U4143 ( .I(n3380), .ZN(n3381) );
  NR2D0BWP12T U4144 ( .A1(n3381), .A2(n3384), .ZN(n3387) );
  CKND0BWP12T U4145 ( .I(n3382), .ZN(n3385) );
  OAI21D0BWP12T U4146 ( .A1(n3385), .A2(n3384), .B(n3383), .ZN(n3386) );
  AOI21D1BWP12T U4147 ( .A1(n3483), .A2(n3387), .B(n3386), .ZN(n3389) );
  XOR2XD1BWP12T U4148 ( .A1(n3389), .A2(n3388), .Z(n4726) );
  INVD1BWP12T U4149 ( .I(n3391), .ZN(n3401) );
  INVD1BWP12T U4150 ( .I(n3394), .ZN(n3404) );
  NR4D0BWP12T U4151 ( .A1(n4837), .A2(n4786), .A3(n4726), .A4(n4720), .ZN(
        n3430) );
  NR2D0BWP12T U4152 ( .A1(n3391), .A2(n3393), .ZN(n3396) );
  TPOAI21D0BWP12T U4153 ( .A1(n3394), .A2(n3393), .B(n3392), .ZN(n3395) );
  AOI21D1BWP12T U4154 ( .A1(n3483), .A2(n3396), .B(n3395), .ZN(n3400) );
  ND2D1BWP12T U4155 ( .A1(n3188), .A2(n3398), .ZN(n3399) );
  XOR2XD1BWP12T U4156 ( .A1(n3400), .A2(n3399), .Z(n5139) );
  CKND2D1BWP12T U4157 ( .A1(n3401), .A2(n3403), .ZN(n3409) );
  INVD0BWP12T U4158 ( .I(n3409), .ZN(n3406) );
  AOI21D1BWP12T U4159 ( .A1(n3404), .A2(n3403), .B(n3402), .ZN(n3412) );
  INVD1BWP12T U4160 ( .I(n3412), .ZN(n3405) );
  AOI21D1BWP12T U4161 ( .A1(n3483), .A2(n3406), .B(n3405), .ZN(n3408) );
  XOR2XD1BWP12T U4162 ( .A1(n3408), .A2(n3407), .Z(n4687) );
  AOI21D1BWP12T U4163 ( .A1(n3483), .A2(n3433), .B(n3415), .ZN(n3418) );
  CKND2D1BWP12T U4164 ( .A1(n3416), .A2(n3432), .ZN(n3417) );
  XOR2XD1BWP12T U4165 ( .A1(n3418), .A2(n3417), .Z(n4911) );
  NR4D0BWP12T U4166 ( .A1(n5139), .A2(n4687), .A3(n4629), .A4(n4911), .ZN(
        n3429) );
  TPOAI21D0BWP12T U4167 ( .A1(n3421), .A2(n3420), .B(n3419), .ZN(n3424) );
  CKND2D1BWP12T U4168 ( .A1(n3242), .A2(n3422), .ZN(n3423) );
  XNR2XD1BWP12T U4169 ( .A1(n3424), .A2(n3423), .ZN(n5095) );
  NR4D0BWP12T U4170 ( .A1(n3427), .A2(n3426), .A3(n3425), .A4(n5095), .ZN(
        n3428) );
  INVD0BWP12T U4171 ( .I(n3442), .ZN(n3437) );
  TPNR2D0BWP12T U4172 ( .A1(n3470), .A2(n3437), .ZN(n3439) );
  INVD1BWP12T U4173 ( .I(n3444), .ZN(n3436) );
  OAI21D1BWP12T U4174 ( .A1(n3480), .A2(n3437), .B(n3436), .ZN(n3438) );
  AOI21D1BWP12T U4175 ( .A1(n3483), .A2(n3439), .B(n3438), .ZN(n3441) );
  CKND2D1BWP12T U4176 ( .A1(n3268), .A2(n3443), .ZN(n3440) );
  XOR2XD1BWP12T U4177 ( .A1(n3441), .A2(n3440), .Z(n4983) );
  CKND2D1BWP12T U4178 ( .A1(n3448), .A2(n3447), .ZN(n3449) );
  XNR2D1BWP12T U4179 ( .A1(n3483), .A2(n3449), .ZN(n4777) );
  INVD1BWP12T U4180 ( .I(n3450), .ZN(n3469) );
  CKND2D1BWP12T U4181 ( .A1(n3469), .A2(n3453), .ZN(n3455) );
  TPNR2D0BWP12T U4182 ( .A1(n3470), .A2(n3455), .ZN(n3457) );
  INVD1BWP12T U4183 ( .I(n3451), .ZN(n3477) );
  AOI21D1BWP12T U4184 ( .A1(n3477), .A2(n3453), .B(n3452), .ZN(n3454) );
  OAI21D1BWP12T U4185 ( .A1(n3480), .A2(n3455), .B(n3454), .ZN(n3456) );
  AOI21D1BWP12T U4186 ( .A1(n3483), .A2(n3457), .B(n3456), .ZN(n3459) );
  XOR2XD1BWP12T U4187 ( .A1(n3459), .A2(n3458), .Z(n4622) );
  CKND2D1BWP12T U4188 ( .A1(n3469), .A2(n3467), .ZN(n3461) );
  TPNR2D0BWP12T U4189 ( .A1(n3470), .A2(n3461), .ZN(n3463) );
  AOI21D1BWP12T U4190 ( .A1(n3477), .A2(n3467), .B(n3471), .ZN(n3460) );
  OAI21D1BWP12T U4191 ( .A1(n3480), .A2(n3461), .B(n3460), .ZN(n3462) );
  AOI21D1BWP12T U4192 ( .A1(n3483), .A2(n3463), .B(n3462), .ZN(n3466) );
  INVD1BWP12T U4193 ( .I(n3473), .ZN(n3464) );
  ND2D1BWP12T U4194 ( .A1(n3464), .A2(n3472), .ZN(n3465) );
  XOR2XD1BWP12T U4195 ( .A1(n3466), .A2(n3465), .Z(n5001) );
  INVD0BWP12T U4196 ( .I(n3467), .ZN(n3468) );
  NR2D1BWP12T U4197 ( .A1(n3468), .A2(n3473), .ZN(n3476) );
  ND2D1BWP12T U4198 ( .A1(n3476), .A2(n3469), .ZN(n3479) );
  TPNR2D0BWP12T U4199 ( .A1(n3470), .A2(n3479), .ZN(n3482) );
  CKND0BWP12T U4200 ( .I(n3471), .ZN(n3474) );
  TPOAI21D0BWP12T U4201 ( .A1(n3474), .A2(n3473), .B(n3472), .ZN(n3475) );
  AOI21D1BWP12T U4202 ( .A1(n3477), .A2(n3476), .B(n3475), .ZN(n3478) );
  OAI21D1BWP12T U4203 ( .A1(n3480), .A2(n3479), .B(n3478), .ZN(n3481) );
  AOI21D1BWP12T U4204 ( .A1(n3483), .A2(n3482), .B(n3481), .ZN(n3485) );
  XOR2XD1BWP12T U4205 ( .A1(n3485), .A2(n3484), .Z(n5174) );
  TPNR2D0BWP12T U4206 ( .A1(n2269), .A2(n3539), .ZN(n3486) );
  ND2D1BWP12T U4207 ( .A1(n3511), .A2(n3486), .ZN(n3490) );
  ND2D1BWP12T U4208 ( .A1(n3488), .A2(n3487), .ZN(n3489) );
  TPOAI21D1BWP12T U4209 ( .A1(n3491), .A2(n3490), .B(n3489), .ZN(n4300) );
  INVD1BWP12T U4210 ( .I(n3544), .ZN(n3493) );
  TPAOI21D0BWP12T U4211 ( .A1(n3493), .A2(n3875), .B(n5214), .ZN(n3508) );
  AOI22D0BWP12T U4212 ( .A1(n3496), .A2(n3495), .B1(n3494), .B2(n4510), .ZN(
        n3500) );
  AOI22D0BWP12T U4213 ( .A1(n3498), .A2(n4891), .B1(n3497), .B2(n4511), .ZN(
        n3499) );
  CKND2D1BWP12T U4214 ( .A1(n3500), .A2(n3499), .ZN(n3514) );
  NR2D1BWP12T U4215 ( .A1(n3514), .A2(n3539), .ZN(n3504) );
  OAI21D0BWP12T U4216 ( .A1(n3594), .A2(n5192), .B(n3905), .ZN(n3501) );
  NR4D1BWP12T U4217 ( .A1(n3504), .A2(n3503), .A3(n3502), .A4(n3501), .ZN(
        n3507) );
  AOI21D0BWP12T U4218 ( .A1(n3515), .A2(n3707), .B(n4301), .ZN(n3505) );
  OAI21D0BWP12T U4219 ( .A1(n3513), .A2(n3609), .B(n3505), .ZN(n3506) );
  TPOAI21D1BWP12T U4220 ( .A1(n3508), .A2(n5211), .B(n3565), .ZN(n5220) );
  MUX2ND0BWP12T U4221 ( .I0(n3509), .I1(n5108), .S(n5196), .ZN(n3525) );
  ND3D1BWP12T U4222 ( .A1(n3512), .A2(n3511), .A3(n3510), .ZN(n3526) );
  AOI22D1BWP12T U4223 ( .A1(n3526), .A2(n4601), .B1(n3527), .B2(n3617), .ZN(
        n3698) );
  TPOAI21D0BWP12T U4224 ( .A1(n3525), .A2(n3905), .B(n3698), .ZN(n3542) );
  INVD1BWP12T U4225 ( .I(n3542), .ZN(n4634) );
  TPOAI21D0BWP12T U4226 ( .A1(n4634), .A2(n3838), .B(n3844), .ZN(n3523) );
  INVD1BWP12T U4227 ( .I(n3513), .ZN(n3530) );
  AOI22D1BWP12T U4228 ( .A1(n4601), .A2(n3514), .B1(n3530), .B2(n3707), .ZN(
        n3522) );
  CKND0BWP12T U4229 ( .I(n3515), .ZN(n3516) );
  TPOAI21D0BWP12T U4230 ( .A1(n3516), .A2(n3607), .B(n3882), .ZN(n3520) );
  NR2D1BWP12T U4231 ( .A1(n3518), .A2(n3517), .ZN(n3529) );
  TPNR2D0BWP12T U4232 ( .A1(n3529), .A2(n3609), .ZN(n3519) );
  NR2D1BWP12T U4233 ( .A1(n3520), .A2(n3519), .ZN(n3521) );
  ND2D1BWP12T U4234 ( .A1(n3522), .A2(n3521), .ZN(n4902) );
  AOI21D1BWP12T U4235 ( .A1(n3523), .A2(n4902), .B(n5323), .ZN(n4903) );
  OAI21D1BWP12T U4236 ( .A1(n3525), .A2(n3948), .B(n3524), .ZN(n3543) );
  INVD1BWP12T U4237 ( .I(n3543), .ZN(n5156) );
  CKMUX2D1BWP12T U4238 ( .I0(n3527), .I1(n3526), .S(n4175), .Z(n3528) );
  OAI21D1BWP12T U4239 ( .A1(n3528), .A2(n4301), .B(n4953), .ZN(n3533) );
  INVD1BWP12T U4240 ( .I(n3529), .ZN(n3531) );
  AOI22D1BWP12T U4241 ( .A1(n3617), .A2(n3531), .B1(n3530), .B2(n4601), .ZN(
        n3532) );
  ND2D1BWP12T U4242 ( .A1(n3533), .A2(n3532), .ZN(n3729) );
  CKND2D0BWP12T U4243 ( .A1(n4903), .A2(n5272), .ZN(n3534) );
  NR2D0BWP12T U4244 ( .A1(n5220), .A2(n3534), .ZN(n3636) );
  AOI21D1BWP12T U4245 ( .A1(n3547), .A2(n3948), .B(n3695), .ZN(n4801) );
  OAI22D1BWP12T U4246 ( .A1(n4176), .A2(n3607), .B1(n3619), .B2(n3730), .ZN(
        n3708) );
  CKND1BWP12T U4247 ( .I(n3537), .ZN(n3540) );
  TPNR2D0BWP12T U4248 ( .A1(n3855), .A2(n3564), .ZN(n3538) );
  AOI21D1BWP12T U4249 ( .A1(n3540), .A2(n3539), .B(n3538), .ZN(n3549) );
  ND4D0BWP12T U4250 ( .A1(n4801), .A2(n4819), .A3(n4678), .A4(n4703), .ZN(
        n3541) );
  OAI31D0BWP12T U4251 ( .A1(n3543), .A2(n3542), .A3(n3541), .B(n4633), .ZN(
        n3546) );
  INVD1BWP12T U4252 ( .I(n4633), .ZN(n3582) );
  TPOAI21D0BWP12T U4253 ( .A1(n3544), .A2(n3582), .B(n3580), .ZN(n4746) );
  INR3XD0BWP12T U4254 ( .A1(n3546), .B1(n3545), .B2(n4746), .ZN(n3635) );
  INVD1BWP12T U4255 ( .I(n3580), .ZN(n4941) );
  TPNR2D1BWP12T U4256 ( .A1(n4941), .A2(n3625), .ZN(n4657) );
  ND2D1BWP12T U4257 ( .A1(n3565), .A2(n3582), .ZN(n3554) );
  OAI21D0BWP12T U4258 ( .A1(n4980), .A2(n4942), .B(n3554), .ZN(n3550) );
  INVD1BWP12T U4259 ( .I(n4657), .ZN(n3552) );
  AOI21D1BWP12T U4260 ( .A1(n3548), .A2(n4633), .B(n3552), .ZN(n4912) );
  INR2D1BWP12T U4261 ( .A1(n3905), .B1(n3549), .ZN(n3626) );
  TPOAI21D0BWP12T U4262 ( .A1(n3552), .A2(n3626), .B(n3554), .ZN(n4997) );
  ND4D0BWP12T U4263 ( .A1(n3551), .A2(n3550), .A3(n4912), .A4(n4997), .ZN(
        n3567) );
  IOA21D0BWP12T U4264 ( .A1(n3580), .A2(n3553), .B(n3552), .ZN(n3556) );
  INVD1BWP12T U4265 ( .I(n5127), .ZN(n3555) );
  INVD1BWP12T U4266 ( .I(n3554), .ZN(n4940) );
  AOI21D1BWP12T U4267 ( .A1(n3556), .A2(n3555), .B(n4940), .ZN(n5115) );
  INVD1BWP12T U4268 ( .I(n3557), .ZN(n3563) );
  CKND0BWP12T U4269 ( .I(n3558), .ZN(n3561) );
  AOI21D1BWP12T U4270 ( .A1(n3559), .A2(n4601), .B(n4301), .ZN(n3560) );
  IOA21D1BWP12T U4271 ( .A1(n3617), .A2(n3561), .B(n3560), .ZN(n3562) );
  AOI21D1BWP12T U4272 ( .A1(n3563), .A2(n3948), .B(n3562), .ZN(n3732) );
  MUX2NXD0BWP12T U4273 ( .I0(n3731), .I1(n3564), .S(n3730), .ZN(n3579) );
  NR4D0BWP12T U4274 ( .A1(n3567), .A2(n3566), .A3(n5115), .A4(n5230), .ZN(
        n3634) );
  NR2D1BWP12T U4275 ( .A1(n4819), .A2(n3882), .ZN(n4210) );
  NR2D1BWP12T U4276 ( .A1(n3571), .A2(n3730), .ZN(n3774) );
  AOI22D1BWP12T U4277 ( .A1(n3875), .A2(n4210), .B1(n5320), .B2(n5214), .ZN(
        n5328) );
  OAI211D0BWP12T U4278 ( .A1(n3583), .A2(n3582), .B(n3581), .C(n5322), .ZN(
        n3584) );
  NR2D0BWP12T U4279 ( .A1(n4614), .A2(n3584), .ZN(n3585) );
  ND4D0BWP12T U4280 ( .A1(n3586), .A2(n5328), .A3(n5078), .A4(n3585), .ZN(
        n3632) );
  OAI22D0BWP12T U4281 ( .A1(n3588), .A2(n5032), .B1(n3587), .B2(n3900), .ZN(
        n3593) );
  OAI22D0BWP12T U4282 ( .A1(n3591), .A2(n437), .B1(n3589), .B2(n3910), .ZN(
        n3592) );
  NR2D1BWP12T U4283 ( .A1(n3593), .A2(n3592), .ZN(n3610) );
  NR2D1BWP12T U4284 ( .A1(n3610), .A2(n3607), .ZN(n3601) );
  IND2D0BWP12T U4285 ( .A1(n3806), .B1(n5192), .ZN(n3598) );
  TPAOI21D1BWP12T U4286 ( .A1(n3603), .A2(n4870), .B(n5323), .ZN(n4866) );
  CKND2D0BWP12T U4287 ( .A1(n3604), .A2(n4866), .ZN(n3631) );
  OAI22D1BWP12T U4288 ( .A1(n3606), .A2(n4953), .B1(n3605), .B2(n3861), .ZN(
        n4764) );
  AOI21D1BWP12T U4289 ( .A1(n4764), .A2(n3875), .B(n4941), .ZN(n4756) );
  OAI22D0BWP12T U4290 ( .A1(n3614), .A2(n3609), .B1(n3608), .B2(n3607), .ZN(
        n3613) );
  TPOAI21D0BWP12T U4291 ( .A1(n3620), .A2(n3618), .B(n3882), .ZN(n3612) );
  NR2D1BWP12T U4292 ( .A1(n3610), .A2(n3730), .ZN(n3611) );
  NR3D1BWP12T U4293 ( .A1(n3613), .A2(n3612), .A3(n3611), .ZN(n5008) );
  NR2D1BWP12T U4294 ( .A1(n5008), .A2(n3838), .ZN(n5035) );
  INVD0BWP12T U4295 ( .I(n3614), .ZN(n3616) );
  AOI22D1BWP12T U4296 ( .A1(n3617), .A2(n3616), .B1(n3615), .B2(n3703), .ZN(
        n3624) );
  OAI21D0BWP12T U4297 ( .A1(n3619), .A2(n3618), .B(n3882), .ZN(n3622) );
  NR2D1BWP12T U4298 ( .A1(n3622), .A2(n3621), .ZN(n3623) );
  ND2D1BWP12T U4299 ( .A1(n3624), .A2(n3623), .ZN(n3734) );
  NR2D0BWP12T U4300 ( .A1(n3626), .A2(n3625), .ZN(n3627) );
  OAI21D0BWP12T U4301 ( .A1(n3627), .A2(n3838), .B(n3844), .ZN(n3628) );
  AOI21D1BWP12T U4302 ( .A1(n3734), .A2(n3628), .B(n5323), .ZN(n5043) );
  ND4D0BWP12T U4303 ( .A1(n3629), .A2(n4756), .A3(n5029), .A4(n5043), .ZN(
        n3630) );
  TPNR3D0BWP12T U4304 ( .A1(n3632), .A2(n3631), .A3(n3630), .ZN(n3633) );
  ND4D1BWP12T U4305 ( .A1(n3636), .A2(n3635), .A3(n3634), .A4(n3633), .ZN(
        n3693) );
  AOI22D1BWP12T U4306 ( .A1(n454), .A2(n3637), .B1(n2250), .B2(n4568), .ZN(
        n3647) );
  AOI22D1BWP12T U4307 ( .A1(n5118), .A2(n3639), .B1(n3638), .B2(n4914), .ZN(
        n3646) );
  AOI22D0BWP12T U4308 ( .A1(a[18]), .A2(n3641), .B1(n3640), .B2(n4672), .ZN(
        n3645) );
  AOI22D0BWP12T U4309 ( .A1(n448), .A2(n3643), .B1(n3642), .B2(n4565), .ZN(
        n3644) );
  ND4D1BWP12T U4310 ( .A1(n3647), .A2(n3646), .A3(n3645), .A4(n3644), .ZN(
        n3678) );
  AOI22D0BWP12T U4311 ( .A1(n5256), .A2(n1222), .B1(n3648), .B2(a[17]), .ZN(
        n3657) );
  AOI22D0BWP12T U4312 ( .A1(n5234), .A2(n3650), .B1(n3649), .B2(n4508), .ZN(
        n3656) );
  AOI22D0BWP12T U4313 ( .A1(n4518), .A2(n3652), .B1(n3651), .B2(n4502), .ZN(
        n3655) );
  AOI22D0BWP12T U4314 ( .A1(n5079), .A2(n2155), .B1(n3653), .B2(n4509), .ZN(
        n3654) );
  ND4D1BWP12T U4315 ( .A1(n3657), .A2(n3656), .A3(n3655), .A4(n3654), .ZN(
        n3677) );
  AOI22D0BWP12T U4316 ( .A1(n4891), .A2(n2227), .B1(n3658), .B2(n4511), .ZN(
        n3665) );
  AOI22D0BWP12T U4317 ( .A1(n4541), .A2(n3882), .B1(n3659), .B2(n4510), .ZN(
        n3664) );
  AOI22D0BWP12T U4318 ( .A1(n5192), .A2(n3906), .B1(n3660), .B2(n5030), .ZN(
        n3663) );
  AOI22D0BWP12T U4319 ( .A1(n480), .A2(n3233), .B1(n3905), .B2(n3661), .ZN(
        n3662) );
  ND4D1BWP12T U4320 ( .A1(n3665), .A2(n3664), .A3(n3663), .A4(n3662), .ZN(
        n3676) );
  AOI22D1BWP12T U4321 ( .A1(n1), .A2(n3667), .B1(n3666), .B2(n5146), .ZN(n3674) );
  AOI22D1BWP12T U4322 ( .A1(n4943), .A2(n689), .B1(n3668), .B2(n4990), .ZN(
        n3673) );
  AOI22D1BWP12T U4323 ( .A1(n4649), .A2(n3670), .B1(n3669), .B2(n2773), .ZN(
        n3672) );
  ND4D1BWP12T U4324 ( .A1(n3674), .A2(n3673), .A3(n3672), .A4(n3671), .ZN(
        n3675) );
  NR4D0BWP12T U4325 ( .A1(n3678), .A2(n3677), .A3(n3676), .A4(n3675), .ZN(
        n3958) );
  CKND2D0BWP12T U4326 ( .A1(n4170), .A2(n5148), .ZN(n3810) );
  NR4D0BWP12T U4327 ( .A1(n4672), .A2(n3679), .A3(n5030), .A4(n4509), .ZN(
        n3683) );
  NR4D0BWP12T U4328 ( .A1(a[18]), .A2(n5118), .A3(n4696), .A4(a[25]), .ZN(
        n3682) );
  NR4D0BWP12T U4329 ( .A1(n2825), .A2(n4649), .A3(n4914), .A4(n4943), .ZN(
        n3681) );
  NR4D0BWP12T U4330 ( .A1(n2773), .A2(n4990), .A3(n1), .A4(n480), .ZN(n3680)
         );
  ND4D1BWP12T U4331 ( .A1(n3683), .A2(n3682), .A3(n3681), .A4(n3680), .ZN(
        n3690) );
  NR4D0BWP12T U4332 ( .A1(n4518), .A2(n4521), .A3(n5192), .A4(n4541), .ZN(
        n3685) );
  ND4D0BWP12T U4333 ( .A1(n3685), .A2(n5296), .A3(n3898), .A4(n410), .ZN(n3689) );
  NR4D0BWP12T U4334 ( .A1(n5256), .A2(n448), .A3(n4508), .A4(n4891), .ZN(n3687) );
  NR4D0BWP12T U4335 ( .A1(n4788), .A2(n5049), .A3(n5234), .A4(n3661), .ZN(
        n3686) );
  CKND2D1BWP12T U4336 ( .A1(n3687), .A2(n3686), .ZN(n3688) );
  NR4D0BWP12T U4337 ( .A1(n3810), .A2(n3690), .A3(n3689), .A4(n3688), .ZN(
        n3691) );
  AOI22D0BWP12T U4338 ( .A1(n3958), .A2(n3925), .B1(n3691), .B2(n3875), .ZN(
        n3692) );
  AOI21D0BWP12T U4339 ( .A1(n3693), .A2(n3692), .B(n5108), .ZN(n4128) );
  AOI21D0BWP12T U4340 ( .A1(n4176), .A2(n3906), .B(n3905), .ZN(n3694) );
  NR2D1BWP12T U4341 ( .A1(n3695), .A2(n3694), .ZN(n3697) );
  INR2D1BWP12T U4342 ( .A1(n3703), .B1(n4995), .ZN(n3696) );
  TPNR2D1BWP12T U4343 ( .A1(n3697), .A2(n3696), .ZN(n4209) );
  CKND1BWP12T U4344 ( .I(n4209), .ZN(n4795) );
  ND4D0BWP12T U4345 ( .A1(n4710), .A2(n4819), .A3(n4978), .A4(n4795), .ZN(
        n3702) );
  INVD1BWP12T U4346 ( .I(n3727), .ZN(n5160) );
  CKND0BWP12T U4347 ( .I(n4995), .ZN(n4177) );
  CKND0BWP12T U4348 ( .I(n3726), .ZN(n3699) );
  ND4D0BWP12T U4349 ( .A1(n4177), .A2(n3731), .A3(n3727), .A4(n3699), .ZN(
        n3700) );
  NR3D0BWP12T U4350 ( .A1(n3717), .A2(n4660), .A3(n3700), .ZN(n3701) );
  CKND2D0BWP12T U4351 ( .A1(n4925), .A2(n3701), .ZN(n4197) );
  NR2D0BWP12T U4352 ( .A1(n3702), .A2(n4197), .ZN(n3712) );
  ND2XD0BWP12T U4353 ( .A1(n3727), .A2(n3703), .ZN(n3706) );
  INVD1BWP12T U4354 ( .I(n3704), .ZN(n3705) );
  INR2XD1BWP12T U4355 ( .A1(n3706), .B1(n3705), .ZN(n4738) );
  CKND0BWP12T U4356 ( .I(n3724), .ZN(n4289) );
  NR3D0BWP12T U4357 ( .A1(n4738), .A2(n4289), .A3(n4945), .ZN(n3711) );
  CKND2D1BWP12T U4358 ( .A1(n4995), .A2(n3707), .ZN(n3710) );
  INVD1BWP12T U4359 ( .I(n3708), .ZN(n3709) );
  NR2D0BWP12T U4360 ( .A1(n5127), .A2(n5009), .ZN(n4291) );
  AOI31D0BWP12T U4361 ( .A1(n3712), .A2(n3711), .A3(n4291), .B(n3844), .ZN(
        n3722) );
  NR2D1BWP12T U4362 ( .A1(n4209), .A2(n3882), .ZN(n4869) );
  CKND0BWP12T U4363 ( .I(n4870), .ZN(n3716) );
  INVD1BWP12T U4364 ( .I(n5009), .ZN(n4681) );
  ND2D1BWP12T U4365 ( .A1(n4681), .A2(n4301), .ZN(n4196) );
  AOI21D0BWP12T U4366 ( .A1(n5035), .A2(n4196), .B(n3713), .ZN(n3715) );
  OAI211D0BWP12T U4367 ( .A1(n4869), .A2(n3716), .B(n3715), .C(n3714), .ZN(
        n3721) );
  CKND1BWP12T U4368 ( .I(n4902), .ZN(n4287) );
  INVD1BWP12T U4369 ( .I(n3717), .ZN(n4890) );
  ND4D0BWP12T U4370 ( .A1(n5328), .A2(n5212), .A3(n4882), .A4(n3718), .ZN(
        n3719) );
  NR4D0BWP12T U4371 ( .A1(n3722), .A2(n3721), .A3(n3720), .A4(n3719), .ZN(
        n3965) );
  NR3D0BWP12T U4372 ( .A1(n3725), .A2(n5073), .A3(n4764), .ZN(n4283) );
  ND2D1BWP12T U4373 ( .A1(n3726), .A2(n4301), .ZN(n4762) );
  OAI21D1BWP12T U4374 ( .A1(n3727), .A2(n3730), .B(n4301), .ZN(n3728) );
  ND2D1BWP12T U4375 ( .A1(n3729), .A2(n3728), .ZN(n5276) );
  AOI31D0BWP12T U4376 ( .A1(n4283), .A2(n4762), .A3(n5276), .B(n3838), .ZN(
        n3741) );
  CKND2D1BWP12T U4377 ( .A1(n4738), .A2(n3875), .ZN(n5210) );
  AOI21D0BWP12T U4378 ( .A1(n5210), .A2(n3844), .B(n5211), .ZN(n3740) );
  OAI21D1BWP12T U4379 ( .A1(n3731), .A2(n3730), .B(n4301), .ZN(n3733) );
  INR2D1BWP12T U4380 ( .A1(n3733), .B1(n3732), .ZN(n5240) );
  INVD1BWP12T U4381 ( .I(n3734), .ZN(n3736) );
  TPAOI21D0BWP12T U4382 ( .A1(n4995), .A2(n4601), .B(n3882), .ZN(n3735) );
  TPNR2D1BWP12T U4383 ( .A1(n3736), .A2(n3735), .ZN(n5048) );
  OAI21D0BWP12T U4384 ( .A1(n5240), .A2(n5048), .B(n3875), .ZN(n3738) );
  CKND2D0BWP12T U4385 ( .A1(n3738), .A2(n3737), .ZN(n3739) );
  TPNR3D0BWP12T U4386 ( .A1(n3741), .A2(n3740), .A3(n3739), .ZN(n3964) );
  OAI22D0BWP12T U4387 ( .A1(n4153), .A2(n3872), .B1(n4131), .B2(n3871), .ZN(
        n3743) );
  OAI22D0BWP12T U4388 ( .A1(n4152), .A2(n3869), .B1(n4140), .B2(n3870), .ZN(
        n3742) );
  NR2D1BWP12T U4389 ( .A1(n3743), .A2(n3742), .ZN(n3767) );
  OAI22D0BWP12T U4390 ( .A1(n4241), .A2(n3872), .B1(n4243), .B2(n3871), .ZN(
        n3745) );
  OAI22D0BWP12T U4391 ( .A1(n4130), .A2(n3869), .B1(n4129), .B2(n3870), .ZN(
        n3744) );
  TPOAI21D0BWP12T U4392 ( .A1(n3745), .A2(n3744), .B(n4178), .ZN(n3746) );
  OAI211D0BWP12T U4393 ( .A1(n3861), .A2(n3767), .B(n3875), .C(n3746), .ZN(
        n3747) );
  AOI21D1BWP12T U4394 ( .A1(n3775), .A2(n4301), .B(n3747), .ZN(n4972) );
  ND3D0BWP12T U4395 ( .A1(n3875), .A2(n3905), .A3(n3748), .ZN(n3752) );
  CKND0BWP12T U4396 ( .I(n3749), .ZN(n3751) );
  AOI222D1BWP12T U4397 ( .A1(n3752), .A2(n3844), .B1(n3751), .B2(n3880), .C1(
        n3750), .C2(n4178), .ZN(n4706) );
  MUX2ND0BWP12T U4398 ( .I0(n5118), .I1(n4565), .S(b[0]), .ZN(n4233) );
  MUX2ND0BWP12T U4399 ( .I0(a[18]), .I1(n4788), .S(b[0]), .ZN(n4232) );
  AOI22D0BWP12T U4400 ( .A1(n3855), .A2(n4233), .B1(n4232), .B2(n3854), .ZN(
        n3754) );
  MUX2ND0BWP12T U4401 ( .I0(a[14]), .I1(n4502), .S(b[0]), .ZN(n4221) );
  MUX2ND0BWP12T U4402 ( .I0(n4822), .I1(n4508), .S(b[0]), .ZN(n4234) );
  AOI22D0BWP12T U4403 ( .A1(n3853), .A2(n4221), .B1(n4234), .B2(n3852), .ZN(
        n3753) );
  ND2D1BWP12T U4404 ( .A1(n3754), .A2(n3753), .ZN(n3789) );
  MUX2ND0BWP12T U4405 ( .I0(n5234), .I1(n5079), .S(b[0]), .ZN(n4227) );
  AOI22D1BWP12T U4406 ( .A1(n3853), .A2(n4216), .B1(n4227), .B2(n3855), .ZN(
        n3756) );
  AOI22D1BWP12T U4407 ( .A1(n3852), .A2(n4228), .B1(n4226), .B2(n3854), .ZN(
        n3755) );
  ND2D1BWP12T U4408 ( .A1(n3756), .A2(n3755), .ZN(n3827) );
  INVD1BWP12T U4409 ( .I(n3817), .ZN(n3849) );
  AOI22D0BWP12T U4410 ( .A1(n3855), .A2(n4166), .B1(n4163), .B2(n3854), .ZN(
        n3759) );
  AOI22D0BWP12T U4411 ( .A1(n3853), .A2(n4150), .B1(n3757), .B2(n3852), .ZN(
        n3758) );
  ND2D1BWP12T U4412 ( .A1(n3759), .A2(n3758), .ZN(n3795) );
  OAI22D1BWP12T U4413 ( .A1(n3761), .A2(n3872), .B1(n3760), .B2(n3870), .ZN(
        n3764) );
  NR2D1BWP12T U4414 ( .A1(n3762), .A2(n3871), .ZN(n3763) );
  NR2D1BWP12T U4415 ( .A1(n3764), .A2(n3763), .ZN(n3831) );
  AOI22D1BWP12T U4416 ( .A1(n3853), .A2(n4139), .B1(n4137), .B2(n3852), .ZN(
        n3766) );
  AOI22D1BWP12T U4417 ( .A1(n3855), .A2(n4151), .B1(n4138), .B2(n3854), .ZN(
        n3765) );
  ND2D1BWP12T U4418 ( .A1(n3766), .A2(n3765), .ZN(n3832) );
  CKND2D0BWP12T U4419 ( .A1(n5116), .A2(n4680), .ZN(n3773) );
  NR2XD0BWP12T U4420 ( .A1(n3767), .A2(n4953), .ZN(n3772) );
  INVD0BWP12T U4421 ( .I(n3768), .ZN(n3769) );
  NR2XD0BWP12T U4422 ( .A1(n3769), .A2(n3861), .ZN(n3771) );
  INVD1BWP12T U4423 ( .I(n3777), .ZN(n4860) );
  NR2D0BWP12T U4424 ( .A1(n4860), .A2(n3882), .ZN(n3770) );
  NR4D0BWP12T U4425 ( .A1(n3772), .A2(n3771), .A3(n3849), .A4(n3770), .ZN(
        n4798) );
  NR4D0BWP12T U4426 ( .A1(n4972), .A2(n4706), .A3(n3773), .A4(n4798), .ZN(
        n3826) );
  INVD1BWP12T U4427 ( .I(n3774), .ZN(n5316) );
  ND4D0BWP12T U4428 ( .A1(n5087), .A2(n5316), .A3(n3867), .A4(n3775), .ZN(
        n3798) );
  CKND0BWP12T U4429 ( .I(n3848), .ZN(n3776) );
  CKND2D0BWP12T U4430 ( .A1(n3776), .A2(n3790), .ZN(n3784) );
  ND3D0BWP12T U4431 ( .A1(n3831), .A2(n3778), .A3(n3777), .ZN(n3783) );
  OAI31D0BWP12T U4432 ( .A1(n3784), .A2(n3783), .A3(n4899), .B(n5214), .ZN(
        n3796) );
  MUX2ND0BWP12T U4433 ( .I0(n4649), .I1(n4914), .S(b[0]), .ZN(n4310) );
  AOI22D0BWP12T U4434 ( .A1(n3854), .A2(n4312), .B1(n4310), .B2(n3852), .ZN(
        n3787) );
  MUX2ND0BWP12T U4435 ( .I0(n1), .I1(n2773), .S(b[0]), .ZN(n4308) );
  CKND2D0BWP12T U4436 ( .A1(n4308), .A2(n3855), .ZN(n3786) );
  MUX2ND4BWP12T U4437 ( .I0(n2825), .I1(n4672), .S(b[0]), .ZN(n4314) );
  CKND2D0BWP12T U4438 ( .A1(n4314), .A2(n3853), .ZN(n3785) );
  AOI31D0BWP12T U4439 ( .A1(n3787), .A2(n3786), .A3(n3785), .B(n4953), .ZN(
        n3788) );
  AOI211D0BWP12T U4440 ( .A1(n3880), .A2(n3789), .B(n3788), .C(n3838), .ZN(
        n3792) );
  AOI22D0BWP12T U4441 ( .A1(n4262), .A2(n3827), .B1(n3790), .B2(n4260), .ZN(
        n3791) );
  ND2D1BWP12T U4442 ( .A1(n3792), .A2(n3791), .ZN(n4600) );
  ND4D0BWP12T U4443 ( .A1(n4772), .A2(n3796), .A3(n4600), .A4(n4996), .ZN(
        n3797) );
  AOI21D0BWP12T U4444 ( .A1(n5214), .A2(n3798), .B(n3797), .ZN(n3825) );
  INVD0BWP12T U4445 ( .I(n4232), .ZN(n3835) );
  INVD1BWP12T U4446 ( .I(n4233), .ZN(n4220) );
  OAI22D0BWP12T U4447 ( .A1(n3835), .A2(n3870), .B1(n4220), .B2(n3871), .ZN(
        n3800) );
  INVD1BWP12T U4448 ( .I(n4234), .ZN(n4182) );
  INVD1BWP12T U4449 ( .I(n4314), .ZN(n4237) );
  OAI22D0BWP12T U4450 ( .A1(n4182), .A2(n3869), .B1(n4237), .B2(n3872), .ZN(
        n3799) );
  NR2D1BWP12T U4451 ( .A1(n3800), .A2(n3799), .ZN(n3812) );
  OAI22D0BWP12T U4452 ( .A1(n4899), .A2(n3882), .B1(n3812), .B2(n4953), .ZN(
        n3804) );
  INVD1BWP12T U4453 ( .I(n4226), .ZN(n3818) );
  INVD1BWP12T U4454 ( .I(n4221), .ZN(n4225) );
  OAI22D1BWP12T U4455 ( .A1(n3818), .A2(n3870), .B1(n4225), .B2(n3872), .ZN(
        n3802) );
  INVD1BWP12T U4456 ( .I(n4227), .ZN(n4219) );
  OAI22D1BWP12T U4457 ( .A1(n4215), .A2(n3869), .B1(n4219), .B2(n3871), .ZN(
        n3801) );
  NR2D1BWP12T U4458 ( .A1(n3802), .A2(n3801), .ZN(n3843) );
  NR2D0BWP12T U4459 ( .A1(n3843), .A2(n3905), .ZN(n3803) );
  NR3D1BWP12T U4460 ( .A1(n3804), .A2(n3803), .A3(n3849), .ZN(n4632) );
  NR2D0BWP12T U4461 ( .A1(n3805), .A2(n4632), .ZN(n3824) );
  INVD1BWP12T U4462 ( .I(n4312), .ZN(n4184) );
  INVD1BWP12T U4463 ( .I(n4310), .ZN(n4183) );
  OAI22D0BWP12T U4464 ( .A1(n4184), .A2(n3870), .B1(n4183), .B2(n3869), .ZN(
        n3809) );
  CKND0BWP12T U4465 ( .I(n4308), .ZN(n3807) );
  OAI22D1BWP12T U4466 ( .A1(n3807), .A2(n3871), .B1(n3806), .B2(n4990), .ZN(
        n3808) );
  OAI21D0BWP12T U4467 ( .A1(n3809), .A2(n3808), .B(n4178), .ZN(n3811) );
  ND3D0BWP12T U4468 ( .A1(n3811), .A2(n3875), .A3(n3810), .ZN(n3816) );
  NR2D0BWP12T U4469 ( .A1(n4899), .A2(n3858), .ZN(n3815) );
  NR2XD0BWP12T U4470 ( .A1(n3812), .A2(n3861), .ZN(n3814) );
  TPNR2D0BWP12T U4471 ( .A1(n3843), .A2(n3859), .ZN(n3813) );
  NR4D0BWP12T U4472 ( .A1(n3816), .A2(n3815), .A3(n3814), .A4(n3813), .ZN(
        n5159) );
  IOA21D1BWP12T U4473 ( .A1(n4301), .A2(n4816), .B(n3817), .ZN(n3820) );
  TPOAI22D0BWP12T U4474 ( .A1(n3860), .A2(n3905), .B1(n3862), .B2(n4953), .ZN(
        n3819) );
  NR2D1BWP12T U4475 ( .A1(n3820), .A2(n3819), .ZN(n4828) );
  INVD1BWP12T U4476 ( .I(n3821), .ZN(n5180) );
  CKND2D1BWP12T U4477 ( .A1(n5180), .A2(n3905), .ZN(n3839) );
  NR2D0BWP12T U4478 ( .A1(n3839), .A2(n3844), .ZN(n3822) );
  NR4D0BWP12T U4479 ( .A1(n5159), .A2(n4828), .A3(n3822), .A4(n5232), .ZN(
        n3823) );
  ND4D1BWP12T U4480 ( .A1(n3826), .A2(n3825), .A3(n3824), .A4(n3823), .ZN(
        n3962) );
  INVD1BWP12T U4481 ( .I(n3827), .ZN(n3829) );
  MUX2D1BWP12T U4482 ( .I0(n3829), .I1(n3828), .S(n3948), .Z(n3830) );
  ND2D1BWP12T U4483 ( .A1(n3830), .A2(n5214), .ZN(n5233) );
  INVD1BWP12T U4484 ( .I(n3831), .ZN(n5022) );
  INVD1BWP12T U4485 ( .I(n3832), .ZN(n3833) );
  MUX2D1BWP12T U4486 ( .I0(n5022), .I1(n3833), .S(n3905), .Z(n3834) );
  CKND2D1BWP12T U4487 ( .A1(n3834), .A2(n5214), .ZN(n5057) );
  OAI22D1BWP12T U4488 ( .A1(n3869), .A2(n4227), .B1(n4221), .B2(n3870), .ZN(
        n3868) );
  NR2D0BWP12T U4489 ( .A1(n3868), .A2(n4953), .ZN(n3836) );
  AOI22D1BWP12T U4490 ( .A1(n3855), .A2(n3835), .B1(n4182), .B2(n3854), .ZN(
        n3879) );
  AOI22D0BWP12T U4491 ( .A1(n3880), .A2(n3837), .B1(n3836), .B2(n3879), .ZN(
        n3841) );
  OAI21D0BWP12T U4492 ( .A1(n3839), .A2(n3838), .B(n3844), .ZN(n3840) );
  ND2D1BWP12T U4493 ( .A1(n3841), .A2(n3840), .ZN(n4734) );
  ND4D0BWP12T U4494 ( .A1(n5233), .A2(n3842), .A3(n5057), .A4(n4734), .ZN(
        n3886) );
  INVD0BWP12T U4495 ( .I(n3845), .ZN(n3847) );
  OAI22D0BWP12T U4496 ( .A1(n3847), .A2(n4953), .B1(n3846), .B2(n3905), .ZN(
        n3851) );
  NR2D0BWP12T U4497 ( .A1(n3848), .A2(n3882), .ZN(n3850) );
  NR3D1BWP12T U4498 ( .A1(n3851), .A2(n3850), .A3(n3849), .ZN(n4922) );
  AOI22D0BWP12T U4499 ( .A1(n3853), .A2(n4232), .B1(n4233), .B2(n3852), .ZN(
        n3857) );
  AOI22D0BWP12T U4500 ( .A1(n3855), .A2(n4310), .B1(n4314), .B2(n3854), .ZN(
        n3856) );
  AOI21D0BWP12T U4501 ( .A1(n3857), .A2(n3856), .B(n4953), .ZN(n3866) );
  OAI21D0BWP12T U4502 ( .A1(n4144), .A2(n3858), .B(n3875), .ZN(n3865) );
  TPNR2D0BWP12T U4503 ( .A1(n3860), .A2(n3859), .ZN(n3864) );
  NR2XD0BWP12T U4504 ( .A1(n3862), .A2(n3861), .ZN(n3863) );
  NR4D0BWP12T U4505 ( .A1(n3866), .A2(n3865), .A3(n3864), .A4(n3863), .ZN(
        n4659) );
  NR3D0BWP12T U4506 ( .A1(n5253), .A2(n4922), .A3(n4659), .ZN(n3885) );
  INVD1BWP12T U4507 ( .I(n3867), .ZN(n3883) );
  INVD1BWP12T U4508 ( .I(n3868), .ZN(n3878) );
  OAI22D0BWP12T U4509 ( .A1(n4237), .A2(n3870), .B1(n4220), .B2(n3869), .ZN(
        n3874) );
  RCOAI22D0BWP12T U4510 ( .A1(n4184), .A2(n3872), .B1(n4183), .B2(n3871), .ZN(
        n3873) );
  TPOAI21D0BWP12T U4511 ( .A1(n3874), .A2(n3873), .B(n4178), .ZN(n3876) );
  TPND2D0BWP12T U4512 ( .A1(n3876), .A2(n3875), .ZN(n3877) );
  AOI31D1BWP12T U4513 ( .A1(n3880), .A2(n3879), .A3(n3878), .B(n3877), .ZN(
        n3881) );
  OAI21D1BWP12T U4514 ( .A1(n3883), .A2(n3882), .B(n3881), .ZN(n4939) );
  IND4D0BWP12T U4515 ( .A1(n3886), .B1(n3885), .B2(n4939), .B3(n3884), .ZN(
        n3961) );
  AOI22D0BWP12T U4516 ( .A1(n4920), .A2(n4916), .B1(n4635), .B2(b[22]), .ZN(
        n3894) );
  AOI22D0BWP12T U4517 ( .A1(n26), .A2(n3888), .B1(n3887), .B2(n17), .ZN(n3893)
         );
  AOI22D0BWP12T U4518 ( .A1(n16), .A2(n3890), .B1(n3889), .B2(n25), .ZN(n3892)
         );
  AOI22D0BWP12T U4519 ( .A1(n4826), .A2(n4578), .B1(n4790), .B2(n4794), .ZN(
        n3891) );
  ND4D1BWP12T U4520 ( .A1(n3894), .A2(n3893), .A3(n3892), .A4(n3891), .ZN(
        n3929) );
  AOI22D0BWP12T U4521 ( .A1(n32), .A2(n3895), .B1(n5260), .B2(n5264), .ZN(
        n3904) );
  AOI22D0BWP12T U4522 ( .A1(n5237), .A2(n5235), .B1(n3896), .B2(n5054), .ZN(
        n3903) );
  AOI22D0BWP12T U4523 ( .A1(n5085), .A2(n5081), .B1(n3897), .B2(n3939), .ZN(
        n3902) );
  AOI22D0BWP12T U4524 ( .A1(n3900), .A2(n3937), .B1(n3930), .B2(n3898), .ZN(
        n3901) );
  ND4D1BWP12T U4525 ( .A1(n3904), .A2(n3903), .A3(n3902), .A4(n3901), .ZN(
        n3928) );
  OAI22D0BWP12T U4526 ( .A1(n5192), .A2(n3906), .B1(n3905), .B2(n3661), .ZN(
        n3907) );
  AOI211D0BWP12T U4527 ( .A1(n3908), .A2(n410), .B(n3907), .C(n5290), .ZN(
        n3924) );
  AOI22D0BWP12T U4528 ( .A1(n4896), .A2(n3910), .B1(n3909), .B2(n3938), .ZN(
        n3923) );
  INVD1BWP12T U4529 ( .I(n3911), .ZN(n5032) );
  AOI22D0BWP12T U4530 ( .A1(n5032), .A2(n5033), .B1(n4301), .B2(n3912), .ZN(
        n3922) );
  AOI22D0BWP12T U4531 ( .A1(n22), .A2(n4607), .B1(n407), .B2(n31), .ZN(n3919)
         );
  AOI22D0BWP12T U4532 ( .A1(n21), .A2(n3914), .B1(n7), .B2(n4944), .ZN(n3918)
         );
  AOI22D0BWP12T U4533 ( .A1(n4655), .A2(n4651), .B1(n3915), .B2(n4977), .ZN(
        n3917) );
  ND4D1BWP12T U4534 ( .A1(n3919), .A2(n3918), .A3(n3917), .A4(n3916), .ZN(
        n3920) );
  NR2D0BWP12T U4535 ( .A1(n3920), .A2(n5106), .ZN(n3921) );
  ND4D1BWP12T U4536 ( .A1(n3924), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(
        n3927) );
  ND2D1BWP12T U4537 ( .A1(n3936), .A2(n3925), .ZN(n3926) );
  OAI31D1BWP12T U4538 ( .A1(n3929), .A2(n3928), .A3(n3927), .B(n3926), .ZN(
        n3959) );
  AOI22D0BWP12T U4539 ( .A1(n4565), .A2(n16), .B1(n4826), .B2(n448), .ZN(n3934) );
  AOI22D0BWP12T U4540 ( .A1(n4788), .A2(n4794), .B1(n5237), .B2(n5234), .ZN(
        n3933) );
  AOI22D0BWP12T U4541 ( .A1(n402), .A2(n480), .B1(n32), .B2(n4508), .ZN(n3932)
         );
  AOI22D0BWP12T U4542 ( .A1(n4990), .A2(n31), .B1(n3930), .B2(n4511), .ZN(
        n3931) );
  ND4D1BWP12T U4543 ( .A1(n3934), .A2(n3933), .A3(n3932), .A4(n3931), .ZN(
        n3956) );
  AOI21D1BWP12T U4544 ( .A1(n25), .A2(a[18]), .B(n5294), .ZN(n3935) );
  CKND2D1BWP12T U4545 ( .A1(n3935), .A2(n4422), .ZN(n3943) );
  AOI22D0BWP12T U4546 ( .A1(n5108), .A2(n3936), .B1(n5085), .B2(n5079), .ZN(
        n3942) );
  AOI22D0BWP12T U4547 ( .A1(n5049), .A2(n5054), .B1(n3937), .B2(n4509), .ZN(
        n3941) );
  AOI22D0BWP12T U4548 ( .A1(n4518), .A2(n3939), .B1(n3938), .B2(n4510), .ZN(
        n3940) );
  IND4D1BWP12T U4549 ( .A1(n3943), .B1(n3942), .B2(n3941), .B3(n3940), .ZN(
        n3955) );
  AOI22D1BWP12T U4550 ( .A1(n5146), .A2(n5153), .B1(n21), .B2(n2773), .ZN(
        n3947) );
  AOI22D0BWP12T U4551 ( .A1(n2825), .A2(b[22]), .B1(n22), .B2(n1), .ZN(n3946)
         );
  AOI22D0BWP12T U4552 ( .A1(n5118), .A2(n26), .B1(n4920), .B2(n4914), .ZN(
        n3945) );
  AOI22D0BWP12T U4553 ( .A1(n4672), .A2(n17), .B1(n4977), .B2(n4568), .ZN(
        n3944) );
  ND4D1BWP12T U4554 ( .A1(n3947), .A2(n3946), .A3(n3945), .A4(n3944), .ZN(
        n3954) );
  AOI22D0BWP12T U4555 ( .A1(n4943), .A2(n4944), .B1(n5033), .B2(n5030), .ZN(
        n3952) );
  AOI22D0BWP12T U4556 ( .A1(n3948), .A2(n436), .B1(n4655), .B2(n4649), .ZN(
        n3951) );
  AOI22D0BWP12T U4557 ( .A1(n4849), .A2(n4501), .B1(n4301), .B2(n4541), .ZN(
        n3950) );
  AOI22D0BWP12T U4558 ( .A1(n5256), .A2(n5264), .B1(n5196), .B2(n5192), .ZN(
        n3949) );
  ND4D1BWP12T U4559 ( .A1(n3952), .A2(n3951), .A3(n3950), .A4(n3949), .ZN(
        n3953) );
  NR4D0BWP12T U4560 ( .A1(n3956), .A2(n3955), .A3(n3954), .A4(n3953), .ZN(
        n3957) );
  AOI21D1BWP12T U4561 ( .A1(n3959), .A2(n3958), .B(n3957), .ZN(n3960) );
  OAI21D1BWP12T U4562 ( .A1(n3962), .A2(n3961), .B(n3960), .ZN(n3963) );
  AOI21D1BWP12T U4563 ( .A1(n3965), .A2(n3964), .B(n3963), .ZN(n4127) );
  INVD1BWP12T U4564 ( .I(n3972), .ZN(n3967) );
  CKND2D1BWP12T U4565 ( .A1(n3985), .A2(n3967), .ZN(n3969) );
  INVD1BWP12T U4566 ( .I(n3975), .ZN(n3966) );
  AOI21D1BWP12T U4567 ( .A1(n3988), .A2(n3967), .B(n3966), .ZN(n3968) );
  OAI21D1BWP12T U4568 ( .A1(n4116), .A2(n3969), .B(n3968), .ZN(n3971) );
  TPND2D0BWP12T U4569 ( .A1(n3970), .A2(n3973), .ZN(n4466) );
  XNR2D1BWP12T U4570 ( .A1(n3971), .A2(n4466), .ZN(n4598) );
  NR2D0BWP12T U4571 ( .A1(n3972), .A2(n3974), .ZN(n3977) );
  TPND2D0BWP12T U4572 ( .A1(n3985), .A2(n3977), .ZN(n3979) );
  OAI21D0BWP12T U4573 ( .A1(n3975), .A2(n3974), .B(n3973), .ZN(n3976) );
  TPAOI21D0BWP12T U4574 ( .A1(n3988), .A2(n3977), .B(n3976), .ZN(n3978) );
  OAI21D1BWP12T U4575 ( .A1(n4116), .A2(n3979), .B(n3978), .ZN(n3981) );
  ND2D1BWP12T U4576 ( .A1(n3980), .A2(n4480), .ZN(n4473) );
  XNR2D1BWP12T U4577 ( .A1(n3981), .A2(n4473), .ZN(n5000) );
  CKND2D1BWP12T U4578 ( .A1(n3983), .A2(n3982), .ZN(n4457) );
  NR4D0BWP12T U4579 ( .A1(n3984), .A2(n4598), .A3(n5000), .A4(n4952), .ZN(
        n4125) );
  TPND2D0BWP12T U4580 ( .A1(n3985), .A2(n3987), .ZN(n3990) );
  TPAOI21D0BWP12T U4581 ( .A1(n3988), .A2(n3987), .B(n3986), .ZN(n3989) );
  OAI21D1BWP12T U4582 ( .A1(n4116), .A2(n3990), .B(n3989), .ZN(n3993) );
  CKND2D1BWP12T U4583 ( .A1(n3992), .A2(n3991), .ZN(n4492) );
  XNR2D1BWP12T U4584 ( .A1(n3993), .A2(n4492), .ZN(n5172) );
  CKND0BWP12T U4585 ( .I(n3998), .ZN(n3995) );
  INVD1BWP12T U4586 ( .I(n4002), .ZN(n3994) );
  OAI21D1BWP12T U4587 ( .A1(n4116), .A2(n3995), .B(n3994), .ZN(n3997) );
  INVD1BWP12T U4588 ( .I(n3996), .ZN(n4001) );
  CKND2D1BWP12T U4589 ( .A1(n4001), .A2(n3999), .ZN(n4338) );
  XNR2D1BWP12T U4590 ( .A1(n3997), .A2(n4338), .ZN(n4744) );
  CKND2D0BWP12T U4591 ( .A1(n3998), .A2(n4001), .ZN(n4004) );
  CKND0BWP12T U4592 ( .I(n3999), .ZN(n4000) );
  TPAOI21D0BWP12T U4593 ( .A1(n4002), .A2(n4001), .B(n4000), .ZN(n4003) );
  OAI21D1BWP12T U4594 ( .A1(n4116), .A2(n4004), .B(n4003), .ZN(n4007) );
  CKND0BWP12T U4595 ( .I(n4005), .ZN(n4006) );
  CKND2D1BWP12T U4596 ( .A1(n4006), .A2(n4342), .ZN(n4340) );
  XNR2D1BWP12T U4597 ( .A1(n4007), .A2(n4340), .ZN(n4712) );
  OAI21D1BWP12T U4598 ( .A1(n4116), .A2(n4010), .B(n4011), .ZN(n4009) );
  INVD1BWP12T U4599 ( .I(n4008), .ZN(n4013) );
  CKND2D1BWP12T U4600 ( .A1(n4013), .A2(n4012), .ZN(n4347) );
  XNR2D1BWP12T U4601 ( .A1(n4009), .A2(n4347), .ZN(n5134) );
  INVD1BWP12T U4602 ( .I(n4010), .ZN(n4103) );
  INVD1BWP12T U4603 ( .I(n4011), .ZN(n4112) );
  OR4D0BWP12T U4604 ( .A1(n4744), .A2(n4712), .A3(n5134), .A4(n4686), .Z(n4035) );
  CKND1BWP12T U4605 ( .I(n4095), .ZN(n4024) );
  INVD1BWP12T U4606 ( .I(n4387), .ZN(n4097) );
  ND2XD0BWP12T U4607 ( .A1(n4024), .A2(n4097), .ZN(n4016) );
  CKND1BWP12T U4608 ( .I(n4094), .ZN(n4028) );
  INVD0BWP12T U4609 ( .I(n4388), .ZN(n4014) );
  AOI21D1BWP12T U4610 ( .A1(n4028), .A2(n4097), .B(n4014), .ZN(n4015) );
  OAI21D1BWP12T U4611 ( .A1(n4096), .A2(n4016), .B(n4015), .ZN(n4018) );
  INVD1BWP12T U4612 ( .I(n4406), .ZN(n4017) );
  CKND2D1BWP12T U4613 ( .A1(n4017), .A2(n4405), .ZN(n4400) );
  XNR2XD1BWP12T U4614 ( .A1(n4018), .A2(n4400), .ZN(n5045) );
  CKND2D0BWP12T U4615 ( .A1(n4024), .A2(n4023), .ZN(n4020) );
  AOI21D0BWP12T U4616 ( .A1(n4028), .A2(n4023), .B(n4025), .ZN(n4019) );
  OAI21D1BWP12T U4617 ( .A1(n4096), .A2(n4020), .B(n4019), .ZN(n4022) );
  INVD1BWP12T U4618 ( .I(n4027), .ZN(n4021) );
  CKND2D1BWP12T U4619 ( .A1(n4021), .A2(n4026), .ZN(n4409) );
  XNR2XD1BWP12T U4620 ( .A1(n4022), .A2(n4409), .ZN(n5278) );
  INVD1BWP12T U4621 ( .I(n4029), .ZN(n4395) );
  CKND2D1BWP12T U4622 ( .A1(n4395), .A2(n4393), .ZN(n4449) );
  OAI21D1BWP12T U4623 ( .A1(n4116), .A2(n4061), .B(n4062), .ZN(n4033) );
  CKND0BWP12T U4624 ( .I(n4030), .ZN(n4329) );
  CKND2D0BWP12T U4625 ( .A1(n4329), .A2(n4031), .ZN(n4032) );
  XNR2D1BWP12T U4626 ( .A1(n4033), .A2(n4032), .ZN(n4805) );
  OR4D1BWP12T U4627 ( .A1(n5045), .A2(n5278), .A3(n4761), .A4(n4805), .Z(n4034) );
  NR4D0BWP12T U4628 ( .A1(n5172), .A2(n4036), .A3(n4035), .A4(n4034), .ZN(
        n4124) );
  INVD1BWP12T U4629 ( .I(n4069), .ZN(n4102) );
  NR2XD0BWP12T U4630 ( .A1(n4102), .A2(n4100), .ZN(n4038) );
  CKND2D0BWP12T U4631 ( .A1(n4038), .A2(n4103), .ZN(n4040) );
  INVD1BWP12T U4632 ( .I(n4068), .ZN(n4109) );
  OAI21D0BWP12T U4633 ( .A1(n4109), .A2(n4100), .B(n4104), .ZN(n4037) );
  AOI21D1BWP12T U4634 ( .A1(n4112), .A2(n4038), .B(n4037), .ZN(n4039) );
  OAI21D1BWP12T U4635 ( .A1(n4116), .A2(n4040), .B(n4039), .ZN(n4042) );
  CKND2D1BWP12T U4636 ( .A1(n4106), .A2(n4374), .ZN(n4041) );
  XNR2D1BWP12T U4637 ( .A1(n4042), .A2(n4041), .ZN(n4662) );
  CKND0BWP12T U4638 ( .I(n4046), .ZN(n4047) );
  AOI21D1BWP12T U4639 ( .A1(n4050), .A2(n4049), .B(n4048), .ZN(n4053) );
  CKND0BWP12T U4640 ( .I(n4051), .ZN(n4423) );
  CKND2D1BWP12T U4641 ( .A1(n4423), .A2(n4422), .ZN(n4052) );
  XOR2XD1BWP12T U4642 ( .A1(n4053), .A2(n4052), .Z(n4880) );
  NR4D0BWP12T U4643 ( .A1(n5011), .A2(n4055), .A3(n4880), .A4(n4054), .ZN(
        n4067) );
  INVD1BWP12T U4644 ( .I(n4056), .ZN(n4430) );
  INVD1BWP12T U4645 ( .I(n4058), .ZN(n4434) );
  OR2XD0BWP12T U4646 ( .A1(n480), .A2(n3016), .Z(n4060) );
  AN2XD1BWP12T U4647 ( .A1(n4060), .A2(n4059), .Z(n5304) );
  NR4D0BWP12T U4648 ( .A1(n5198), .A2(n4844), .A3(n5304), .A4(n4970), .ZN(
        n4065) );
  XOR2XD1BWP12T U4649 ( .A1(n4116), .A2(n4396), .Z(n4818) );
  INR4D0BWP12T U4650 ( .A1(n4065), .B1(n4064), .B2(n4063), .B3(n4818), .ZN(
        n4066) );
  IND3D1BWP12T U4651 ( .A1(n4662), .B1(n4067), .B2(n4066), .ZN(n4083) );
  CKND2D0BWP12T U4652 ( .A1(n4103), .A2(n4069), .ZN(n4071) );
  AOI21D0BWP12T U4653 ( .A1(n4112), .A2(n4069), .B(n4068), .ZN(n4070) );
  OAI21D1BWP12T U4654 ( .A1(n4116), .A2(n4071), .B(n4070), .ZN(n4074) );
  TPND2D0BWP12T U4655 ( .A1(n4072), .A2(n4361), .ZN(n4073) );
  XNR2D1BWP12T U4656 ( .A1(n4074), .A2(n4073), .ZN(n4630) );
  NR2D1BWP12T U4657 ( .A1(n4102), .A2(n4075), .ZN(n4077) );
  CKND2D1BWP12T U4658 ( .A1(n4077), .A2(n4103), .ZN(n4079) );
  OAI21D1BWP12T U4659 ( .A1(n4109), .A2(n4075), .B(n4361), .ZN(n4076) );
  AOI21D1BWP12T U4660 ( .A1(n4112), .A2(n4077), .B(n4076), .ZN(n4078) );
  OAI21D1BWP12T U4661 ( .A1(n4116), .A2(n4079), .B(n4078), .ZN(n4082) );
  ND2D1BWP12T U4662 ( .A1(n4366), .A2(n4080), .ZN(n4081) );
  XNR2D1BWP12T U4663 ( .A1(n4082), .A2(n4081), .ZN(n4929) );
  NR3XD0BWP12T U4664 ( .A1(n4083), .A2(n4630), .A3(n4929), .ZN(n4123) );
  TPND2D0BWP12T U4665 ( .A1(n4084), .A2(n4087), .ZN(n4090) );
  INVD0BWP12T U4666 ( .I(n4085), .ZN(n4086) );
  TPAOI21D0BWP12T U4667 ( .A1(n4088), .A2(n4087), .B(n4086), .ZN(n4089) );
  OAI21D1BWP12T U4668 ( .A1(n4096), .A2(n4090), .B(n4089), .ZN(n4093) );
  CKND2D1BWP12T U4669 ( .A1(n4384), .A2(n4382), .ZN(n4092) );
  XNR2XD1BWP12T U4670 ( .A1(n4093), .A2(n4092), .ZN(n5077) );
  OR4D1BWP12T U4671 ( .A1(n4099), .A2(n4098), .A3(n5077), .A4(n5242), .Z(n4121) );
  INVD0BWP12T U4672 ( .I(n4100), .ZN(n4101) );
  ND2D1BWP12T U4673 ( .A1(n4101), .A2(n4106), .ZN(n4110) );
  NR2D1BWP12T U4674 ( .A1(n4110), .A2(n4102), .ZN(n4113) );
  CKND2D1BWP12T U4675 ( .A1(n4113), .A2(n4103), .ZN(n4115) );
  INVD0BWP12T U4676 ( .I(n4104), .ZN(n4107) );
  TPAOI21D0BWP12T U4677 ( .A1(n4107), .A2(n4106), .B(n4105), .ZN(n4108) );
  OAI21D1BWP12T U4678 ( .A1(n4110), .A2(n4109), .B(n4108), .ZN(n4111) );
  AOI21D1BWP12T U4679 ( .A1(n4113), .A2(n4112), .B(n4111), .ZN(n4114) );
  OAI21D1BWP12T U4680 ( .A1(n4116), .A2(n4115), .B(n4114), .ZN(n4120) );
  ND2D1BWP12T U4681 ( .A1(n4118), .A2(n4117), .ZN(n4119) );
  XNR2D1BWP12T U4682 ( .A1(n4120), .A2(n4119), .ZN(n4971) );
  NR2D0BWP12T U4683 ( .A1(n4121), .A2(n4971), .ZN(n4122) );
  ND4D1BWP12T U4684 ( .A1(n4125), .A2(n4124), .A3(n4123), .A4(n4122), .ZN(
        n4126) );
  AOI22D1BWP12T U4685 ( .A1(n4242), .A2(n4133), .B1(n4132), .B2(n4245), .ZN(
        n4136) );
  CKND2D1BWP12T U4686 ( .A1(n2839), .A2(n4134), .ZN(n4135) );
  ND2D1BWP12T U4687 ( .A1(n4136), .A2(n4135), .ZN(n5019) );
  INVD1BWP12T U4688 ( .I(n5019), .ZN(n4275) );
  INVD1BWP12T U4689 ( .I(n4253), .ZN(n4278) );
  ND2D1BWP12T U4690 ( .A1(n5162), .A2(n4185), .ZN(n4298) );
  ND3XD0BWP12T U4691 ( .A1(n4814), .A2(n4299), .A3(n4277), .ZN(n4149) );
  CKND2D0BWP12T U4692 ( .A1(n4242), .A2(n4233), .ZN(n4143) );
  AOI22D0BWP12T U4693 ( .A1(n4245), .A2(n4314), .B1(n4244), .B2(n4232), .ZN(
        n4142) );
  CKND2D0BWP12T U4694 ( .A1(n2839), .A2(n4310), .ZN(n4141) );
  TPAOI31D0BWP12T U4695 ( .A1(n4143), .A2(n4142), .A3(n4141), .B(n5183), .ZN(
        n4146) );
  OAI21D0BWP12T U4696 ( .A1(n5162), .A2(n4144), .B(n4185), .ZN(n4145) );
  NR2D1BWP12T U4697 ( .A1(n4146), .A2(n4145), .ZN(n4148) );
  ND2XD0BWP12T U4698 ( .A1(n4813), .A2(n4267), .ZN(n4147) );
  ND3D1BWP12T U4699 ( .A1(n4149), .A2(n4148), .A3(n4147), .ZN(n4646) );
  OAI22D1BWP12T U4700 ( .A1(n4311), .A2(n4151), .B1(n4150), .B2(n4313), .ZN(
        n4161) );
  INVD0BWP12T U4701 ( .I(n4161), .ZN(n4154) );
  AOI22D1BWP12T U4702 ( .A1(n2839), .A2(n4153), .B1(n4244), .B2(n4152), .ZN(
        n4160) );
  TPAOI21D0BWP12T U4703 ( .A1(n4154), .A2(n4160), .B(n5183), .ZN(n4157) );
  CKND0BWP12T U4704 ( .I(n4207), .ZN(n4155) );
  TPNR2D0BWP12T U4705 ( .A1(n4817), .A2(n4155), .ZN(n4156) );
  AOI211D1BWP12T U4706 ( .A1(n4158), .A2(n4267), .B(n4157), .C(n4156), .ZN(
        n4803) );
  ND4D0BWP12T U4707 ( .A1(n4684), .A2(n4646), .A3(n4159), .A4(n4803), .ZN(
        n4259) );
  CKND2D0BWP12T U4708 ( .A1(n4160), .A2(n4267), .ZN(n4162) );
  NR2XD0BWP12T U4709 ( .A1(n4162), .A2(n4161), .ZN(n4172) );
  AOI22D0BWP12T U4710 ( .A1(n4245), .A2(n4164), .B1(n4244), .B2(n4163), .ZN(
        n4169) );
  CKND2D0BWP12T U4711 ( .A1(n2839), .A2(n4165), .ZN(n4168) );
  CKND2D0BWP12T U4712 ( .A1(n4242), .A2(n4166), .ZN(n4167) );
  TPAOI31D0BWP12T U4713 ( .A1(n4169), .A2(n4168), .A3(n4167), .B(n5183), .ZN(
        n4171) );
  NR3XD0BWP12T U4714 ( .A1(n4172), .A2(n4171), .A3(n4170), .ZN(n4173) );
  OAI21D1BWP12T U4715 ( .A1(n4174), .A2(n4281), .B(n4173), .ZN(n4181) );
  MUX2ND0BWP12T U4716 ( .I0(n4177), .I1(n4176), .S(n4175), .ZN(n4179) );
  CKND2D1BWP12T U4717 ( .A1(n4179), .A2(n4178), .ZN(n4180) );
  ND2D1BWP12T U4718 ( .A1(n4181), .A2(n4180), .ZN(n4982) );
  NR3D0BWP12T U4719 ( .A1(n4982), .A2(n4956), .A3(n4186), .ZN(n4258) );
  INR2D1BWP12T U4720 ( .A1(n4208), .B1(n4187), .ZN(n4188) );
  AOI21D0BWP12T U4721 ( .A1(n4189), .A2(n4297), .B(n4188), .ZN(n4191) );
  AOI21D0BWP12T U4722 ( .A1(n4202), .A2(n4299), .B(n4298), .ZN(n4190) );
  CKND2D1BWP12T U4723 ( .A1(n4191), .A2(n4190), .ZN(n4708) );
  AOI22D1BWP12T U4724 ( .A1(n4192), .A2(n4208), .B1(n4266), .B2(n4297), .ZN(
        n4194) );
  TPAOI21D0BWP12T U4725 ( .A1(n4203), .A2(n4299), .B(n4298), .ZN(n4193) );
  ND2D1BWP12T U4726 ( .A1(n4194), .A2(n4193), .ZN(n4913) );
  ND4D0BWP12T U4727 ( .A1(n4708), .A2(n5071), .A3(n4195), .A4(n4913), .ZN(
        n4214) );
  INVD1BWP12T U4728 ( .I(n4196), .ZN(n5034) );
  INVD0BWP12T U4729 ( .I(n4197), .ZN(n4206) );
  IND3D0BWP12T U4730 ( .A1(n5312), .B1(n4202), .B2(n5163), .ZN(n4204) );
  CKND0BWP12T U4731 ( .I(n4203), .ZN(n4268) );
  NR3D0BWP12T U4732 ( .A1(n4204), .A2(n4268), .A3(n5019), .ZN(n4205) );
  OAI211D0BWP12T U4733 ( .A1(n5008), .A2(n5034), .B(n4206), .C(n4205), .ZN(
        n4213) );
  AOI22D1BWP12T U4734 ( .A1(n4209), .A2(n4301), .B1(n4208), .B2(n4207), .ZN(
        n4871) );
  CKND0BWP12T U4735 ( .I(n5320), .ZN(n4211) );
  INVD0BWP12T U4736 ( .I(n4210), .ZN(n5311) );
  ND4D0BWP12T U4737 ( .A1(n4871), .A2(n4211), .A3(n4954), .A4(n5311), .ZN(
        n4212) );
  TPNR3D0BWP12T U4738 ( .A1(n4214), .A2(n4213), .A3(n4212), .ZN(n4257) );
  INR2D1BWP12T U4739 ( .A1(n4215), .B1(n4311), .ZN(n4218) );
  OAI22D1BWP12T U4740 ( .A1(n4315), .A2(n4216), .B1(n4313), .B2(n4226), .ZN(
        n4217) );
  AOI211XD1BWP12T U4741 ( .A1(n2839), .A2(n4219), .B(n4218), .C(n4217), .ZN(
        n4307) );
  INR2D0BWP12T U4742 ( .A1(n4220), .B1(n4309), .ZN(n4224) );
  TPNR2D0BWP12T U4743 ( .A1(n4311), .A2(n4234), .ZN(n4223) );
  OAI22D0BWP12T U4744 ( .A1(n4315), .A2(n4221), .B1(n4313), .B2(n4232), .ZN(
        n4222) );
  NR3D1BWP12T U4745 ( .A1(n4224), .A2(n4223), .A3(n4222), .ZN(n4306) );
  INR2D0BWP12T U4746 ( .A1(n4225), .B1(n4309), .ZN(n4231) );
  NR2D1BWP12T U4747 ( .A1(n4311), .A2(n4226), .ZN(n4230) );
  OAI22D1BWP12T U4748 ( .A1(n4315), .A2(n4228), .B1(n4313), .B2(n4227), .ZN(
        n4229) );
  NR3D1BWP12T U4749 ( .A1(n4231), .A2(n4230), .A3(n4229), .ZN(n4271) );
  TPNR2D0BWP12T U4750 ( .A1(n4311), .A2(n4232), .ZN(n4236) );
  OAI22D0BWP12T U4751 ( .A1(n4315), .A2(n4234), .B1(n4313), .B2(n4233), .ZN(
        n4235) );
  AOI211XD0BWP12T U4752 ( .A1(n2839), .A2(n4237), .B(n4236), .C(n4235), .ZN(
        n4238) );
  OAI222D1BWP12T U4753 ( .A1(n4817), .A2(n5163), .B1(n4815), .B2(n4271), .C1(
        n5183), .C2(n4238), .ZN(n4637) );
  CKND0BWP12T U4754 ( .I(n5162), .ZN(n4240) );
  RCAOI22D0BWP12T U4755 ( .A1(n4240), .A2(n5019), .B1(n4239), .B2(n4267), .ZN(
        n4255) );
  CKND0BWP12T U4756 ( .I(n4817), .ZN(n4252) );
  CKND2D0BWP12T U4757 ( .A1(n4242), .A2(n4241), .ZN(n4250) );
  AOI22D0BWP12T U4758 ( .A1(n4246), .A2(n4245), .B1(n4244), .B2(n4243), .ZN(
        n4249) );
  TPND2D0BWP12T U4759 ( .A1(n2839), .A2(n4247), .ZN(n4248) );
  TPAOI31D0BWP12T U4760 ( .A1(n4250), .A2(n4249), .A3(n4248), .B(n5183), .ZN(
        n4251) );
  RCAOI21D0BWP12T U4761 ( .A1(n4253), .A2(n4252), .B(n4251), .ZN(n4254) );
  CKND2D1BWP12T U4762 ( .A1(n4255), .A2(n4254), .ZN(n4998) );
  NR4D0BWP12T U4763 ( .A1(n5130), .A2(n4637), .A3(n5165), .A4(n4998), .ZN(
        n4256) );
  IND4D1BWP12T U4764 ( .A1(n4259), .B1(n4258), .B2(n4257), .B3(n4256), .ZN(
        n4328) );
  CKND2D2BWP12T U4765 ( .A1(n4954), .A2(n4260), .ZN(n5185) );
  INVD0BWP12T U4766 ( .I(n4261), .ZN(n4263) );
  CKND2D1BWP12T U4767 ( .A1(n4263), .A2(n4262), .ZN(n5186) );
  AN2XD0BWP12T U4768 ( .A1(n5185), .A2(n5186), .Z(n4265) );
  INVD1BWP12T U4769 ( .I(n5211), .ZN(n5184) );
  CKND0BWP12T U4770 ( .I(n5182), .ZN(n4264) );
  AOI21D0BWP12T U4771 ( .A1(n4265), .A2(n5184), .B(n4264), .ZN(n4269) );
  OAI211D0BWP12T U4772 ( .A1(n4301), .A2(n4270), .B(n4269), .C(n4766), .ZN(
        n4272) );
  INR3XD0BWP12T U4773 ( .A1(n4273), .B1(n4272), .B2(n5280), .ZN(n4284) );
  CKND2D1BWP12T U4774 ( .A1(n4275), .A2(n4274), .ZN(n4280) );
  INVD0BWP12T U4775 ( .I(n4281), .ZN(n4276) );
  TPAOI21D0BWP12T U4776 ( .A1(n4278), .A2(n4277), .B(n4276), .ZN(n4279) );
  AOI21D1BWP12T U4777 ( .A1(n4280), .A2(n4279), .B(n5048), .ZN(n5047) );
  MUX2NXD0BWP12T U4778 ( .I0(n4307), .I1(n4319), .S(n4297), .ZN(n4282) );
  ND4D0BWP12T U4779 ( .A1(n4284), .A2(n4283), .A3(n5047), .A4(n5227), .ZN(
        n4327) );
  CKND0BWP12T U4780 ( .I(n4710), .ZN(n4286) );
  NR2D0BWP12T U4781 ( .A1(n4286), .A2(n4285), .ZN(n4293) );
  ND4D0BWP12T U4782 ( .A1(n4288), .A2(n4861), .A3(n4287), .A4(n4819), .ZN(
        n4290) );
  INR3XD0BWP12T U4783 ( .A1(n4795), .B1(n4290), .B2(n4289), .ZN(n4292) );
  AOI31D0BWP12T U4784 ( .A1(n4293), .A2(n4292), .A3(n4291), .B(n4301), .ZN(
        n4326) );
  INVD1BWP12T U4785 ( .I(n4294), .ZN(n4295) );
  AOI22D1BWP12T U4786 ( .A1(n4297), .A2(n4296), .B1(n4295), .B2(n4208), .ZN(
        n4305) );
  AOI21D0BWP12T U4787 ( .A1(n4299), .A2(n5182), .B(n4298), .ZN(n4304) );
  INVD1BWP12T U4788 ( .I(n4300), .ZN(n4303) );
  OAI21D0BWP12T U4789 ( .A1(n4954), .A2(n4301), .B(n4953), .ZN(n4302) );
  AOI22D1BWP12T U4790 ( .A1(n4305), .A2(n4304), .B1(n4303), .B2(n4302), .ZN(
        n4739) );
  OAI22D0BWP12T U4791 ( .A1(n4307), .A2(n4817), .B1(n4306), .B2(n4815), .ZN(
        n4322) );
  NR2D0BWP12T U4792 ( .A1(n4309), .A2(n4308), .ZN(n4318) );
  NR2D0BWP12T U4793 ( .A1(n4311), .A2(n4310), .ZN(n4317) );
  OAI22D0BWP12T U4794 ( .A1(n4315), .A2(n4314), .B1(n4313), .B2(n4312), .ZN(
        n4316) );
  NR3XD0BWP12T U4795 ( .A1(n4318), .A2(n4317), .A3(n4316), .ZN(n4320) );
  OAI22D0BWP12T U4796 ( .A1(n4320), .A2(n5183), .B1(n4319), .B2(n5162), .ZN(
        n4321) );
  NR2D1BWP12T U4797 ( .A1(n4322), .A2(n4321), .ZN(n4605) );
  IND4D0BWP12T U4798 ( .A1(n4324), .B1(n4323), .B2(n4739), .B3(n4605), .ZN(
        n4325) );
  NR4D0BWP12T U4799 ( .A1(n4328), .A2(n4327), .A3(n4326), .A4(n4325), .ZN(
        n4592) );
  CKND0BWP12T U4800 ( .I(n4330), .ZN(n4331) );
  NR2D0BWP12T U4801 ( .A1(n4331), .A2(n4334), .ZN(n4337) );
  CKND0BWP12T U4802 ( .I(n4332), .ZN(n4335) );
  OAI21D0BWP12T U4803 ( .A1(n4335), .A2(n4334), .B(n4333), .ZN(n4336) );
  AOI21D1BWP12T U4804 ( .A1(n4491), .A2(n4337), .B(n4336), .ZN(n4339) );
  XOR2XD1BWP12T U4805 ( .A1(n4339), .A2(n4338), .Z(n4727) );
  INVD1BWP12T U4806 ( .I(n4341), .ZN(n4349) );
  INVD1BWP12T U4807 ( .I(n4344), .ZN(n4352) );
  TPNR2D0BWP12T U4808 ( .A1(n4341), .A2(n4343), .ZN(n4346) );
  OAI21D1BWP12T U4809 ( .A1(n4344), .A2(n4343), .B(n4342), .ZN(n4345) );
  AOI21D1BWP12T U4810 ( .A1(n4491), .A2(n4346), .B(n4345), .ZN(n4348) );
  XOR2XD1BWP12T U4811 ( .A1(n4348), .A2(n4347), .Z(n5114) );
  NR4D0BWP12T U4812 ( .A1(n4787), .A2(n4727), .A3(n4694), .A4(n5114), .ZN(
        n4448) );
  CKND2D1BWP12T U4813 ( .A1(n4349), .A2(n4351), .ZN(n4354) );
  AOI21D1BWP12T U4814 ( .A1(n4352), .A2(n4351), .B(n4350), .ZN(n4357) );
  NR2D0BWP12T U4815 ( .A1(n4354), .A2(n4356), .ZN(n4359) );
  TPOAI21D0BWP12T U4816 ( .A1(n4357), .A2(n4356), .B(n4355), .ZN(n4358) );
  AOI21D1BWP12T U4817 ( .A1(n4491), .A2(n4359), .B(n4358), .ZN(n4363) );
  CKND2D1BWP12T U4818 ( .A1(n4072), .A2(n4361), .ZN(n4362) );
  XOR2XD1BWP12T U4819 ( .A1(n4363), .A2(n4362), .Z(n4631) );
  AOI21D1BWP12T U4820 ( .A1(n4491), .A2(n4365), .B(n4364), .ZN(n4368) );
  ND2D1BWP12T U4821 ( .A1(n4366), .A2(n4369), .ZN(n4367) );
  XOR2XD1BWP12T U4822 ( .A1(n4368), .A2(n4367), .Z(n4930) );
  NR2D0BWP12T U4823 ( .A1(n4478), .A2(n4370), .ZN(n4372) );
  TPOAI21D0BWP12T U4824 ( .A1(n4488), .A2(n4370), .B(n4369), .ZN(n4371) );
  AOI21D1BWP12T U4825 ( .A1(n4491), .A2(n4372), .B(n4371), .ZN(n4376) );
  CKND2D1BWP12T U4826 ( .A1(n4106), .A2(n4374), .ZN(n4375) );
  XOR2XD1BWP12T U4827 ( .A1(n4376), .A2(n4375), .Z(n4663) );
  NR4D0BWP12T U4828 ( .A1(n4670), .A2(n4631), .A3(n4930), .A4(n4663), .ZN(
        n4447) );
  OAI21D1BWP12T U4829 ( .A1(n4408), .A2(n4380), .B(n4381), .ZN(n4379) );
  INVD1BWP12T U4830 ( .I(n4377), .ZN(n4384) );
  CKND2D1BWP12T U4831 ( .A1(n4384), .A2(n4382), .ZN(n4378) );
  XNR2XD1BWP12T U4832 ( .A1(n4379), .A2(n4378), .ZN(n5092) );
  INVD1BWP12T U4833 ( .I(n4380), .ZN(n4403) );
  TPND2D0BWP12T U4834 ( .A1(n4403), .A2(n4384), .ZN(n4386) );
  INVD1BWP12T U4835 ( .I(n4381), .ZN(n4407) );
  INVD1BWP12T U4836 ( .I(n4382), .ZN(n4383) );
  AOI21D1BWP12T U4837 ( .A1(n4407), .A2(n4384), .B(n4383), .ZN(n4385) );
  OAI21D1BWP12T U4838 ( .A1(n4408), .A2(n4386), .B(n4385), .ZN(n4390) );
  CKND2D1BWP12T U4839 ( .A1(n4097), .A2(n4388), .ZN(n4389) );
  XNR2XD1BWP12T U4840 ( .A1(n4390), .A2(n4389), .ZN(n5229) );
  NR4D0BWP12T U4841 ( .A1(n4392), .A2(n4391), .A3(n5092), .A4(n5229), .ZN(
        n4446) );
  INVD1BWP12T U4842 ( .I(n4393), .ZN(n4394) );
  AOI21D1BWP12T U4843 ( .A1(n4491), .A2(n4395), .B(n4394), .ZN(n4397) );
  XOR2XD1BWP12T U4844 ( .A1(n4397), .A2(n4396), .Z(n4812) );
  ND2XD0BWP12T U4845 ( .A1(n4403), .A2(n4402), .ZN(n4399) );
  AOI21D1BWP12T U4846 ( .A1(n4407), .A2(n4402), .B(n4404), .ZN(n4398) );
  OAI21D1BWP12T U4847 ( .A1(n4408), .A2(n4399), .B(n4398), .ZN(n4401) );
  XNR2XD1BWP12T U4848 ( .A1(n4401), .A2(n4400), .ZN(n5060) );
  AOI21D1BWP12T U4849 ( .A1(n4421), .A2(n4413), .B(n4415), .ZN(n4411) );
  CKND2D1BWP12T U4850 ( .A1(n4047), .A2(n4416), .ZN(n4410) );
  XOR2XD1BWP12T U4851 ( .A1(n4411), .A2(n4410), .Z(n5007) );
  NR2D0BWP12T U4852 ( .A1(n4412), .A2(n5007), .ZN(n4442) );
  CKND0BWP12T U4853 ( .I(n4413), .ZN(n4414) );
  NR2XD0BWP12T U4854 ( .A1(n4414), .A2(n4417), .ZN(n4420) );
  CKND0BWP12T U4855 ( .I(n4415), .ZN(n4418) );
  OAI21D0BWP12T U4856 ( .A1(n4418), .A2(n4417), .B(n4416), .ZN(n4419) );
  AOI21D1BWP12T U4857 ( .A1(n4421), .A2(n4420), .B(n4419), .ZN(n4425) );
  TPND2D0BWP12T U4858 ( .A1(n4423), .A2(n4422), .ZN(n4424) );
  XOR2XD1BWP12T U4859 ( .A1(n4425), .A2(n4424), .Z(n4881) );
  NR2D0BWP12T U4860 ( .A1(n4426), .A2(n4881), .ZN(n4441) );
  INVD1BWP12T U4861 ( .I(n4427), .ZN(n4435) );
  OAI21D1BWP12T U4862 ( .A1(n4435), .A2(n4428), .B(n4433), .ZN(n4432) );
  ND2XD0BWP12T U4863 ( .A1(n4430), .A2(n4429), .ZN(n4431) );
  XNR2XD1BWP12T U4864 ( .A1(n4432), .A2(n4431), .ZN(n5190) );
  ND2D1BWP12T U4865 ( .A1(n4437), .A2(n4436), .ZN(n4438) );
  XNR2D1BWP12T U4866 ( .A1(n3016), .A2(n4438), .ZN(n5314) );
  OR3D0BWP12T U4867 ( .A1(n4965), .A2(n4843), .A3(n5314), .Z(n4439) );
  NR2D0BWP12T U4868 ( .A1(n5190), .A2(n4439), .ZN(n4440) );
  IND4D1BWP12T U4869 ( .A1(n4443), .B1(n4442), .B2(n4441), .B3(n4440), .ZN(
        n4444) );
  NR4D0BWP12T U4870 ( .A1(n4812), .A2(n5060), .A3(n5270), .A4(n4444), .ZN(
        n4445) );
  ND4D1BWP12T U4871 ( .A1(n4448), .A2(n4447), .A3(n4446), .A4(n4445), .ZN(
        n4499) );
  XNR2XD1BWP12T U4872 ( .A1(n4491), .A2(n4449), .ZN(n4760) );
  NR3D0BWP12T U4873 ( .A1(n4760), .A2(n4451), .A3(n4450), .ZN(n4497) );
  INVD1BWP12T U4874 ( .I(n4452), .ZN(n4455) );
  NR2D0BWP12T U4875 ( .A1(n4981), .A2(n4937), .ZN(n4496) );
  INVD1BWP12T U4876 ( .I(n4458), .ZN(n4477) );
  ND2D1BWP12T U4877 ( .A1(n4477), .A2(n4461), .ZN(n4463) );
  TPNR2D0BWP12T U4878 ( .A1(n4478), .A2(n4463), .ZN(n4465) );
  INVD1BWP12T U4879 ( .I(n4459), .ZN(n4485) );
  AOI21D1BWP12T U4880 ( .A1(n4485), .A2(n4461), .B(n4460), .ZN(n4462) );
  OAI21D1BWP12T U4881 ( .A1(n4488), .A2(n4463), .B(n4462), .ZN(n4464) );
  AOI21D1BWP12T U4882 ( .A1(n4491), .A2(n4465), .B(n4464), .ZN(n4467) );
  XOR2XD1BWP12T U4883 ( .A1(n4467), .A2(n4466), .Z(n4599) );
  NR2D0BWP12T U4884 ( .A1(n4468), .A2(n4599), .ZN(n4495) );
  CKND2D1BWP12T U4885 ( .A1(n4477), .A2(n4475), .ZN(n4470) );
  TPNR2D0BWP12T U4886 ( .A1(n4478), .A2(n4470), .ZN(n4472) );
  AOI21D1BWP12T U4887 ( .A1(n4485), .A2(n4475), .B(n4479), .ZN(n4469) );
  OAI21D1BWP12T U4888 ( .A1(n4488), .A2(n4470), .B(n4469), .ZN(n4471) );
  AOI21D1BWP12T U4889 ( .A1(n4491), .A2(n4472), .B(n4471), .ZN(n4474) );
  XOR2XD1BWP12T U4890 ( .A1(n4474), .A2(n4473), .Z(n4999) );
  INVD0BWP12T U4891 ( .I(n4475), .ZN(n4476) );
  NR2XD0BWP12T U4892 ( .A1(n4476), .A2(n4481), .ZN(n4484) );
  ND2D1BWP12T U4893 ( .A1(n4484), .A2(n4477), .ZN(n4487) );
  TPNR2D0BWP12T U4894 ( .A1(n4478), .A2(n4487), .ZN(n4490) );
  CKND0BWP12T U4895 ( .I(n4479), .ZN(n4482) );
  TPOAI21D0BWP12T U4896 ( .A1(n4482), .A2(n4481), .B(n4480), .ZN(n4483) );
  AOI21D1BWP12T U4897 ( .A1(n4485), .A2(n4484), .B(n4483), .ZN(n4486) );
  OAI21D1BWP12T U4898 ( .A1(n4488), .A2(n4487), .B(n4486), .ZN(n4489) );
  AOI21D1BWP12T U4899 ( .A1(n4491), .A2(n4490), .B(n4489), .ZN(n4493) );
  XOR2XD1BWP12T U4900 ( .A1(n4493), .A2(n4492), .Z(n5170) );
  NR2D0BWP12T U4901 ( .A1(n4999), .A2(n5170), .ZN(n4494) );
  ND4D1BWP12T U4902 ( .A1(n4497), .A2(n4496), .A3(n4495), .A4(n4494), .ZN(
        n4498) );
  ND4D0BWP12T U4903 ( .A1(n4500), .A2(a[18]), .A3(n5118), .A4(n4565), .ZN(
        n4507) );
  ND4D0BWP12T U4904 ( .A1(n4568), .A2(n454), .A3(n4649), .A4(n4914), .ZN(n4506) );
  ND4D0BWP12T U4905 ( .A1(n4502), .A2(n5234), .A3(n5030), .A4(n4501), .ZN(
        n4505) );
  ND4D1BWP12T U4906 ( .A1(n1), .A2(n4503), .A3(n4943), .A4(n4990), .ZN(n4504)
         );
  NR4D0BWP12T U4907 ( .A1(n4507), .A2(n4506), .A3(n4505), .A4(n4504), .ZN(
        n4517) );
  ND4D0BWP12T U4908 ( .A1(n4788), .A2(n5256), .A3(n448), .A4(n4508), .ZN(n4515) );
  ND4D0BWP12T U4909 ( .A1(n5146), .A2(n4510), .A3(n4891), .A4(n4509), .ZN(
        n4514) );
  ND4D0BWP12T U4910 ( .A1(n5079), .A2(n4511), .A3(n4541), .A4(n5236), .ZN(
        n4513) );
  ND4D0BWP12T U4911 ( .A1(n5108), .A2(n4518), .A3(n5192), .A4(n436), .ZN(n4512) );
  NR4D0BWP12T U4912 ( .A1(n4515), .A2(n4514), .A3(n4513), .A4(n4512), .ZN(
        n4516) );
  AN2D0BWP12T U4913 ( .A1(n4517), .A2(n4516), .Z(n4591) );
  TPNR2D0BWP12T U4914 ( .A1(n4519), .A2(n4518), .ZN(n4520) );
  CKND2D1BWP12T U4915 ( .A1(n4577), .A2(n4520), .ZN(n4522) );
  XOR2XD1BWP12T U4916 ( .A1(n4522), .A2(n4521), .Z(n5090) );
  NR4D0BWP12T U4917 ( .A1(n4524), .A2(n4523), .A3(n5090), .A4(n5231), .ZN(
        n4550) );
  INVD1BWP12T U4918 ( .I(n4572), .ZN(n4532) );
  NR2D0BWP12T U4919 ( .A1(n4532), .A2(n5118), .ZN(n4525) );
  CKND2D1BWP12T U4920 ( .A1(n4582), .A2(n4525), .ZN(n4526) );
  XOR2XD1BWP12T U4921 ( .A1(n4526), .A2(n4672), .Z(n4685) );
  NR2XD0BWP12T U4922 ( .A1(n4532), .A2(n4529), .ZN(n4527) );
  CKND2D1BWP12T U4923 ( .A1(n4582), .A2(n4527), .ZN(n4528) );
  XOR2D1BWP12T U4924 ( .A1(n4528), .A2(n2825), .Z(n4638) );
  CKND0BWP12T U4925 ( .I(n4529), .ZN(n4530) );
  CKND2D0BWP12T U4926 ( .A1(n4530), .A2(n4635), .ZN(n4531) );
  NR2D1BWP12T U4927 ( .A1(n4532), .A2(n4531), .ZN(n4533) );
  CKND2D1BWP12T U4928 ( .A1(n4582), .A2(n4533), .ZN(n4534) );
  XOR2D1BWP12T U4929 ( .A1(n4534), .A2(n4914), .Z(n4928) );
  NR4D0BWP12T U4930 ( .A1(n4535), .A2(n4685), .A3(n4638), .A4(n4928), .ZN(
        n4549) );
  XNR2XD1BWP12T U4931 ( .A1(n4501), .A2(n3015), .ZN(n4850) );
  XNR2D0BWP12T U4932 ( .A1(n4536), .A2(n5192), .ZN(n5199) );
  OR4D0BWP12T U4933 ( .A1(n4850), .A2(n5104), .A3(n4537), .A4(n5199), .Z(n4538) );
  NR4D0BWP12T U4934 ( .A1(n4540), .A2(n5102), .A3(n4539), .A4(n4538), .ZN(
        n4548) );
  NR2XD0BWP12T U4935 ( .A1(n4543), .A2(n4542), .ZN(n4544) );
  XNR2D1BWP12T U4936 ( .A1(n4544), .A2(n4891), .ZN(n4878) );
  XNR2XD1BWP12T U4937 ( .A1(n4582), .A2(n448), .ZN(n4832) );
  CKND0BWP12T U4938 ( .I(n4571), .ZN(n4545) );
  TPND2D0BWP12T U4939 ( .A1(n4582), .A2(n4545), .ZN(n4546) );
  XOR2D1BWP12T U4940 ( .A1(n4546), .A2(n4649), .Z(n4648) );
  NR4D0BWP12T U4941 ( .A1(n5020), .A2(n4878), .A3(n4832), .A4(n4648), .ZN(
        n4547) );
  ND4D1BWP12T U4942 ( .A1(n4550), .A2(n4549), .A3(n4548), .A4(n4547), .ZN(
        n4589) );
  INVD0BWP12T U4943 ( .I(n4559), .ZN(n4551) );
  NR2D1BWP12T U4944 ( .A1(n4571), .A2(n4551), .ZN(n4552) );
  CKND2D1BWP12T U4945 ( .A1(n4552), .A2(n4582), .ZN(n4553) );
  XOR2D1BWP12T U4946 ( .A1(n4553), .A2(n1), .Z(n4617) );
  CKND2D1BWP12T U4947 ( .A1(n4559), .A2(n4607), .ZN(n4554) );
  NR2D1BWP12T U4948 ( .A1(n4571), .A2(n4554), .ZN(n4555) );
  CKND2D1BWP12T U4949 ( .A1(n4555), .A2(n4582), .ZN(n4556) );
  XOR2D1BWP12T U4950 ( .A1(n4556), .A2(n2255), .Z(n4989) );
  INVD0BWP12T U4951 ( .I(n4557), .ZN(n4558) );
  TPND2D0BWP12T U4952 ( .A1(n4559), .A2(n4558), .ZN(n4560) );
  TPNR2D0BWP12T U4953 ( .A1(n4571), .A2(n4560), .ZN(n4561) );
  TPND2D0BWP12T U4954 ( .A1(n4561), .A2(n4582), .ZN(n4562) );
  XOR2XD1BWP12T U4955 ( .A1(n4562), .A2(n5146), .Z(n5158) );
  NR4D0BWP12T U4956 ( .A1(n4563), .A2(n4617), .A3(n4989), .A4(n5158), .ZN(
        n4587) );
  NR2D1BWP12T U4957 ( .A1(n4580), .A2(a[18]), .ZN(n4564) );
  CKND2D1BWP12T U4958 ( .A1(n4582), .A2(n4564), .ZN(n4566) );
  XOR2XD1BWP12T U4959 ( .A1(n4566), .A2(n4696), .Z(n4709) );
  NR2D1BWP12T U4960 ( .A1(n4571), .A2(n4649), .ZN(n4567) );
  CKND2D1BWP12T U4961 ( .A1(n4567), .A2(n4582), .ZN(n4569) );
  XOR2D1BWP12T U4962 ( .A1(n4569), .A2(n4568), .Z(n4973) );
  CKND2D1BWP12T U4963 ( .A1(n4582), .A2(n4572), .ZN(n4573) );
  XOR2D1BWP12T U4964 ( .A1(n4573), .A2(n5118), .Z(n5128) );
  NR4D0BWP12T U4965 ( .A1(n4709), .A2(n4973), .A3(n4951), .A4(n5128), .ZN(
        n4586) );
  INVD0BWP12T U4966 ( .I(n4574), .ZN(n4576) );
  NR2D0BWP12T U4967 ( .A1(n5059), .A2(n5268), .ZN(n4585) );
  CKND2D1BWP12T U4968 ( .A1(n4582), .A2(n4578), .ZN(n4579) );
  XOR2XD1BWP12T U4969 ( .A1(n4579), .A2(n4788), .Z(n4802) );
  CKND0BWP12T U4970 ( .I(n4580), .ZN(n4581) );
  CKND2D1BWP12T U4971 ( .A1(n4582), .A2(n4581), .ZN(n4583) );
  XOR2XD1BWP12T U4972 ( .A1(n4583), .A2(a[18]), .Z(n4736) );
  NR3D0BWP12T U4973 ( .A1(n4758), .A2(n4802), .A3(n4736), .ZN(n4584) );
  ND4D1BWP12T U4974 ( .A1(n4587), .A2(n4586), .A3(n4585), .A4(n4584), .ZN(
        n4588) );
  NR2D1BWP12T U4975 ( .A1(n4589), .A2(n4588), .ZN(n4590) );
  INR2D1BWP12T U4976 ( .A1(n4594), .B1(n4593), .ZN(n4595) );
  ND2D4BWP12T U4977 ( .A1(n4597), .A2(n5292), .ZN(n4627) );
  INR2D1BWP12T U4978 ( .A1(n4598), .B1(n4970), .ZN(n4621) );
  INVD1BWP12T U4979 ( .I(n4599), .ZN(n4619) );
  INVD1BWP12T U4980 ( .I(n4600), .ZN(n4603) );
  INR2D1BWP12T U4981 ( .A1(n4601), .B1(n4924), .ZN(n5161) );
  AOI22D1BWP12T U4982 ( .A1(n4603), .A2(n5252), .B1(n5161), .B2(n4602), .ZN(
        n4604) );
  OAI21D1BWP12T U4983 ( .A1(n4605), .A2(n5312), .B(n4604), .ZN(n4616) );
  CKMUX2D1BWP12T U4984 ( .I0(n5258), .I1(n5257), .S(n22), .Z(n4606) );
  NR2D0BWP12T U4985 ( .A1(n4606), .A2(n5296), .ZN(n4608) );
  OA21D0BWP12T U4986 ( .A1(n4611), .A2(n5296), .B(n22), .Z(n4612) );
  AO211D1BWP12T U4987 ( .A1(n4614), .A2(n5322), .B(n4613), .C(n4612), .Z(n4615) );
  AOI211D1BWP12T U4988 ( .A1(n5297), .A2(n4617), .B(n4616), .C(n4615), .ZN(
        n4618) );
  OAI21D1BWP12T U4989 ( .A1(n4619), .A2(n4965), .B(n4618), .ZN(n4620) );
  AOI211XD1BWP12T U4990 ( .A1(n4622), .A2(n5308), .B(n4621), .C(n4620), .ZN(
        n4623) );
  IOA21D2BWP12T U4991 ( .A1(n4624), .A2(n5305), .B(n4623), .ZN(n4625) );
  INVD3BWP12T U4992 ( .I(n4625), .ZN(n4626) );
  CKND2D4BWP12T U4993 ( .A1(n4628), .A2(n5292), .ZN(n4643) );
  INR2D1BWP12T U4994 ( .A1(n4629), .B1(n5105), .ZN(n4640) );
  ND2D1BWP12T U4995 ( .A1(n4633), .A2(n5322), .ZN(n5155) );
  AOI211XD1BWP12T U4996 ( .A1(n4641), .A2(n5305), .B(n4640), .C(n4639), .ZN(
        n4642) );
  TPND2D8BWP12T U4997 ( .A1(n4643), .A2(n4642), .ZN(result[22]) );
  NR2XD0BWP12T U4998 ( .A1(n4646), .A2(n5312), .ZN(n4647) );
  AOI21D1BWP12T U4999 ( .A1(n4648), .A2(n5297), .B(n4647), .ZN(n4661) );
  OAI21D1BWP12T U5000 ( .A1(n4649), .A2(n5255), .B(n5254), .ZN(n4654) );
  CKMUX2D1BWP12T U5001 ( .I0(n5258), .I1(n5257), .S(n4655), .Z(n4650) );
  NR2D0BWP12T U5002 ( .A1(n4650), .A2(n5296), .ZN(n4652) );
  MUX2ND0BWP12T U5003 ( .I0(n4652), .I1(n5299), .S(n4651), .ZN(n4653) );
  RCAOI21D0BWP12T U5004 ( .A1(n4655), .A2(n4654), .B(n4653), .ZN(n4656) );
  TPOAI21D0BWP12T U5005 ( .A1(n4657), .A2(n5271), .B(n4656), .ZN(n4658) );
  CKND2D1BWP12T U5006 ( .A1(n4924), .A2(n5155), .ZN(n4821) );
  TPAOI21D2BWP12T U5007 ( .A1(n4665), .A2(n5305), .B(n4664), .ZN(n4666) );
  CKND2D4BWP12T U5008 ( .A1(n4668), .A2(n5292), .ZN(n4691) );
  CKND2D1BWP12T U5009 ( .A1(n4669), .A2(n5305), .ZN(n4689) );
  OAI21D0BWP12T U5010 ( .A1(n4672), .A2(n5255), .B(n5254), .ZN(n4675) );
  MUX2D1BWP12T U5011 ( .I0(n5295), .I1(n5294), .S(n17), .Z(n4671) );
  CKND2D0BWP12T U5012 ( .A1(n4671), .A2(n5254), .ZN(n4673) );
  MUX2XD0BWP12T U5013 ( .I0(n5236), .I1(n4673), .S(n4672), .Z(n4674) );
  AOI21D1BWP12T U5014 ( .A1(n17), .A2(n4675), .B(n4674), .ZN(n4677) );
  OA21D0BWP12T U5015 ( .A1(n4678), .A2(n5155), .B(n4677), .Z(n4679) );
  TPOAI21D0BWP12T U5016 ( .A1(n5232), .A2(n4680), .B(n4679), .ZN(n4683) );
  INVD1BWP12T U5017 ( .I(n5151), .ZN(n4702) );
  TPOAI21D0BWP12T U5018 ( .A1(n4681), .A2(n4924), .B(n4702), .ZN(n4682) );
  AN2XD2BWP12T U5019 ( .A1(n4689), .A2(n4688), .Z(n4690) );
  TPND2D8BWP12T U5020 ( .A1(n4691), .A2(n4690), .ZN(result[21]) );
  INVD1BWP12T U5021 ( .I(n4693), .ZN(n4722) );
  INVD1BWP12T U5022 ( .I(n4694), .ZN(n4718) );
  OAI21D0BWP12T U5023 ( .A1(n4696), .A2(n5255), .B(n5254), .ZN(n4699) );
  MUX2XD0BWP12T U5024 ( .I0(n5295), .I1(n5294), .S(n16), .Z(n4695) );
  ND2XD0BWP12T U5025 ( .A1(n4695), .A2(n5254), .ZN(n4697) );
  MUX2D0BWP12T U5026 ( .I0(n5236), .I1(n4697), .S(n4696), .Z(n4698) );
  AOI21D1BWP12T U5027 ( .A1(n16), .A2(n4699), .B(n4698), .ZN(n4701) );
  ND2D1BWP12T U5028 ( .A1(n4702), .A2(n4701), .ZN(n4705) );
  NR2D1BWP12T U5029 ( .A1(n4703), .A2(n5155), .ZN(n4704) );
  AOI211D1BWP12T U5030 ( .A1(n4706), .A2(n5252), .B(n4705), .C(n4704), .ZN(
        n4707) );
  TPOAI21D0BWP12T U5031 ( .A1(n5312), .A2(n4708), .B(n4707), .ZN(n4716) );
  INVD1BWP12T U5032 ( .I(n4709), .ZN(n4711) );
  OAI22D1BWP12T U5033 ( .A1(n4711), .A2(n5104), .B1(n4924), .B2(n4710), .ZN(
        n4714) );
  CKND2D1BWP12T U5034 ( .A1(n4712), .A2(n5303), .ZN(n4713) );
  IND2XD1BWP12T U5035 ( .A1(n4714), .B1(n4713), .ZN(n4715) );
  NR2D1BWP12T U5036 ( .A1(n4716), .A2(n4715), .ZN(n4717) );
  OAI21D1BWP12T U5037 ( .A1(n4718), .A2(n4965), .B(n4717), .ZN(n4719) );
  AOI21D1BWP12T U5038 ( .A1(n4720), .A2(n5308), .B(n4719), .ZN(n4721) );
  OA21D2BWP12T U5039 ( .A1(n4722), .A2(n5203), .B(n4721), .Z(n4723) );
  INVD1BWP12T U5040 ( .I(n4726), .ZN(n4750) );
  INVD1BWP12T U5041 ( .I(n4727), .ZN(n4743) );
  OAI21D1BWP12T U5042 ( .A1(a[18]), .A2(n5255), .B(n5254), .ZN(n4731) );
  MUX2XD0BWP12T U5043 ( .I0(n5295), .I1(n5294), .S(n25), .Z(n4728) );
  ND2XD0BWP12T U5044 ( .A1(n4728), .A2(n5254), .ZN(n4729) );
  MUX2XD0BWP12T U5045 ( .I0(n5236), .I1(n4729), .S(a[18]), .Z(n4730) );
  AOI21D1BWP12T U5046 ( .A1(n25), .A2(n4731), .B(n4730), .ZN(n4733) );
  OAI21D1BWP12T U5047 ( .A1(n4734), .A2(n5232), .B(n4733), .ZN(n4735) );
  AOI21D1BWP12T U5048 ( .A1(n4736), .A2(n5297), .B(n4735), .ZN(n4737) );
  IOA21D1BWP12T U5049 ( .A1(n4738), .A2(n4974), .B(n4737), .ZN(n4741) );
  NR2D1BWP12T U5050 ( .A1(n4739), .A2(n5312), .ZN(n4740) );
  NR2D1BWP12T U5051 ( .A1(n4741), .A2(n4740), .ZN(n4742) );
  OAI21D1BWP12T U5052 ( .A1(n4743), .A2(n4965), .B(n4742), .ZN(n4748) );
  ND2D1BWP12T U5053 ( .A1(n4744), .A2(n5303), .ZN(n4745) );
  IOA21D1BWP12T U5054 ( .A1(n5322), .A2(n4746), .B(n4745), .ZN(n4747) );
  TPNR2D1BWP12T U5055 ( .A1(n4748), .A2(n4747), .ZN(n4749) );
  OAI21D1BWP12T U5056 ( .A1(n4750), .A2(n5105), .B(n4749), .ZN(n4751) );
  TPAOI21D2BWP12T U5057 ( .A1(n4752), .A2(n5305), .B(n4751), .ZN(n4753) );
  ND2XD3BWP12T U5058 ( .A1(n4755), .A2(n5292), .ZN(n4784) );
  NR2D1BWP12T U5059 ( .A1(n4756), .A2(n5271), .ZN(n4757) );
  AO21D1BWP12T U5060 ( .A1(n4758), .A2(n5297), .B(n4757), .Z(n4759) );
  AOI21D1BWP12T U5061 ( .A1(n4760), .A2(n5313), .B(n4759), .ZN(n4782) );
  ND2D1BWP12T U5062 ( .A1(n4761), .A2(n5303), .ZN(n4776) );
  INVD1BWP12T U5063 ( .I(n4762), .ZN(n4763) );
  TPOAI21D0BWP12T U5064 ( .A1(n4764), .A2(n4763), .B(n5072), .ZN(n4765) );
  OAI21D1BWP12T U5065 ( .A1(n4766), .A2(n5312), .B(n4765), .ZN(n4774) );
  OAI21D0BWP12T U5066 ( .A1(n4508), .A2(n5255), .B(n5254), .ZN(n4769) );
  CKMUX2D1BWP12T U5067 ( .I0(n5236), .I1(n4767), .S(n4508), .Z(n4768) );
  AOI21D1BWP12T U5068 ( .A1(n32), .A2(n4769), .B(n4768), .ZN(n4771) );
  OAI21D1BWP12T U5069 ( .A1(n4772), .A2(n5232), .B(n4771), .ZN(n4773) );
  NR2D1BWP12T U5070 ( .A1(n4774), .A2(n4773), .ZN(n4775) );
  ND2D1BWP12T U5071 ( .A1(n4776), .A2(n4775), .ZN(n4781) );
  CKND2D1BWP12T U5072 ( .A1(n4777), .A2(n5308), .ZN(n4778) );
  IOA21D1BWP12T U5073 ( .A1(n4779), .A2(n5305), .B(n4778), .ZN(n4780) );
  INR3D2BWP12T U5074 ( .A1(n4782), .B1(n4781), .B2(n4780), .ZN(n4783) );
  ND2D4BWP12T U5075 ( .A1(n4784), .A2(n4783), .ZN(result[15]) );
  INR2D1BWP12T U5076 ( .A1(n4786), .B1(n5105), .ZN(n4807) );
  OAI21D0BWP12T U5077 ( .A1(n4788), .A2(n5255), .B(n5254), .ZN(n4793) );
  MUX2XD0BWP12T U5078 ( .I0(n5258), .I1(n5257), .S(n4794), .Z(n4789) );
  NR2D0BWP12T U5079 ( .A1(n4789), .A2(n5296), .ZN(n4791) );
  MUX2NXD0BWP12T U5080 ( .I0(n4791), .I1(n5299), .S(n4790), .ZN(n4792) );
  TPAOI21D1BWP12T U5081 ( .A1(n4794), .A2(n4793), .B(n4792), .ZN(n4797) );
  NR2D0BWP12T U5082 ( .A1(n4795), .A2(n4924), .ZN(n4796) );
  INR3D0BWP12T U5083 ( .A1(n4797), .B1(n5151), .B2(n4796), .ZN(n4800) );
  CKND2D1BWP12T U5084 ( .A1(n4798), .A2(n5252), .ZN(n4799) );
  INVD1BWP12T U5085 ( .I(n4802), .ZN(n4804) );
  AOI211XD1BWP12T U5086 ( .A1(n4808), .A2(n5305), .B(n4807), .C(n4806), .ZN(
        n4809) );
  TPND2D2BWP12T U5087 ( .A1(n4811), .A2(n5292), .ZN(n4842) );
  INVD1BWP12T U5088 ( .I(n4812), .ZN(n4835) );
  INVD0BWP12T U5089 ( .I(n4819), .ZN(n4820) );
  CKND2D1BWP12T U5090 ( .A1(n4821), .A2(n4820), .ZN(n4830) );
  OAI21D1BWP12T U5091 ( .A1(n4822), .A2(n5255), .B(n5254), .ZN(n4825) );
  MUX2XD0BWP12T U5092 ( .I0(n5299), .I1(n4823), .S(n448), .Z(n4824) );
  IOA21D1BWP12T U5093 ( .A1(n4826), .A2(n4825), .B(n4824), .ZN(n4827) );
  AOI211D1BWP12T U5094 ( .A1(n5252), .A2(n4828), .B(n5151), .C(n4827), .ZN(
        n4829) );
  CKND2D1BWP12T U5095 ( .A1(n4830), .A2(n4829), .ZN(n4831) );
  AOI21D1BWP12T U5096 ( .A1(n4832), .A2(n5297), .B(n4831), .ZN(n4833) );
  OAI211D1BWP12T U5097 ( .A1(n4965), .A2(n4835), .B(n4834), .C(n4833), .ZN(
        n4836) );
  AOI21D1BWP12T U5098 ( .A1(n5308), .A2(n4837), .B(n4836), .ZN(n4838) );
  IOA21D1BWP12T U5099 ( .A1(n4839), .A2(n5305), .B(n4838), .ZN(n4840) );
  INVD1P75BWP12T U5100 ( .I(n4840), .ZN(n4841) );
  ND2D4BWP12T U5101 ( .A1(n4842), .A2(n4841), .ZN(result[16]) );
  AOI22D1BWP12T U5102 ( .A1(n4844), .A2(n5303), .B1(n4843), .B2(n5313), .ZN(
        n4857) );
  OAI21D0BWP12T U5103 ( .A1(n3684), .A2(n5255), .B(n5254), .ZN(n4848) );
  MUX2XD0BWP12T U5104 ( .I0(n5258), .I1(n5257), .S(n4849), .Z(n4845) );
  NR2XD0BWP12T U5105 ( .A1(n4845), .A2(n5296), .ZN(n4846) );
  MUX2D1BWP12T U5106 ( .I0(n5299), .I1(n4846), .S(n4501), .Z(n4847) );
  IOA21D1BWP12T U5107 ( .A1(n4849), .A2(n4848), .B(n4847), .ZN(n4852) );
  CKAN2D1BWP12T U5108 ( .A1(n4850), .A2(n5297), .Z(n4851) );
  NR2XD0BWP12T U5109 ( .A1(n4852), .A2(n4851), .ZN(n4856) );
  AOI22D1BWP12T U5110 ( .A1(n4854), .A2(n5308), .B1(n4853), .B2(n5305), .ZN(
        n4855) );
  ND3D1BWP12T U5111 ( .A1(n4857), .A2(n4856), .A3(n4855), .ZN(n4858) );
  RCAOI21D0BWP12T U5112 ( .A1(n5292), .A2(n4859), .B(n4858), .ZN(n4865) );
  ND2D1BWP12T U5113 ( .A1(n5181), .A2(n4860), .ZN(n4864) );
  INVD1BWP12T U5114 ( .I(n4861), .ZN(n4862) );
  ND2D1BWP12T U5115 ( .A1(n4862), .A2(n5321), .ZN(n4863) );
  ND3D1BWP12T U5116 ( .A1(n4865), .A2(n4864), .A3(n4863), .ZN(n4868) );
  INR2D2BWP12T U5117 ( .A1(n5322), .B1(n4866), .ZN(n4867) );
  NR2D2BWP12T U5118 ( .A1(n4868), .A2(n4867), .ZN(n4875) );
  INR3XD1BWP12T U5119 ( .A1(n4870), .B1(n5327), .B2(n4869), .ZN(n4873) );
  TPNR2D1BWP12T U5120 ( .A1(n4871), .A2(n5312), .ZN(n4872) );
  ND2D4BWP12T U5121 ( .A1(n4875), .A2(n4874), .ZN(result[1]) );
  INVD1P75BWP12T U5122 ( .I(n4876), .ZN(n4877) );
  TPNR2D2BWP12T U5123 ( .A1(n4877), .A2(n5112), .ZN(n4908) );
  AOI22D1BWP12T U5124 ( .A1(n5308), .A2(n4879), .B1(n4878), .B2(n5297), .ZN(
        n4888) );
  AOI22D1BWP12T U5125 ( .A1(n5313), .A2(n4881), .B1(n4880), .B2(n5303), .ZN(
        n4887) );
  INVD1BWP12T U5126 ( .I(n4882), .ZN(n4883) );
  ND2XD0BWP12T U5127 ( .A1(n4883), .A2(n5212), .ZN(n4886) );
  CKND2D1BWP12T U5128 ( .A1(n4884), .A2(n5305), .ZN(n4885) );
  AN4D2BWP12T U5129 ( .A1(n4888), .A2(n4887), .A3(n4886), .A4(n4885), .Z(n4907) );
  OAI21D0BWP12T U5130 ( .A1(n4890), .A2(n5312), .B(n4889), .ZN(n4901) );
  OAI21D0BWP12T U5131 ( .A1(n4891), .A2(n5255), .B(n5254), .ZN(n4895) );
  MUX2D1BWP12T U5132 ( .I0(n5236), .I1(n4893), .S(n4891), .Z(n4894) );
  OAI21D1BWP12T U5133 ( .A1(n5163), .A2(n5017), .B(n4897), .ZN(n4898) );
  AOI21D1BWP12T U5134 ( .A1(n4899), .A2(n5181), .B(n4898), .ZN(n4900) );
  IOA21D1BWP12T U5135 ( .A1(n4902), .A2(n4901), .B(n4900), .ZN(n4905) );
  TPNR2D1BWP12T U5136 ( .A1(n4903), .A2(n5271), .ZN(n4904) );
  NR2D2BWP12T U5137 ( .A1(n4905), .A2(n4904), .ZN(n4906) );
  IND3D4BWP12T U5138 ( .A1(n4908), .B1(n4907), .B2(n4906), .ZN(result[6]) );
  AOI22D1BWP12T U5139 ( .A1(n5308), .A2(n4911), .B1(n4910), .B2(n5305), .ZN(
        n4933) );
  OAI22D1BWP12T U5140 ( .A1(n4913), .A2(n5312), .B1(n4912), .B2(n5271), .ZN(
        n4927) );
  TPOAI21D0BWP12T U5141 ( .A1(n4914), .A2(n5255), .B(n5254), .ZN(n4919) );
  MUX2D1BWP12T U5142 ( .I0(n5295), .I1(n5294), .S(n4920), .Z(n4915) );
  CKND2D1BWP12T U5143 ( .A1(n4915), .A2(n5254), .ZN(n4917) );
  MUX2ND0BWP12T U5144 ( .I0(n4917), .I1(n5236), .S(n4916), .ZN(n4918) );
  IOA21D1BWP12T U5145 ( .A1(n4920), .A2(n4919), .B(n4918), .ZN(n4921) );
  AOI21D1BWP12T U5146 ( .A1(n4922), .A2(n5252), .B(n4921), .ZN(n4923) );
  OAI21D1BWP12T U5147 ( .A1(n4925), .A2(n4924), .B(n4923), .ZN(n4926) );
  AOI211D1BWP12T U5148 ( .A1(n4928), .A2(n5297), .B(n4927), .C(n4926), .ZN(
        n4932) );
  AOI22D1BWP12T U5149 ( .A1(n4930), .A2(n5313), .B1(n4929), .B2(n5303), .ZN(
        n4931) );
  INVD1BWP12T U5150 ( .I(n4937), .ZN(n4966) );
  INVD1BWP12T U5151 ( .I(n4938), .ZN(n4961) );
  NR2D1BWP12T U5152 ( .A1(n4939), .A2(n5232), .ZN(n4950) );
  INR2D1BWP12T U5153 ( .A1(n5322), .B1(n4940), .ZN(n4979) );
  INVD1BWP12T U5154 ( .I(n4979), .ZN(n4948) );
  NR2XD0BWP12T U5155 ( .A1(n4942), .A2(n4941), .ZN(n4947) );
  OAI21D1BWP12T U5156 ( .A1(n4948), .A2(n4947), .B(n4946), .ZN(n4949) );
  AOI211XD0BWP12T U5157 ( .A1(n4951), .A2(n5297), .B(n4950), .C(n4949), .ZN(
        n4959) );
  INR2D0BWP12T U5158 ( .A1(n4952), .B1(n4970), .ZN(n4958) );
  NR2D1BWP12T U5159 ( .A1(n4954), .A2(n4953), .ZN(n4955) );
  OA21D1BWP12T U5160 ( .A1(n4956), .A2(n4955), .B(n5281), .Z(n4957) );
  INR3XD0BWP12T U5161 ( .A1(n4959), .B1(n4958), .B2(n4957), .ZN(n4960) );
  OAI21D1BWP12T U5162 ( .A1(n4961), .A2(n5203), .B(n4960), .ZN(n4962) );
  AOI21D1BWP12T U5163 ( .A1(n5308), .A2(n4963), .B(n4962), .ZN(n4964) );
  OA21XD2BWP12T U5164 ( .A1(n4966), .A2(n4965), .B(n4964), .Z(n4967) );
  TPND2D8BWP12T U5165 ( .A1(n4968), .A2(n4967), .ZN(result[26]) );
  ND2XD8BWP12T U5166 ( .A1(n4969), .A2(n5292), .ZN(n4987) );
  INVD3BWP12T U5167 ( .I(n4985), .ZN(n4986) );
  TPND2D8BWP12T U5168 ( .A1(n4987), .A2(n4986), .ZN(result[25]) );
  TPND2D8BWP12T U5169 ( .A1(n4988), .A2(n5292), .ZN(n5006) );
  MUX2ND0BWP12T U5170 ( .I0(n5295), .I1(n5294), .S(n31), .ZN(n4992) );
  NR2D0BWP12T U5171 ( .A1(n4992), .A2(n5296), .ZN(n4994) );
  CKND2D2BWP12T U5172 ( .A1(n5002), .A2(n5305), .ZN(n5003) );
  AN2D4BWP12T U5173 ( .A1(n5004), .A2(n5003), .Z(n5005) );
  ND2XD16BWP12T U5174 ( .A1(n5006), .A2(n5005), .ZN(result[29]) );
  ND2D1BWP12T U5175 ( .A1(n5007), .A2(n5313), .ZN(n5028) );
  INVD0BWP12T U5176 ( .I(n5008), .ZN(n5013) );
  TPND2D0BWP12T U5177 ( .A1(n5009), .A2(n5281), .ZN(n5010) );
  CKND2D1BWP12T U5178 ( .A1(n5010), .A2(n4889), .ZN(n5012) );
  AOI22D1BWP12T U5179 ( .A1(n5013), .A2(n5012), .B1(n5011), .B2(n5303), .ZN(
        n5016) );
  CKND2D1BWP12T U5180 ( .A1(n5014), .A2(n5308), .ZN(n5015) );
  ND2D1BWP12T U5181 ( .A1(n5016), .A2(n5015), .ZN(n5027) );
  CKND0BWP12T U5182 ( .I(n5017), .ZN(n5018) );
  ND2D1BWP12T U5183 ( .A1(n5019), .A2(n5018), .ZN(n5025) );
  AOI22D1BWP12T U5184 ( .A1(n5021), .A2(n5305), .B1(n5020), .B2(n5297), .ZN(
        n5024) );
  ND2D1BWP12T U5185 ( .A1(n5181), .A2(n5022), .ZN(n5023) );
  ND3D1BWP12T U5186 ( .A1(n5025), .A2(n5024), .A3(n5023), .ZN(n5026) );
  INR3XD1BWP12T U5187 ( .A1(n5028), .B1(n5027), .B2(n5026), .ZN(n5042) );
  CKMUX2D1BWP12T U5188 ( .I0(n5295), .I1(n5294), .S(n2190), .Z(n5031) );
  NR2D1BWP12T U5189 ( .A1(n5034), .A2(n5327), .ZN(n5036) );
  AN2XD2BWP12T U5190 ( .A1(n5036), .A2(n5035), .Z(n5037) );
  NR2D2BWP12T U5191 ( .A1(n5038), .A2(n5037), .ZN(n5041) );
  CKND2D2BWP12T U5192 ( .A1(n5039), .A2(n5292), .ZN(n5040) );
  ND3D4BWP12T U5193 ( .A1(n5042), .A2(n5041), .A3(n5040), .ZN(result[5]) );
  NR2D1BWP12T U5194 ( .A1(n5043), .A2(n5271), .ZN(n5044) );
  AOI21D1BWP12T U5195 ( .A1(n5045), .A2(n5303), .B(n5044), .ZN(n5046) );
  OAI21D1BWP12T U5196 ( .A1(n5047), .A2(n5312), .B(n5046), .ZN(n5068) );
  INVD1BWP12T U5197 ( .I(n5275), .ZN(n5241) );
  TPND2D1BWP12T U5198 ( .A1(n5048), .A2(n5241), .ZN(n5056) );
  OAI21D0BWP12T U5199 ( .A1(n5049), .A2(n5255), .B(n5254), .ZN(n5053) );
  MUX2D1BWP12T U5200 ( .I0(n5295), .I1(n5294), .S(n5054), .Z(n5050) );
  ND2XD0BWP12T U5201 ( .A1(n5050), .A2(n5254), .ZN(n5051) );
  CKMUX2D1BWP12T U5202 ( .I0(n5236), .I1(n5051), .S(n5049), .Z(n5052) );
  AOI21D1BWP12T U5203 ( .A1(n5054), .A2(n5053), .B(n5052), .ZN(n5055) );
  OAI211D1BWP12T U5204 ( .A1(n5232), .A2(n5057), .B(n5056), .C(n5055), .ZN(
        n5058) );
  AOI21D1BWP12T U5205 ( .A1(n5059), .A2(n5297), .B(n5058), .ZN(n5064) );
  ND2D1BWP12T U5206 ( .A1(n5060), .A2(n5313), .ZN(n5063) );
  CKND2D1BWP12T U5207 ( .A1(n5061), .A2(n5305), .ZN(n5062) );
  ND3D1BWP12T U5208 ( .A1(n5064), .A2(n5063), .A3(n5062), .ZN(n5067) );
  AN2XD2BWP12T U5209 ( .A1(n5065), .A2(n5308), .Z(n5066) );
  TPNR3D1BWP12T U5210 ( .A1(n5068), .A2(n5067), .A3(n5066), .ZN(n5069) );
  RCOAI21D2BWP12T U5211 ( .A1(n5070), .A2(n5112), .B(n5069), .ZN(result[13])
         );
  INVD1BWP12T U5212 ( .I(n5071), .ZN(n5075) );
  AOI22D1BWP12T U5213 ( .A1(n5075), .A2(n5074), .B1(n5073), .B2(n5072), .ZN(
        n5076) );
  IOA21D1BWP12T U5214 ( .A1(n5077), .A2(n5303), .B(n5076), .ZN(n5094) );
  NR2D1BWP12T U5215 ( .A1(n5078), .A2(n5271), .ZN(n5089) );
  OAI21D0BWP12T U5216 ( .A1(n5079), .A2(n5255), .B(n5254), .ZN(n5084) );
  MUX2XD0BWP12T U5217 ( .I0(n5258), .I1(n5257), .S(n5085), .Z(n5080) );
  NR2D0BWP12T U5218 ( .A1(n5080), .A2(n5296), .ZN(n5082) );
  MUX2NXD0BWP12T U5219 ( .I0(n5082), .I1(n5299), .S(n5081), .ZN(n5083) );
  AOI21D1BWP12T U5220 ( .A1(n5085), .A2(n5084), .B(n5083), .ZN(n5086) );
  OAI21D1BWP12T U5221 ( .A1(n5087), .A2(n5317), .B(n5086), .ZN(n5088) );
  AOI211D1BWP12T U5222 ( .A1(n5090), .A2(n5297), .B(n5089), .C(n5088), .ZN(
        n5091) );
  IOA21D1BWP12T U5223 ( .A1(n5092), .A2(n5313), .B(n5091), .ZN(n5093) );
  AOI211XD1BWP12T U5224 ( .A1(n5095), .A2(n5308), .B(n5094), .C(n5093), .ZN(
        n5096) );
  IOA21D2BWP12T U5225 ( .A1(n5305), .A2(n5097), .B(n5096), .ZN(n5098) );
  AO21D4BWP12T U5226 ( .A1(n5099), .A2(n5292), .B(n5098), .Z(result[11]) );
  XNR2D1BWP12T U5227 ( .A1(n5101), .A2(n5100), .ZN(n5113) );
  NR2D1BWP12T U5228 ( .A1(n5110), .A2(n5109), .ZN(n5111) );
  TPOAI21D1BWP12T U5229 ( .A1(n5113), .A2(n5112), .B(n5111), .ZN(v) );
  ND2D1BWP12T U5230 ( .A1(n5114), .A2(n5313), .ZN(n5137) );
  CKND2D1BWP12T U5231 ( .A1(n5115), .A2(n5322), .ZN(n5133) );
  NR2XD0BWP12T U5232 ( .A1(n5116), .A2(n5232), .ZN(n5124) );
  OAI21D0BWP12T U5233 ( .A1(n5118), .A2(n5255), .B(n5254), .ZN(n5121) );
  MUX2D1BWP12T U5234 ( .I0(n5258), .I1(n5257), .S(n26), .Z(n5117) );
  NR2D0BWP12T U5235 ( .A1(n5117), .A2(n5296), .ZN(n5119) );
  MUX2D0BWP12T U5236 ( .I0(n5299), .I1(n5119), .S(n5118), .Z(n5120) );
  IOA21D1BWP12T U5237 ( .A1(n26), .A2(n5121), .B(n5120), .ZN(n5123) );
  NR2D1BWP12T U5238 ( .A1(n5124), .A2(n5123), .ZN(n5125) );
  IOA21D1BWP12T U5239 ( .A1(n5127), .A2(n5126), .B(n5125), .ZN(n5132) );
  CKND2D1BWP12T U5240 ( .A1(n5128), .A2(n5297), .ZN(n5129) );
  IOA21D1BWP12T U5241 ( .A1(n5281), .A2(n5130), .B(n5129), .ZN(n5131) );
  INR3XD0BWP12T U5242 ( .A1(n5133), .B1(n5132), .B2(n5131), .ZN(n5136) );
  CKND2D1BWP12T U5243 ( .A1(n5134), .A2(n5303), .ZN(n5135) );
  ND3D1BWP12T U5244 ( .A1(n5137), .A2(n5136), .A3(n5135), .ZN(n5138) );
  AOI21D1BWP12T U5245 ( .A1(n5308), .A2(n5139), .B(n5138), .ZN(n5140) );
  INVD1P75BWP12T U5246 ( .I(n5142), .ZN(n5143) );
  RCOAI21D2BWP12T U5247 ( .A1(n5144), .A2(n5112), .B(n5143), .ZN(result[20])
         );
  OAI21D1BWP12T U5248 ( .A1(n5146), .A2(n5255), .B(n5254), .ZN(n5152) );
  NR2D0BWP12T U5249 ( .A1(n5147), .A2(n5296), .ZN(n5149) );
  MUX2ND0BWP12T U5250 ( .I0(n5149), .I1(n5299), .S(n5148), .ZN(n5150) );
  AOI211XD0BWP12T U5251 ( .A1(n5153), .A2(n5152), .B(n5151), .C(n5150), .ZN(
        n5154) );
  TPOAI21D0BWP12T U5252 ( .A1(n5156), .A2(n5155), .B(n5154), .ZN(n5157) );
  AOI21D1BWP12T U5253 ( .A1(n5158), .A2(n5297), .B(n5157), .ZN(n5168) );
  AOI22D1BWP12T U5254 ( .A1(n5161), .A2(n5160), .B1(n5159), .B2(n5252), .ZN(
        n5167) );
  NR2D1BWP12T U5255 ( .A1(n5163), .A2(n5162), .ZN(n5164) );
  OAI21D1BWP12T U5256 ( .A1(n5165), .A2(n5164), .B(n5281), .ZN(n5166) );
  ND3D1BWP12T U5257 ( .A1(n5168), .A2(n5167), .A3(n5166), .ZN(n5169) );
  AOI21D1BWP12T U5258 ( .A1(n5170), .A2(n5313), .B(n5169), .ZN(n5171) );
  IOA21D1BWP12T U5259 ( .A1(n5172), .A2(n5303), .B(n5171), .ZN(n5173) );
  AOI21D1BWP12T U5260 ( .A1(n5308), .A2(n5174), .B(n5173), .ZN(n5177) );
  ND2D1BWP12T U5261 ( .A1(n5175), .A2(n5305), .ZN(n5176) );
  AN2XD2BWP12T U5262 ( .A1(n5177), .A2(n5176), .Z(n5178) );
  ND2XD3BWP12T U5263 ( .A1(n5179), .A2(n5178), .ZN(result[30]) );
  ND2D1BWP12T U5264 ( .A1(n5181), .A2(n5180), .ZN(n5189) );
  NR3D1BWP12T U5265 ( .A1(n5183), .A2(n5182), .A3(n5312), .ZN(n5188) );
  INR3D2BWP12T U5266 ( .A1(n5189), .B1(n5188), .B2(n5187), .ZN(n5219) );
  ND2XD0BWP12T U5267 ( .A1(n5190), .A2(n5313), .ZN(n5202) );
  OAI21D0BWP12T U5268 ( .A1(n5192), .A2(n5255), .B(n5254), .ZN(n5195) );
  MUX2D1BWP12T U5269 ( .I0(n5258), .I1(n5257), .S(n5196), .Z(n5191) );
  NR2XD0BWP12T U5270 ( .A1(n5191), .A2(n5296), .ZN(n5193) );
  MUX2XD0BWP12T U5271 ( .I0(n5299), .I1(n5193), .S(n5192), .Z(n5194) );
  IOA21D1BWP12T U5272 ( .A1(n5196), .A2(n5195), .B(n5194), .ZN(n5197) );
  TPAOI21D0BWP12T U5273 ( .A1(n5198), .A2(n5303), .B(n5197), .ZN(n5201) );
  ND2D0BWP12T U5274 ( .A1(n5199), .A2(n5297), .ZN(n5200) );
  ND3D1BWP12T U5275 ( .A1(n5202), .A2(n5201), .A3(n5200), .ZN(n5209) );
  OR2D0BWP12T U5276 ( .A1(n5204), .A2(n5203), .Z(n5207) );
  ND2XD0BWP12T U5277 ( .A1(n5205), .A2(n5308), .ZN(n5206) );
  CKND2D1BWP12T U5278 ( .A1(n5207), .A2(n5206), .ZN(n5208) );
  NR2D1BWP12T U5279 ( .A1(n5209), .A2(n5208), .ZN(n5217) );
  INVD1BWP12T U5280 ( .I(n5210), .ZN(n5215) );
  INR2D1BWP12T U5281 ( .A1(n5212), .B1(n5211), .ZN(n5213) );
  OA21D1BWP12T U5282 ( .A1(n5215), .A2(n5214), .B(n5213), .Z(n5216) );
  INR2D2BWP12T U5283 ( .A1(n5217), .B1(n5216), .ZN(n5218) );
  CKND2D2BWP12T U5284 ( .A1(n5219), .A2(n5218), .ZN(n5224) );
  AOI22D1BWP12T U5285 ( .A1(n5226), .A2(n5305), .B1(n5225), .B2(n5308), .ZN(
        n5248) );
  INVD1BWP12T U5286 ( .I(n5227), .ZN(n5228) );
  AOI22D1BWP12T U5287 ( .A1(n5229), .A2(n5313), .B1(n5281), .B2(n5228), .ZN(
        n5246) );
  AOI22D1BWP12T U5288 ( .A1(n5231), .A2(n5297), .B1(n5322), .B2(n5230), .ZN(
        n5245) );
  NR2D1BWP12T U5289 ( .A1(n5233), .A2(n5232), .ZN(n5239) );
  AOI211D1BWP12T U5290 ( .A1(n5241), .A2(n5240), .B(n5239), .C(n5238), .ZN(
        n5244) );
  CKND2D1BWP12T U5291 ( .A1(n5242), .A2(n5303), .ZN(n5243) );
  AN4XD1BWP12T U5292 ( .A1(n5246), .A2(n5245), .A3(n5244), .A4(n5243), .Z(
        n5247) );
  AO21D4BWP12T U5293 ( .A1(n5250), .A2(n5292), .B(n5249), .Z(result[12]) );
  CKND2D1BWP12T U5294 ( .A1(n5251), .A2(n5305), .ZN(n5286) );
  CKND2D1BWP12T U5295 ( .A1(n5253), .A2(n5252), .ZN(n5266) );
  OAI21D1BWP12T U5296 ( .A1(a[14]), .A2(n5255), .B(n5254), .ZN(n5263) );
  MUX2XD0BWP12T U5297 ( .I0(n5258), .I1(n5257), .S(n5264), .Z(n5259) );
  NR2D0BWP12T U5298 ( .A1(n5259), .A2(n5296), .ZN(n5261) );
  MUX2NXD0BWP12T U5299 ( .I0(n5261), .I1(n5299), .S(n5260), .ZN(n5262) );
  AOI21D1BWP12T U5300 ( .A1(n5264), .A2(n5263), .B(n5262), .ZN(n5265) );
  ND2D1BWP12T U5301 ( .A1(n5266), .A2(n5265), .ZN(n5267) );
  AOI21D1BWP12T U5302 ( .A1(n5268), .A2(n5297), .B(n5267), .ZN(n5269) );
  IOA21D1BWP12T U5303 ( .A1(n5270), .A2(n5313), .B(n5269), .ZN(n5274) );
  NR2D1BWP12T U5304 ( .A1(n5272), .A2(n5271), .ZN(n5273) );
  TPNR2D1BWP12T U5305 ( .A1(n5274), .A2(n5273), .ZN(n5285) );
  NR2D1BWP12T U5306 ( .A1(n5276), .A2(n5275), .ZN(n5277) );
  AOI21D1BWP12T U5307 ( .A1(n5278), .A2(n5303), .B(n5277), .ZN(n5279) );
  IOA21D1BWP12T U5308 ( .A1(n5281), .A2(n5280), .B(n5279), .ZN(n5282) );
  AOI21D1BWP12T U5309 ( .A1(n5283), .A2(n5308), .B(n5282), .ZN(n5284) );
  ND3D1BWP12T U5310 ( .A1(n5286), .A2(n5285), .A3(n5284), .ZN(n5287) );
  AO21D4BWP12T U5311 ( .A1(n5288), .A2(n5292), .B(n5287), .Z(result[14]) );
  AOI22D0BWP12T U5312 ( .A1(n5290), .A2(n5289), .B1(n402), .B2(n5296), .ZN(
        n5291) );
  IOA21D1BWP12T U5313 ( .A1(n5293), .A2(n5292), .B(n5291), .ZN(n5302) );
  MUX2ND0BWP12T U5314 ( .I0(n5295), .I1(n5294), .S(n402), .ZN(n5298) );
  NR3D0BWP12T U5315 ( .A1(n5298), .A2(n5297), .A3(n5296), .ZN(n5300) );
  MUX2ND0BWP12T U5316 ( .I0(n5300), .I1(n5299), .S(n3015), .ZN(n5301) );
  RCAOI211D0BWP12T U5317 ( .A1(n5304), .A2(n5303), .B(n5302), .C(n5301), .ZN(
        n5310) );
  RCAOI22D0BWP12T U5318 ( .A1(n5308), .A2(n5307), .B1(n5306), .B2(n5305), .ZN(
        n5309) );
  OAI211D1BWP12T U5319 ( .A1(n5312), .A2(n5311), .B(n5310), .C(n5309), .ZN(
        n5319) );
  CKND2D1BWP12T U5320 ( .A1(n5314), .A2(n5313), .ZN(n5315) );
  OAI21D1BWP12T U5321 ( .A1(n5317), .A2(n5316), .B(n5315), .ZN(n5318) );
  AOI211XD0BWP12T U5322 ( .A1(n5321), .A2(n5320), .B(n5319), .C(n5318), .ZN(
        n5326) );
  INVD1BWP12T U5323 ( .I(n5328), .ZN(n5324) );
  OAI21D1BWP12T U5324 ( .A1(n5324), .A2(n5323), .B(n5322), .ZN(n5325) );
  OAI211D1BWP12T U5325 ( .A1(n5328), .A2(n5327), .B(n5326), .C(n5325), .ZN(
        result[0]) );
endmodule


module top7 ( clk, reset, MEM_MEMCTRL_from_mem_data, 
        MEMCTRL_MEM_to_mem_read_enable, MEMCTRL_MEM_to_mem_write_enable, 
        MEMCTRL_MEM_to_mem_mem_enable, MEMCTRL_MEM_to_mem_address, 
        MEMCTRL_MEM_to_mem_data );
  input [15:0] MEM_MEMCTRL_from_mem_data;
  output [11:0] MEMCTRL_MEM_to_mem_address;
  output [15:0] MEMCTRL_MEM_to_mem_data;
  input clk, reset;
  output MEMCTRL_MEM_to_mem_read_enable, MEMCTRL_MEM_to_mem_write_enable,
         MEMCTRL_MEM_to_mem_mem_enable;
  wire   DEC_CPSR_update_flag_n, new_n, ALU_OUT_n, RF_OUT_n,
         DEC_CPSR_update_flag_c, new_c, ALU_OUT_c, RF_OUT_c,
         DEC_CPSR_update_flag_z, new_z, ALU_OUT_z, RF_OUT_z,
         DEC_CPSR_update_flag_v, new_v, ALU_OUT_v, RF_OUT_v,
         DEC_RF_alu_write_to_reg_enable, DEC_RF_memory_write_to_reg_enable,
         DEC_MISC_OUT_memory_address_source_is_reg,
         DEC_MEMCTRL_memorycontroller_sign_extend,
         DEC_MEMCTRL_memory_load_request, DEC_MEMCTRL_memory_store_request,
         DEC_IF_stall_to_instructionfetch, ALU_IN_c, irdecode_inst1_N912,
         irdecode_inst1_N911, irdecode_inst1_N907, irdecode_inst1_N906,
         irdecode_inst1_N707, irdecode_inst1_N706, irdecode_inst1_N705,
         irdecode_inst1_N704, irdecode_inst1_N703, irdecode_inst1_N702,
         irdecode_inst1_N701, irdecode_inst1_N546, irdecode_inst1_N545,
         irdecode_inst1_N544, irdecode_inst1_N543, irdecode_inst1_N542,
         irdecode_inst1_N541, irdecode_inst1_N540, irdecode_inst1_N539,
         irdecode_inst1_split_instruction, irdecode_inst1_next_step_0_,
         irdecode_inst1_next_step_2_, irdecode_inst1_next_step_3_,
         irdecode_inst1_next_step_4_, irdecode_inst1_next_step_5_,
         irdecode_inst1_next_step_6_, irdecode_inst1_next_step_7_,
         irdecode_inst1_itstate_0_, irdecode_inst1_itstate_1_,
         irdecode_inst1_itstate_2_, irdecode_inst1_itstate_3_,
         irdecode_inst1_itstate_4_, irdecode_inst1_itstate_5_,
         irdecode_inst1_itstate_6_, irdecode_inst1_itstate_7_,
         irdecode_inst1_next_alu_write_to_reg_enable,
         irdecode_inst1_next_update_flag_v, irdecode_inst1_next_update_flag_c,
         irdecode_inst1_next_update_flag_n,
         memory_interface_inst1_delayed_is_signed, Instruction_Fetch_inst1_N98,
         Instruction_Fetch_inst1_N97, Instruction_Fetch_inst1_N96,
         Instruction_Fetch_inst1_N95, Instruction_Fetch_inst1_N94,
         Instruction_Fetch_inst1_N93, Instruction_Fetch_inst1_N92,
         Instruction_Fetch_inst1_N91, Instruction_Fetch_inst1_N90,
         Instruction_Fetch_inst1_N89, Instruction_Fetch_inst1_N88,
         Instruction_Fetch_inst1_N87, Instruction_Fetch_inst1_N86,
         Instruction_Fetch_inst1_N85, Instruction_Fetch_inst1_N84,
         Instruction_Fetch_inst1_N83, Instruction_Fetch_inst1_N80,
         Instruction_Fetch_inst1_N79,
         Instruction_Fetch_inst1_first_instruction_fetched,
         Instruction_Fetch_inst1_fetched_instruction_reg_0_,
         Instruction_Fetch_inst1_fetched_instruction_reg_1_,
         Instruction_Fetch_inst1_fetched_instruction_reg_2_,
         Instruction_Fetch_inst1_fetched_instruction_reg_3_,
         Instruction_Fetch_inst1_fetched_instruction_reg_4_,
         Instruction_Fetch_inst1_fetched_instruction_reg_5_,
         Instruction_Fetch_inst1_fetched_instruction_reg_6_,
         Instruction_Fetch_inst1_fetched_instruction_reg_7_,
         Instruction_Fetch_inst1_fetched_instruction_reg_8_,
         Instruction_Fetch_inst1_fetched_instruction_reg_9_,
         Instruction_Fetch_inst1_fetched_instruction_reg_10_,
         Instruction_Fetch_inst1_fetched_instruction_reg_11_,
         Instruction_Fetch_inst1_fetched_instruction_reg_12_,
         Instruction_Fetch_inst1_fetched_instruction_reg_13_,
         Instruction_Fetch_inst1_fetched_instruction_reg_14_,
         Instruction_Fetch_inst1_fetched_instruction_reg_15_,
         Instruction_Fetch_inst1_currentState_0_,
         Instruction_Fetch_inst1_currentState_1_,
         memory_interface_inst1_fsm_N35, memory_interface_inst1_fsm_N34,
         memory_interface_inst1_fsm_N33, memory_interface_inst1_fsm_N32,
         memory_interface_inst1_fsm_state_0_,
         memory_interface_inst1_fsm_state_1_,
         memory_interface_inst1_fsm_state_2_,
         memory_interface_inst1_fsm_state_3_, n754, n777, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53;
  wire   [7:0] IF_DEC_instruction;
  wire   [4:0] DEC_RF_operand_a;
  wire   [4:0] DEC_RF_operand_b;
  wire   [31:0] DEC_RF_offset_b;
  wire   [4:0] DEC_ALU_alu_opcode;
  wire   [4:0] DEC_RF_alu_write_to_reg;
  wire   [4:0] DEC_RF_memory_write_to_reg;
  wire   [4:0] DEC_RF_memory_store_data_reg;
  wire   [4:0] DEC_RF_memory_store_address_reg;
  wire   [1:0] DEC_MEMCTRL_load_store_width;
  wire   [31:0] ALU_MISC_OUT_result;
  wire   [31:0] MEMCTRL_RF_IF_data_in;
  wire   [31:0] IF_RF_incremented_pc_out;
  wire   [31:0] RF_ALU_operand_a;
  wire   [31:0] RF_ALU_operand_b;
  wire   [31:0] RF_MEMCTRL_data_reg;
  wire   [12:2] RF_MEMCTRL_address_reg;
  wire   [31:0] RF_pc_out;
  wire   [11:0] MEMCTRL_IN_address;
  wire   [7:0] irdecode_inst1_step;
  wire   [15:0] memory_interface_inst1_delay_first_two_bytes_out;
  wire   [31:0] memory_interface_inst1_delay_data_in32;
  wire   [11:0] memory_interface_inst1_delay_addr_for_adder;

  register_file register_file_inst1 ( .readA_sel(DEC_RF_operand_a), 
        .readB_sel(DEC_RF_operand_b), .readC_sel(DEC_RF_memory_store_data_reg), 
        .readD_sel(DEC_RF_memory_store_address_reg), .write1_sel(
        DEC_RF_alu_write_to_reg), .write2_sel(DEC_RF_memory_write_to_reg), 
        .write1_en(DEC_RF_alu_write_to_reg_enable), .write2_en(
        DEC_RF_memory_write_to_reg_enable), .write1_in(ALU_MISC_OUT_result), 
        .write2_in(MEMCTRL_RF_IF_data_in), .immediate1_in({n864, n864, n864, 
        n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, 
        n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, 
        n864, n864, n864, n864, n864}), .immediate2_in(DEC_RF_offset_b), 
        .next_pc_in({IF_RF_incremented_pc_out[31:28], n1843, 
        IF_RF_incremented_pc_out[26], n1842, IF_RF_incremented_pc_out[24:2], 
        MEMCTRL_IN_address[0], IF_RF_incremented_pc_out[0]}), .next_cpsr_in({
        new_n, new_c, new_z, new_v}), .next_sp_in({n864, n864, n864, n864, 
        n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, 
        n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, 
        n864, n864, n864, n864}), .clk(clk), .reset(reset), .regA_out(
        RF_ALU_operand_a), .regB_out(RF_ALU_operand_b), .regC_out(
        RF_MEMCTRL_data_reg), .regD_out({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        RF_MEMCTRL_address_reg, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21}), .pc_out(RF_pc_out), .cpsr_out({RF_OUT_n, 
        RF_OUT_c, RF_OUT_z, RF_OUT_v}), .sp_out({SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53}), .next_pc_en_BAR(n754) );
  ALU_VARIABLE ALU_VARIABLE_inst1 ( .a({RF_ALU_operand_a[31:18], n1853, 
        RF_ALU_operand_a[16:5], n1852, RF_ALU_operand_a[3:2], n1851, 
        RF_ALU_operand_a[0]}), .b({RF_ALU_operand_b[31:2], n1850, n1849}), 
        .op(DEC_ALU_alu_opcode[3:0]), .c_in(ALU_IN_c), .result(
        ALU_MISC_OUT_result), .c_out(ALU_OUT_c), .z(ALU_OUT_z), .n(ALU_OUT_n), 
        .v(ALU_OUT_v) );
  CKAN2D2BWP12T irdecode_inst1_C5193 ( .A1(irdecode_inst1_next_step_7_), .A2(
        IF_DEC_instruction[7]), .Z(irdecode_inst1_N539) );
  CKAN2D2BWP12T irdecode_inst1_C5194 ( .A1(irdecode_inst1_next_step_6_), .A2(
        IF_DEC_instruction[6]), .Z(irdecode_inst1_N540) );
  CKAN2D2BWP12T irdecode_inst1_C5195 ( .A1(irdecode_inst1_next_step_5_), .A2(
        IF_DEC_instruction[5]), .Z(irdecode_inst1_N541) );
  CKAN2D2BWP12T irdecode_inst1_C5196 ( .A1(irdecode_inst1_next_step_4_), .A2(
        IF_DEC_instruction[4]), .Z(irdecode_inst1_N542) );
  CKAN2D2BWP12T irdecode_inst1_C5197 ( .A1(irdecode_inst1_next_step_3_), .A2(
        IF_DEC_instruction[3]), .Z(irdecode_inst1_N543) );
  CKAN2D2BWP12T irdecode_inst1_C5198 ( .A1(irdecode_inst1_next_step_2_), .A2(
        IF_DEC_instruction[2]), .Z(irdecode_inst1_N544) );
  CKAN2D2BWP12T irdecode_inst1_C5199 ( .A1(n1841), .A2(IF_DEC_instruction[1]), 
        .Z(irdecode_inst1_N545) );
  CKAN2D2BWP12T irdecode_inst1_C5200 ( .A1(irdecode_inst1_next_step_0_), .A2(
        IF_DEC_instruction[0]), .Z(irdecode_inst1_N546) );
  CKAN2D2BWP12T irdecode_inst1_C5280 ( .A1(irdecode_inst1_next_step_6_), .A2(
        IF_DEC_instruction[6]), .Z(irdecode_inst1_N701) );
  CKAN2D2BWP12T irdecode_inst1_C5281 ( .A1(irdecode_inst1_next_step_5_), .A2(
        IF_DEC_instruction[5]), .Z(irdecode_inst1_N702) );
  CKAN2D2BWP12T irdecode_inst1_C5282 ( .A1(irdecode_inst1_next_step_4_), .A2(
        IF_DEC_instruction[4]), .Z(irdecode_inst1_N703) );
  CKAN2D2BWP12T irdecode_inst1_C5283 ( .A1(irdecode_inst1_next_step_3_), .A2(
        IF_DEC_instruction[3]), .Z(irdecode_inst1_N704) );
  CKAN2D2BWP12T irdecode_inst1_C5284 ( .A1(irdecode_inst1_next_step_2_), .A2(
        IF_DEC_instruction[2]), .Z(irdecode_inst1_N705) );
  CKAN2D2BWP12T irdecode_inst1_C5285 ( .A1(n1841), .A2(IF_DEC_instruction[1]), 
        .Z(irdecode_inst1_N706) );
  CKAN2D2BWP12T irdecode_inst1_C5286 ( .A1(irdecode_inst1_next_step_0_), .A2(
        IF_DEC_instruction[0]), .Z(irdecode_inst1_N707) );
  CKAN2D2BWP12T irdecode_inst1_C2476 ( .A1(n1841), .A2(
        irdecode_inst1_next_step_0_), .Z(irdecode_inst1_N906) );
  CKAN2D2BWP12T irdecode_inst1_C2482 ( .A1(irdecode_inst1_N907), .A2(n1854), 
        .Z(irdecode_inst1_N911) );
  OR2XD4BWP12T irdecode_inst1_C2484 ( .A1(n1841), .A2(n1854), .Z(
        irdecode_inst1_N912) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_0_ ( .D(
        MEM_MEMCTRL_from_mem_data[8]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[0]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_1_ ( .D(
        MEM_MEMCTRL_from_mem_data[9]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[1]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_2_ ( .D(
        MEM_MEMCTRL_from_mem_data[10]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_3_ ( .D(
        MEM_MEMCTRL_from_mem_data[11]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_4_ ( .D(
        MEM_MEMCTRL_from_mem_data[12]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[4]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_5_ ( .D(
        MEM_MEMCTRL_from_mem_data[13]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[5]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_6_ ( .D(
        MEM_MEMCTRL_from_mem_data[14]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_7_ ( .D(
        MEM_MEMCTRL_from_mem_data[15]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_8_ ( .D(
        MEM_MEMCTRL_from_mem_data[0]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_9_ ( .D(
        MEM_MEMCTRL_from_mem_data[1]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_10_ ( .D(
        MEM_MEMCTRL_from_mem_data[2]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_11_ ( .D(
        MEM_MEMCTRL_from_mem_data[3]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[11]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_12_ ( .D(
        MEM_MEMCTRL_from_mem_data[4]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[12]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_13_ ( .D(
        MEM_MEMCTRL_from_mem_data[5]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[13]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_14_ ( .D(
        MEM_MEMCTRL_from_mem_data[6]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[14]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_15_ ( .D(
        MEM_MEMCTRL_from_mem_data[7]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[15]) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_1_ ( .D(
        memory_interface_inst1_fsm_N33), .CP(clk), .Q(
        memory_interface_inst1_fsm_state_1_) );
  DFQD1BWP12T irdecode_inst1_load_store_width_reg_1_ ( .D(n837), .CP(clk), .Q(
        DEC_MEMCTRL_load_store_width[1]) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_0_ ( .D(
        memory_interface_inst1_fsm_N32), .CP(clk), .Q(
        memory_interface_inst1_fsm_state_0_) );
  DFQD1BWP12T irdecode_inst1_memory_load_request_reg ( .D(n861), .CP(clk), .Q(
        DEC_MEMCTRL_memory_load_request) );
  DFQD1BWP12T Instruction_Fetch_inst1_currentState_reg_1_ ( .D(
        Instruction_Fetch_inst1_N80), .CP(clk), .Q(
        Instruction_Fetch_inst1_currentState_1_) );
  DFQD1BWP12T Instruction_Fetch_inst1_currentState_reg_0_ ( .D(
        Instruction_Fetch_inst1_N79), .CP(clk), .Q(
        Instruction_Fetch_inst1_currentState_0_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_0_ ( .D(
        Instruction_Fetch_inst1_N83), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_0_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_1_ ( .D(
        Instruction_Fetch_inst1_N84), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_1_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_2_ ( .D(
        Instruction_Fetch_inst1_N85), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_2_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_3_ ( .D(
        Instruction_Fetch_inst1_N86), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_3_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_4_ ( .D(
        Instruction_Fetch_inst1_N87), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_4_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_5_ ( .D(
        Instruction_Fetch_inst1_N88), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_5_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_6_ ( .D(
        Instruction_Fetch_inst1_N89), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_6_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_7_ ( .D(
        Instruction_Fetch_inst1_N90), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_7_) );
  DFQD1BWP12T memory_interface_inst1_delayed_is_signed_reg ( .D(
        DEC_MEMCTRL_memorycontroller_sign_extend), .CP(clk), .Q(
        memory_interface_inst1_delayed_is_signed) );
  DFQD1BWP12T irdecode_inst1_step_reg_1_ ( .D(n1841), .CP(clk), .Q(
        irdecode_inst1_step[1]) );
  DFQD1BWP12T irdecode_inst1_split_instruction_reg ( .D(n847), .CP(clk), .Q(
        irdecode_inst1_split_instruction) );
  DFQD1BWP12T irdecode_inst1_step_reg_6_ ( .D(irdecode_inst1_next_step_6_), 
        .CP(clk), .Q(irdecode_inst1_step[6]) );
  DFQD1BWP12T irdecode_inst1_step_reg_5_ ( .D(irdecode_inst1_next_step_5_), 
        .CP(clk), .Q(irdecode_inst1_step[5]) );
  DFQD1BWP12T irdecode_inst1_step_reg_0_ ( .D(irdecode_inst1_next_step_0_), 
        .CP(clk), .Q(irdecode_inst1_step[0]) );
  DFQD1BWP12T irdecode_inst1_step_reg_2_ ( .D(irdecode_inst1_next_step_2_), 
        .CP(clk), .Q(irdecode_inst1_step[2]) );
  DFQD1BWP12T irdecode_inst1_step_reg_3_ ( .D(irdecode_inst1_next_step_3_), 
        .CP(clk), .Q(irdecode_inst1_step[3]) );
  DFQD1BWP12T irdecode_inst1_step_reg_4_ ( .D(irdecode_inst1_next_step_4_), 
        .CP(clk), .Q(irdecode_inst1_step[4]) );
  DFQD1BWP12T irdecode_inst1_step_reg_7_ ( .D(irdecode_inst1_next_step_7_), 
        .CP(clk), .Q(irdecode_inst1_step[7]) );
  DFQD1BWP12T irdecode_inst1_memory_store_request_reg ( .D(n852), .CP(clk), 
        .Q(DEC_MEMCTRL_memory_store_request) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_6_ ( .D(n854), .CP(clk), .Q(
        irdecode_inst1_itstate_6_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_7_ ( .D(n853), .CP(clk), .Q(
        irdecode_inst1_itstate_7_) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_0_ ( .D(n830), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[0]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_2_ ( .D(n828), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[2]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_3_ ( .D(n827), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[3]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_4_ ( .D(n826), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[4]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_0_ ( .D(n824), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[0]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_2_ ( .D(n822), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[2]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_4_ ( .D(n848), .CP(clk), .Q(
        DEC_ALU_alu_opcode[4]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_3_ ( .D(n821), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[3]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_4_ ( .D(n820), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[4]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_1_ ( .D(n850), .CP(clk), .Q(
        DEC_ALU_alu_opcode[1]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_2_ ( .D(n846), .CP(clk), .Q(
        DEC_ALU_alu_opcode[2]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_0_ ( .D(n851), .CP(clk), .Q(
        DEC_ALU_alu_opcode[0]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_3_ ( .D(n849), .CP(clk), .Q(
        DEC_ALU_alu_opcode[3]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_2_ ( .D(n818), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[2]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_3_ ( .D(n817), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[3]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_4_ ( .D(n815), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[4]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_0_ ( .D(n816), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[0]) );
  DFQD1BWP12T irdecode_inst1_memory_address_source_is_reg_reg ( .D(n836), .CP(
        clk), .Q(DEC_MISC_OUT_memory_address_source_is_reg) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_1_ ( .D(n829), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[1]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_enable_reg ( .D(n825), .CP(
        clk), .Q(DEC_RF_memory_write_to_reg_enable) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_1_ ( .D(n823), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[1]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_0_ ( .D(n809), .CP(clk), .Q(
        DEC_RF_offset_b[0]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_1_ ( .D(n808), .CP(clk), .Q(
        DEC_RF_offset_b[1]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_2_ ( .D(n807), .CP(clk), .Q(
        DEC_RF_offset_b[2]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_3_ ( .D(n806), .CP(clk), .Q(
        DEC_RF_offset_b[3]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_4_ ( .D(n805), .CP(clk), .Q(
        DEC_RF_offset_b[4]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_5_ ( .D(n804), .CP(clk), .Q(
        DEC_RF_offset_b[5]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_6_ ( .D(n803), .CP(clk), .Q(
        DEC_RF_offset_b[6]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_8_ ( .D(n801), .CP(clk), .Q(
        DEC_RF_offset_b[8]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_9_ ( .D(n800), .CP(clk), .Q(
        DEC_RF_offset_b[9]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_10_ ( .D(n799), .CP(clk), .Q(
        DEC_RF_offset_b[10]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_11_ ( .D(n798), .CP(clk), .Q(
        DEC_RF_offset_b[11]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_12_ ( .D(n797), .CP(clk), .Q(
        DEC_RF_offset_b[12]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_13_ ( .D(n796), .CP(clk), .Q(
        DEC_RF_offset_b[13]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_14_ ( .D(n795), .CP(clk), .Q(
        DEC_RF_offset_b[14]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_15_ ( .D(n794), .CP(clk), .Q(
        DEC_RF_offset_b[15]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_16_ ( .D(n793), .CP(clk), .Q(
        DEC_RF_offset_b[16]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_17_ ( .D(n792), .CP(clk), .Q(
        DEC_RF_offset_b[17]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_18_ ( .D(n791), .CP(clk), .Q(
        DEC_RF_offset_b[18]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_19_ ( .D(n790), .CP(clk), .Q(
        DEC_RF_offset_b[19]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_20_ ( .D(n789), .CP(clk), .Q(
        DEC_RF_offset_b[20]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_21_ ( .D(n788), .CP(clk), .Q(
        DEC_RF_offset_b[21]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_22_ ( .D(n787), .CP(clk), .Q(
        DEC_RF_offset_b[22]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_23_ ( .D(n786), .CP(clk), .Q(
        DEC_RF_offset_b[23]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_24_ ( .D(n785), .CP(clk), .Q(
        DEC_RF_offset_b[24]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_25_ ( .D(n784), .CP(clk), .Q(
        DEC_RF_offset_b[25]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_26_ ( .D(n783), .CP(clk), .Q(
        DEC_RF_offset_b[26]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_27_ ( .D(n782), .CP(clk), .Q(
        DEC_RF_offset_b[27]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_28_ ( .D(n781), .CP(clk), .Q(
        DEC_RF_offset_b[28]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_29_ ( .D(n780), .CP(clk), .Q(
        DEC_RF_offset_b[29]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_30_ ( .D(n779), .CP(clk), .Q(
        DEC_RF_offset_b[30]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_3_ ( .D(
        MEMCTRL_IN_address[3]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_6_ ( .D(
        MEMCTRL_IN_address[6]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_7_ ( .D(
        MEMCTRL_IN_address[7]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_8_ ( .D(
        MEMCTRL_IN_address[8]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_9_ ( .D(
        MEMCTRL_IN_address[9]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_10_ ( .D(
        MEMCTRL_IN_address[10]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_11_ ( .D(
        MEMCTRL_IN_address[11]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[11]) );
  DFQD4BWP12T memory_interface_inst1_fsm_state_reg_3_ ( .D(
        memory_interface_inst1_fsm_N35), .CP(clk), .Q(
        memory_interface_inst1_fsm_state_3_) );
  DFD4BWP12T irdecode_inst1_operand_a_reg_2_ ( .D(n813), .CP(clk), .Q(
        DEC_RF_operand_a[2]), .QN(n1000) );
  DFD4BWP12T irdecode_inst1_operand_a_reg_1_ ( .D(n814), .CP(clk), .Q(
        DEC_RF_operand_a[1]), .QN(n998) );
  DFD4BWP12T irdecode_inst1_operand_a_reg_3_ ( .D(n812), .CP(clk), .Q(
        DEC_RF_operand_a[3]), .QN(n1004) );
  DFD4BWP12T irdecode_inst1_operand_b_reg_0_ ( .D(n844), .CP(clk), .Q(
        DEC_RF_operand_b[0]) );
  DFD4BWP12T irdecode_inst1_operand_a_reg_4_ ( .D(n810), .CP(clk), .Q(
        DEC_RF_operand_a[4]), .QN(n1840) );
  DFD4BWP12T irdecode_inst1_operand_b_reg_2_ ( .D(n842), .CP(clk), .Q(
        DEC_RF_operand_b[2]), .QN(n1002) );
  DFD4BWP12T irdecode_inst1_operand_b_reg_4_ ( .D(n840), .CP(clk), .Q(
        DEC_RF_operand_b[4]), .QN(n868) );
  DFD4BWP12T irdecode_inst1_operand_b_reg_1_ ( .D(n843), .CP(clk), .Q(
        DEC_RF_operand_b[1]), .QN(n866) );
  DFD4BWP12T irdecode_inst1_operand_b_reg_3_ ( .D(n841), .CP(clk), .Q(
        DEC_RF_operand_b[3]) );
  DFXD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_0_ ( .D(
        MEMCTRL_IN_address[0]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[0]), .QN(n1847) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_21_ ( .D(
        RF_MEMCTRL_data_reg[21]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[21]) );
  DFXD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_12_ ( .D(
        Instruction_Fetch_inst1_N95), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_12_) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_5_ ( .D(
        RF_MEMCTRL_data_reg[5]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[5]) );
  DFXD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_11_ ( .D(
        Instruction_Fetch_inst1_N94), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_11_) );
  DFXD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_15_ ( .D(
        Instruction_Fetch_inst1_N98), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_15_) );
  DFXD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_13_ ( .D(
        Instruction_Fetch_inst1_N96), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_13_) );
  DFXD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_9_ ( .D(
        Instruction_Fetch_inst1_N92), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_9_) );
  DFXD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_14_ ( .D(
        Instruction_Fetch_inst1_N97), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_14_) );
  DFXD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_10_ ( .D(
        Instruction_Fetch_inst1_N93), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_10_) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_4_ ( .D(
        RF_MEMCTRL_data_reg[4]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[4]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_11_ ( .D(
        RF_MEMCTRL_data_reg[11]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[11]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_7_ ( .D(
        RF_MEMCTRL_data_reg[7]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[7]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_1_ ( .D(
        RF_MEMCTRL_data_reg[1]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[1]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_28_ ( .D(
        RF_MEMCTRL_data_reg[28]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[28]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_31_ ( .D(
        RF_MEMCTRL_data_reg[31]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[31]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_27_ ( .D(
        RF_MEMCTRL_data_reg[27]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[27]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_29_ ( .D(
        RF_MEMCTRL_data_reg[29]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[29]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_26_ ( .D(
        RF_MEMCTRL_data_reg[26]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[26]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_25_ ( .D(
        RF_MEMCTRL_data_reg[25]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[25]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_30_ ( .D(
        RF_MEMCTRL_data_reg[30]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[30]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_24_ ( .D(
        RF_MEMCTRL_data_reg[24]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[24]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_0_ ( .D(
        RF_MEMCTRL_data_reg[0]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[0]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_9_ ( .D(
        RF_MEMCTRL_data_reg[9]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[9]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_20_ ( .D(
        RF_MEMCTRL_data_reg[20]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[20]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_19_ ( .D(
        RF_MEMCTRL_data_reg[19]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[19]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_6_ ( .D(
        RF_MEMCTRL_data_reg[6]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[6]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_18_ ( .D(
        RF_MEMCTRL_data_reg[18]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[18]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_8_ ( .D(
        RF_MEMCTRL_data_reg[8]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[8]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_15_ ( .D(
        RF_MEMCTRL_data_reg[15]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[15]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_12_ ( .D(
        RF_MEMCTRL_data_reg[12]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[12]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_17_ ( .D(
        RF_MEMCTRL_data_reg[17]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[17]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_22_ ( .D(
        RF_MEMCTRL_data_reg[22]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[22]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_14_ ( .D(
        RF_MEMCTRL_data_reg[14]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[14]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_16_ ( .D(
        RF_MEMCTRL_data_reg[16]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[16]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_23_ ( .D(
        RF_MEMCTRL_data_reg[23]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[23]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_13_ ( .D(
        RF_MEMCTRL_data_reg[13]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[13]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_3_ ( .D(
        RF_MEMCTRL_data_reg[3]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[3]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_2_ ( .D(
        RF_MEMCTRL_data_reg[2]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[2]) );
  DFXD1BWP12T memory_interface_inst1_delay_data_in32_reg_10_ ( .D(
        RF_MEMCTRL_data_reg[10]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[10]) );
  DFXD1BWP12T irdecode_inst1_memory_store_address_reg_reg_1_ ( .D(n834), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[1]) );
  DFXD1BWP12T Instruction_Fetch_inst1_first_instruction_fetched_reg ( .D(n862), 
        .CP(clk), .Q(Instruction_Fetch_inst1_first_instruction_fetched) );
  DFXD1BWP12T irdecode_inst1_memorycontroller_sign_extend_reg ( .D(n839), .CP(
        clk), .Q(DEC_MEMCTRL_memorycontroller_sign_extend) );
  DFXD1BWP12T irdecode_inst1_load_store_width_reg_0_ ( .D(n838), .CP(clk), .Q(
        DEC_MEMCTRL_load_store_width[0]), .QN(n1846) );
  DFXD1BWP12T irdecode_inst1_itstate_reg_0_ ( .D(n860), .CP(clk), .Q(
        irdecode_inst1_itstate_0_) );
  DFXD1BWP12T irdecode_inst1_stall_to_instructionfetch_reg ( .D(n845), .CP(clk), .Q(DEC_IF_stall_to_instructionfetch) );
  DFXD1BWP12T irdecode_inst1_itstate_reg_5_ ( .D(n855), .CP(clk), .Q(
        irdecode_inst1_itstate_5_), .QN(n1845) );
  DFXD1BWP12T irdecode_inst1_itstate_reg_4_ ( .D(n856), .CP(clk), .Q(
        irdecode_inst1_itstate_4_) );
  DFXD1BWP12T irdecode_inst1_itstate_reg_3_ ( .D(n857), .CP(clk), .Q(
        irdecode_inst1_itstate_3_) );
  DFXD1BWP12T irdecode_inst1_itstate_reg_2_ ( .D(n858), .CP(clk), .Q(
        irdecode_inst1_itstate_2_) );
  DFXD1BWP12T irdecode_inst1_itstate_reg_1_ ( .D(n859), .CP(clk), .Q(
        irdecode_inst1_itstate_1_) );
  DFXD1BWP12T irdecode_inst1_update_flag_v_reg ( .D(
        irdecode_inst1_next_update_flag_v), .CP(clk), .Q(
        DEC_CPSR_update_flag_v), .QN(n1844) );
  DFXD1BWP12T irdecode_inst1_update_flag_c_reg ( .D(
        irdecode_inst1_next_update_flag_c), .CP(clk), .Q(
        DEC_CPSR_update_flag_c) );
  DFXD1BWP12T irdecode_inst1_alu_write_to_reg_enable_reg ( .D(
        irdecode_inst1_next_alu_write_to_reg_enable), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg_enable) );
  DFXD1BWP12T irdecode_inst1_memory_store_address_reg_reg_3_ ( .D(n832), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[3]) );
  DFXD1BWP12T irdecode_inst1_update_flag_z_reg ( .D(
        irdecode_inst1_next_update_flag_n), .CP(clk), .Q(
        DEC_CPSR_update_flag_z), .QN(n1839) );
  DFXD1BWP12T irdecode_inst1_update_flag_n_reg ( .D(
        irdecode_inst1_next_update_flag_n), .CP(clk), .Q(
        DEC_CPSR_update_flag_n), .QN(n1838) );
  DFXD1BWP12T irdecode_inst1_memory_store_address_reg_reg_2_ ( .D(n833), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[2]) );
  DFXD1BWP12T irdecode_inst1_memory_store_address_reg_reg_0_ ( .D(n835), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[0]) );
  DFXD1BWP12T irdecode_inst1_memory_store_address_reg_reg_4_ ( .D(n831), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[4]) );
  DFXD1BWP12T irdecode_inst1_alu_write_to_reg_reg_1_ ( .D(n819), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[1]) );
  DFXD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_1_ ( .D(
        MEMCTRL_IN_address[1]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[1]) );
  DFXD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_2_ ( .D(
        MEMCTRL_IN_address[2]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[2]), .QN(n1848) );
  DFXD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_4_ ( .D(
        MEMCTRL_IN_address[4]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[4]) );
  DFXD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_5_ ( .D(
        MEMCTRL_IN_address[5]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[5]) );
  DFCNQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_8_ ( .D(
        Instruction_Fetch_inst1_N91), .CP(clk), .CDN(n1837), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_8_) );
  DFMQD4BWP12T irdecode_inst1_offset_b_reg_31_ ( .DB(n864), .DA(n777), .SA(
        n1837), .CP(clk), .Q(DEC_RF_offset_b[31]) );
  DFMQD4BWP12T irdecode_inst1_operand_a_reg_0_ ( .DB(n864), .DA(n811), .SA(
        n1837), .CP(clk), .Q(DEC_RF_operand_a[0]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_7_ ( .D(n802), .CP(clk), .Q(
        DEC_RF_offset_b[7]) );
  DFQD4BWP12T memory_interface_inst1_fsm_state_reg_2_ ( .D(
        memory_interface_inst1_fsm_N34), .CP(clk), .Q(
        memory_interface_inst1_fsm_state_2_) );
  TIELBWP12T U1022 ( .ZN(n864) );
  INVD1BWP12T U1023 ( .I(n864), .ZN(MEMCTRL_MEM_to_mem_mem_enable) );
  AO21D4BWP12T U1024 ( .A1(ALU_OUT_c), .A2(DEC_CPSR_update_flag_c), .B(n1464), 
        .Z(new_c) );
  ND2XD8BWP12T U1025 ( .A1(n1013), .A2(n1017), .ZN(n1730) );
  TPND2D2BWP12T U1026 ( .A1(n1005), .A2(irdecode_inst1_N912), .ZN(n1321) );
  DCCKND4BWP12T U1027 ( .I(irdecode_inst1_N906), .ZN(n1005) );
  AO22D4BWP12T U1028 ( .A1(n1731), .A2(MEMCTRL_RF_IF_data_in[2]), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_2_), .B2(n1257), .Z(
        IF_DEC_instruction[2]) );
  AO22D4BWP12T U1029 ( .A1(n1731), .A2(MEMCTRL_RF_IF_data_in[3]), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_3_), .B2(n1257), .Z(
        IF_DEC_instruction[3]) );
  AO22XD2BWP12T U1030 ( .A1(n1731), .A2(MEMCTRL_RF_IF_data_in[6]), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_6_), .B2(n1257), .Z(
        IF_DEC_instruction[6]) );
  AO22XD2BWP12T U1031 ( .A1(n1731), .A2(MEMCTRL_RF_IF_data_in[5]), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_5_), .B2(n1257), .Z(
        IF_DEC_instruction[5]) );
  AO22D4BWP12T U1032 ( .A1(n1731), .A2(MEMCTRL_RF_IF_data_in[4]), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_4_), .B2(n1257), .Z(
        IF_DEC_instruction[4]) );
  MUX2D4BWP12T U1033 ( .I0(memory_interface_inst1_delay_first_two_bytes_out[0]), .I1(MEM_MEMCTRL_from_mem_data[8]), .S(n1730), .Z(MEMCTRL_RF_IF_data_in[0])
         );
  NR2XD3BWP12T U1034 ( .A1(irdecode_inst1_N539), .A2(irdecode_inst1_N540), 
        .ZN(n1328) );
  TPNR2D1BWP12T U1035 ( .A1(n1082), .A2(n1081), .ZN(n1630) );
  TPNR2D1BWP12T U1036 ( .A1(n1082), .A2(n1070), .ZN(n1071) );
  INVD3BWP12T U1037 ( .I(memory_interface_inst1_fsm_state_2_), .ZN(n1011) );
  AO22D4BWP12T U1038 ( .A1(n1731), .A2(MEMCTRL_RF_IF_data_in[7]), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_7_), .B2(n1257), .Z(
        IF_DEC_instruction[7]) );
  DCCKND4BWP12T U1039 ( .I(irdecode_inst1_N546), .ZN(n1632) );
  TPNR2D2BWP12T U1040 ( .A1(n1333), .A2(n1327), .ZN(n1351) );
  CKND2D2BWP12T U1041 ( .A1(n960), .A2(n1332), .ZN(n1333) );
  NR2D2BWP12T U1042 ( .A1(n1342), .A2(irdecode_inst1_N707), .ZN(n865) );
  TPNR2D1BWP12T U1043 ( .A1(n1342), .A2(irdecode_inst1_N707), .ZN(n1640) );
  CKND2D2BWP12T U1044 ( .A1(n1640), .A2(n1102), .ZN(n1642) );
  TPND2D1BWP12T U1045 ( .A1(n865), .A2(n1346), .ZN(n1641) );
  NR2D2BWP12T U1046 ( .A1(n1767), .A2(n1103), .ZN(n1370) );
  TPOAI21D1BWP12T U1047 ( .A1(n1661), .A2(n1642), .B(n1692), .ZN(n1103) );
  INR2D2BWP12T U1048 ( .A1(n1079), .B1(n1714), .ZN(n1772) );
  TPNR3D2BWP12T U1049 ( .A1(n1657), .A2(irdecode_inst1_N539), .A3(
        irdecode_inst1_N541), .ZN(n1079) );
  TPND2D2BWP12T U1050 ( .A1(n1685), .A2(n1790), .ZN(n1256) );
  NR3D2BWP12T U1051 ( .A1(n1075), .A2(n1074), .A3(n1353), .ZN(n1076) );
  INR2D2BWP12T U1052 ( .A1(n1073), .B1(n1684), .ZN(n1353) );
  TPOAI22D1BWP12T U1053 ( .A1(n1720), .A2(n1823), .B1(n1710), .B2(n1709), .ZN(
        n1711) );
  ND2D4BWP12T U1054 ( .A1(n1256), .A2(n1255), .ZN(n1841) );
  INR2D1BWP12T U1055 ( .A1(n1841), .B1(n1253), .ZN(n1248) );
  INVD3BWP12T U1056 ( .I(n1679), .ZN(n1720) );
  TPAOI21D2BWP12T U1057 ( .A1(n1256), .A2(n1255), .B(n1254), .ZN(n1679) );
  TPOAI21D1BWP12T U1058 ( .A1(n1248), .A2(n1247), .B(n1809), .ZN(n1697) );
  RCAOI211D1BWP12T U1059 ( .A1(IF_DEC_instruction[3]), .A2(n1691), .B(n1690), 
        .C(n1689), .ZN(n1695) );
  TPNR3D2BWP12T U1060 ( .A1(n1639), .A2(n1100), .A3(n1099), .ZN(n1104) );
  BUFFD6BWP12T U1061 ( .I(RF_ALU_operand_a[4]), .Z(n1852) );
  CKND0BWP12T U1062 ( .I(n866), .ZN(n867) );
  INVD1BWP12T U1063 ( .I(n868), .ZN(n869) );
  MUX2NXD1BWP12T U1064 ( .I0(MEM_MEMCTRL_from_mem_data[15]), .I1(n1225), .S(
        n1224), .ZN(n1833) );
  AN3XD0BWP12T U1065 ( .A1(n1220), .A2(MEM_MEMCTRL_from_mem_data[7]), .A3(
        memory_interface_inst1_delayed_is_signed), .Z(n1225) );
  NR2D0BWP12T U1066 ( .A1(n1223), .A2(n1222), .ZN(n1224) );
  INR2D1BWP12T U1067 ( .A1(memory_interface_inst1_delayed_is_signed), .B1(
        n1221), .ZN(n1222) );
  INR2D1BWP12T U1068 ( .A1(n1152), .B1(n1056), .ZN(n1210) );
  TPND2D1BWP12T U1069 ( .A1(n1011), .A2(n1010), .ZN(n1483) );
  INR2D1BWP12T U1070 ( .A1(n1210), .B1(n1209), .ZN(n1214) );
  IOA21D1BWP12T U1071 ( .A1(n1834), .A2(MEM_MEMCTRL_from_mem_data[0]), .B(
        n1833), .ZN(MEMCTRL_RF_IF_data_in[24]) );
  IOA21D1BWP12T U1072 ( .A1(n1834), .A2(MEM_MEMCTRL_from_mem_data[2]), .B(
        n1833), .ZN(MEMCTRL_RF_IF_data_in[26]) );
  IOA21D1BWP12T U1073 ( .A1(n1834), .A2(MEM_MEMCTRL_from_mem_data[3]), .B(
        n1833), .ZN(MEMCTRL_RF_IF_data_in[27]) );
  INVD1BWP12T U1074 ( .I(reset), .ZN(n1435) );
  AN2D1BWP12T U1075 ( .A1(n1253), .A2(n1740), .Z(n1254) );
  INR2D1BWP12T U1076 ( .A1(IF_DEC_instruction[7]), .B1(n1832), .ZN(n1723) );
  NR2D1BWP12T U1077 ( .A1(n1154), .A2(n1153), .ZN(n1779) );
  CKND0BWP12T U1078 ( .I(IF_DEC_instruction[6]), .ZN(n1823) );
  INVD1BWP12T U1079 ( .I(n1809), .ZN(n1832) );
  TPND2D1BWP12T U1080 ( .A1(n1731), .A2(n1435), .ZN(n1733) );
  INVD1BWP12T U1081 ( .I(DEC_MEMCTRL_memory_store_request), .ZN(n1580) );
  ND2D1BWP12T U1082 ( .A1(n1046), .A2(n1435), .ZN(n1364) );
  CKND0BWP12T U1083 ( .I(n1661), .ZN(n1656) );
  INVD1BWP12T U1084 ( .I(n1364), .ZN(n1836) );
  NR2D2BWP12T U1085 ( .A1(n1021), .A2(n1834), .ZN(n1109) );
  ND2D1BWP12T U1086 ( .A1(MEMCTRL_RF_IF_data_in[0]), .A2(n1731), .ZN(n1203) );
  ND2D1BWP12T U1087 ( .A1(MEMCTRL_RF_IF_data_in[1]), .A2(n1731), .ZN(n1207) );
  NR2D2BWP12T U1088 ( .A1(n1343), .A2(irdecode_inst1_N707), .ZN(n870) );
  TPND2D2BWP12T U1089 ( .A1(n870), .A2(n1102), .ZN(n1773) );
  IND2D0BWP12T U1090 ( .A1(n1492), .B1(n1534), .ZN(n1493) );
  IND2XD2BWP12T U1091 ( .A1(irdecode_inst1_N545), .B1(n1632), .ZN(n1615) );
  NR2D0BWP12T U1092 ( .A1(RF_pc_out[9]), .A2(n1286), .ZN(n871) );
  MAOI22D0BWP12T U1093 ( .A1(n871), .A2(RF_pc_out[10]), .B1(n871), .B2(
        RF_pc_out[10]), .ZN(n1513) );
  OAI21D0BWP12T U1094 ( .A1(n1441), .A2(n1281), .B(n1458), .ZN(n872) );
  AOI21D0BWP12T U1095 ( .A1(n1441), .A2(n1281), .B(n872), .ZN(
        IF_RF_incremented_pc_out[11]) );
  AO222D0BWP12T U1096 ( .A1(ALU_MISC_OUT_result[2]), .A2(n1566), .B1(n1568), 
        .B2(n1567), .C1(n1569), .C2(RF_MEMCTRL_address_reg[2]), .Z(
        MEMCTRL_IN_address[1]) );
  CKND2D0BWP12T U1097 ( .A1(DEC_RF_offset_b[15]), .A2(n1836), .ZN(n873) );
  OAI211D0BWP12T U1098 ( .A1(n1396), .A2(n1469), .B(n1696), .C(n873), .ZN(n794) );
  OAI22D0BWP12T U1099 ( .A1(n1787), .A2(n1786), .B1(n1789), .B2(n1788), .ZN(
        n874) );
  AOI22D1BWP12T U1100 ( .A1(DEC_RF_memory_write_to_reg[2]), .A2(n1836), .B1(
        n1790), .B2(n874), .ZN(n875) );
  IND3D1BWP12T U1101 ( .A1(n1792), .B1(n1791), .B2(n875), .ZN(n822) );
  ND2D1BWP12T U1102 ( .A1(n1329), .A2(irdecode_inst1_N544), .ZN(n876) );
  NR2D1BWP12T U1103 ( .A1(n1616), .A2(n876), .ZN(n1617) );
  ND3D1BWP12T U1104 ( .A1(irdecode_inst1_N703), .A2(n1349), .A3(n865), .ZN(
        n1802) );
  CKND0BWP12T U1105 ( .I(n1578), .ZN(n877) );
  AOI222D0BWP12T U1106 ( .A1(n877), .A2(RF_MEMCTRL_data_reg[22]), .B1(n1575), 
        .B2(memory_interface_inst1_delay_data_in32[6]), .C1(n1576), .C2(
        memory_interface_inst1_delay_data_in32[22]), .ZN(n878) );
  IOA21D0BWP12T U1107 ( .A1(RF_MEMCTRL_data_reg[6]), .A2(n1577), .B(n878), 
        .ZN(MEMCTRL_MEM_to_mem_data[14]) );
  AN2D0BWP12T U1108 ( .A1(n1310), .A2(n1458), .Z(IF_RF_incremented_pc_out[15])
         );
  CKND2D0BWP12T U1109 ( .A1(DEC_RF_operand_b[3]), .A2(n1836), .ZN(n879) );
  OAI211D0BWP12T U1110 ( .A1(n1823), .A2(n1613), .B(n1755), .C(n879), .ZN(n841) );
  AO222D0BWP12T U1111 ( .A1(ALU_MISC_OUT_result[12]), .A2(n1566), .B1(n1568), 
        .B2(n1482), .C1(n1569), .C2(RF_MEMCTRL_address_reg[12]), .Z(
        MEMCTRL_IN_address[11]) );
  CKND2D0BWP12T U1112 ( .A1(n1836), .A2(DEC_RF_offset_b[13]), .ZN(n880) );
  OAI211D0BWP12T U1113 ( .A1(n1783), .A2(n1469), .B(n1696), .C(n880), .ZN(n796) );
  CKND0BWP12T U1114 ( .I(MEMCTRL_RF_IF_data_in[7]), .ZN(n881) );
  MOAI22D0BWP12T U1115 ( .A1(n1733), .A2(n881), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_7_), .B2(n1732), .ZN(
        Instruction_Fetch_inst1_N90) );
  AN4D0BWP12T U1116 ( .A1(n1388), .A2(n1710), .A3(n1387), .A4(n1692), .Z(n1390) );
  TPNR2D1BWP12T U1117 ( .A1(irdecode_inst1_N543), .A2(irdecode_inst1_N542), 
        .ZN(n882) );
  TPND2D1BWP12T U1118 ( .A1(n882), .A2(n1088), .ZN(n1082) );
  INVD1BWP12T U1119 ( .I(n1372), .ZN(n883) );
  AOI21D0BWP12T U1120 ( .A1(n1718), .A2(n1162), .B(n883), .ZN(n1760) );
  MAOI22D0BWP12T U1121 ( .A1(n1836), .A2(irdecode_inst1_step[1]), .B1(n1661), 
        .B2(n1094), .ZN(n884) );
  CKND0BWP12T U1122 ( .I(n1160), .ZN(n885) );
  OA211D1BWP12T U1123 ( .A1(n1632), .A2(n1693), .B(n884), .C(n885), .Z(n1255)
         );
  CKND0BWP12T U1124 ( .I(n1509), .ZN(n886) );
  AOI222D0BWP12T U1125 ( .A1(n886), .A2(RF_MEMCTRL_data_reg[9]), .B1(
        MEM_MEMCTRL_from_mem_data[1]), .B2(n1551), .C1(n1576), .C2(
        memory_interface_inst1_delay_data_in32[25]), .ZN(n887) );
  IOA21D0BWP12T U1126 ( .A1(memory_interface_inst1_delay_data_in32[9]), .A2(
        n1506), .B(n887), .ZN(MEMCTRL_MEM_to_mem_data[1]) );
  NR2D0BWP12T U1127 ( .A1(n1287), .A2(n1457), .ZN(n888) );
  OAI21D0BWP12T U1128 ( .A1(n888), .A2(RF_pc_out[6]), .B(n1458), .ZN(n889) );
  AOI21D0BWP12T U1129 ( .A1(n888), .A2(RF_pc_out[6]), .B(n889), .ZN(
        IF_RF_incremented_pc_out[6]) );
  AO222D0BWP12T U1130 ( .A1(ALU_MISC_OUT_result[11]), .A2(n1566), .B1(n1568), 
        .B2(n1511), .C1(n1569), .C2(RF_MEMCTRL_address_reg[11]), .Z(
        MEMCTRL_IN_address[10]) );
  CKND0BWP12T U1131 ( .I(MEMCTRL_RF_IF_data_in[6]), .ZN(n890) );
  MOAI22D0BWP12T U1132 ( .A1(n1733), .A2(n890), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_6_), .B2(n1732), .ZN(
        Instruction_Fetch_inst1_N89) );
  IIND4D1BWP12T U1133 ( .A1(irdecode_inst1_N706), .A2(n1105), .B1(
        irdecode_inst1_N704), .B2(n1095), .ZN(n1774) );
  CKND2D0BWP12T U1134 ( .A1(n1625), .A2(n1633), .ZN(n891) );
  AOI21D1BWP12T U1135 ( .A1(n891), .A2(n1648), .B(n1626), .ZN(n1654) );
  CKND0BWP12T U1136 ( .I(n1578), .ZN(n892) );
  AOI222D0BWP12T U1137 ( .A1(n892), .A2(RF_MEMCTRL_data_reg[17]), .B1(n1575), 
        .B2(memory_interface_inst1_delay_data_in32[1]), .C1(n1576), .C2(
        memory_interface_inst1_delay_data_in32[17]), .ZN(n893) );
  IOA21D0BWP12T U1138 ( .A1(RF_MEMCTRL_data_reg[1]), .A2(n1577), .B(n893), 
        .ZN(MEMCTRL_MEM_to_mem_data[9]) );
  OAI21D0BWP12T U1139 ( .A1(n1457), .A2(n1287), .B(n1458), .ZN(n894) );
  AOI21D0BWP12T U1140 ( .A1(n1457), .A2(n1287), .B(n894), .ZN(
        IF_RF_incremented_pc_out[5]) );
  OAI21D0BWP12T U1141 ( .A1(n1442), .A2(RF_pc_out[12]), .B(n1458), .ZN(n895)
         );
  AOI21D0BWP12T U1142 ( .A1(n1442), .A2(RF_pc_out[12]), .B(n895), .ZN(
        IF_RF_incremented_pc_out[12]) );
  IND2D0BWP12T U1143 ( .A1(n1004), .B1(n1836), .ZN(n896) );
  OAI211D0BWP12T U1144 ( .A1(n1757), .A2(n1614), .B(n1622), .C(n896), .ZN(n812) );
  AO222D0BWP12T U1145 ( .A1(ALU_MISC_OUT_result[10]), .A2(n1566), .B1(n1568), 
        .B2(n1513), .C1(n1569), .C2(RF_MEMCTRL_address_reg[10]), .Z(
        MEMCTRL_IN_address[9]) );
  CKND2D0BWP12T U1146 ( .A1(n1836), .A2(DEC_RF_offset_b[12]), .ZN(n897) );
  OAI211D0BWP12T U1147 ( .A1(n1721), .A2(n1469), .B(n1696), .C(n897), .ZN(n797) );
  CKND0BWP12T U1148 ( .I(MEMCTRL_RF_IF_data_in[5]), .ZN(n898) );
  MOAI22D0BWP12T U1149 ( .A1(n1733), .A2(n898), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_5_), .B2(n1732), .ZN(
        Instruction_Fetch_inst1_N88) );
  IND4D0BWP12T U1150 ( .A1(n1775), .B1(n1774), .B2(n1773), .B3(n1776), .ZN(
        n899) );
  NR2D1BWP12T U1151 ( .A1(n1777), .A2(n899), .ZN(n1803) );
  NR2D0BWP12T U1152 ( .A1(RF_pc_out[3]), .A2(n1291), .ZN(n900) );
  MAOI22D0BWP12T U1153 ( .A1(RF_pc_out[4]), .A2(n900), .B1(RF_pc_out[4]), .B2(
        n900), .ZN(n1563) );
  CKND0BWP12T U1154 ( .I(n1509), .ZN(n901) );
  AOI222D0BWP12T U1155 ( .A1(n901), .A2(RF_MEMCTRL_data_reg[11]), .B1(
        MEM_MEMCTRL_from_mem_data[3]), .B2(n1551), .C1(n1576), .C2(
        memory_interface_inst1_delay_data_in32[27]), .ZN(n902) );
  IOA21D0BWP12T U1156 ( .A1(memory_interface_inst1_delay_data_in32[11]), .A2(
        n1506), .B(n902), .ZN(MEMCTRL_MEM_to_mem_data[3]) );
  AO222D0BWP12T U1157 ( .A1(ALU_MISC_OUT_result[9]), .A2(n1566), .B1(n1568), 
        .B2(n1516), .C1(n1569), .C2(RF_MEMCTRL_address_reg[9]), .Z(
        MEMCTRL_IN_address[8]) );
  OAI22D0BWP12T U1158 ( .A1(n1713), .A2(n1788), .B1(n1712), .B2(n1823), .ZN(
        n903) );
  AOI21D0BWP12T U1159 ( .A1(n1722), .A2(n1714), .B(n903), .ZN(n904) );
  CKND2D0BWP12T U1160 ( .A1(n1715), .A2(IF_DEC_instruction[0]), .ZN(n905) );
  OAI211D1BWP12T U1161 ( .A1(n1783), .A2(n1720), .B(n904), .C(n905), .ZN(n906)
         );
  AO222D1BWP12T U1162 ( .A1(n906), .A2(n1809), .B1(n1735), .B2(n1723), .C1(
        n1836), .C2(DEC_RF_offset_b[2]), .Z(n807) );
  CKND0BWP12T U1163 ( .I(MEMCTRL_RF_IF_data_in[4]), .ZN(n907) );
  MOAI22D0BWP12T U1164 ( .A1(n1733), .A2(n907), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_4_), .B2(n1732), .ZN(
        Instruction_Fetch_inst1_N87) );
  IND4D1BWP12T U1165 ( .A1(n1105), .B1(irdecode_inst1_N706), .B2(n1344), .B3(
        n1095), .ZN(n1799) );
  IND3D0BWP12T U1166 ( .A1(n1801), .B1(n1618), .B2(n1642), .ZN(n1624) );
  NR2D0BWP12T U1167 ( .A1(n1361), .A2(n1669), .ZN(n908) );
  CKND2D0BWP12T U1168 ( .A1(n908), .A2(n1151), .ZN(n1191) );
  IND2D1BWP12T U1169 ( .A1(n1082), .B1(irdecode_inst1_N540), .ZN(n1657) );
  CKND0BWP12T U1170 ( .I(n1578), .ZN(n909) );
  AOI222D0BWP12T U1171 ( .A1(n909), .A2(RF_MEMCTRL_data_reg[19]), .B1(n1575), 
        .B2(memory_interface_inst1_delay_data_in32[3]), .C1(n1576), .C2(
        memory_interface_inst1_delay_data_in32[19]), .ZN(n910) );
  IOA21D0BWP12T U1172 ( .A1(RF_MEMCTRL_data_reg[3]), .A2(n1577), .B(n910), 
        .ZN(MEMCTRL_MEM_to_mem_data[11]) );
  OAI21D0BWP12T U1173 ( .A1(n1314), .A2(RF_pc_out[3]), .B(n1458), .ZN(n911) );
  AOI21D0BWP12T U1174 ( .A1(n1314), .A2(RF_pc_out[3]), .B(n911), .ZN(
        IF_RF_incremented_pc_out[3]) );
  NR2D0BWP12T U1175 ( .A1(n1446), .A2(n1447), .ZN(n912) );
  OAI21D0BWP12T U1176 ( .A1(n912), .A2(RF_pc_out[14]), .B(n1458), .ZN(n913) );
  AOI21D0BWP12T U1177 ( .A1(n912), .A2(RF_pc_out[14]), .B(n913), .ZN(
        IF_RF_incremented_pc_out[14]) );
  AO222D0BWP12T U1178 ( .A1(ALU_MISC_OUT_result[8]), .A2(n1566), .B1(n1568), 
        .B2(n1521), .C1(n1569), .C2(RF_MEMCTRL_address_reg[8]), .Z(
        MEMCTRL_IN_address[7]) );
  CKND2D0BWP12T U1179 ( .A1(DEC_RF_alu_write_to_reg[3]), .A2(n1836), .ZN(n914)
         );
  OAI211D0BWP12T U1180 ( .A1(n1757), .A2(n1623), .B(n1622), .C(n914), .ZN(n817) );
  CKND0BWP12T U1181 ( .I(MEMCTRL_RF_IF_data_in[3]), .ZN(n915) );
  MOAI22D0BWP12T U1182 ( .A1(n1733), .A2(n915), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_3_), .B2(n1732), .ZN(
        Instruction_Fetch_inst1_N86) );
  INR3D0BWP12T U1183 ( .A1(irdecode_inst1_N701), .B1(irdecode_inst1_N702), 
        .B2(n1347), .ZN(n1348) );
  AN2D0BWP12T U1184 ( .A1(n1458), .A2(n1427), .Z(IF_RF_incremented_pc_out[26])
         );
  NR2D0BWP12T U1185 ( .A1(n1616), .A2(n1615), .ZN(n916) );
  CKND2D0BWP12T U1186 ( .A1(n1636), .A2(n916), .ZN(n1620) );
  CKND0BWP12T U1187 ( .I(n1509), .ZN(n917) );
  AOI222D0BWP12T U1188 ( .A1(n917), .A2(RF_MEMCTRL_data_reg[10]), .B1(
        MEM_MEMCTRL_from_mem_data[2]), .B2(n1551), .C1(n1576), .C2(
        memory_interface_inst1_delay_data_in32[26]), .ZN(n918) );
  IOA21D0BWP12T U1189 ( .A1(memory_interface_inst1_delay_data_in32[10]), .A2(
        n1506), .B(n918), .ZN(MEMCTRL_MEM_to_mem_data[2]) );
  CKND2D0BWP12T U1190 ( .A1(n1836), .A2(DEC_RF_offset_b[11]), .ZN(n919) );
  OAI211D1BWP12T U1191 ( .A1(n1787), .A2(n1697), .B(n1696), .C(n919), .ZN(n798) );
  CKND2D0BWP12T U1192 ( .A1(n1402), .A2(n1384), .ZN(n920) );
  AOI211D0BWP12T U1193 ( .A1(n1714), .A2(n1406), .B(n1597), .C(n920), .ZN(n921) );
  AOI31D0BWP12T U1194 ( .A1(n921), .A2(n1386), .A3(n1385), .B(n1757), .ZN(n922) );
  AO211D1BWP12T U1195 ( .A1(DEC_ALU_alu_opcode[2]), .A2(n1836), .B(n922), .C(
        n1761), .Z(n846) );
  AN2D0BWP12T U1196 ( .A1(n1568), .A2(n1428), .Z(n1842) );
  CKND0BWP12T U1197 ( .I(n1669), .ZN(n923) );
  ND4D1BWP12T U1198 ( .A1(n1687), .A2(n1672), .A3(n1671), .A4(n1778), .ZN(n924) );
  AOI211D0BWP12T U1199 ( .A1(n1745), .A2(n923), .B(n1744), .C(n924), .ZN(n1828) );
  AN3XD1BWP12T U1200 ( .A1(n925), .A2(n865), .A3(irdecode_inst1_N702), .Z(
        n1658) );
  CKND0BWP12T U1201 ( .I(n1347), .ZN(n925) );
  CKND0BWP12T U1202 ( .I(n1578), .ZN(n926) );
  AOI222D0BWP12T U1203 ( .A1(n926), .A2(RF_MEMCTRL_data_reg[18]), .B1(n1575), 
        .B2(memory_interface_inst1_delay_data_in32[2]), .C1(n1576), .C2(
        memory_interface_inst1_delay_data_in32[18]), .ZN(n927) );
  IOA21D0BWP12T U1204 ( .A1(RF_MEMCTRL_data_reg[2]), .A2(n1577), .B(n927), 
        .ZN(MEMCTRL_MEM_to_mem_data[10]) );
  MAOI22D0BWP12T U1205 ( .A1(memory_interface_inst1_delay_addr_for_adder[9]), 
        .A2(n1515), .B1(memory_interface_inst1_delay_addr_for_adder[9]), .B2(
        n1514), .ZN(n928) );
  AO21D0BWP12T U1206 ( .A1(MEMCTRL_IN_address[9]), .A2(n1574), .B(n928), .Z(
        MEMCTRL_MEM_to_mem_address[9]) );
  AO222D0BWP12T U1207 ( .A1(ALU_MISC_OUT_result[7]), .A2(n1566), .B1(n1568), 
        .B2(n1527), .C1(n1569), .C2(RF_MEMCTRL_address_reg[7]), .Z(
        MEMCTRL_IN_address[6]) );
  CKND0BWP12T U1208 ( .I(MEMCTRL_RF_IF_data_in[2]), .ZN(n929) );
  MOAI22D0BWP12T U1209 ( .A1(n1733), .A2(n929), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_2_), .B2(n1732), .ZN(
        Instruction_Fetch_inst1_N85) );
  CKND0BWP12T U1210 ( .I(n1620), .ZN(n930) );
  CKND2D0BWP12T U1211 ( .A1(irdecode_inst1_step[2]), .A2(n1836), .ZN(n931) );
  OAI211D0BWP12T U1212 ( .A1(n1693), .A2(n930), .B(n1621), .C(n931), .ZN(
        irdecode_inst1_next_step_2_) );
  IND4D0BWP12T U1213 ( .A1(n1306), .B1(RF_pc_out[16]), .B2(RF_pc_out[15]), 
        .B3(n1305), .ZN(n932) );
  NR2D1BWP12T U1214 ( .A1(n1239), .A2(n932), .ZN(n1230) );
  IND2XD2BWP12T U1215 ( .A1(n1355), .B1(n1799), .ZN(n1639) );
  IND2D0BWP12T U1216 ( .A1(n1534), .B1(n1492), .ZN(n1578) );
  AN2D0BWP12T U1217 ( .A1(n1458), .A2(n1219), .Z(IF_RF_incremented_pc_out[28])
         );
  AO222D1BWP12T U1218 ( .A1(ALU_MISC_OUT_result[4]), .A2(n1566), .B1(n1568), 
        .B2(n1563), .C1(n1569), .C2(RF_MEMCTRL_address_reg[4]), .Z(
        MEMCTRL_IN_address[3]) );
  CKND2D0BWP12T U1219 ( .A1(n1836), .A2(DEC_RF_offset_b[10]), .ZN(n933) );
  OAI211D1BWP12T U1220 ( .A1(n1822), .A2(n1697), .B(n1696), .C(n933), .ZN(n799) );
  CKND0BWP12T U1221 ( .I(MEMCTRL_RF_IF_data_in[1]), .ZN(n934) );
  MOAI22D0BWP12T U1222 ( .A1(n1733), .A2(n934), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_1_), .B2(n1732), .ZN(
        Instruction_Fetch_inst1_N84) );
  MAOI22D0BWP12T U1223 ( .A1(n1836), .A2(irdecode_inst1_step[3]), .B1(n1661), 
        .B2(n1619), .ZN(n935) );
  OAI211D0BWP12T U1224 ( .A1(n1693), .A2(n1625), .B(n935), .C(n1621), .ZN(
        irdecode_inst1_next_step_3_) );
  NR2D0BWP12T U1225 ( .A1(n1331), .A2(n1330), .ZN(n936) );
  CKND2D0BWP12T U1226 ( .A1(n936), .A2(n1332), .ZN(n1633) );
  NR2D1BWP12T U1227 ( .A1(n1343), .A2(irdecode_inst1_N706), .ZN(n937) );
  ND2D1BWP12T U1228 ( .A1(n937), .A2(n865), .ZN(n1619) );
  CKND0BWP12T U1229 ( .I(n1578), .ZN(n938) );
  AOI222D0BWP12T U1230 ( .A1(n938), .A2(RF_MEMCTRL_data_reg[21]), .B1(n1575), 
        .B2(memory_interface_inst1_delay_data_in32[5]), .C1(n1576), .C2(
        memory_interface_inst1_delay_data_in32[21]), .ZN(n939) );
  IOA21D0BWP12T U1231 ( .A1(n1577), .A2(RF_MEMCTRL_data_reg[5]), .B(n939), 
        .ZN(MEMCTRL_MEM_to_mem_data[13]) );
  AN2D0BWP12T U1232 ( .A1(RF_pc_out[3]), .A2(n1314), .Z(n940) );
  OAI21D0BWP12T U1233 ( .A1(n940), .A2(RF_pc_out[4]), .B(n1458), .ZN(n941) );
  AOI21D0BWP12T U1234 ( .A1(n940), .A2(RF_pc_out[4]), .B(n941), .ZN(
        IF_RF_incremented_pc_out[4]) );
  NR2D0BWP12T U1235 ( .A1(n1832), .A2(n1823), .ZN(n942) );
  AOI22D0BWP12T U1236 ( .A1(n942), .A2(n1715), .B1(n1836), .B2(
        DEC_RF_offset_b[8]), .ZN(n943) );
  OAI21D0BWP12T U1237 ( .A1(n1720), .A2(n1674), .B(n943), .ZN(n801) );
  CKND0BWP12T U1238 ( .I(DEC_RF_memory_store_data_reg[2]), .ZN(n944) );
  CKND2D0BWP12T U1239 ( .A1(n1779), .A2(n1361), .ZN(n945) );
  OAI211D0BWP12T U1240 ( .A1(n1788), .A2(n1362), .B(n1830), .C(n945), .ZN(n946) );
  OAI31D0BWP12T U1241 ( .A1(n1367), .A2(n1810), .A3(n946), .B(n1790), .ZN(n947) );
  OAI211D1BWP12T U1242 ( .A1(n1364), .A2(n944), .B(n1791), .C(n947), .ZN(n828)
         );
  IND4D0BWP12T U1243 ( .A1(n1449), .B1(n1448), .B2(RF_pc_out[8]), .B3(
        RF_pc_out[7]), .ZN(n1239) );
  CKND0BWP12T U1244 ( .I(n1328), .ZN(n948) );
  INVD1BWP12T U1245 ( .I(n1633), .ZN(n949) );
  AOI211D0BWP12T U1246 ( .A1(n1351), .A2(n948), .B(n1617), .C(n949), .ZN(n1769) );
  CKND2D0BWP12T U1247 ( .A1(n1586), .A2(n1579), .ZN(n950) );
  NR2D0BWP12T U1248 ( .A1(n1484), .A2(n950), .ZN(n1562) );
  AN2D0BWP12T U1249 ( .A1(n1568), .A2(n1425), .Z(n1843) );
  INR2D1BWP12T U1250 ( .A1(n1188), .B1(n1320), .ZN(n1794) );
  OAI21D0BWP12T U1251 ( .A1(DEC_IF_stall_to_instructionfetch), .A2(
        Instruction_Fetch_inst1_currentState_1_), .B(
        Instruction_Fetch_inst1_currentState_0_), .ZN(n951) );
  AOI32D0BWP12T U1252 ( .A1(n1302), .A2(n1733), .A3(n951), .B1(reset), .B2(
        n1733), .ZN(Instruction_Fetch_inst1_N79) );
  AOI22D0BWP12T U1253 ( .A1(n1659), .A2(n1656), .B1(n1836), .B2(
        irdecode_inst1_step[5]), .ZN(n952) );
  OAI211D0BWP12T U1254 ( .A1(n1693), .A2(n1628), .B(n952), .C(n1654), .ZN(
        irdecode_inst1_next_step_5_) );
  IND2D1BWP12T U1255 ( .A1(n1306), .B1(n1443), .ZN(n1309) );
  OR2D0BWP12T U1256 ( .A1(n1231), .A2(n1237), .Z(n953) );
  OAI21D0BWP12T U1257 ( .A1(n1232), .A2(n953), .B(n1458), .ZN(n954) );
  AOI21D0BWP12T U1258 ( .A1(n1232), .A2(n953), .B(n954), .ZN(
        IF_RF_incremented_pc_out[19]) );
  INR2D1BWP12T U1259 ( .A1(n1740), .B1(n1670), .ZN(n1687) );
  NR2D0BWP12T U1260 ( .A1(n1814), .A2(n1320), .ZN(n955) );
  OAI21D0BWP12T U1261 ( .A1(n955), .A2(n1683), .B(n1470), .ZN(n1748) );
  CKND2D0BWP12T U1262 ( .A1(n1615), .A2(n1332), .ZN(n956) );
  OAI211D1BWP12T U1263 ( .A1(n1655), .A2(n1333), .B(n1769), .C(n956), .ZN(
        n1818) );
  IND3D1BWP12T U1264 ( .A1(n1011), .B1(memory_interface_inst1_fsm_state_3_), 
        .B2(n1015), .ZN(n1485) );
  OAI21D0BWP12T U1265 ( .A1(n1456), .A2(RF_pc_out[7]), .B(n1458), .ZN(n957) );
  AOI21D0BWP12T U1266 ( .A1(n1456), .A2(RF_pc_out[7]), .B(n957), .ZN(
        IF_RF_incremented_pc_out[7]) );
  CKND0BWP12T U1267 ( .I(MEMCTRL_RF_IF_data_in[0]), .ZN(n958) );
  MOAI22D0BWP12T U1268 ( .A1(n1733), .A2(n958), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_0_), .B2(n1732), .ZN(
        Instruction_Fetch_inst1_N83) );
  OA211D0BWP12T U1269 ( .A1(n1301), .A2(DEC_IF_stall_to_instructionfetch), .B(
        n1300), .C(n1302), .Z(n959) );
  NR2D0BWP12T U1270 ( .A1(reset), .A2(n959), .ZN(Instruction_Fetch_inst1_N80)
         );
  TPNR2D2BWP12T U1271 ( .A1(n1331), .A2(irdecode_inst1_N543), .ZN(n960) );
  NR2D1BWP12T U1272 ( .A1(n1094), .A2(irdecode_inst1_N705), .ZN(n961) );
  ND2D1BWP12T U1273 ( .A1(n961), .A2(n1102), .ZN(n1798) );
  OAI21D1BWP12T U1274 ( .A1(n1266), .A2(RF_pc_out[31]), .B(n1458), .ZN(n962)
         );
  AOI21D1BWP12T U1275 ( .A1(n1266), .A2(RF_pc_out[31]), .B(n962), .ZN(
        IF_RF_incremented_pc_out[31]) );
  NR3D0BWP12T U1276 ( .A1(n1197), .A2(n1826), .A3(n1163), .ZN(n963) );
  ND4D1BWP12T U1277 ( .A1(n1603), .A2(n1470), .A3(n1378), .A4(n963), .ZN(n1367) );
  CKND0BWP12T U1278 ( .I(n1578), .ZN(n964) );
  AOI222D0BWP12T U1279 ( .A1(n964), .A2(RF_MEMCTRL_data_reg[16]), .B1(n1575), 
        .B2(memory_interface_inst1_delay_data_in32[0]), .C1(n1576), .C2(
        memory_interface_inst1_delay_data_in32[16]), .ZN(n965) );
  IOA21D0BWP12T U1280 ( .A1(RF_MEMCTRL_data_reg[0]), .A2(n1577), .B(n965), 
        .ZN(MEMCTRL_MEM_to_mem_data[8]) );
  NR2D0BWP12T U1281 ( .A1(n1572), .A2(
        memory_interface_inst1_delay_addr_for_adder[3]), .ZN(n966) );
  AO222D0BWP12T U1282 ( .A1(n1564), .A2(n966), .B1(MEMCTRL_IN_address[3]), 
        .B2(n1574), .C1(n1565), .C2(
        memory_interface_inst1_delay_addr_for_adder[3]), .Z(
        MEMCTRL_MEM_to_mem_address[3]) );
  CKND0BWP12T U1283 ( .I(n1446), .ZN(n967) );
  OAI21D0BWP12T U1284 ( .A1(n1443), .A2(n967), .B(n1458), .ZN(n968) );
  AOI21D0BWP12T U1285 ( .A1(n1443), .A2(n967), .B(n968), .ZN(
        IF_RF_incremented_pc_out[13]) );
  CKND2D0BWP12T U1286 ( .A1(irdecode_inst1_step[4]), .A2(n1836), .ZN(n969) );
  OAI211D0BWP12T U1287 ( .A1(n1627), .A2(n1661), .B(n1654), .C(n969), .ZN(
        irdecode_inst1_next_step_4_) );
  OAI21D0BWP12T U1288 ( .A1(n1304), .A2(n1303), .B(n1458), .ZN(n970) );
  AOI21D0BWP12T U1289 ( .A1(n1304), .A2(n1303), .B(n970), .ZN(
        IF_RF_incremented_pc_out[24]) );
  CKND0BWP12T U1290 ( .I(n1578), .ZN(n971) );
  AOI222D0BWP12T U1291 ( .A1(n971), .A2(RF_MEMCTRL_data_reg[20]), .B1(n1575), 
        .B2(memory_interface_inst1_delay_data_in32[4]), .C1(n1576), .C2(
        memory_interface_inst1_delay_data_in32[20]), .ZN(n972) );
  IOA21D0BWP12T U1292 ( .A1(RF_MEMCTRL_data_reg[4]), .A2(n1577), .B(n972), 
        .ZN(MEMCTRL_MEM_to_mem_data[12]) );
  OAI21D0BWP12T U1293 ( .A1(n1307), .A2(RF_pc_out[16]), .B(n1458), .ZN(n973)
         );
  AOI21D0BWP12T U1294 ( .A1(n1307), .A2(RF_pc_out[16]), .B(n973), .ZN(
        IF_RF_incremented_pc_out[16]) );
  AOI21D0BWP12T U1295 ( .A1(n1822), .A2(n1821), .B(n1820), .ZN(n974) );
  OAI22D0BWP12T U1296 ( .A1(n1824), .A2(n1823), .B1(n1825), .B2(n974), .ZN(
        n975) );
  AOI21D0BWP12T U1297 ( .A1(n1826), .A2(n1827), .B(n975), .ZN(n976) );
  OAI211D0BWP12T U1298 ( .A1(n1830), .A2(n1829), .B(n1828), .C(n976), .ZN(n977) );
  AOI31D0BWP12T U1299 ( .A1(n1831), .A2(n1841), .A3(n1854), .B(n977), .ZN(n978) );
  MOAI22D0BWP12T U1300 ( .A1(n1832), .A2(n978), .B1(DEC_ALU_alu_opcode[0]), 
        .B2(n1836), .ZN(n851) );
  NR2D0BWP12T U1301 ( .A1(n1659), .A2(n1658), .ZN(n979) );
  CKND2D0BWP12T U1302 ( .A1(irdecode_inst1_step[6]), .A2(n1836), .ZN(n980) );
  OAI211D1BWP12T U1303 ( .A1(n979), .A2(n1661), .B(n1660), .C(n980), .ZN(
        irdecode_inst1_next_step_6_) );
  TPNR2D1BWP12T U1304 ( .A1(n1304), .A2(n1303), .ZN(n981) );
  ND2D1BWP12T U1305 ( .A1(n981), .A2(RF_pc_out[25]), .ZN(n1426) );
  MAOI22D0BWP12T U1306 ( .A1(n981), .A2(RF_pc_out[25]), .B1(n981), .B2(
        RF_pc_out[25]), .ZN(n1428) );
  IND2D1BWP12T U1307 ( .A1(n1240), .B1(n1454), .ZN(n1441) );
  OAI21D0BWP12T U1308 ( .A1(n1227), .A2(n1226), .B(n1458), .ZN(n982) );
  AOI21D0BWP12T U1309 ( .A1(n1227), .A2(n1226), .B(n982), .ZN(
        IF_RF_incremented_pc_out[22]) );
  TPNR2D1BWP12T U1310 ( .A1(n1078), .A2(irdecode_inst1_N543), .ZN(n983) );
  TPND2D1BWP12T U1311 ( .A1(n983), .A2(n1088), .ZN(n1628) );
  CKND0BWP12T U1312 ( .I(n1578), .ZN(n984) );
  AOI222D0BWP12T U1313 ( .A1(n984), .A2(RF_MEMCTRL_data_reg[23]), .B1(n1575), 
        .B2(memory_interface_inst1_delay_data_in32[7]), .C1(n1576), .C2(
        memory_interface_inst1_delay_data_in32[23]), .ZN(n985) );
  IOA21D0BWP12T U1314 ( .A1(RF_MEMCTRL_data_reg[7]), .A2(n1577), .B(n985), 
        .ZN(MEMCTRL_MEM_to_mem_data[15]) );
  CKND0BWP12T U1315 ( .I(MEMCTRL_IN_address[10]), .ZN(n986) );
  CKND2D0BWP12T U1316 ( .A1(memory_interface_inst1_delay_addr_for_adder[9]), 
        .A2(n1514), .ZN(n987) );
  OAI22D0BWP12T U1317 ( .A1(n1562), .A2(n986), .B1(
        memory_interface_inst1_delay_addr_for_adder[10]), .B2(n987), .ZN(n988)
         );
  AO21D0BWP12T U1318 ( .A1(memory_interface_inst1_delay_addr_for_adder[10]), 
        .A2(n1512), .B(n988), .Z(MEMCTRL_MEM_to_mem_address[10]) );
  CKND2D0BWP12T U1319 ( .A1(n1828), .A2(n1829), .ZN(n989) );
  NR4D0BWP12T U1320 ( .A1(n1673), .A2(n1826), .A3(n1685), .A4(n989), .ZN(n990)
         );
  MOAI22D0BWP12T U1321 ( .A1(n990), .A2(n1832), .B1(n1836), .B2(
        DEC_ALU_alu_opcode[4]), .ZN(n848) );
  NR2D0BWP12T U1322 ( .A1(n1572), .A2(n1486), .ZN(n1514) );
  OAI21D0BWP12T U1323 ( .A1(n1437), .A2(RF_pc_out[23]), .B(n1458), .ZN(n991)
         );
  AOI21D0BWP12T U1324 ( .A1(n1437), .A2(RF_pc_out[23]), .B(n991), .ZN(
        IF_RF_incremented_pc_out[23]) );
  MAOI22D0BWP12T U1325 ( .A1(n1228), .A2(RF_pc_out[21]), .B1(n1228), .B2(
        RF_pc_out[21]), .ZN(n1229) );
  CKND0BWP12T U1326 ( .I(n1745), .ZN(n992) );
  OAI21D0BWP12T U1327 ( .A1(n1714), .A2(n992), .B(n1596), .ZN(n1753) );
  IND2D0BWP12T U1328 ( .A1(n1794), .B1(n1789), .ZN(n1810) );
  INR2D0BWP12T U1329 ( .A1(n1459), .B1(n1460), .ZN(MEMCTRL_IN_address[0]) );
  CKND0BWP12T U1330 ( .I(n1836), .ZN(n993) );
  OAI21D0BWP12T U1331 ( .A1(n1840), .A2(n993), .B(n1835), .ZN(n810) );
  AOI211D0BWP12T U1332 ( .A1(n1350), .A2(n1830), .B(n1775), .C(n1815), .ZN(
        n994) );
  NR2D0BWP12T U1333 ( .A1(n1778), .A2(n994), .ZN(n995) );
  NR4D0BWP12T U1334 ( .A1(n1363), .A2(n1366), .A3(n995), .A4(n1784), .ZN(n996)
         );
  OAI22D0BWP12T U1335 ( .A1(n1580), .A2(n1364), .B1(n996), .B2(n1832), .ZN(
        n852) );
  AOI21D0BWP12T U1336 ( .A1(n1836), .A2(irdecode_inst1_step[7]), .B(n1656), 
        .ZN(n997) );
  OAI211D0BWP12T U1337 ( .A1(n1693), .A2(n1657), .B(n1660), .C(n997), .ZN(
        irdecode_inst1_next_step_7_) );
  AOI22D0BWP12T U1338 ( .A1(n1200), .A2(n1790), .B1(n1836), .B2(
        DEC_RF_operand_b[0]), .ZN(n1201) );
  INVD1BWP12T U1339 ( .I(n998), .ZN(n999) );
  INVD1BWP12T U1340 ( .I(n1000), .ZN(n1001) );
  INVD1BWP12T U1341 ( .I(n1002), .ZN(n1003) );
  BUFFXD12BWP12T U1342 ( .I(RF_ALU_operand_a[17]), .Z(n1853) );
  TPNR2D2BWP12T U1343 ( .A1(n1247), .A2(n1249), .ZN(n1740) );
  TPNR2D3BWP12T U1344 ( .A1(n1160), .A2(n1159), .ZN(n1854) );
  IOA21D2BWP12T U1345 ( .A1(RF_OUT_n), .A2(n1838), .B(n1465), .ZN(new_n) );
  TPND2D2BWP12T U1346 ( .A1(ALU_OUT_n), .A2(DEC_CPSR_update_flag_n), .ZN(n1465) );
  TIEHBWP12T U1347 ( .Z(n1837) );
  BUFFXD16BWP12T U1348 ( .I(RF_ALU_operand_a[1]), .Z(n1851) );
  INR2D1BWP12T U1349 ( .A1(memory_interface_inst1_fsm_state_0_), .B1(
        memory_interface_inst1_fsm_state_1_), .ZN(n1015) );
  INR2D1BWP12T U1350 ( .A1(memory_interface_inst1_fsm_state_3_), .B1(n1015), 
        .ZN(n1008) );
  INR2D2BWP12T U1351 ( .A1(memory_interface_inst1_fsm_state_2_), .B1(
        memory_interface_inst1_fsm_state_1_), .ZN(n1013) );
  INR2D2BWP12T U1352 ( .A1(memory_interface_inst1_fsm_state_1_), .B1(
        memory_interface_inst1_fsm_state_2_), .ZN(n1018) );
  TPNR2D0BWP12T U1353 ( .A1(n1013), .A2(n1018), .ZN(n1006) );
  INVD1BWP12T U1354 ( .I(memory_interface_inst1_fsm_state_0_), .ZN(n1012) );
  MUX2D1BWP12T U1355 ( .I0(n1011), .I1(n1006), .S(n1012), .Z(n1007) );
  INR2D2BWP12T U1356 ( .A1(n1008), .B1(n1007), .ZN(n1484) );
  CKND2D1BWP12T U1357 ( .A1(n1018), .A2(memory_interface_inst1_fsm_state_0_), 
        .ZN(n1444) );
  CKND2D2BWP12T U1358 ( .A1(n1485), .A2(n1444), .ZN(n1009) );
  TPNR2D2BWP12T U1359 ( .A1(n1484), .A2(n1009), .ZN(n1478) );
  INVD1P75BWP12T U1360 ( .I(memory_interface_inst1_fsm_state_3_), .ZN(n1010)
         );
  INVD1P75BWP12T U1361 ( .I(n1483), .ZN(n1014) );
  INR2D2BWP12T U1362 ( .A1(n1014), .B1(memory_interface_inst1_fsm_state_1_), 
        .ZN(n1220) );
  CKND2D2BWP12T U1363 ( .A1(n1220), .A2(n1012), .ZN(n1579) );
  TPND2D2BWP12T U1364 ( .A1(n1478), .A2(n1579), .ZN(n1223) );
  TPNR2D3BWP12T U1365 ( .A1(memory_interface_inst1_fsm_state_0_), .A2(
        memory_interface_inst1_fsm_state_3_), .ZN(n1017) );
  ND2D1BWP12T U1366 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  ND2D2BWP12T U1367 ( .A1(n1730), .A2(n1016), .ZN(n1025) );
  TPNR2D1BWP12T U1368 ( .A1(n1223), .A2(n1025), .ZN(n1021) );
  INVD4BWP12T U1369 ( .I(n1730), .ZN(n1834) );
  TPND2D0BWP12T U1370 ( .A1(n1109), .A2(MEM_MEMCTRL_from_mem_data[7]), .ZN(
        n1023) );
  TPND2D0BWP12T U1371 ( .A1(n1834), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[15]), .ZN(n1022) );
  CKND2D2BWP12T U1372 ( .A1(n1018), .A2(n1017), .ZN(n1221) );
  TPNR2D0BWP12T U1373 ( .A1(n1221), .A2(
        memory_interface_inst1_delayed_is_signed), .ZN(n1019) );
  TPNR2D1BWP12T U1374 ( .A1(n1019), .A2(MEM_MEMCTRL_from_mem_data[15]), .ZN(
        n1020) );
  TPND2D2BWP12T U1375 ( .A1(n1021), .A2(n1020), .ZN(n1111) );
  ND3D1BWP12T U1376 ( .A1(n1023), .A2(n1022), .A3(n1111), .ZN(
        MEMCTRL_RF_IF_data_in[15]) );
  INVD1P75BWP12T U1377 ( .I(Instruction_Fetch_inst1_currentState_1_), .ZN(
        n1024) );
  OR2XD4BWP12T U1378 ( .A1(n1024), .A2(Instruction_Fetch_inst1_currentState_0_), .Z(n1026) );
  INVD3BWP12T U1379 ( .I(n1026), .ZN(n1568) );
  INVD1P75BWP12T U1380 ( .I(n1568), .ZN(n1460) );
  INVD4BWP12T U1381 ( .I(n1460), .ZN(n1458) );
  INR2D4BWP12T U1382 ( .A1(Instruction_Fetch_inst1_currentState_0_), .B1(
        Instruction_Fetch_inst1_currentState_1_), .ZN(n1257) );
  INR2D4BWP12T U1383 ( .A1(n1221), .B1(n1025), .ZN(n1586) );
  TPNR2D8BWP12T U1384 ( .A1(n1586), .A2(n1026), .ZN(n1731) );
  INVD6BWP12T U1385 ( .I(n1731), .ZN(n754) );
  INVD3BWP12T U1386 ( .I(n1257), .ZN(n1301) );
  ND2D4BWP12T U1387 ( .A1(n754), .A2(n1301), .ZN(n1300) );
  IOA21D1BWP12T U1388 ( .A1(n1257), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_15_), .B(n1300), .ZN(
        n1027) );
  AO21D2BWP12T U1389 ( .A1(MEMCTRL_RF_IF_data_in[15]), .A2(n1458), .B(n1027), 
        .Z(n1149) );
  TPND2D0BWP12T U1390 ( .A1(n1109), .A2(MEM_MEMCTRL_from_mem_data[5]), .ZN(
        n1029) );
  CKND2D1BWP12T U1391 ( .A1(n1834), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[13]), .ZN(n1028) );
  ND3D1BWP12T U1392 ( .A1(n1029), .A2(n1111), .A3(n1028), .ZN(
        MEMCTRL_RF_IF_data_in[13]) );
  ND2D1BWP12T U1393 ( .A1(MEMCTRL_RF_IF_data_in[13]), .A2(n1568), .ZN(n1032)
         );
  INVD1P75BWP12T U1394 ( .I(n1300), .ZN(n1050) );
  INR2D1BWP12T U1395 ( .A1(Instruction_Fetch_inst1_fetched_instruction_reg_13_), .B1(n1301), .ZN(n1030) );
  TPNR2D1BWP12T U1396 ( .A1(n1050), .A2(n1030), .ZN(n1031) );
  TPND2D2BWP12T U1397 ( .A1(n1032), .A2(n1031), .ZN(n1161) );
  ND2D1BWP12T U1398 ( .A1(n1149), .A2(n1161), .ZN(n1056) );
  INVD1BWP12T U1399 ( .I(n1056), .ZN(n1036) );
  TPND2D0BWP12T U1400 ( .A1(n1109), .A2(MEM_MEMCTRL_from_mem_data[6]), .ZN(
        n1034) );
  CKND2D1BWP12T U1401 ( .A1(n1834), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[14]), .ZN(n1033) );
  ND3D1BWP12T U1402 ( .A1(n1034), .A2(n1111), .A3(n1033), .ZN(
        MEMCTRL_RF_IF_data_in[14]) );
  INR2D2BWP12T U1403 ( .A1(Instruction_Fetch_inst1_fetched_instruction_reg_14_), .B1(n1301), .ZN(n1035) );
  TPAOI21D2BWP12T U1404 ( .A1(MEMCTRL_RF_IF_data_in[14]), .A2(n1731), .B(n1035), .ZN(n1152) );
  INVD1BWP12T U1405 ( .I(n1152), .ZN(n1044) );
  ND2D1BWP12T U1406 ( .A1(n1036), .A2(n1044), .ZN(n1115) );
  INVD1BWP12T U1407 ( .I(n1115), .ZN(n1144) );
  CKND2D1BWP12T U1408 ( .A1(n1109), .A2(MEM_MEMCTRL_from_mem_data[4]), .ZN(
        n1038) );
  CKND2D1BWP12T U1409 ( .A1(n1834), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[12]), .ZN(n1037) );
  ND3D1BWP12T U1410 ( .A1(n1038), .A2(n1111), .A3(n1037), .ZN(
        MEMCTRL_RF_IF_data_in[12]) );
  ND2D1BWP12T U1411 ( .A1(MEMCTRL_RF_IF_data_in[12]), .A2(n1568), .ZN(n1041)
         );
  INR2D1BWP12T U1412 ( .A1(Instruction_Fetch_inst1_fetched_instruction_reg_12_), .B1(n1301), .ZN(n1039) );
  NR2D2BWP12T U1413 ( .A1(n1050), .A2(n1039), .ZN(n1040) );
  TPND2D3BWP12T U1414 ( .A1(n1041), .A2(n1040), .ZN(n1410) );
  CKND2D2BWP12T U1415 ( .A1(n1144), .A2(n1410), .ZN(n1387) );
  INR2D2BWP12T U1416 ( .A1(n1321), .B1(n1387), .ZN(n1685) );
  ND3D1BWP12T U1417 ( .A1(DEC_IF_stall_to_instructionfetch), .A2(
        irdecode_inst1_split_instruction), .A3(n1435), .ZN(n1043) );
  TPND2D2BWP12T U1418 ( .A1(n1586), .A2(DEC_MEMCTRL_memory_load_request), .ZN(
        n1042) );
  TPOAI21D2BWP12T U1419 ( .A1(n1484), .A2(n1580), .B(n1042), .ZN(n1046) );
  TPAOI21D4BWP12T U1420 ( .A1(n1733), .A2(n1043), .B(n1046), .ZN(n1790) );
  INVD1P75BWP12T U1421 ( .I(n1161), .ZN(n1148) );
  TPND2D2BWP12T U1422 ( .A1(n1149), .A2(n1148), .ZN(n1154) );
  INVD3BWP12T U1423 ( .I(n1410), .ZN(n1402) );
  ND2D1BWP12T U1424 ( .A1(n1044), .A2(n1402), .ZN(n1045) );
  NR2D2BWP12T U1425 ( .A1(n1154), .A2(n1045), .ZN(n1814) );
  CKND2D2BWP12T U1426 ( .A1(n1814), .A2(n1790), .ZN(n1661) );
  INVD1BWP12T U1427 ( .I(irdecode_inst1_N707), .ZN(n1094) );
  TPND2D0BWP12T U1428 ( .A1(n1109), .A2(MEM_MEMCTRL_from_mem_data[1]), .ZN(
        n1048) );
  TPND2D0BWP12T U1429 ( .A1(n1834), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[9]), .ZN(n1047) );
  ND3D1BWP12T U1430 ( .A1(n1048), .A2(n1111), .A3(n1047), .ZN(
        MEMCTRL_RF_IF_data_in[9]) );
  ND2D1BWP12T U1431 ( .A1(MEMCTRL_RF_IF_data_in[9]), .A2(n1568), .ZN(n1052) );
  INR2XD0BWP12T U1432 ( .A1(Instruction_Fetch_inst1_fetched_instruction_reg_9_), .B1(n1301), .ZN(n1049) );
  NR2D1BWP12T U1433 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  ND2D3BWP12T U1434 ( .A1(n1052), .A2(n1051), .ZN(n1795) );
  TPND2D0BWP12T U1435 ( .A1(n1109), .A2(MEM_MEMCTRL_from_mem_data[2]), .ZN(
        n1054) );
  TPND2D0BWP12T U1436 ( .A1(n1834), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[10]), .ZN(n1053) );
  ND3D1BWP12T U1437 ( .A1(n1054), .A2(n1111), .A3(n1053), .ZN(
        MEMCTRL_RF_IF_data_in[10]) );
  IOA21D1BWP12T U1438 ( .A1(n1257), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_10_), .B(n1300), .ZN(
        n1055) );
  TPAOI21D2BWP12T U1439 ( .A1(MEMCTRL_RF_IF_data_in[10]), .A2(n1568), .B(n1055), .ZN(n1787) );
  NR2D1BWP12T U1440 ( .A1(n1795), .A2(n1787), .ZN(n1057) );
  ND2D1BWP12T U1441 ( .A1(n1210), .A2(n1410), .ZN(n1119) );
  INR2D2BWP12T U1442 ( .A1(n1057), .B1(n1119), .ZN(n1817) );
  CKND2D2BWP12T U1443 ( .A1(n1817), .A2(n1790), .ZN(n1693) );
  TPNR3D0BWP12T U1444 ( .A1(irdecode_inst1_N544), .A2(irdecode_inst1_N542), 
        .A3(irdecode_inst1_N541), .ZN(n1061) );
  CKND2D1BWP12T U1445 ( .A1(n1109), .A2(MEM_MEMCTRL_from_mem_data[0]), .ZN(
        n1059) );
  TPND2D0BWP12T U1446 ( .A1(n1834), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[8]), .ZN(n1058) );
  ND3D1BWP12T U1447 ( .A1(n1059), .A2(n1111), .A3(n1058), .ZN(
        MEMCTRL_RF_IF_data_in[8]) );
  IOA21D1BWP12T U1448 ( .A1(n1257), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_8_), .B(n1300), .ZN(
        n1060) );
  AOI21D2BWP12T U1449 ( .A1(MEMCTRL_RF_IF_data_in[8]), .A2(n1568), .B(n1060), 
        .ZN(n1684) );
  ND2D1BWP12T U1450 ( .A1(n1684), .A2(n1328), .ZN(n1077) );
  INR2D1BWP12T U1451 ( .A1(n1061), .B1(n1077), .ZN(n1066) );
  INVD1BWP12T U1452 ( .I(irdecode_inst1_N543), .ZN(n1330) );
  TPND3D0BWP12T U1453 ( .A1(n1066), .A2(irdecode_inst1_N545), .A3(n1330), .ZN(
        n1064) );
  TPNR2D0BWP12T U1454 ( .A1(irdecode_inst1_N545), .A2(irdecode_inst1_N543), 
        .ZN(n1062) );
  TPND2D0BWP12T U1455 ( .A1(n1066), .A2(n1062), .ZN(n1063) );
  MUX2NXD0BWP12T U1456 ( .I0(n1064), .I1(n1063), .S(irdecode_inst1_N546), .ZN(
        n1087) );
  NR2D1BWP12T U1457 ( .A1(n1615), .A2(n1330), .ZN(n1065) );
  ND2D1BWP12T U1458 ( .A1(n1066), .A2(n1065), .ZN(n1634) );
  INVD0BWP12T U1459 ( .I(n1615), .ZN(n1329) );
  NR2D0BWP12T U1460 ( .A1(irdecode_inst1_N543), .A2(irdecode_inst1_N541), .ZN(
        n1067) );
  INVD1BWP12T U1461 ( .I(irdecode_inst1_N542), .ZN(n1078) );
  ND4D0BWP12T U1462 ( .A1(n1329), .A2(n1067), .A3(n1078), .A4(
        irdecode_inst1_N544), .ZN(n1068) );
  TPNR2D0BWP12T U1463 ( .A1(n1077), .A2(n1068), .ZN(n1075) );
  INVD1P75BWP12T U1464 ( .I(n1684), .ZN(n1714) );
  NR2D2BWP12T U1465 ( .A1(n1615), .A2(irdecode_inst1_N544), .ZN(n1088) );
  CKND0BWP12T U1466 ( .I(irdecode_inst1_N540), .ZN(n1069) );
  INVD1BWP12T U1467 ( .I(irdecode_inst1_N541), .ZN(n1081) );
  CKND2D1BWP12T U1468 ( .A1(n1069), .A2(n1081), .ZN(n1070) );
  CKND2D1BWP12T U1469 ( .A1(n1071), .A2(irdecode_inst1_N539), .ZN(n1629) );
  TPNR2D0BWP12T U1470 ( .A1(n1714), .A2(n1629), .ZN(n1074) );
  INVD1BWP12T U1471 ( .I(n1071), .ZN(n1072) );
  NR2D1BWP12T U1472 ( .A1(n1072), .A2(irdecode_inst1_N539), .ZN(n1073) );
  ND2D1BWP12T U1473 ( .A1(n1634), .A2(n1076), .ZN(n1771) );
  INVD1BWP12T U1474 ( .I(n1077), .ZN(n1083) );
  NR2D0BWP12T U1475 ( .A1(n1628), .A2(irdecode_inst1_N541), .ZN(n1080) );
  AOI21D1BWP12T U1476 ( .A1(n1083), .A2(n1080), .B(n1772), .ZN(n1085) );
  CKND2D1BWP12T U1477 ( .A1(n1083), .A2(n1630), .ZN(n1084) );
  ND2D1BWP12T U1478 ( .A1(n1085), .A2(n1084), .ZN(n1086) );
  TPNR3D2BWP12T U1479 ( .A1(n1087), .A2(n1771), .A3(n1086), .ZN(n1332) );
  INVD1BWP12T U1480 ( .I(n1088), .ZN(n1331) );
  INVD1BWP12T U1481 ( .I(n1630), .ZN(n1089) );
  ND2D1BWP12T U1482 ( .A1(n1089), .A2(n1628), .ZN(n1327) );
  TPND2D1BWP12T U1483 ( .A1(n1351), .A2(n1328), .ZN(n1636) );
  TPNR2D1BWP12T U1484 ( .A1(n1636), .A2(n1693), .ZN(n1767) );
  TPNR2D0BWP12T U1485 ( .A1(irdecode_inst1_N707), .A2(irdecode_inst1_N705), 
        .ZN(n1090) );
  MUX2XD2BWP12T U1486 ( .I0(
        memory_interface_inst1_delay_first_two_bytes_out[7]), .I1(
        MEM_MEMCTRL_from_mem_data[15]), .S(n1730), .Z(MEMCTRL_RF_IF_data_in[7]) );
  INR2D0BWP12T U1487 ( .A1(n1090), .B1(IF_DEC_instruction[7]), .ZN(n1095) );
  NR2D1BWP12T U1488 ( .A1(irdecode_inst1_N702), .A2(irdecode_inst1_N701), .ZN(
        n1096) );
  INVD1BWP12T U1489 ( .I(irdecode_inst1_N703), .ZN(n1091) );
  ND2D1BWP12T U1490 ( .A1(n1096), .A2(n1091), .ZN(n1105) );
  INVD1BWP12T U1491 ( .I(irdecode_inst1_N704), .ZN(n1344) );
  NR2D1BWP12T U1492 ( .A1(irdecode_inst1_N706), .A2(irdecode_inst1_N707), .ZN(
        n1341) );
  INVD1BWP12T U1493 ( .I(irdecode_inst1_N705), .ZN(n1343) );
  ND2D1BWP12T U1494 ( .A1(n1341), .A2(n1343), .ZN(n1345) );
  NR2D1BWP12T U1495 ( .A1(n1345), .A2(irdecode_inst1_N704), .ZN(n1349) );
  ND2D1BWP12T U1496 ( .A1(n1349), .A2(n1091), .ZN(n1347) );
  INR3XD0BWP12T U1497 ( .A1(irdecode_inst1_N702), .B1(irdecode_inst1_N701), 
        .B2(n1347), .ZN(n1092) );
  INR2D1BWP12T U1498 ( .A1(n1092), .B1(IF_DEC_instruction[7]), .ZN(n1355) );
  NR3XD0BWP12T U1499 ( .A1(n1105), .A2(irdecode_inst1_N706), .A3(
        irdecode_inst1_N704), .ZN(n1093) );
  INR2D1BWP12T U1500 ( .A1(n1093), .B1(IF_DEC_instruction[7]), .ZN(n1102) );
  ND2D1BWP12T U1501 ( .A1(n1798), .A2(n1773), .ZN(n1100) );
  ND3XD0BWP12T U1502 ( .A1(n1349), .A2(n1096), .A3(irdecode_inst1_N703), .ZN(
        n1097) );
  TPNR2D0BWP12T U1503 ( .A1(IF_DEC_instruction[7]), .A2(n1097), .ZN(n1354) );
  INVD1BWP12T U1504 ( .I(n1354), .ZN(n1098) );
  ND2D1BWP12T U1505 ( .A1(n1774), .A2(n1098), .ZN(n1099) );
  INR2XD0BWP12T U1506 ( .A1(n1348), .B1(IF_DEC_instruction[7]), .ZN(n1101) );
  INVD1BWP12T U1507 ( .I(n1101), .ZN(n1108) );
  ND2D1BWP12T U1508 ( .A1(n1104), .A2(n1108), .ZN(n1342) );
  INVD6BWP12T U1509 ( .I(n1790), .ZN(n1757) );
  ND2D2BWP12T U1510 ( .A1(n1757), .A2(n1364), .ZN(n1692) );
  INVD1BWP12T U1511 ( .I(n1104), .ZN(n1350) );
  CKND0BWP12T U1512 ( .I(n1349), .ZN(n1106) );
  TPNR2D0BWP12T U1513 ( .A1(n1106), .A2(n1105), .ZN(n1107) );
  TPND2D0BWP12T U1514 ( .A1(IF_DEC_instruction[7]), .A2(n1107), .ZN(n1637) );
  ND2D1BWP12T U1515 ( .A1(n1108), .A2(n1637), .ZN(n1775) );
  NR2D1BWP12T U1516 ( .A1(n1350), .A2(n1775), .ZN(n1618) );
  OAI22D1BWP12T U1517 ( .A1(n1332), .A2(n1693), .B1(n1618), .B2(n1661), .ZN(
        n1157) );
  TPND2D0BWP12T U1518 ( .A1(n1109), .A2(MEM_MEMCTRL_from_mem_data[3]), .ZN(
        n1112) );
  TPND2D0BWP12T U1519 ( .A1(n1834), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[11]), .ZN(n1110) );
  ND3D1BWP12T U1520 ( .A1(n1112), .A2(n1111), .A3(n1110), .ZN(
        MEMCTRL_RF_IF_data_in[11]) );
  IOA21D1BWP12T U1521 ( .A1(n1257), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_11_), .B(n1300), .ZN(
        n1113) );
  TPAOI21D1BWP12T U1522 ( .A1(MEMCTRL_RF_IF_data_in[11]), .A2(n1568), .B(n1113), .ZN(n1114) );
  BUFFXD4BWP12T U1523 ( .I(n1114), .Z(n1830) );
  ND2D1BWP12T U1524 ( .A1(n1402), .A2(n1830), .ZN(n1118) );
  NR2D1BWP12T U1525 ( .A1(n1115), .A2(n1118), .ZN(n1247) );
  NR2D1BWP12T U1526 ( .A1(n1402), .A2(n1152), .ZN(n1116) );
  INR2D2BWP12T U1527 ( .A1(n1116), .B1(n1154), .ZN(n1249) );
  INVD1BWP12T U1528 ( .I(n1149), .ZN(n1117) );
  ND2D1BWP12T U1529 ( .A1(n1117), .A2(n1152), .ZN(n1378) );
  NR3D1BWP12T U1530 ( .A1(n1161), .A2(n1149), .A3(n1152), .ZN(n1188) );
  INVD1BWP12T U1531 ( .I(n1118), .ZN(n1162) );
  CKND2D1BWP12T U1532 ( .A1(n1188), .A2(n1162), .ZN(n1603) );
  ND3XD0BWP12T U1533 ( .A1(n1740), .A2(n1378), .A3(n1603), .ZN(n1150) );
  AOI21D0BWP12T U1534 ( .A1(n1714), .A2(n1787), .B(n1795), .ZN(n1120) );
  INVD2BWP12T U1535 ( .I(n1830), .ZN(n1821) );
  CKND2D1BWP12T U1536 ( .A1(n1821), .A2(n1787), .ZN(n1736) );
  INVD1BWP12T U1537 ( .I(n1119), .ZN(n1151) );
  IOA21D0BWP12T U1538 ( .A1(n1120), .A2(n1736), .B(n1151), .ZN(n1146) );
  INR2D2BWP12T U1539 ( .A1(n1402), .B1(n1830), .ZN(n1820) );
  NR3D1BWP12T U1540 ( .A1(irdecode_inst1_itstate_0_), .A2(
        irdecode_inst1_itstate_2_), .A3(irdecode_inst1_itstate_1_), .ZN(n1215)
         );
  NR3XD0BWP12T U1541 ( .A1(irdecode_inst1_itstate_4_), .A2(
        irdecode_inst1_itstate_3_), .A3(irdecode_inst1_itstate_5_), .ZN(n1121)
         );
  NR2D1BWP12T U1542 ( .A1(irdecode_inst1_itstate_7_), .A2(
        irdecode_inst1_itstate_6_), .ZN(n1132) );
  ND3D1BWP12T U1543 ( .A1(n1215), .A2(n1121), .A3(n1132), .ZN(n1407) );
  CKND2D0BWP12T U1544 ( .A1(irdecode_inst1_itstate_6_), .A2(RF_OUT_n), .ZN(
        n1123) );
  INR2XD0BWP12T U1545 ( .A1(RF_OUT_c), .B1(RF_OUT_z), .ZN(n1173) );
  INVD0BWP12T U1546 ( .I(irdecode_inst1_itstate_6_), .ZN(n1592) );
  ND2XD0BWP12T U1547 ( .A1(n1173), .A2(n1592), .ZN(n1122) );
  MUX2ND0BWP12T U1548 ( .I0(n1123), .I1(n1122), .S(irdecode_inst1_itstate_7_), 
        .ZN(n1124) );
  AOI21D0BWP12T U1549 ( .A1(RF_OUT_z), .A2(n1132), .B(n1124), .ZN(n1131) );
  INVD1BWP12T U1550 ( .I(RF_OUT_z), .ZN(n1170) );
  XOR2D1BWP12T U1551 ( .A1(RF_OUT_v), .A2(RF_OUT_n), .Z(n1171) );
  INR2D1BWP12T U1552 ( .A1(n1170), .B1(n1171), .ZN(n1168) );
  CKND2D1BWP12T U1553 ( .A1(irdecode_inst1_itstate_7_), .A2(
        irdecode_inst1_itstate_6_), .ZN(n1125) );
  INVD1BWP12T U1554 ( .I(n1125), .ZN(n1133) );
  ND2D1BWP12T U1555 ( .A1(n1168), .A2(n1133), .ZN(n1130) );
  INR2D1BWP12T U1556 ( .A1(irdecode_inst1_itstate_7_), .B1(n1171), .ZN(n1129)
         );
  INVD1BWP12T U1557 ( .I(RF_OUT_c), .ZN(n1463) );
  CKND0BWP12T U1558 ( .I(n1132), .ZN(n1127) );
  TPND2D0BWP12T U1559 ( .A1(irdecode_inst1_itstate_6_), .A2(RF_OUT_v), .ZN(
        n1126) );
  OAI211D1BWP12T U1560 ( .A1(n1463), .A2(n1127), .B(n1126), .C(n1125), .ZN(
        n1128) );
  OAI21D1BWP12T U1561 ( .A1(n1129), .A2(n1128), .B(irdecode_inst1_itstate_5_), 
        .ZN(n1136) );
  OAI211D1BWP12T U1562 ( .A1(irdecode_inst1_itstate_5_), .A2(n1131), .B(n1130), 
        .C(n1136), .ZN(n1142) );
  AOI21D0BWP12T U1563 ( .A1(n1132), .A2(n1170), .B(irdecode_inst1_itstate_5_), 
        .ZN(n1140) );
  INVD0BWP12T U1564 ( .I(n1168), .ZN(n1174) );
  CKND2D1BWP12T U1565 ( .A1(n1174), .A2(n1133), .ZN(n1139) );
  NR2D0BWP12T U1566 ( .A1(n1592), .A2(RF_OUT_n), .ZN(n1135) );
  NR2D0BWP12T U1567 ( .A1(n1173), .A2(irdecode_inst1_itstate_6_), .ZN(n1134)
         );
  MUX2NXD0BWP12T U1568 ( .I0(n1135), .I1(n1134), .S(irdecode_inst1_itstate_7_), 
        .ZN(n1138) );
  INVD1BWP12T U1569 ( .I(n1136), .ZN(n1137) );
  AOI31D1BWP12T U1570 ( .A1(n1140), .A2(n1139), .A3(n1138), .B(n1137), .ZN(
        n1141) );
  MUX2D1BWP12T U1571 ( .I0(n1142), .I1(n1141), .S(irdecode_inst1_itstate_4_), 
        .Z(n1143) );
  INR2D2BWP12T U1572 ( .A1(n1407), .B1(n1143), .ZN(n1195) );
  AOI21D0BWP12T U1573 ( .A1(n1144), .A2(n1820), .B(n1195), .ZN(n1145) );
  ND2D1BWP12T U1574 ( .A1(n1146), .A2(n1145), .ZN(n1197) );
  CKND2D0BWP12T U1575 ( .A1(n1402), .A2(n1152), .ZN(n1147) );
  NR2D1BWP12T U1576 ( .A1(n1154), .A2(n1147), .ZN(n1735) );
  NR3D1BWP12T U1577 ( .A1(n1149), .A2(n1148), .A3(n1152), .ZN(n1703) );
  TPNR2D1BWP12T U1578 ( .A1(n1735), .A2(n1703), .ZN(n1384) );
  CKND2D1BWP12T U1579 ( .A1(n1188), .A2(n1410), .ZN(n1338) );
  ND2D1BWP12T U1580 ( .A1(n1384), .A2(n1338), .ZN(n1743) );
  NR3D1BWP12T U1581 ( .A1(n1150), .A2(n1197), .A3(n1743), .ZN(n1388) );
  CKND2D1BWP12T U1582 ( .A1(n1830), .A2(n1787), .ZN(n1361) );
  INVD1P75BWP12T U1583 ( .I(n1795), .ZN(n1822) );
  CKND2D1BWP12T U1584 ( .A1(n1822), .A2(n1684), .ZN(n1669) );
  INVD1BWP12T U1585 ( .I(n1820), .ZN(n1320) );
  CKND2D0BWP12T U1586 ( .A1(n1410), .A2(n1152), .ZN(n1153) );
  TPNR2D1BWP12T U1587 ( .A1(n1794), .A2(n1779), .ZN(n1786) );
  ND2D1BWP12T U1588 ( .A1(n1210), .A2(n1402), .ZN(n1470) );
  CKND2D2BWP12T U1589 ( .A1(n1786), .A2(n1470), .ZN(n1744) );
  INR2D2BWP12T U1590 ( .A1(n1191), .B1(n1744), .ZN(n1710) );
  INVD0BWP12T U1591 ( .I(n1387), .ZN(n1831) );
  INR2D1BWP12T U1592 ( .A1(n1830), .B1(n1387), .ZN(n1670) );
  AOI21D0BWP12T U1593 ( .A1(n1831), .A2(irdecode_inst1_N911), .B(n1670), .ZN(
        n1155) );
  TPAOI31D0BWP12T U1594 ( .A1(n1388), .A2(n1710), .A3(n1155), .B(n1757), .ZN(
        n1156) );
  NR2D1BWP12T U1595 ( .A1(n1157), .A2(n1156), .ZN(n1158) );
  TPND2D2BWP12T U1596 ( .A1(n1370), .A2(n1158), .ZN(n1160) );
  INR2D1BWP12T U1597 ( .A1(irdecode_inst1_step[0]), .B1(n1364), .ZN(n1159) );
  INVD2BWP12T U1598 ( .I(n1854), .ZN(irdecode_inst1_next_step_0_) );
  INR2D1BWP12T U1599 ( .A1(n1795), .B1(n1338), .ZN(n1737) );
  CKND2D1BWP12T U1600 ( .A1(n1737), .A2(n1361), .ZN(n1789) );
  CKND2D1BWP12T U1601 ( .A1(n1740), .A2(n1387), .ZN(n1163) );
  INVD1BWP12T U1602 ( .I(n1191), .ZN(n1826) );
  TPOAI31D0BWP12T U1603 ( .A1(n1810), .A2(n1821), .A3(n1367), .B(n1790), .ZN(
        n1666) );
  CKND2D1BWP12T U1604 ( .A1(n1370), .A2(n1666), .ZN(n1263) );
  AO21D1BWP12T U1605 ( .A1(n1836), .A2(DEC_RF_memory_store_data_reg[4]), .B(
        n1263), .Z(n826) );
  MUX2D1BWP12T U1606 ( .I0(memory_interface_inst1_delay_first_two_bytes_out[5]), .I1(MEM_MEMCTRL_from_mem_data[13]), .S(n1730), .Z(MEMCTRL_RF_IF_data_in[5])
         );
  NR2D1BWP12T U1607 ( .A1(n1378), .A2(n1161), .ZN(n1403) );
  INR2D1BWP12T U1608 ( .A1(n1338), .B1(n1403), .ZN(n1612) );
  CKND2D1BWP12T U1609 ( .A1(n1612), .A2(n1384), .ZN(n1691) );
  INVD1P75BWP12T U1610 ( .I(n1710), .ZN(n1715) );
  NR2XD0BWP12T U1611 ( .A1(n1715), .A2(n1197), .ZN(n1377) );
  INVD1BWP12T U1612 ( .I(n1787), .ZN(n1675) );
  INR2D2BWP12T U1613 ( .A1(n1675), .B1(n1603), .ZN(n1745) );
  CKND2D1BWP12T U1614 ( .A1(n1745), .A2(n1795), .ZN(n1372) );
  INR2D2BWP12T U1615 ( .A1(n1161), .B1(n1378), .ZN(n1718) );
  ND2D1BWP12T U1616 ( .A1(n1377), .A2(n1760), .ZN(n1690) );
  INVD1BWP12T U1617 ( .I(n1163), .ZN(n1749) );
  INVD1BWP12T U1618 ( .I(n1817), .ZN(n1742) );
  ND2D1BWP12T U1619 ( .A1(n1749), .A2(n1742), .ZN(n1606) );
  NR2XD0BWP12T U1620 ( .A1(n1690), .A2(n1606), .ZN(n1614) );
  INVD0BWP12T U1621 ( .I(n1614), .ZN(n1165) );
  NR2D1BWP12T U1622 ( .A1(n1814), .A2(n1718), .ZN(n1683) );
  MUX2D1BWP12T U1623 ( .I0(memory_interface_inst1_delay_first_two_bytes_out[2]), .I1(MEM_MEMCTRL_from_mem_data[10]), .S(n1730), .Z(MEMCTRL_RF_IF_data_in[2])
         );
  INVD1BWP12T U1624 ( .I(IF_DEC_instruction[2]), .ZN(n1788) );
  OAI22D0BWP12T U1625 ( .A1(n1683), .A2(n1787), .B1(n1603), .B2(n1788), .ZN(
        n1164) );
  AOI211XD0BWP12T U1626 ( .A1(IF_DEC_instruction[5]), .A2(n1691), .B(n1165), 
        .C(n1164), .ZN(n1167) );
  ND2D1BWP12T U1627 ( .A1(n1836), .A2(n1001), .ZN(n1166) );
  OAI211D1BWP12T U1628 ( .A1(n1757), .A2(n1167), .B(n1692), .C(n1166), .ZN(
        n813) );
  INVD1BWP12T U1629 ( .I(n1361), .ZN(n1340) );
  NR2D0BWP12T U1630 ( .A1(n1787), .A2(n1168), .ZN(n1169) );
  AOI22D0BWP12T U1631 ( .A1(n1340), .A2(n1170), .B1(n1169), .B2(n1821), .ZN(
        n1187) );
  NR2D1BWP12T U1632 ( .A1(n1795), .A2(n1684), .ZN(n1319) );
  INVD1BWP12T U1633 ( .I(n1319), .ZN(n1412) );
  CKND0BWP12T U1634 ( .I(n1171), .ZN(n1172) );
  MUX2ND0BWP12T U1635 ( .I0(n1173), .I1(n1172), .S(n1795), .ZN(n1178) );
  MUX2XD0BWP12T U1636 ( .I0(RF_OUT_n), .I1(RF_OUT_v), .S(n1795), .Z(n1179) );
  NR2D0BWP12T U1637 ( .A1(n1795), .A2(n1174), .ZN(n1175) );
  MUX2ND0BWP12T U1638 ( .I0(n1179), .I1(n1175), .S(n1821), .ZN(n1177) );
  MUX2ND0BWP12T U1639 ( .I0(RF_OUT_z), .I1(RF_OUT_c), .S(n1795), .ZN(n1176) );
  OAI222D0BWP12T U1640 ( .A1(n1736), .A2(n1178), .B1(n1787), .B2(n1177), .C1(
        n1361), .C2(n1176), .ZN(n1185) );
  CKND0BWP12T U1641 ( .I(n1178), .ZN(n1183) );
  INVD0BWP12T U1642 ( .I(n1179), .ZN(n1180) );
  ND3D0BWP12T U1643 ( .A1(n1180), .A2(n1830), .A3(n1675), .ZN(n1182) );
  ND3D0BWP12T U1644 ( .A1(n1340), .A2(n1463), .A3(n1795), .ZN(n1181) );
  OAI211D0BWP12T U1645 ( .A1(n1183), .A2(n1736), .B(n1182), .C(n1181), .ZN(
        n1184) );
  MUX2ND0BWP12T U1646 ( .I0(n1185), .I1(n1184), .S(n1714), .ZN(n1186) );
  OAI21D0BWP12T U1647 ( .A1(n1187), .A2(n1412), .B(n1186), .ZN(n1194) );
  NR4D0BWP12T U1648 ( .A1(n1748), .A2(n1817), .A3(n1247), .A4(n1831), .ZN(
        n1192) );
  INVD1BWP12T U1649 ( .I(IF_DEC_instruction[7]), .ZN(n1827) );
  MUX2D1BWP12T U1650 ( .I0(memory_interface_inst1_delay_first_two_bytes_out[6]), .I1(MEM_MEMCTRL_from_mem_data[14]), .S(n1730), .Z(MEMCTRL_RF_IF_data_in[6])
         );
  ND2XD0BWP12T U1651 ( .A1(n1827), .A2(IF_DEC_instruction[6]), .ZN(n1414) );
  NR2D0BWP12T U1652 ( .A1(n1361), .A2(n1410), .ZN(n1189) );
  CKND2D1BWP12T U1653 ( .A1(n1189), .A2(n1188), .ZN(n1824) );
  AOI31D0BWP12T U1654 ( .A1(n1684), .A2(n1795), .A3(n1414), .B(n1824), .ZN(
        n1190) );
  NR2D1BWP12T U1655 ( .A1(n1190), .A2(n1403), .ZN(n1596) );
  CKND2D1BWP12T U1656 ( .A1(n1745), .A2(n1412), .ZN(n1385) );
  ND4D0BWP12T U1657 ( .A1(n1192), .A2(n1596), .A3(n1191), .A4(n1385), .ZN(
        n1193) );
  AOI21D0BWP12T U1658 ( .A1(n1194), .A2(n1249), .B(n1193), .ZN(n1196) );
  NR2D4BWP12T U1659 ( .A1(n1195), .A2(n1757), .ZN(n1809) );
  NR2XD0BWP12T U1660 ( .A1(n1196), .A2(n1832), .ZN(
        irdecode_inst1_next_alu_write_to_reg_enable) );
  INVD1BWP12T U1661 ( .I(n1197), .ZN(n1759) );
  INR2D1BWP12T U1662 ( .A1(n1410), .B1(n1830), .ZN(n1699) );
  INVD1BWP12T U1663 ( .I(n1403), .ZN(n1825) );
  AOI21D1BWP12T U1664 ( .A1(n1787), .A2(n1699), .B(n1825), .ZN(n1722) );
  INVD0BWP12T U1665 ( .I(n1722), .ZN(n1602) );
  ND4D0BWP12T U1666 ( .A1(n1759), .A2(n1683), .A3(n1692), .A4(n1602), .ZN(
        n1199) );
  TPND2D0BWP12T U1667 ( .A1(n1710), .A2(n1384), .ZN(n1605) );
  INR2D1BWP12T U1668 ( .A1(n1692), .B1(n1790), .ZN(n1389) );
  INVD1BWP12T U1669 ( .I(n1389), .ZN(n1198) );
  OAI31D1BWP12T U1670 ( .A1(n1199), .A2(n1606), .A3(n1605), .B(n1198), .ZN(
        n1755) );
  MUX2D1BWP12T U1671 ( .I0(memory_interface_inst1_delay_first_two_bytes_out[3]), .I1(MEM_MEMCTRL_from_mem_data[11]), .S(n1730), .Z(MEMCTRL_RF_IF_data_in[3])
         );
  CKND0BWP12T U1672 ( .I(IF_DEC_instruction[3]), .ZN(n1396) );
  OAI22D0BWP12T U1673 ( .A1(n1612), .A2(n1823), .B1(n1396), .B2(n1603), .ZN(
        n1200) );
  TPND2D0BWP12T U1674 ( .A1(n1755), .A2(n1201), .ZN(n844) );
  CKND2D1BWP12T U1675 ( .A1(n1257), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_0_), .ZN(n1202) );
  TPND2D2BWP12T U1676 ( .A1(n1203), .A2(n1202), .ZN(IF_DEC_instruction[0]) );
  AOI22D0BWP12T U1677 ( .A1(n1722), .A2(IF_DEC_instruction[6]), .B1(n1718), 
        .B2(IF_DEC_instruction[0]), .ZN(n1204) );
  INR2D1BWP12T U1678 ( .A1(n1821), .B1(n1387), .ZN(n1739) );
  TPND2D0BWP12T U1679 ( .A1(n1739), .A2(irdecode_inst1_N911), .ZN(n1758) );
  TPAOI21D0BWP12T U1680 ( .A1(n1204), .A2(n1758), .B(n1832), .ZN(n1205) );
  AO21D1BWP12T U1681 ( .A1(DEC_RF_offset_b[0]), .A2(n1836), .B(n1205), .Z(n809) );
  MUX2D1BWP12T U1682 ( .I0(memory_interface_inst1_delay_first_two_bytes_out[1]), .I1(MEM_MEMCTRL_from_mem_data[9]), .S(n1730), .Z(MEMCTRL_RF_IF_data_in[1])
         );
  TPND2D0BWP12T U1683 ( .A1(n1257), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_1_), .ZN(n1206) );
  ND2D2BWP12T U1684 ( .A1(n1207), .A2(n1206), .ZN(IF_DEC_instruction[1]) );
  NR3XD0BWP12T U1685 ( .A1(n1822), .A2(n1787), .A3(n1684), .ZN(n1208) );
  ND2D1BWP12T U1686 ( .A1(n1208), .A2(n1699), .ZN(n1209) );
  NR4D0BWP12T U1687 ( .A1(IF_DEC_instruction[3]), .A2(IF_DEC_instruction[2]), 
        .A3(IF_DEC_instruction[1]), .A4(IF_DEC_instruction[0]), .ZN(n1212) );
  NR2D1BWP12T U1688 ( .A1(n1212), .A2(n1757), .ZN(n1211) );
  ND2D1BWP12T U1689 ( .A1(n1214), .A2(n1211), .ZN(n1593) );
  INVD1BWP12T U1690 ( .I(n1593), .ZN(n1264) );
  CKND2D1BWP12T U1691 ( .A1(n1214), .A2(n1212), .ZN(n1213) );
  AOI21D1BWP12T U1692 ( .A1(n1213), .A2(n1790), .B(reset), .ZN(n1590) );
  AOI211D1BWP12T U1693 ( .A1(n1215), .A2(irdecode_inst1_itstate_3_), .B(n1214), 
        .C(n1757), .ZN(n1591) );
  AO222D0BWP12T U1694 ( .A1(IF_DEC_instruction[1]), .A2(n1264), .B1(n1590), 
        .B2(irdecode_inst1_itstate_1_), .C1(irdecode_inst1_itstate_0_), .C2(
        n1591), .Z(n859) );
  AO222D0BWP12T U1695 ( .A1(IF_DEC_instruction[2]), .A2(n1264), .B1(n1590), 
        .B2(irdecode_inst1_itstate_2_), .C1(irdecode_inst1_itstate_1_), .C2(
        n1591), .Z(n858) );
  CKND2D1BWP12T U1696 ( .A1(RF_pc_out[9]), .A2(RF_pc_out[10]), .ZN(n1240) );
  CKND2D0BWP12T U1697 ( .A1(RF_pc_out[11]), .A2(RF_pc_out[12]), .ZN(n1216) );
  NR2D1BWP12T U1698 ( .A1(n1240), .A2(n1216), .ZN(n1305) );
  CKND2D0BWP12T U1699 ( .A1(RF_pc_out[13]), .A2(RF_pc_out[14]), .ZN(n1306) );
  ND2XD0BWP12T U1700 ( .A1(RF_pc_out[5]), .A2(RF_pc_out[6]), .ZN(n1449) );
  CKND2D0BWP12T U1701 ( .A1(RF_pc_out[3]), .A2(RF_pc_out[4]), .ZN(n1217) );
  ND2XD0BWP12T U1702 ( .A1(RF_pc_out[2]), .A2(RF_pc_out[1]), .ZN(n1313) );
  NR2D1BWP12T U1703 ( .A1(n1217), .A2(n1313), .ZN(n1448) );
  CKND2D0BWP12T U1704 ( .A1(RF_pc_out[17]), .A2(RF_pc_out[18]), .ZN(n1231) );
  INVD1BWP12T U1705 ( .I(RF_pc_out[19]), .ZN(n1232) );
  NR2XD0BWP12T U1706 ( .A1(n1231), .A2(n1232), .ZN(n1218) );
  ND2D1BWP12T U1707 ( .A1(n1230), .A2(n1218), .ZN(n1245) );
  INVD1BWP12T U1708 ( .I(RF_pc_out[20]), .ZN(n1244) );
  NR2D1BWP12T U1709 ( .A1(n1245), .A2(n1244), .ZN(n1228) );
  CKND2D1BWP12T U1710 ( .A1(n1228), .A2(RF_pc_out[21]), .ZN(n1227) );
  INVD1BWP12T U1711 ( .I(RF_pc_out[22]), .ZN(n1226) );
  NR2D1BWP12T U1712 ( .A1(n1227), .A2(n1226), .ZN(n1437) );
  CKND2D1BWP12T U1713 ( .A1(n1437), .A2(RF_pc_out[23]), .ZN(n1304) );
  INVD1BWP12T U1714 ( .I(RF_pc_out[24]), .ZN(n1303) );
  AN2XD1BWP12T U1715 ( .A1(n1229), .A2(n1458), .Z(IF_RF_incremented_pc_out[21]) );
  INVD1BWP12T U1716 ( .I(n1230), .ZN(n1237) );
  INVD0BWP12T U1717 ( .I(RF_pc_out[17]), .ZN(n1236) );
  NR2D1BWP12T U1718 ( .A1(n1237), .A2(n1236), .ZN(n1234) );
  CKND0BWP12T U1719 ( .I(RF_pc_out[18]), .ZN(n1233) );
  XNR2D1BWP12T U1720 ( .A1(n1234), .A2(n1233), .ZN(n1235) );
  AN2XD1BWP12T U1721 ( .A1(n1235), .A2(n1458), .Z(IF_RF_incremented_pc_out[18]) );
  CKXOR2D1BWP12T U1722 ( .A1(n1237), .A2(n1236), .Z(n1238) );
  AN2D0BWP12T U1723 ( .A1(n1238), .A2(n1458), .Z(IF_RF_incremented_pc_out[17])
         );
  INVD1BWP12T U1724 ( .I(n1239), .ZN(n1454) );
  CKND2D1BWP12T U1725 ( .A1(n1454), .A2(RF_pc_out[9]), .ZN(n1242) );
  CKND0BWP12T U1726 ( .I(RF_pc_out[10]), .ZN(n1241) );
  XOR2D1BWP12T U1727 ( .A1(n1242), .A2(n1241), .Z(n1243) );
  AN2D0BWP12T U1728 ( .A1(n1243), .A2(n1458), .Z(IF_RF_incremented_pc_out[10])
         );
  CKXOR2D1BWP12T U1729 ( .A1(n1245), .A2(n1244), .Z(n1246) );
  AN2D0BWP12T U1730 ( .A1(n1246), .A2(n1458), .Z(IF_RF_incremented_pc_out[20])
         );
  AN2D0BWP12T U1731 ( .A1(n1458), .A2(RF_pc_out[0]), .Z(
        IF_RF_incremented_pc_out[0]) );
  MUX2D1BWP12T U1732 ( .I0(memory_interface_inst1_delay_first_two_bytes_out[4]), .I1(MEM_MEMCTRL_from_mem_data[12]), .S(n1730), .Z(MEMCTRL_RF_IF_data_in[4])
         );
  ND2D1BWP12T U1733 ( .A1(n1854), .A2(n1739), .ZN(n1253) );
  ND2D3BWP12T U1734 ( .A1(n1249), .A2(n1723), .ZN(n1696) );
  CKND0BWP12T U1735 ( .I(n1696), .ZN(n1250) );
  TPAOI21D0BWP12T U1736 ( .A1(n1836), .A2(DEC_RF_offset_b[9]), .B(n1250), .ZN(
        n1252) );
  TPND2D0BWP12T U1737 ( .A1(n1744), .A2(n1723), .ZN(n1251) );
  OAI211D1BWP12T U1738 ( .A1(n1684), .A2(n1697), .B(n1252), .C(n1251), .ZN(
        n800) );
  AOI22D0BWP12T U1739 ( .A1(n1735), .A2(n1795), .B1(n1703), .B2(n1714), .ZN(
        n1260) );
  NR2D0BWP12T U1740 ( .A1(n1699), .A2(n1787), .ZN(n1258) );
  AOI22D0BWP12T U1741 ( .A1(n1258), .A2(n1403), .B1(n1718), .B2(
        IF_DEC_instruction[4]), .ZN(n1259) );
  OAI211D1BWP12T U1742 ( .A1(n1788), .A2(n1710), .B(n1260), .C(n1259), .ZN(
        n1261) );
  TPAOI21D0BWP12T U1743 ( .A1(IF_DEC_instruction[3]), .A2(n1679), .B(n1261), 
        .ZN(n1262) );
  MOAI22D1BWP12T U1744 ( .A1(n1262), .A2(n1832), .B1(n1836), .B2(
        DEC_RF_offset_b[4]), .ZN(n805) );
  INR2D1BWP12T U1745 ( .A1(n1353), .B1(n1693), .ZN(n1651) );
  AO211D1BWP12T U1746 ( .A1(n1836), .A2(DEC_RF_memory_store_data_reg[3]), .B(
        n1263), .C(n1651), .Z(n827) );
  AO222D0BWP12T U1747 ( .A1(IF_DEC_instruction[4]), .A2(n1264), .B1(n1591), 
        .B2(irdecode_inst1_itstate_3_), .C1(irdecode_inst1_itstate_4_), .C2(
        n1590), .Z(n856) );
  AO222D0BWP12T U1748 ( .A1(IF_DEC_instruction[3]), .A2(n1264), .B1(n1591), 
        .B2(irdecode_inst1_itstate_2_), .C1(n1590), .C2(
        irdecode_inst1_itstate_3_), .Z(n857) );
  INVD1BWP12T U1749 ( .I(IF_DEC_instruction[0]), .ZN(n1721) );
  MOAI22D0BWP12T U1750 ( .A1(n1721), .A2(n1593), .B1(n1590), .B2(
        irdecode_inst1_itstate_0_), .ZN(n860) );
  HICIND1BWP12T U1751 ( .A(RF_pc_out[28]), .CIN(n1265), .CO(n1269), .S(n1219)
         );
  HICIND1BWP12T U1752 ( .A(RF_pc_out[30]), .CIN(n1267), .CO(n1266), .S(n1268)
         );
  AN2D0BWP12T U1753 ( .A1(n1268), .A2(n1458), .Z(IF_RF_incremented_pc_out[30])
         );
  HICOND1BWP12T U1754 ( .A(RF_pc_out[29]), .CI(n1269), .CON(n1267), .S(n1270)
         );
  AN2D0BWP12T U1755 ( .A1(n1270), .A2(n1458), .Z(IF_RF_incremented_pc_out[29])
         );
  NR4D0BWP12T U1756 ( .A1(RF_pc_out[16]), .A2(RF_pc_out[31]), .A3(
        RF_pc_out[22]), .A4(RF_pc_out[26]), .ZN(n1299) );
  NR2D0BWP12T U1757 ( .A1(RF_pc_out[2]), .A2(RF_pc_out[1]), .ZN(n1290) );
  NR2D0BWP12T U1758 ( .A1(RF_pc_out[3]), .A2(RF_pc_out[4]), .ZN(n1271) );
  CKND2D1BWP12T U1759 ( .A1(n1290), .A2(n1271), .ZN(n1275) );
  NR2D0BWP12T U1760 ( .A1(RF_pc_out[5]), .A2(RF_pc_out[6]), .ZN(n1276) );
  NR2D0BWP12T U1761 ( .A1(RF_pc_out[7]), .A2(RF_pc_out[8]), .ZN(n1272) );
  TPND2D0BWP12T U1762 ( .A1(n1276), .A2(n1272), .ZN(n1273) );
  OR2XD1BWP12T U1763 ( .A1(n1275), .A2(n1273), .Z(n1286) );
  OR2XD0BWP12T U1764 ( .A1(RF_pc_out[9]), .A2(RF_pc_out[10]), .Z(n1274) );
  NR2D1BWP12T U1765 ( .A1(n1286), .A2(n1274), .ZN(n1282) );
  CKXOR2D0BWP12T U1766 ( .A1(n1282), .A2(RF_pc_out[11]), .Z(n1511) );
  INVD1BWP12T U1767 ( .I(n1275), .ZN(n1289) );
  ND2D1BWP12T U1768 ( .A1(n1289), .A2(n1276), .ZN(n1278) );
  NR2XD0BWP12T U1769 ( .A1(n1278), .A2(RF_pc_out[7]), .ZN(n1277) );
  CKXOR2D0BWP12T U1770 ( .A1(n1277), .A2(RF_pc_out[8]), .Z(n1521) );
  NR4D0BWP12T U1771 ( .A1(RF_pc_out[14]), .A2(n1511), .A3(n1521), .A4(
        RF_pc_out[28]), .ZN(n1280) );
  XNR2D0BWP12T U1772 ( .A1(n1278), .A2(RF_pc_out[7]), .ZN(n1527) );
  NR4D0BWP12T U1773 ( .A1(n1513), .A2(RF_pc_out[17]), .A3(n1527), .A4(
        RF_pc_out[29]), .ZN(n1279) );
  CKND2D1BWP12T U1774 ( .A1(n1280), .A2(n1279), .ZN(n1284) );
  CKND0BWP12T U1775 ( .I(RF_pc_out[11]), .ZN(n1281) );
  CKND2D1BWP12T U1776 ( .A1(n1282), .A2(n1281), .ZN(n1283) );
  XNR2D0BWP12T U1777 ( .A1(n1283), .A2(RF_pc_out[12]), .ZN(n1482) );
  NR4D0BWP12T U1778 ( .A1(RF_pc_out[23]), .A2(n1284), .A3(n1482), .A4(
        RF_pc_out[20]), .ZN(n1298) );
  OR3XD0BWP12T U1779 ( .A1(RF_pc_out[18]), .A2(RF_pc_out[30]), .A3(
        RF_pc_out[13]), .Z(n1285) );
  NR4D0BWP12T U1780 ( .A1(RF_pc_out[24]), .A2(n1285), .A3(RF_pc_out[21]), .A4(
        RF_pc_out[25]), .ZN(n1297) );
  XNR2D1BWP12T U1781 ( .A1(n1286), .A2(RF_pc_out[9]), .ZN(n1516) );
  CKND1BWP12T U1782 ( .I(n1516), .ZN(n1294) );
  CKND0BWP12T U1783 ( .I(RF_pc_out[5]), .ZN(n1287) );
  ND2D1BWP12T U1784 ( .A1(n1289), .A2(n1287), .ZN(n1288) );
  XNR2D0BWP12T U1785 ( .A1(n1288), .A2(RF_pc_out[6]), .ZN(n1543) );
  CKXOR2D0BWP12T U1786 ( .A1(n1289), .A2(RF_pc_out[5]), .Z(n1553) );
  INVD0BWP12T U1787 ( .I(n1290), .ZN(n1291) );
  XNR2D0BWP12T U1788 ( .A1(n1291), .A2(RF_pc_out[3]), .ZN(n1536) );
  XNR2XD0BWP12T U1789 ( .A1(RF_pc_out[2]), .A2(RF_pc_out[1]), .ZN(n1567) );
  CKND0BWP12T U1790 ( .I(RF_pc_out[1]), .ZN(n1459) );
  OR3D0BWP12T U1791 ( .A1(n1567), .A2(n1459), .A3(n1563), .Z(n1292) );
  NR4D0BWP12T U1792 ( .A1(n1543), .A2(n1553), .A3(n1536), .A4(n1292), .ZN(
        n1293) );
  CKND2D1BWP12T U1793 ( .A1(n1294), .A2(n1293), .ZN(n1295) );
  NR4D0BWP12T U1794 ( .A1(RF_pc_out[27]), .A2(RF_pc_out[15]), .A3(
        RF_pc_out[19]), .A4(n1295), .ZN(n1296) );
  AN4XD1BWP12T U1795 ( .A1(n1299), .A2(n1298), .A3(n1297), .A4(n1296), .Z(
        n1587) );
  ND3XD0BWP12T U1796 ( .A1(n1587), .A2(n1568), .A3(
        Instruction_Fetch_inst1_first_instruction_fetched), .ZN(n1302) );
  ND2D1BWP12T U1797 ( .A1(n1454), .A2(n1305), .ZN(n1447) );
  INVD1BWP12T U1798 ( .I(n1447), .ZN(n1443) );
  CKND0BWP12T U1799 ( .I(RF_pc_out[15]), .ZN(n1308) );
  NR2D1BWP12T U1800 ( .A1(n1309), .A2(n1308), .ZN(n1307) );
  CKXOR2D1BWP12T U1801 ( .A1(n1309), .A2(n1308), .Z(n1310) );
  CKND0BWP12T U1802 ( .I(RF_pc_out[2]), .ZN(n1311) );
  XNR2XD0BWP12T U1803 ( .A1(n1311), .A2(RF_pc_out[1]), .ZN(n1312) );
  AN2D0BWP12T U1804 ( .A1(n1312), .A2(n1458), .Z(IF_RF_incremented_pc_out[2])
         );
  INVD0BWP12T U1805 ( .I(n1313), .ZN(n1314) );
  INVD1BWP12T U1806 ( .I(IF_DEC_instruction[5]), .ZN(n1709) );
  NR2D1BWP12T U1807 ( .A1(n1720), .A2(n1709), .ZN(n1316) );
  INVD1BWP12T U1808 ( .I(n1718), .ZN(n1713) );
  CKND0BWP12T U1809 ( .I(n1703), .ZN(n1712) );
  OAI22D0BWP12T U1810 ( .A1(n1713), .A2(n1823), .B1(n1712), .B2(n1787), .ZN(
        n1315) );
  AOI211D1BWP12T U1811 ( .A1(n1715), .A2(IF_DEC_instruction[4]), .B(n1316), 
        .C(n1315), .ZN(n1317) );
  MOAI22D1BWP12T U1812 ( .A1(n1317), .A2(n1832), .B1(n1836), .B2(
        DEC_RF_offset_b[6]), .ZN(n803) );
  CKND0BWP12T U1813 ( .I(DEC_RF_alu_write_to_reg[4]), .ZN(n1324) );
  CKND2D0BWP12T U1814 ( .A1(n1795), .A2(n1684), .ZN(n1318) );
  NR2D1BWP12T U1815 ( .A1(n1824), .A2(n1318), .ZN(n1418) );
  MOAI22D1BWP12T U1816 ( .A1(n1320), .A2(n1713), .B1(n1745), .B2(n1319), .ZN(
        n1763) );
  AOI21D1BWP12T U1817 ( .A1(n1418), .A2(n1414), .B(n1763), .ZN(n1601) );
  INVD1BWP12T U1818 ( .I(n1743), .ZN(n1672) );
  ND4D1BWP12T U1819 ( .A1(n1601), .A2(n1672), .A3(n1759), .A4(n1786), .ZN(
        n1373) );
  ND2D1BWP12T U1820 ( .A1(n1739), .A2(n1321), .ZN(n1813) );
  INVD0BWP12T U1821 ( .I(n1813), .ZN(n1322) );
  OAI21D0BWP12T U1822 ( .A1(n1373), .A2(n1322), .B(n1790), .ZN(n1323) );
  OAI211D0BWP12T U1823 ( .A1(n1364), .A2(n1324), .B(n1323), .C(n1692), .ZN(
        n815) );
  CKND0BWP12T U1824 ( .I(DEC_ALU_alu_opcode[1]), .ZN(n1337) );
  CKND0BWP12T U1825 ( .I(n1699), .ZN(n1326) );
  NR2D0BWP12T U1826 ( .A1(n1326), .A2(n1378), .ZN(n1673) );
  AOI22D0BWP12T U1827 ( .A1(n1673), .A2(n1795), .B1(n1402), .B2(n1403), .ZN(
        n1325) );
  OAI211D1BWP12T U1828 ( .A1(n1713), .A2(n1326), .B(n1813), .C(n1325), .ZN(
        n1334) );
  INVD1BWP12T U1829 ( .I(n1327), .ZN(n1655) );
  INVD1BWP12T U1830 ( .I(n1332), .ZN(n1616) );
  OAI21D1BWP12T U1831 ( .A1(n1818), .A2(n1616), .B(n1817), .ZN(n1829) );
  NR2D1BWP12T U1832 ( .A1(n1829), .A2(n1821), .ZN(n1363) );
  TPOAI31D0BWP12T U1833 ( .A1(n1334), .A2(n1763), .A3(n1363), .B(n1809), .ZN(
        n1336) );
  INVD0BWP12T U1834 ( .I(n1824), .ZN(n1406) );
  OAI21D0BWP12T U1835 ( .A1(n1826), .A2(n1406), .B(n1723), .ZN(n1335) );
  OAI211D0BWP12T U1836 ( .A1(n1364), .A2(n1337), .B(n1336), .C(n1335), .ZN(
        n850) );
  NR2D0BWP12T U1837 ( .A1(n1338), .A2(n1795), .ZN(n1381) );
  INVD1BWP12T U1838 ( .I(n1381), .ZN(n1339) );
  CKND2D1BWP12T U1839 ( .A1(n1339), .A2(n1384), .ZN(n1768) );
  NR2XD0BWP12T U1840 ( .A1(n1768), .A2(n1779), .ZN(n1808) );
  NR2D1BWP12T U1841 ( .A1(n1808), .A2(n1821), .ZN(n1366) );
  ND2D1BWP12T U1842 ( .A1(n1737), .A2(n1340), .ZN(n1362) );
  INVD1BWP12T U1843 ( .I(n1362), .ZN(n1784) );
  TPNR2D0BWP12T U1844 ( .A1(n1342), .A2(n1341), .ZN(n1801) );
  TPNR2D0BWP12T U1845 ( .A1(n1345), .A2(n1344), .ZN(n1346) );
  ND2D1BWP12T U1846 ( .A1(n1619), .A2(n1641), .ZN(n1777) );
  INVD1BWP12T U1847 ( .I(n1658), .ZN(n1804) );
  ND2D0BWP12T U1848 ( .A1(n865), .A2(n1348), .ZN(n1776) );
  ND3D1BWP12T U1849 ( .A1(n1804), .A2(n1776), .A3(n1802), .ZN(n1356) );
  OR3D1BWP12T U1850 ( .A1(n1801), .A2(n1777), .A3(n1356), .Z(n1815) );
  INVD1BWP12T U1851 ( .I(n1814), .ZN(n1778) );
  INVD1BWP12T U1852 ( .I(n1693), .ZN(n1648) );
  CKND2D0BWP12T U1853 ( .A1(n1655), .A2(n1629), .ZN(n1352) );
  OR4D0BWP12T U1854 ( .A1(n1353), .A2(n1772), .A3(n1352), .A4(n1351), .Z(n1360) );
  CKND0BWP12T U1855 ( .I(n1370), .ZN(n1359) );
  CKND2D0BWP12T U1856 ( .A1(n1768), .A2(n1790), .ZN(n1646) );
  NR2XD0BWP12T U1857 ( .A1(n1355), .A2(n1354), .ZN(n1800) );
  INR3XD0BWP12T U1858 ( .A1(n1800), .B1(n1775), .B2(n1356), .ZN(n1357) );
  OAI22D1BWP12T U1859 ( .A1(n1646), .A2(n1788), .B1(n1357), .B2(n1661), .ZN(
        n1358) );
  AOI211D1BWP12T U1860 ( .A1(n1648), .A2(n1360), .B(n1359), .C(n1358), .ZN(
        n1791) );
  TPNR2D0BWP12T U1861 ( .A1(n1363), .A2(n1814), .ZN(n1365) );
  INVD1BWP12T U1862 ( .I(DEC_MISC_OUT_memory_address_source_is_reg), .ZN(n1481) );
  OAI22D0BWP12T U1863 ( .A1(n1365), .A2(n1832), .B1(n1481), .B2(n1364), .ZN(
        n836) );
  TPOAI31D0BWP12T U1864 ( .A1(n1784), .A2(n1367), .A3(n1366), .B(n1790), .ZN(
        n1369) );
  TPOAI21D0BWP12T U1865 ( .A1(n1648), .A2(n1656), .B(n1830), .ZN(n1368) );
  CKND2D1BWP12T U1866 ( .A1(n1369), .A2(n1368), .ZN(n1792) );
  INVD1BWP12T U1867 ( .I(n1792), .ZN(n1653) );
  CKND2D1BWP12T U1868 ( .A1(n1370), .A2(n1653), .ZN(n1371) );
  AO21D0BWP12T U1869 ( .A1(n1836), .A2(DEC_RF_memory_write_to_reg[4]), .B(
        n1371), .Z(n820) );
  AO211D0BWP12T U1870 ( .A1(n1836), .A2(DEC_RF_memory_write_to_reg[3]), .B(
        n1371), .C(n1651), .Z(n821) );
  NR2XD0BWP12T U1871 ( .A1(n1372), .A2(n1684), .ZN(n1751) );
  NR3XD0BWP12T U1872 ( .A1(n1373), .A2(n1826), .A3(n1751), .ZN(n1706) );
  INVD0BWP12T U1873 ( .I(n1706), .ZN(n1374) );
  NR2D1BWP12T U1874 ( .A1(n1374), .A2(n1606), .ZN(n1623) );
  AOI22D0BWP12T U1875 ( .A1(n1753), .A2(IF_DEC_instruction[2]), .B1(n1675), 
        .B2(n1748), .ZN(n1375) );
  TPAOI21D0BWP12T U1876 ( .A1(n1623), .A2(n1375), .B(n1757), .ZN(n1376) );
  INVD1BWP12T U1877 ( .I(n1692), .ZN(n1761) );
  AO211D0BWP12T U1878 ( .A1(n1836), .A2(DEC_RF_alu_write_to_reg[2]), .B(n1376), 
        .C(n1761), .Z(n818) );
  INR3XD0BWP12T U1879 ( .A1(n1377), .B1(n1814), .B2(n1606), .ZN(n1386) );
  INVD0BWP12T U1880 ( .I(n1386), .ZN(n1380) );
  OAI211D0BWP12T U1881 ( .A1(n1410), .A2(n1712), .B(n1603), .C(n1378), .ZN(
        n1379) );
  AOI211D0BWP12T U1882 ( .A1(n1787), .A2(n1381), .B(n1380), .C(n1379), .ZN(
        n1383) );
  TPND2D0BWP12T U1883 ( .A1(n1836), .A2(DEC_MEMCTRL_load_store_width[1]), .ZN(
        n1382) );
  OAI211D0BWP12T U1884 ( .A1(n1757), .A2(n1383), .B(n1692), .C(n1382), .ZN(
        n837) );
  NR2XD0BWP12T U1885 ( .A1(n1713), .A2(n1820), .ZN(n1597) );
  NR2D1BWP12T U1886 ( .A1(n1390), .A2(n1389), .ZN(n1626) );
  AO21D0BWP12T U1887 ( .A1(n1836), .A2(DEC_RF_memory_store_address_reg[4]), 
        .B(n1626), .Z(n831) );
  AO21D1BWP12T U1888 ( .A1(n1390), .A2(n1742), .B(n1389), .Z(n1756) );
  AOI22D0BWP12T U1889 ( .A1(n1656), .A2(n1675), .B1(n1836), .B2(
        DEC_RF_memory_store_address_reg[2]), .ZN(n1391) );
  CKND2D1BWP12T U1890 ( .A1(n1756), .A2(n1391), .ZN(n833) );
  AOI22D0BWP12T U1891 ( .A1(n1656), .A2(n1714), .B1(n1836), .B2(
        DEC_RF_memory_store_address_reg[0]), .ZN(n1392) );
  CKND2D1BWP12T U1892 ( .A1(n1756), .A2(n1392), .ZN(n835) );
  ND2D1BWP12T U1893 ( .A1(n1670), .A2(n1809), .ZN(n1469) );
  TPND2D0BWP12T U1894 ( .A1(n1836), .A2(DEC_RF_offset_b[18]), .ZN(n1393) );
  OAI211D0BWP12T U1895 ( .A1(n1823), .A2(n1469), .B(n1393), .C(n1696), .ZN(
        n791) );
  INVD1BWP12T U1896 ( .I(IF_DEC_instruction[1]), .ZN(n1783) );
  TPND2D0BWP12T U1897 ( .A1(n1836), .A2(DEC_RF_offset_b[17]), .ZN(n1394) );
  OAI211D0BWP12T U1898 ( .A1(n1709), .A2(n1469), .B(n1394), .C(n1696), .ZN(
        n792) );
  CKND0BWP12T U1899 ( .I(IF_DEC_instruction[4]), .ZN(n1604) );
  TPND2D0BWP12T U1900 ( .A1(n1836), .A2(DEC_RF_offset_b[16]), .ZN(n1395) );
  OAI211D0BWP12T U1901 ( .A1(n1604), .A2(n1469), .B(n1395), .C(n1696), .ZN(
        n793) );
  TPND2D0BWP12T U1902 ( .A1(n1836), .A2(DEC_RF_offset_b[14]), .ZN(n1397) );
  OAI211D0BWP12T U1903 ( .A1(n1788), .A2(n1469), .B(n1397), .C(n1696), .ZN(
        n795) );
  TPND2D0BWP12T U1904 ( .A1(n1836), .A2(DEC_RF_offset_b[22]), .ZN(n1398) );
  OAI211D0BWP12T U1905 ( .A1(n1787), .A2(n1469), .B(n1398), .C(n1696), .ZN(
        n787) );
  TPND2D0BWP12T U1906 ( .A1(n1836), .A2(DEC_RF_offset_b[21]), .ZN(n1399) );
  OAI211D0BWP12T U1907 ( .A1(n1822), .A2(n1469), .B(n1399), .C(n1696), .ZN(
        n788) );
  TPND2D0BWP12T U1908 ( .A1(n1836), .A2(DEC_RF_offset_b[19]), .ZN(n1400) );
  OAI211D0BWP12T U1909 ( .A1(n1827), .A2(n1469), .B(n1400), .C(n1696), .ZN(
        n790) );
  CKND0BWP12T U1910 ( .I(n1414), .ZN(n1417) );
  CKND2D0BWP12T U1911 ( .A1(n1684), .A2(n1417), .ZN(n1401) );
  OAI211D0BWP12T U1912 ( .A1(n1827), .A2(n1669), .B(n1412), .C(n1401), .ZN(
        n1405) );
  NR2D0BWP12T U1913 ( .A1(n1713), .A2(n1402), .ZN(n1404) );
  AOI211D0BWP12T U1914 ( .A1(n1406), .A2(n1405), .B(n1404), .C(n1403), .ZN(
        n1409) );
  CKND0BWP12T U1915 ( .I(n1407), .ZN(n1408) );
  TPND2D0BWP12T U1916 ( .A1(n1790), .A2(n1408), .ZN(n1599) );
  AOI22D0BWP12T U1917 ( .A1(n1763), .A2(n1809), .B1(n1723), .B2(n1418), .ZN(
        n1419) );
  OAI21D0BWP12T U1918 ( .A1(n1409), .A2(n1599), .B(n1419), .ZN(
        irdecode_inst1_next_update_flag_c) );
  CKND0BWP12T U1919 ( .I(n1673), .ZN(n1411) );
  ND3D0BWP12T U1920 ( .A1(n1718), .A2(n1830), .A3(n1410), .ZN(n1671) );
  CKND2D0BWP12T U1921 ( .A1(n1411), .A2(n1671), .ZN(n1416) );
  CKND2D0BWP12T U1922 ( .A1(n1823), .A2(IF_DEC_instruction[7]), .ZN(n1413) );
  AOI211D0BWP12T U1923 ( .A1(n1414), .A2(n1413), .B(n1824), .C(n1412), .ZN(
        n1415) );
  AOI211D0BWP12T U1924 ( .A1(n1418), .A2(n1417), .B(n1416), .C(n1415), .ZN(
        n1420) );
  OAI21D0BWP12T U1925 ( .A1(n1420), .A2(n1599), .B(n1419), .ZN(
        irdecode_inst1_next_update_flag_v) );
  IOA21D0BWP12T U1926 ( .A1(n1836), .A2(DEC_RF_offset_b[23]), .B(n1696), .ZN(
        n786) );
  IOA21D0BWP12T U1927 ( .A1(n1836), .A2(DEC_RF_offset_b[30]), .B(n1696), .ZN(
        n779) );
  IOA21D0BWP12T U1928 ( .A1(n1836), .A2(DEC_RF_offset_b[29]), .B(n1696), .ZN(
        n780) );
  IOA21D0BWP12T U1929 ( .A1(n1836), .A2(DEC_RF_offset_b[31]), .B(n1696), .ZN(
        n777) );
  IOA21D0BWP12T U1930 ( .A1(n1836), .A2(DEC_RF_offset_b[28]), .B(n1696), .ZN(
        n781) );
  TPND2D0BWP12T U1931 ( .A1(n1836), .A2(DEC_RF_memory_store_address_reg[1]), 
        .ZN(n1421) );
  TPOAI31D0BWP12T U1932 ( .A1(n1822), .A2(n1832), .A3(n1778), .B(n1421), .ZN(
        n834) );
  IOA21D0BWP12T U1933 ( .A1(n1836), .A2(DEC_RF_offset_b[27]), .B(n1696), .ZN(
        n782) );
  IOA21D0BWP12T U1934 ( .A1(n1836), .A2(DEC_RF_offset_b[26]), .B(n1696), .ZN(
        n783) );
  IOA21D0BWP12T U1935 ( .A1(n1836), .A2(DEC_RF_offset_b[25]), .B(n1696), .ZN(
        n784) );
  CKND0BWP12T U1936 ( .I(n1737), .ZN(n1423) );
  TPND2D0BWP12T U1937 ( .A1(n1836), .A2(
        DEC_MEMCTRL_memorycontroller_sign_extend), .ZN(n1422) );
  TPOAI31D0BWP12T U1938 ( .A1(n1830), .A2(n1832), .A3(n1423), .B(n1422), .ZN(
        n839) );
  IOA21D0BWP12T U1939 ( .A1(n1836), .A2(DEC_RF_offset_b[24]), .B(n1696), .ZN(
        n785) );
  HICOND1BWP12T U1940 ( .A(RF_pc_out[27]), .CI(n1424), .CON(n1265), .S(n1425)
         );
  HICIND1BWP12T U1941 ( .A(RF_pc_out[26]), .CIN(n1426), .CO(n1424), .S(n1427)
         );
  MUX2NXD0BWP12T U1942 ( .I0(MEMCTRL_RF_IF_data_in[13]), .I1(
        Instruction_Fetch_inst1_fetched_instruction_reg_13_), .S(n754), .ZN(
        n1429) );
  CKND2D1BWP12T U1943 ( .A1(n1429), .A2(n1435), .ZN(
        Instruction_Fetch_inst1_N96) );
  MUX2NXD0BWP12T U1944 ( .I0(MEMCTRL_RF_IF_data_in[10]), .I1(
        Instruction_Fetch_inst1_fetched_instruction_reg_10_), .S(n754), .ZN(
        n1430) );
  CKND2D1BWP12T U1945 ( .A1(n1430), .A2(n1435), .ZN(
        Instruction_Fetch_inst1_N93) );
  MUX2NXD0BWP12T U1946 ( .I0(MEMCTRL_RF_IF_data_in[11]), .I1(
        Instruction_Fetch_inst1_fetched_instruction_reg_11_), .S(n754), .ZN(
        n1431) );
  CKND2D1BWP12T U1947 ( .A1(n1431), .A2(n1435), .ZN(
        Instruction_Fetch_inst1_N94) );
  MUX2NXD0BWP12T U1948 ( .I0(MEMCTRL_RF_IF_data_in[9]), .I1(
        Instruction_Fetch_inst1_fetched_instruction_reg_9_), .S(n754), .ZN(
        n1432) );
  CKND2D1BWP12T U1949 ( .A1(n1432), .A2(n1435), .ZN(
        Instruction_Fetch_inst1_N92) );
  MUX2NXD0BWP12T U1950 ( .I0(MEMCTRL_RF_IF_data_in[8]), .I1(
        Instruction_Fetch_inst1_fetched_instruction_reg_8_), .S(n754), .ZN(
        n1433) );
  CKND2D1BWP12T U1951 ( .A1(n1433), .A2(n1435), .ZN(
        Instruction_Fetch_inst1_N91) );
  MUX2NXD0BWP12T U1952 ( .I0(MEMCTRL_RF_IF_data_in[15]), .I1(
        Instruction_Fetch_inst1_fetched_instruction_reg_15_), .S(n754), .ZN(
        n1434) );
  CKND2D1BWP12T U1953 ( .A1(n1434), .A2(n1435), .ZN(
        Instruction_Fetch_inst1_N98) );
  MUX2NXD0BWP12T U1954 ( .I0(MEMCTRL_RF_IF_data_in[12]), .I1(
        Instruction_Fetch_inst1_fetched_instruction_reg_12_), .S(n754), .ZN(
        n1436) );
  CKND2D1BWP12T U1955 ( .A1(n1436), .A2(n1435), .ZN(
        Instruction_Fetch_inst1_N95) );
  BUFFD12BWP12T U1956 ( .I(RF_ALU_operand_b[1]), .Z(n1850) );
  AOI211D0BWP12T U1957 ( .A1(DEC_MEMCTRL_load_store_width[1]), .A2(
        DEC_MEMCTRL_load_store_width[0]), .B(n1579), .C(reset), .ZN(n1439) );
  NR2D0BWP12T U1958 ( .A1(DEC_MEMCTRL_memory_load_request), .A2(
        Instruction_Fetch_inst1_currentState_1_), .ZN(n1583) );
  ND3XD0BWP12T U1959 ( .A1(n1439), .A2(DEC_MEMCTRL_memory_store_request), .A3(
        n1583), .ZN(n1445) );
  OR2XD1BWP12T U1960 ( .A1(DEC_MEMCTRL_load_store_width[1]), .A2(
        DEC_MEMCTRL_load_store_width[0]), .Z(n1532) );
  INVD1BWP12T U1961 ( .I(n1532), .ZN(n1480) );
  OA21XD0BWP12T U1962 ( .A1(memory_interface_inst1_fsm_state_3_), .A2(n1444), 
        .B(n1485), .Z(n1438) );
  TPOAI22D0BWP12T U1963 ( .A1(n1445), .A2(n1480), .B1(reset), .B2(n1438), .ZN(
        memory_interface_inst1_fsm_N34) );
  CKND0BWP12T U1964 ( .I(n1439), .ZN(n1440) );
  OAI31D0BWP12T U1965 ( .A1(n1480), .A2(n1583), .A3(n1440), .B(n1445), .ZN(
        memory_interface_inst1_fsm_N32) );
  NR2D1BWP12T U1966 ( .A1(n1441), .A2(n1281), .ZN(n1442) );
  CKND0BWP12T U1967 ( .I(RF_pc_out[13]), .ZN(n1446) );
  INR2D0BWP12T U1968 ( .A1(memory_interface_inst1_fsm_state_3_), .B1(n1444), 
        .ZN(n1491) );
  CKND1BWP12T U1969 ( .I(n1485), .ZN(n1576) );
  NR2D1BWP12T U1970 ( .A1(n1491), .A2(n1576), .ZN(n1479) );
  OAI21D0BWP12T U1971 ( .A1(reset), .A2(n1479), .B(n1445), .ZN(
        memory_interface_inst1_fsm_N35) );
  INVD1BWP12T U1972 ( .I(n1448), .ZN(n1457) );
  NR2D1BWP12T U1973 ( .A1(n1457), .A2(n1449), .ZN(n1456) );
  CKND2D1BWP12T U1974 ( .A1(n1456), .A2(RF_pc_out[7]), .ZN(n1451) );
  CKND0BWP12T U1975 ( .I(RF_pc_out[8]), .ZN(n1450) );
  XOR2D1BWP12T U1976 ( .A1(n1451), .A2(n1450), .Z(n1452) );
  AN2D0BWP12T U1977 ( .A1(n1452), .A2(n1458), .Z(IF_RF_incremented_pc_out[8])
         );
  INVD0BWP12T U1978 ( .I(RF_pc_out[9]), .ZN(n1453) );
  XNR2XD1BWP12T U1979 ( .A1(n1454), .A2(n1453), .ZN(n1455) );
  AN2D0BWP12T U1980 ( .A1(n1455), .A2(n1458), .Z(IF_RF_incremented_pc_out[9])
         );
  NR2D0BWP12T U1981 ( .A1(DEC_ALU_alu_opcode[3]), .A2(DEC_ALU_alu_opcode[0]), 
        .ZN(n1461) );
  ND3D0BWP12T U1982 ( .A1(n1461), .A2(DEC_ALU_alu_opcode[1]), .A3(
        DEC_ALU_alu_opcode[2]), .ZN(n1462) );
  MUX2NXD0BWP12T U1983 ( .I0(n1463), .I1(n1462), .S(DEC_ALU_alu_opcode[4]), 
        .ZN(ALU_IN_c) );
  INR2D1BWP12T U1984 ( .A1(RF_OUT_c), .B1(DEC_CPSR_update_flag_c), .ZN(n1464)
         );
  TPND2D2BWP12T U1985 ( .A1(ALU_OUT_z), .A2(DEC_CPSR_update_flag_z), .ZN(n1467) );
  ND2D1BWP12T U1986 ( .A1(n1839), .A2(RF_OUT_z), .ZN(n1466) );
  ND2D2BWP12T U1987 ( .A1(n1467), .A2(n1466), .ZN(new_z) );
  TPND2D0BWP12T U1988 ( .A1(n1836), .A2(DEC_RF_offset_b[20]), .ZN(n1468) );
  OAI211D0BWP12T U1989 ( .A1(n1684), .A2(n1469), .B(n1468), .C(n1696), .ZN(
        n789) );
  CKND2D0BWP12T U1990 ( .A1(n1691), .A2(IF_DEC_instruction[4]), .ZN(n1473) );
  INVD0BWP12T U1991 ( .I(n1603), .ZN(n1682) );
  OAI22D0BWP12T U1992 ( .A1(n1822), .A2(n1683), .B1(n1470), .B2(n1821), .ZN(
        n1471) );
  AOI211D0BWP12T U1993 ( .A1(n1682), .A2(IF_DEC_instruction[1]), .B(n1471), 
        .C(n1794), .ZN(n1472) );
  ND4D1BWP12T U1994 ( .A1(n1760), .A2(n1473), .A3(n1472), .A4(n1749), .ZN(
        n1474) );
  AO22XD0BWP12T U1995 ( .A1(n1474), .A2(n1809), .B1(n1836), .B2(n999), .Z(n814) );
  BUFFXD16BWP12T U1996 ( .I(RF_ALU_operand_b[0]), .Z(n1849) );
  INVD1BWP12T U1997 ( .I(ALU_OUT_v), .ZN(n1477) );
  INR2D1BWP12T U1998 ( .A1(RF_OUT_v), .B1(DEC_CPSR_update_flag_v), .ZN(n1475)
         );
  INVD1BWP12T U1999 ( .I(n1475), .ZN(n1476) );
  TPOAI21D1BWP12T U2000 ( .A1(n1477), .A2(n1844), .B(n1476), .ZN(new_v) );
  INVD1BWP12T U2001 ( .I(n1841), .ZN(irdecode_inst1_N907) );
  CKND2D0BWP12T U2002 ( .A1(n1478), .A2(n1586), .ZN(n1534) );
  OAI31D1BWP12T U2003 ( .A1(n1480), .A2(n1580), .A3(n1534), .B(n1479), .ZN(
        MEMCTRL_MEM_to_mem_write_enable) );
  NR2D1BWP12T U2004 ( .A1(DEC_MISC_OUT_memory_address_source_is_reg), .A2(
        Instruction_Fetch_inst1_currentState_1_), .ZN(n1566) );
  NR2XD0BWP12T U2005 ( .A1(n1481), .A2(Instruction_Fetch_inst1_currentState_1_), .ZN(n1569) );
  INVD1BWP12T U2006 ( .I(MEMCTRL_IN_address[11]), .ZN(n1490) );
  ND2D1BWP12T U2007 ( .A1(memory_interface_inst1_delay_addr_for_adder[0]), 
        .A2(memory_interface_inst1_delay_addr_for_adder[1]), .ZN(n1541) );
  NR2D1BWP12T U2008 ( .A1(n1541), .A2(n1848), .ZN(n1564) );
  AN3XD1BWP12T U2009 ( .A1(n1564), .A2(
        memory_interface_inst1_delay_addr_for_adder[3]), .A3(
        memory_interface_inst1_delay_addr_for_adder[4]), .Z(n1546) );
  AN3XD1BWP12T U2010 ( .A1(n1546), .A2(
        memory_interface_inst1_delay_addr_for_adder[5]), .A3(
        memory_interface_inst1_delay_addr_for_adder[6]), .Z(n1522) );
  ND3D1BWP12T U2011 ( .A1(n1522), .A2(
        memory_interface_inst1_delay_addr_for_adder[7]), .A3(
        memory_interface_inst1_delay_addr_for_adder[8]), .ZN(n1486) );
  CKND2D0BWP12T U2012 ( .A1(n1730), .A2(n1483), .ZN(n1535) );
  NR2D1BWP12T U2013 ( .A1(n1484), .A2(n1535), .ZN(n1492) );
  ND2D1BWP12T U2014 ( .A1(n1492), .A2(n1485), .ZN(n1557) );
  ND2D1BWP12T U2015 ( .A1(n1557), .A2(n1562), .ZN(n1572) );
  IND4D1BWP12T U2016 ( .A1(memory_interface_inst1_delay_addr_for_adder[11]), 
        .B1(memory_interface_inst1_delay_addr_for_adder[10]), .B2(n1514), .B3(
        memory_interface_inst1_delay_addr_for_adder[9]), .ZN(n1489) );
  NR2D1BWP12T U2017 ( .A1(memory_interface_inst1_delay_addr_for_adder[10]), 
        .A2(n1572), .ZN(n1487) );
  INVD1BWP12T U2018 ( .I(n1572), .ZN(n1556) );
  INVD1BWP12T U2019 ( .I(n1557), .ZN(n1551) );
  AOI21D1BWP12T U2020 ( .A1(n1556), .A2(n1486), .B(n1551), .ZN(n1515) );
  OAI21D1BWP12T U2021 ( .A1(memory_interface_inst1_delay_addr_for_adder[9]), 
        .A2(n1572), .B(n1515), .ZN(n1512) );
  OAI21D1BWP12T U2022 ( .A1(n1487), .A2(n1512), .B(
        memory_interface_inst1_delay_addr_for_adder[11]), .ZN(n1488) );
  OAI211D1BWP12T U2023 ( .A1(n1490), .A2(n1562), .B(n1489), .C(n1488), .ZN(
        MEMCTRL_MEM_to_mem_address[11]) );
  INVD1BWP12T U2024 ( .I(n1491), .ZN(n1584) );
  ND2D1BWP12T U2025 ( .A1(n1584), .A2(n1493), .ZN(n1575) );
  NR2D1BWP12T U2026 ( .A1(n1492), .A2(n1534), .ZN(n1577) );
  INVD1BWP12T U2027 ( .I(RF_MEMCTRL_data_reg[15]), .ZN(n1496) );
  INVD1BWP12T U2028 ( .I(n1577), .ZN(n1509) );
  INVD1BWP12T U2029 ( .I(MEM_MEMCTRL_from_mem_data[7]), .ZN(n1727) );
  MAOI22D0BWP12T U2030 ( .A1(n1576), .A2(
        memory_interface_inst1_delay_data_in32[31]), .B1(n1727), .B2(n1557), 
        .ZN(n1495) );
  INVD1BWP12T U2031 ( .I(n1493), .ZN(n1506) );
  ND2D1BWP12T U2032 ( .A1(n1506), .A2(
        memory_interface_inst1_delay_data_in32[15]), .ZN(n1494) );
  OAI211D1BWP12T U2033 ( .A1(n1496), .A2(n1509), .B(n1495), .C(n1494), .ZN(
        MEMCTRL_MEM_to_mem_data[7]) );
  INVD1BWP12T U2034 ( .I(RF_MEMCTRL_data_reg[14]), .ZN(n1499) );
  INVD1BWP12T U2035 ( .I(MEM_MEMCTRL_from_mem_data[6]), .ZN(n1728) );
  MAOI22D0BWP12T U2036 ( .A1(n1576), .A2(
        memory_interface_inst1_delay_data_in32[30]), .B1(n1728), .B2(n1557), 
        .ZN(n1498) );
  ND2D1BWP12T U2037 ( .A1(n1506), .A2(
        memory_interface_inst1_delay_data_in32[14]), .ZN(n1497) );
  OAI211D1BWP12T U2038 ( .A1(n1499), .A2(n1509), .B(n1498), .C(n1497), .ZN(
        MEMCTRL_MEM_to_mem_data[6]) );
  INVD1BWP12T U2039 ( .I(RF_MEMCTRL_data_reg[13]), .ZN(n1502) );
  INVD1BWP12T U2040 ( .I(MEM_MEMCTRL_from_mem_data[5]), .ZN(n1726) );
  MAOI22D0BWP12T U2041 ( .A1(n1576), .A2(
        memory_interface_inst1_delay_data_in32[29]), .B1(n1726), .B2(n1557), 
        .ZN(n1501) );
  ND2D1BWP12T U2042 ( .A1(n1506), .A2(
        memory_interface_inst1_delay_data_in32[13]), .ZN(n1500) );
  OAI211D1BWP12T U2043 ( .A1(n1502), .A2(n1509), .B(n1501), .C(n1500), .ZN(
        MEMCTRL_MEM_to_mem_data[5]) );
  INVD1BWP12T U2044 ( .I(RF_MEMCTRL_data_reg[12]), .ZN(n1505) );
  INVD1BWP12T U2045 ( .I(MEM_MEMCTRL_from_mem_data[4]), .ZN(n1725) );
  MAOI22D0BWP12T U2046 ( .A1(n1576), .A2(
        memory_interface_inst1_delay_data_in32[28]), .B1(n1725), .B2(n1557), 
        .ZN(n1504) );
  ND2D1BWP12T U2047 ( .A1(n1506), .A2(
        memory_interface_inst1_delay_data_in32[12]), .ZN(n1503) );
  OAI211D1BWP12T U2048 ( .A1(n1505), .A2(n1509), .B(n1504), .C(n1503), .ZN(
        MEMCTRL_MEM_to_mem_data[4]) );
  INVD1BWP12T U2049 ( .I(RF_MEMCTRL_data_reg[8]), .ZN(n1510) );
  AOI22D1BWP12T U2050 ( .A1(n1576), .A2(
        memory_interface_inst1_delay_data_in32[24]), .B1(n1551), .B2(
        MEM_MEMCTRL_from_mem_data[0]), .ZN(n1508) );
  ND2D1BWP12T U2051 ( .A1(n1506), .A2(
        memory_interface_inst1_delay_data_in32[8]), .ZN(n1507) );
  OAI211D1BWP12T U2052 ( .A1(n1510), .A2(n1509), .B(n1508), .C(n1507), .ZN(
        MEMCTRL_MEM_to_mem_data[0]) );
  INVD1BWP12T U2053 ( .I(n1562), .ZN(n1574) );
  INVD1BWP12T U2054 ( .I(MEMCTRL_IN_address[8]), .ZN(n1520) );
  IND4D1BWP12T U2055 ( .A1(memory_interface_inst1_delay_addr_for_adder[8]), 
        .B1(n1522), .B2(n1556), .B3(
        memory_interface_inst1_delay_addr_for_adder[7]), .ZN(n1519) );
  NR2D1BWP12T U2056 ( .A1(memory_interface_inst1_delay_addr_for_adder[7]), 
        .A2(n1574), .ZN(n1517) );
  OAI21D1BWP12T U2057 ( .A1(n1522), .A2(n1574), .B(n1557), .ZN(n1523) );
  OAI21D1BWP12T U2058 ( .A1(n1517), .A2(n1523), .B(
        memory_interface_inst1_delay_addr_for_adder[8]), .ZN(n1518) );
  OAI211D1BWP12T U2059 ( .A1(n1562), .A2(n1520), .B(n1519), .C(n1518), .ZN(
        MEMCTRL_MEM_to_mem_address[8]) );
  INVD1BWP12T U2060 ( .I(n1522), .ZN(n1525) );
  ND2D1BWP12T U2061 ( .A1(memory_interface_inst1_delay_addr_for_adder[7]), 
        .A2(n1523), .ZN(n1524) );
  OAI31D1BWP12T U2062 ( .A1(memory_interface_inst1_delay_addr_for_adder[7]), 
        .A2(n1525), .A3(n1572), .B(n1524), .ZN(n1526) );
  AO21D1BWP12T U2063 ( .A1(n1574), .A2(MEMCTRL_IN_address[7]), .B(n1526), .Z(
        MEMCTRL_MEM_to_mem_address[7]) );
  INVD1BWP12T U2064 ( .I(MEMCTRL_IN_address[6]), .ZN(n1531) );
  IND4D1BWP12T U2065 ( .A1(memory_interface_inst1_delay_addr_for_adder[6]), 
        .B1(n1546), .B2(n1556), .B3(
        memory_interface_inst1_delay_addr_for_adder[5]), .ZN(n1530) );
  NR2D1BWP12T U2066 ( .A1(memory_interface_inst1_delay_addr_for_adder[5]), 
        .A2(n1574), .ZN(n1528) );
  OAI21D1BWP12T U2067 ( .A1(n1546), .A2(n1574), .B(n1557), .ZN(n1547) );
  OAI21D1BWP12T U2068 ( .A1(n1528), .A2(n1547), .B(
        memory_interface_inst1_delay_addr_for_adder[6]), .ZN(n1529) );
  OAI211D1BWP12T U2069 ( .A1(n1562), .A2(n1531), .B(n1530), .C(n1529), .ZN(
        MEMCTRL_MEM_to_mem_address[6]) );
  AOI21D1BWP12T U2070 ( .A1(n1583), .A2(n1532), .B(n1534), .ZN(n1533) );
  AO21D1BWP12T U2071 ( .A1(n1535), .A2(n1534), .B(n1533), .Z(
        MEMCTRL_MEM_to_mem_read_enable) );
  TPND2D0BWP12T U2072 ( .A1(ALU_MISC_OUT_result[3]), .A2(n1566), .ZN(n1538) );
  AOI22D0BWP12T U2073 ( .A1(RF_MEMCTRL_address_reg[3]), .A2(n1569), .B1(n1568), 
        .B2(n1536), .ZN(n1537) );
  ND2D1BWP12T U2074 ( .A1(n1538), .A2(n1537), .ZN(MEMCTRL_IN_address[2]) );
  NR2D1BWP12T U2075 ( .A1(memory_interface_inst1_delay_addr_for_adder[1]), 
        .A2(n1574), .ZN(n1539) );
  OAI21D1BWP12T U2076 ( .A1(memory_interface_inst1_delay_addr_for_adder[0]), 
        .A2(n1574), .B(n1557), .ZN(n1570) );
  OAI21D1BWP12T U2077 ( .A1(n1539), .A2(n1570), .B(
        memory_interface_inst1_delay_addr_for_adder[2]), .ZN(n1540) );
  OAI31D1BWP12T U2078 ( .A1(memory_interface_inst1_delay_addr_for_adder[2]), 
        .A2(n1541), .A3(n1572), .B(n1540), .ZN(n1542) );
  AO21D1BWP12T U2079 ( .A1(n1574), .A2(MEMCTRL_IN_address[2]), .B(n1542), .Z(
        MEMCTRL_MEM_to_mem_address[2]) );
  TPND2D0BWP12T U2080 ( .A1(ALU_MISC_OUT_result[6]), .A2(n1566), .ZN(n1545) );
  AOI22D0BWP12T U2081 ( .A1(RF_MEMCTRL_address_reg[6]), .A2(n1569), .B1(n1568), 
        .B2(n1543), .ZN(n1544) );
  ND2D1BWP12T U2082 ( .A1(n1545), .A2(n1544), .ZN(MEMCTRL_IN_address[5]) );
  INVD1BWP12T U2083 ( .I(n1546), .ZN(n1549) );
  ND2D1BWP12T U2084 ( .A1(memory_interface_inst1_delay_addr_for_adder[5]), 
        .A2(n1547), .ZN(n1548) );
  OAI31D1BWP12T U2085 ( .A1(memory_interface_inst1_delay_addr_for_adder[5]), 
        .A2(n1549), .A3(n1572), .B(n1548), .ZN(n1550) );
  AO21D1BWP12T U2086 ( .A1(n1574), .A2(MEMCTRL_IN_address[5]), .B(n1550), .Z(
        MEMCTRL_MEM_to_mem_address[5]) );
  AOI22D1BWP12T U2087 ( .A1(memory_interface_inst1_delay_addr_for_adder[0]), 
        .A2(n1551), .B1(MEMCTRL_IN_address[0]), .B2(n1574), .ZN(n1552) );
  OAI21D1BWP12T U2088 ( .A1(memory_interface_inst1_delay_addr_for_adder[0]), 
        .A2(n1572), .B(n1552), .ZN(MEMCTRL_MEM_to_mem_address[0]) );
  TPND2D0BWP12T U2089 ( .A1(ALU_MISC_OUT_result[5]), .A2(n1566), .ZN(n1555) );
  AOI22D0BWP12T U2090 ( .A1(RF_MEMCTRL_address_reg[5]), .A2(n1569), .B1(n1568), 
        .B2(n1553), .ZN(n1554) );
  ND2D1BWP12T U2091 ( .A1(n1555), .A2(n1554), .ZN(MEMCTRL_IN_address[4]) );
  INVD1BWP12T U2092 ( .I(MEMCTRL_IN_address[4]), .ZN(n1561) );
  IND4D1BWP12T U2093 ( .A1(memory_interface_inst1_delay_addr_for_adder[4]), 
        .B1(n1564), .B2(n1556), .B3(
        memory_interface_inst1_delay_addr_for_adder[3]), .ZN(n1560) );
  NR2D1BWP12T U2094 ( .A1(memory_interface_inst1_delay_addr_for_adder[3]), 
        .A2(n1574), .ZN(n1558) );
  OAI21D1BWP12T U2095 ( .A1(n1564), .A2(n1574), .B(n1557), .ZN(n1565) );
  OAI21D1BWP12T U2096 ( .A1(n1558), .A2(n1565), .B(
        memory_interface_inst1_delay_addr_for_adder[4]), .ZN(n1559) );
  OAI211D1BWP12T U2097 ( .A1(n1562), .A2(n1561), .B(n1560), .C(n1559), .ZN(
        MEMCTRL_MEM_to_mem_address[4]) );
  ND2D1BWP12T U2098 ( .A1(memory_interface_inst1_delay_addr_for_adder[1]), 
        .A2(n1570), .ZN(n1571) );
  OAI31D1BWP12T U2099 ( .A1(memory_interface_inst1_delay_addr_for_adder[1]), 
        .A2(n1847), .A3(n1572), .B(n1571), .ZN(n1573) );
  AO21D1BWP12T U2100 ( .A1(n1574), .A2(MEMCTRL_IN_address[1]), .B(n1573), .Z(
        MEMCTRL_MEM_to_mem_address[1]) );
  CKND0BWP12T U2101 ( .I(n1579), .ZN(n1582) );
  OAI21D0BWP12T U2102 ( .A1(DEC_MEMCTRL_load_store_width[1]), .A2(n1580), .B(
        n1583), .ZN(n1581) );
  OAI211D0BWP12T U2103 ( .A1(n1583), .A2(n1846), .B(n1582), .C(n1581), .ZN(
        n1585) );
  AOI21D1BWP12T U2104 ( .A1(n1585), .A2(n1584), .B(reset), .ZN(
        memory_interface_inst1_fsm_N33) );
  CKND0BWP12T U2105 ( .I(n1586), .ZN(n1588) );
  AOI21D1BWP12T U2106 ( .A1(n1588), .A2(n1587), .B(
        Instruction_Fetch_inst1_first_instruction_fetched), .ZN(n1589) );
  NR2D1BWP12T U2107 ( .A1(n1589), .A2(reset), .ZN(n862) );
  NR2D1BWP12T U2108 ( .A1(n1591), .A2(n1590), .ZN(n1595) );
  OAI22D1BWP12T U2109 ( .A1(n1595), .A2(n1592), .B1(n1823), .B2(n1593), .ZN(
        n854) );
  OAI22D1BWP12T U2110 ( .A1(n1595), .A2(n1845), .B1(n1709), .B2(n1593), .ZN(
        n855) );
  CKND0BWP12T U2111 ( .I(irdecode_inst1_itstate_7_), .ZN(n1594) );
  OAI22D1BWP12T U2112 ( .A1(n1595), .A2(n1594), .B1(n1827), .B2(n1593), .ZN(
        n853) );
  INVD1BWP12T U2113 ( .I(n1596), .ZN(n1598) );
  NR2D1BWP12T U2114 ( .A1(n1598), .A2(n1597), .ZN(n1600) );
  OAI22D1BWP12T U2115 ( .A1(n1601), .A2(n1832), .B1(n1600), .B2(n1599), .ZN(
        irdecode_inst1_next_update_flag_n) );
  INVD0BWP12T U2116 ( .I(n1723), .ZN(n1674) );
  OAI211D0BWP12T U2117 ( .A1(n1604), .A2(n1603), .B(n1602), .C(n1683), .ZN(
        n1607) );
  OAI31D0BWP12T U2118 ( .A1(n1607), .A2(n1606), .A3(n1605), .B(n1809), .ZN(
        n1609) );
  CKND2D0BWP12T U2119 ( .A1(n1836), .A2(n867), .ZN(n1608) );
  OAI211D1BWP12T U2120 ( .A1(n1612), .A2(n1674), .B(n1609), .C(n1608), .ZN(
        n843) );
  CKND2D0BWP12T U2121 ( .A1(n1745), .A2(n1790), .ZN(n1613) );
  CKND2D0BWP12T U2122 ( .A1(n1714), .A2(n1790), .ZN(n1662) );
  NR2D0BWP12T U2123 ( .A1(n1757), .A2(n1709), .ZN(n1610) );
  AOI22D1BWP12T U2124 ( .A1(n1682), .A2(n1610), .B1(n1836), .B2(n1003), .ZN(
        n1611) );
  OAI211D1BWP12T U2125 ( .A1(n1612), .A2(n1662), .B(n1755), .C(n1611), .ZN(
        n842) );
  OA21D1BWP12T U2126 ( .A1(n1613), .A2(n1827), .B(n1692), .Z(n1622) );
  NR2D1BWP12T U2127 ( .A1(n1620), .A2(n1617), .ZN(n1625) );
  AOI21D1BWP12T U2128 ( .A1(n1656), .A2(n1624), .B(n1626), .ZN(n1621) );
  NR2D1BWP12T U2129 ( .A1(n1624), .A2(n1777), .ZN(n1627) );
  CKND2D1BWP12T U2130 ( .A1(n1627), .A2(n1802), .ZN(n1659) );
  CKND0BWP12T U2131 ( .I(n1629), .ZN(n1631) );
  AOI211D0BWP12T U2132 ( .A1(irdecode_inst1_N545), .A2(n1632), .B(n1631), .C(
        n1630), .ZN(n1635) );
  ND4D0BWP12T U2133 ( .A1(n1636), .A2(n1635), .A3(n1634), .A4(n1633), .ZN(
        n1649) );
  CKND2D0BWP12T U2134 ( .A1(n1774), .A2(n1637), .ZN(n1638) );
  AOI211D0BWP12T U2135 ( .A1(n865), .A2(irdecode_inst1_N706), .B(n1639), .C(
        n1638), .ZN(n1643) );
  ND4D0BWP12T U2136 ( .A1(n1804), .A2(n1643), .A3(n1642), .A4(n1641), .ZN(
        n1644) );
  TPND2D0BWP12T U2137 ( .A1(n1644), .A2(n1656), .ZN(n1645) );
  OAI211D0BWP12T U2138 ( .A1(n1721), .A2(n1646), .B(n1692), .C(n1645), .ZN(
        n1647) );
  AOI21D1BWP12T U2139 ( .A1(n1649), .A2(n1648), .B(n1647), .ZN(n1668) );
  INVD1BWP12T U2140 ( .I(n1789), .ZN(n1793) );
  TPNR2D0BWP12T U2141 ( .A1(n1757), .A2(n1721), .ZN(n1664) );
  MOAI22D0BWP12T U2142 ( .A1(n1786), .A2(n1662), .B1(n1836), .B2(
        DEC_RF_memory_write_to_reg[0]), .ZN(n1650) );
  AOI211XD0BWP12T U2143 ( .A1(n1793), .A2(n1664), .B(n1651), .C(n1650), .ZN(
        n1652) );
  ND3D1BWP12T U2144 ( .A1(n1668), .A2(n1653), .A3(n1652), .ZN(n824) );
  OA21D1BWP12T U2145 ( .A1(n1655), .A2(n1693), .B(n1654), .Z(n1660) );
  CKND0BWP12T U2146 ( .I(n1662), .ZN(n1663) );
  AOI22D0BWP12T U2147 ( .A1(n1663), .A2(n1779), .B1(n1836), .B2(
        DEC_RF_memory_store_data_reg[0]), .ZN(n1667) );
  CKND2D1BWP12T U2148 ( .A1(n1784), .A2(n1664), .ZN(n1665) );
  ND4D1BWP12T U2149 ( .A1(n1668), .A2(n1667), .A3(n1666), .A4(n1665), .ZN(n830) );
  TPND2D0BWP12T U2150 ( .A1(n1715), .A2(IF_DEC_instruction[3]), .ZN(n1677) );
  AOI22D0BWP12T U2151 ( .A1(n1735), .A2(n1675), .B1(n1703), .B2(n1795), .ZN(
        n1676) );
  OAI211D1BWP12T U2152 ( .A1(n1709), .A2(n1713), .B(n1677), .C(n1676), .ZN(
        n1678) );
  TPAOI21D0BWP12T U2153 ( .A1(IF_DEC_instruction[4]), .A2(n1679), .B(n1678), 
        .ZN(n1681) );
  CKND2D1BWP12T U2154 ( .A1(n1836), .A2(DEC_RF_offset_b[5]), .ZN(n1680) );
  OAI21D1BWP12T U2155 ( .A1(n1681), .A2(n1832), .B(n1680), .ZN(n804) );
  MOAI22D0BWP12T U2156 ( .A1(n1684), .A2(n1683), .B1(n1682), .B2(
        IF_DEC_instruction[0]), .ZN(n1686) );
  INR3XD0BWP12T U2157 ( .A1(n1687), .B1(n1686), .B2(n1685), .ZN(n1688) );
  INVD1BWP12T U2158 ( .I(n1688), .ZN(n1689) );
  CKND2D1BWP12T U2159 ( .A1(n1693), .A2(n1692), .ZN(n1707) );
  AOI21D0BWP12T U2160 ( .A1(n1836), .A2(DEC_RF_operand_a[0]), .B(n1707), .ZN(
        n1694) );
  OAI21D1BWP12T U2161 ( .A1(n1695), .A2(n1757), .B(n1694), .ZN(n811) );
  TPNR2D0BWP12T U2162 ( .A1(n1710), .A2(n1783), .ZN(n1701) );
  TPND2D0BWP12T U2163 ( .A1(n1735), .A2(n1714), .ZN(n1698) );
  TPOAI31D0BWP12T U2164 ( .A1(n1822), .A2(n1699), .A3(n1825), .B(n1698), .ZN(
        n1700) );
  RCAOI211D0BWP12T U2165 ( .A1(n1718), .A2(IF_DEC_instruction[3]), .B(n1701), 
        .C(n1700), .ZN(n1702) );
  OAI21D1BWP12T U2166 ( .A1(n1720), .A2(n1788), .B(n1702), .ZN(n1704) );
  AO222D1BWP12T U2167 ( .A1(n1704), .A2(n1809), .B1(n1703), .B2(n1723), .C1(
        n1836), .C2(DEC_RF_offset_b[3]), .Z(n806) );
  AOI22D0BWP12T U2168 ( .A1(n1753), .A2(IF_DEC_instruction[0]), .B1(n1714), 
        .B2(n1748), .ZN(n1705) );
  TPAOI31D0BWP12T U2169 ( .A1(n1720), .A2(n1706), .A3(n1705), .B(n1757), .ZN(
        n1708) );
  AO211D1BWP12T U2170 ( .A1(n1836), .A2(DEC_RF_alu_write_to_reg[0]), .B(n1708), 
        .C(n1707), .Z(n816) );
  AO222D1BWP12T U2171 ( .A1(n1711), .A2(n1809), .B1(n1718), .B2(n1723), .C1(
        n1836), .C2(DEC_RF_offset_b[7]), .Z(n802) );
  CKND0BWP12T U2172 ( .I(n1735), .ZN(n1716) );
  TPOAI21D0BWP12T U2173 ( .A1(n1716), .A2(n1823), .B(n1778), .ZN(n1717) );
  AOI211D0BWP12T U2174 ( .A1(n1718), .A2(IF_DEC_instruction[1]), .B(n1817), 
        .C(n1717), .ZN(n1719) );
  OAI211D1BWP12T U2175 ( .A1(n1721), .A2(n1720), .B(n1719), .C(n1813), .ZN(
        n1724) );
  AO222D1BWP12T U2176 ( .A1(n1724), .A2(n1809), .B1(n1723), .B2(n1722), .C1(
        n1836), .C2(DEC_RF_offset_b[1]), .Z(n808) );
  OAI21D1BWP12T U2177 ( .A1(n1725), .A2(n1730), .B(n1833), .ZN(
        MEMCTRL_RF_IF_data_in[28]) );
  OAI21D1BWP12T U2178 ( .A1(n1726), .A2(n1730), .B(n1833), .ZN(
        MEMCTRL_RF_IF_data_in[29]) );
  OAI21D1BWP12T U2179 ( .A1(n1727), .A2(n1730), .B(n1833), .ZN(
        MEMCTRL_RF_IF_data_in[31]) );
  OAI21D1BWP12T U2180 ( .A1(n1728), .A2(n1730), .B(n1833), .ZN(
        MEMCTRL_RF_IF_data_in[30]) );
  INVD1BWP12T U2181 ( .I(MEM_MEMCTRL_from_mem_data[15]), .ZN(n1729) );
  OAI21D1BWP12T U2182 ( .A1(n1730), .A2(n1729), .B(n1833), .ZN(
        MEMCTRL_RF_IF_data_in[23]) );
  NR2D1BWP12T U2183 ( .A1(n1731), .A2(reset), .ZN(n1732) );
  CKND0BWP12T U2184 ( .I(MEMCTRL_RF_IF_data_in[14]), .ZN(n1734) );
  MOAI22D0BWP12T U2185 ( .A1(n1734), .A2(n1733), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_14_), .B2(n1732), .ZN(
        Instruction_Fetch_inst1_N97) );
  AOI21D0BWP12T U2186 ( .A1(n1737), .A2(n1736), .B(n1735), .ZN(n1738) );
  MOAI22D0BWP12T U2187 ( .A1(n1738), .A2(n1832), .B1(n1836), .B2(
        DEC_MEMCTRL_load_store_width[0]), .ZN(n838) );
  CKND0BWP12T U2188 ( .I(n1739), .ZN(n1741) );
  ND4D0BWP12T U2189 ( .A1(n1742), .A2(n1741), .A3(n1740), .A4(n1778), .ZN(
        n1746) );
  NR4D0BWP12T U2190 ( .A1(n1746), .A2(n1745), .A3(n1744), .A4(n1743), .ZN(
        n1747) );
  MOAI22D0BWP12T U2191 ( .A1(n1747), .A2(n1832), .B1(n1836), .B2(
        DEC_IF_stall_to_instructionfetch), .ZN(n845) );
  CKND0BWP12T U2192 ( .I(n1748), .ZN(n1750) );
  OAI21D0BWP12T U2193 ( .A1(n1750), .A2(n1822), .B(n1749), .ZN(n1752) );
  RCAOI211D0BWP12T U2194 ( .A1(IF_DEC_instruction[1]), .A2(n1753), .B(n1752), 
        .C(n1751), .ZN(n1754) );
  MOAI22D0BWP12T U2195 ( .A1(n1754), .A2(n1832), .B1(n1836), .B2(
        DEC_RF_alu_write_to_reg[1]), .ZN(n819) );
  IOA21D1BWP12T U2196 ( .A1(n1836), .A2(n869), .B(n1755), .ZN(n840) );
  IOA21D1BWP12T U2197 ( .A1(n1836), .A2(DEC_RF_memory_store_address_reg[3]), 
        .B(n1756), .ZN(n832) );
  TPAOI31D0BWP12T U2198 ( .A1(n1760), .A2(n1759), .A3(n1758), .B(n1757), .ZN(
        n1762) );
  NR2D1BWP12T U2199 ( .A1(n1762), .A2(n1761), .ZN(n1835) );
  CKND0BWP12T U2200 ( .I(n1763), .ZN(n1764) );
  OAI21D0BWP12T U2201 ( .A1(n1822), .A2(n1824), .B(n1764), .ZN(n1765) );
  AOI22D0BWP12T U2202 ( .A1(n1765), .A2(n1790), .B1(n1836), .B2(
        DEC_ALU_alu_opcode[3]), .ZN(n1766) );
  IND3D1BWP12T U2203 ( .A1(n1767), .B1(n1835), .B2(n1766), .ZN(n849) );
  CKND0BWP12T U2204 ( .I(n1768), .ZN(n1782) );
  CKND0BWP12T U2205 ( .I(n1769), .ZN(n1770) );
  OAI31D0BWP12T U2206 ( .A1(n1772), .A2(n1771), .A3(n1770), .B(n1817), .ZN(
        n1781) );
  MAOI22D0BWP12T U2207 ( .A1(n1779), .A2(n1795), .B1(n1803), .B2(n1778), .ZN(
        n1780) );
  OAI211D1BWP12T U2208 ( .A1(n1783), .A2(n1782), .B(n1781), .C(n1780), .ZN(
        n1796) );
  AOI22D0BWP12T U2209 ( .A1(n1796), .A2(n1830), .B1(n1784), .B2(
        IF_DEC_instruction[1]), .ZN(n1785) );
  MOAI22D0BWP12T U2210 ( .A1(n1785), .A2(n1832), .B1(n1836), .B2(
        DEC_RF_memory_store_data_reg[1]), .ZN(n829) );
  AOI222D0BWP12T U2211 ( .A1(n1796), .A2(n1821), .B1(n1795), .B2(n1794), .C1(
        IF_DEC_instruction[1]), .C2(n1793), .ZN(n1797) );
  MOAI22D0BWP12T U2212 ( .A1(n1797), .A2(n1832), .B1(n1836), .B2(
        DEC_RF_memory_write_to_reg[1]), .ZN(n823) );
  IND4D0BWP12T U2213 ( .A1(n1801), .B1(n1800), .B2(n1799), .B3(n1798), .ZN(
        n1805) );
  IND4D0BWP12T U2214 ( .A1(n1805), .B1(n1804), .B2(n1803), .B3(n1802), .ZN(
        n1806) );
  CKND2D0BWP12T U2215 ( .A1(n1806), .A2(n1814), .ZN(n1807) );
  TPAOI31D0BWP12T U2216 ( .A1(n1829), .A2(n1808), .A3(n1807), .B(n1830), .ZN(
        n1811) );
  OAI21D1BWP12T U2217 ( .A1(n1811), .A2(n1810), .B(n1809), .ZN(n1812) );
  IOA21D1BWP12T U2218 ( .A1(n1836), .A2(DEC_MEMCTRL_memory_load_request), .B(
        n1812), .ZN(n861) );
  IOA21D1BWP12T U2219 ( .A1(n1836), .A2(DEC_RF_memory_write_to_reg_enable), 
        .B(n1812), .ZN(n825) );
  IOA21D0BWP12T U2220 ( .A1(n1815), .A2(n1814), .B(n1813), .ZN(n1816) );
  AOI21D0BWP12T U2221 ( .A1(n1818), .A2(n1817), .B(n1816), .ZN(n1819) );
  MOAI22D0BWP12T U2222 ( .A1(n1819), .A2(n1832), .B1(n1836), .B2(
        irdecode_inst1_split_instruction), .ZN(n847) );
  IOA21D1BWP12T U2223 ( .A1(n1834), .A2(MEM_MEMCTRL_from_mem_data[1]), .B(
        n1833), .ZN(MEMCTRL_RF_IF_data_in[25]) );
  IOA21D1BWP12T U2224 ( .A1(n1834), .A2(MEM_MEMCTRL_from_mem_data[14]), .B(
        n1833), .ZN(MEMCTRL_RF_IF_data_in[22]) );
  IOA21D1BWP12T U2225 ( .A1(n1834), .A2(MEM_MEMCTRL_from_mem_data[13]), .B(
        n1833), .ZN(MEMCTRL_RF_IF_data_in[21]) );
  IOA21D1BWP12T U2226 ( .A1(n1834), .A2(MEM_MEMCTRL_from_mem_data[11]), .B(
        n1833), .ZN(MEMCTRL_RF_IF_data_in[19]) );
  IOA21D1BWP12T U2227 ( .A1(n1834), .A2(MEM_MEMCTRL_from_mem_data[8]), .B(
        n1833), .ZN(MEMCTRL_RF_IF_data_in[16]) );
  IOA21D1BWP12T U2228 ( .A1(n1834), .A2(MEM_MEMCTRL_from_mem_data[9]), .B(
        n1833), .ZN(MEMCTRL_RF_IF_data_in[17]) );
  IOA21D1BWP12T U2229 ( .A1(n1834), .A2(MEM_MEMCTRL_from_mem_data[10]), .B(
        n1833), .ZN(MEMCTRL_RF_IF_data_in[18]) );
  IOA21D1BWP12T U2230 ( .A1(n1834), .A2(MEM_MEMCTRL_from_mem_data[12]), .B(
        n1833), .ZN(MEMCTRL_RF_IF_data_in[20]) );
endmodule

