
module irdecode ( clk, reset, instruction, instruction_valid, flag_n, flag_z, 
        flag_c, flag_v, memory_write_finished, memory_read_finished, operand_a, 
        operand_b, offset_a, offset_b, alu_opcode, pc_mask_bit, update_flag_n, 
        update_flag_z, update_flag_c, update_flag_v, alu_write_to_reg, 
        alu_write_to_reg_enable, memory_write_to_reg, 
        memory_write_to_reg_enable, memory_store_data_reg, 
        memory_store_address_reg, memory_address_source_is_reg, 
        load_store_width, memorycontroller_sign_extend, memory_load_request, 
        stall_to_instructionfetch, memory_store_request_BAR );
  input [15:0] instruction;
  output [4:0] operand_a;
  output [4:0] operand_b;
  output [31:0] offset_a;
  output [31:0] offset_b;
  output [4:0] alu_opcode;
  output [4:0] alu_write_to_reg;
  output [4:0] memory_write_to_reg;
  output [4:0] memory_store_data_reg;
  output [4:0] memory_store_address_reg;
  output [1:0] load_store_width;
  input clk, reset, instruction_valid, flag_n, flag_z, flag_c, flag_v,
         memory_write_finished, memory_read_finished;
  output pc_mask_bit, update_flag_n, update_flag_z, update_flag_c,
         update_flag_v, alu_write_to_reg_enable, memory_write_to_reg_enable,
         memory_address_source_is_reg, memorycontroller_sign_extend,
         memory_load_request, stall_to_instructionfetch,
         memory_store_request_BAR;
  wire   memory_store_request, next_update_flag_n, next_update_flag_c,
         next_update_flag_v, next_alu_write_to_reg_enable, split_instruction,
         N539, N540, N541, N542, N543, N544, N545, N546, N701, N702, N703,
         N704, N705, N706, N707, N906, N907, N910, N911, N912, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n2, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512;
  wire   [7:0] itstate;
  wire   [7:0] step;
  wire   [7:0] next_step;
  tri   clk;
  tri   reset;
  tri   flag_n;
  tri   flag_z;
  tri   flag_c;
  tri   flag_v;
  tri   [4:0] operand_a;
  tri   [4:0] operand_b;
  tri   [31:0] offset_b;
  tri   [4:0] alu_write_to_reg;
  tri   alu_write_to_reg_enable;
  tri   [4:0] memory_write_to_reg;
  tri   memory_write_to_reg_enable;
  tri   [4:0] memory_store_data_reg;
  tri   [4:0] memory_store_address_reg;
  tri   [31:0] offset_a;

  OR2XD4BWP12T C2484 ( .A1(next_step[1]), .A2(N910), .Z(N912) );
  CKAN2D2BWP12T C2482 ( .A1(N907), .A2(N910), .Z(N911) );
  CKAN2D2BWP12T C2476 ( .A1(next_step[1]), .A2(next_step[0]), .Z(N906) );
  CKAN2D2BWP12T C5286 ( .A1(next_step[0]), .A2(instruction[0]), .Z(N707) );
  CKAN2D2BWP12T C5285 ( .A1(next_step[1]), .A2(instruction[1]), .Z(N706) );
  CKAN2D2BWP12T C5284 ( .A1(next_step[2]), .A2(instruction[2]), .Z(N705) );
  CKAN2D2BWP12T C5283 ( .A1(next_step[3]), .A2(instruction[3]), .Z(N704) );
  CKAN2D2BWP12T C5282 ( .A1(next_step[4]), .A2(instruction[4]), .Z(N703) );
  CKAN2D2BWP12T C5281 ( .A1(next_step[5]), .A2(instruction[5]), .Z(N702) );
  CKAN2D2BWP12T C5280 ( .A1(next_step[6]), .A2(instruction[6]), .Z(N701) );
  CKAN2D2BWP12T C5200 ( .A1(next_step[0]), .A2(instruction[0]), .Z(N546) );
  CKAN2D2BWP12T C5199 ( .A1(next_step[1]), .A2(instruction[1]), .Z(N545) );
  CKAN2D2BWP12T C5198 ( .A1(next_step[2]), .A2(instruction[2]), .Z(N544) );
  CKAN2D2BWP12T C5197 ( .A1(next_step[3]), .A2(instruction[3]), .Z(N543) );
  CKAN2D2BWP12T C5196 ( .A1(next_step[4]), .A2(instruction[4]), .Z(N542) );
  CKAN2D2BWP12T C5195 ( .A1(next_step[5]), .A2(instruction[5]), .Z(N541) );
  CKAN2D2BWP12T C5194 ( .A1(next_step[6]), .A2(instruction[6]), .Z(N540) );
  CKAN2D2BWP12T C5193 ( .A1(next_step[7]), .A2(instruction[7]), .Z(N539) );
  DFQD1BWP12T split_instruction_reg ( .D(n693), .CP(clk), .Q(split_instruction) );
  DFQD1BWP12T itstate_reg_0_ ( .D(n691), .CP(clk), .Q(itstate[0]) );
  DFQD1BWP12T itstate_reg_1_ ( .D(n690), .CP(clk), .Q(itstate[1]) );
  DFQD1BWP12T itstate_reg_2_ ( .D(n689), .CP(clk), .Q(itstate[2]) );
  DFQD1BWP12T itstate_reg_3_ ( .D(n688), .CP(clk), .Q(itstate[3]) );
  DFQD1BWP12T itstate_reg_4_ ( .D(n687), .CP(clk), .Q(itstate[4]) );
  DFQD1BWP12T itstate_reg_5_ ( .D(n686), .CP(clk), .Q(itstate[5]) );
  DFQD1BWP12T itstate_reg_6_ ( .D(n685), .CP(clk), .Q(itstate[6]) );
  DFQD1BWP12T itstate_reg_7_ ( .D(n684), .CP(clk), .Q(itstate[7]) );
  DFQD1BWP12T update_flag_v_reg ( .D(next_update_flag_v), .CP(clk), .Q(
        update_flag_v) );
  DFQD1BWP12T update_flag_c_reg ( .D(next_update_flag_c), .CP(clk), .Q(
        update_flag_c) );
  DFQD1BWP12T alu_write_to_reg_enable_reg ( .D(next_alu_write_to_reg_enable), 
        .CP(clk), .Q(alu_write_to_reg_enable) );
  DFQD1BWP12T update_flag_n_reg ( .D(next_update_flag_n), .CP(clk), .Q(
        update_flag_n) );
  DFQD1BWP12T update_flag_z_reg ( .D(next_update_flag_n), .CP(clk), .Q(
        update_flag_z) );
  DFQD1BWP12T memory_store_request_reg ( .D(n665), .CP(clk), .Q(
        memory_store_request) );
  DFQD1BWP12T alu_write_to_reg_reg_3_ ( .D(n642), .CP(clk), .Q(
        alu_write_to_reg[3]) );
  DFQD1BWP12T operand_b_reg_0_ ( .D(n633), .CP(clk), .Q(operand_b[0]) );
  DFQD1BWP12T operand_b_reg_2_ ( .D(n631), .CP(clk), .Q(operand_b[2]) );
  DFQD1BWP12T operand_b_reg_4_ ( .D(n629), .CP(clk), .Q(operand_b[4]) );
  DFQD1BWP12T stall_to_instructionfetch_reg ( .D(n692), .CP(clk), .Q(
        stall_to_instructionfetch) );
  DFQD1BWP12T alu_opcode_reg_2_ ( .D(n668), .CP(clk), .Q(alu_opcode[2]) );
  DFQD1BWP12T load_store_width_reg_1_ ( .D(n662), .CP(clk), .Q(
        load_store_width[1]) );
  DFQD1BWP12T memory_store_address_reg_reg_0_ ( .D(n660), .CP(clk), .Q(
        memory_store_address_reg[0]) );
  DFQD1BWP12T memory_store_address_reg_reg_2_ ( .D(n658), .CP(clk), .Q(
        memory_store_address_reg[2]) );
  DFQD1BWP12T memory_store_address_reg_reg_3_ ( .D(n657), .CP(clk), .Q(
        memory_store_address_reg[3]) );
  DFQD1BWP12T memory_store_address_reg_reg_4_ ( .D(n656), .CP(clk), .Q(
        memory_store_address_reg[4]) );
  DFQD1BWP12T step_reg_6_ ( .D(next_step[6]), .CP(clk), .Q(step[6]) );
  DFQD1BWP12T step_reg_1_ ( .D(next_step[1]), .CP(clk), .Q(step[1]) );
  DFQD1BWP12T step_reg_0_ ( .D(next_step[0]), .CP(clk), .Q(step[0]) );
  DFQD1BWP12T step_reg_7_ ( .D(next_step[7]), .CP(clk), .Q(step[7]) );
  DFQD1BWP12T step_reg_2_ ( .D(next_step[2]), .CP(clk), .Q(step[2]) );
  DFQD1BWP12T step_reg_3_ ( .D(next_step[3]), .CP(clk), .Q(step[3]) );
  DFQD1BWP12T step_reg_4_ ( .D(next_step[4]), .CP(clk), .Q(step[4]) );
  DFQD1BWP12T step_reg_5_ ( .D(next_step[5]), .CP(clk), .Q(step[5]) );
  DFQD1BWP12T memory_store_data_reg_reg_0_ ( .D(n655), .CP(clk), .Q(
        memory_store_data_reg[0]) );
  DFQD1BWP12T memory_write_to_reg_reg_0_ ( .D(n649), .CP(clk), .Q(
        memory_write_to_reg[0]) );
  DFQD1BWP12T memory_store_data_reg_reg_2_ ( .D(n653), .CP(clk), .Q(
        memory_store_data_reg[2]) );
  DFQD1BWP12T memory_write_to_reg_reg_2_ ( .D(n647), .CP(clk), .Q(
        memory_write_to_reg[2]) );
  DFQD1BWP12T offset_b_reg_8_ ( .D(n679), .CP(clk), .Q(offset_b[8]) );
  DFQD1BWP12T offset_b_reg_7_ ( .D(n678), .CP(clk), .Q(offset_b[7]) );
  DFQD1BWP12T offset_b_reg_6_ ( .D(n677), .CP(clk), .Q(offset_b[6]) );
  DFQD1BWP12T offset_b_reg_5_ ( .D(n676), .CP(clk), .Q(offset_b[5]) );
  DFQD1BWP12T offset_b_reg_4_ ( .D(n675), .CP(clk), .Q(offset_b[4]) );
  DFQD1BWP12T offset_b_reg_3_ ( .D(n674), .CP(clk), .Q(offset_b[3]) );
  DFQD1BWP12T offset_b_reg_2_ ( .D(n673), .CP(clk), .Q(offset_b[2]) );
  DFQD1BWP12T offset_b_reg_1_ ( .D(n672), .CP(clk), .Q(offset_b[1]) );
  DFQD1BWP12T offset_b_reg_0_ ( .D(n671), .CP(clk), .Q(offset_b[0]) );
  DFQD1BWP12T alu_opcode_reg_3_ ( .D(n669), .CP(clk), .Q(alu_opcode[3]) );
  DFQD1BWP12T memory_store_data_reg_reg_3_ ( .D(n652), .CP(clk), .Q(
        memory_store_data_reg[3]) );
  DFQD1BWP12T memory_write_to_reg_reg_3_ ( .D(n646), .CP(clk), .Q(
        memory_write_to_reg[3]) );
  DFQD1BWP12T alu_opcode_reg_4_ ( .D(n670), .CP(clk), .Q(alu_opcode[4]) );
  DFQD1BWP12T memory_store_data_reg_reg_4_ ( .D(n651), .CP(clk), .Q(
        memory_store_data_reg[4]) );
  DFQD1BWP12T alu_opcode_reg_0_ ( .D(n666), .CP(clk), .Q(alu_opcode[0]) );
  DFQD1BWP12T memory_load_request_reg ( .D(n683), .CP(clk), .Q(
        memory_load_request) );
  DFQD1BWP12T alu_opcode_reg_1_ ( .D(n667), .CP(clk), .Q(alu_opcode[1]) );
  DFQD1BWP12T memory_write_to_reg_reg_4_ ( .D(n645), .CP(clk), .Q(
        memory_write_to_reg[4]) );
  DFQD1BWP12T alu_write_to_reg_reg_2_ ( .D(n643), .CP(clk), .Q(
        alu_write_to_reg[2]) );
  DFQD1BWP12T alu_write_to_reg_reg_0_ ( .D(n641), .CP(clk), .Q(
        alu_write_to_reg[0]) );
  DFQD1BWP12T alu_write_to_reg_reg_4_ ( .D(n640), .CP(clk), .Q(
        alu_write_to_reg[4]) );
  DFQD1BWP12T operand_a_reg_2_ ( .D(n637), .CP(clk), .Q(operand_a[2]) );
  DFQD1BWP12T operand_a_reg_3_ ( .D(n636), .CP(clk), .Q(operand_a[3]) );
  DFQD1BWP12T operand_a_reg_0_ ( .D(n635), .CP(clk), .Q(operand_a[0]) );
  DFQD1BWP12T operand_a_reg_4_ ( .D(n634), .CP(clk), .Q(operand_a[4]) );
  DFQD1BWP12T operand_b_reg_3_ ( .D(n630), .CP(clk), .Q(operand_b[3]) );
  DFQD1BWP12T memorycontroller_sign_extend_reg ( .D(n664), .CP(clk), .Q(
        memorycontroller_sign_extend) );
  DFQD1BWP12T load_store_width_reg_0_ ( .D(n663), .CP(clk), .Q(
        load_store_width[0]) );
  DFQD1BWP12T memory_address_source_is_reg_reg ( .D(n661), .CP(clk), .Q(
        memory_address_source_is_reg) );
  DFQD1BWP12T memory_store_address_reg_reg_1_ ( .D(n659), .CP(clk), .Q(
        memory_store_address_reg[1]) );
  DFQD1BWP12T memory_store_data_reg_reg_1_ ( .D(n654), .CP(clk), .Q(
        memory_store_data_reg[1]) );
  DFQD1BWP12T memory_write_to_reg_enable_reg ( .D(n650), .CP(clk), .Q(
        memory_write_to_reg_enable) );
  DFQD1BWP12T memory_write_to_reg_reg_1_ ( .D(n648), .CP(clk), .Q(
        memory_write_to_reg[1]) );
  DFQD1BWP12T alu_write_to_reg_reg_1_ ( .D(n644), .CP(clk), .Q(
        alu_write_to_reg[1]) );
  DFQD1BWP12T operand_a_reg_1_ ( .D(n638), .CP(clk), .Q(operand_a[1]) );
  DFQD1BWP12T operand_b_reg_1_ ( .D(n632), .CP(clk), .Q(operand_b[1]) );
  DFQD1BWP12T offset_b_reg_11_ ( .D(n682), .CP(clk), .Q(offset_b[11]) );
  DFQD1BWP12T offset_b_reg_10_ ( .D(n681), .CP(clk), .Q(offset_b[10]) );
  DFQD1BWP12T offset_b_reg_9_ ( .D(n680), .CP(clk), .Q(offset_b[9]) );
  DFQD1BWP12T offset_b_reg_12_ ( .D(n628), .CP(clk), .Q(offset_b[12]) );
  DFQD1BWP12T offset_b_reg_13_ ( .D(n627), .CP(clk), .Q(offset_b[13]) );
  DFQD1BWP12T offset_b_reg_14_ ( .D(n626), .CP(clk), .Q(offset_b[14]) );
  DFQD1BWP12T offset_b_reg_15_ ( .D(n625), .CP(clk), .Q(offset_b[15]) );
  DFQD1BWP12T offset_b_reg_16_ ( .D(n624), .CP(clk), .Q(offset_b[16]) );
  DFQD1BWP12T offset_b_reg_17_ ( .D(n623), .CP(clk), .Q(offset_b[17]) );
  DFQD1BWP12T offset_b_reg_18_ ( .D(n622), .CP(clk), .Q(offset_b[18]) );
  DFQD1BWP12T offset_b_reg_19_ ( .D(n621), .CP(clk), .Q(offset_b[19]) );
  DFQD1BWP12T offset_b_reg_20_ ( .D(n620), .CP(clk), .Q(offset_b[20]) );
  DFQD1BWP12T offset_b_reg_21_ ( .D(n619), .CP(clk), .Q(offset_b[21]) );
  DFQD1BWP12T offset_b_reg_22_ ( .D(n618), .CP(clk), .Q(offset_b[22]) );
  DFQD1BWP12T offset_b_reg_23_ ( .D(n617), .CP(clk), .Q(offset_b[23]) );
  DFQD1BWP12T offset_b_reg_24_ ( .D(n616), .CP(clk), .Q(offset_b[24]) );
  DFQD1BWP12T offset_b_reg_25_ ( .D(n615), .CP(clk), .Q(offset_b[25]) );
  DFQD1BWP12T offset_b_reg_26_ ( .D(n614), .CP(clk), .Q(offset_b[26]) );
  DFQD1BWP12T offset_b_reg_27_ ( .D(n613), .CP(clk), .Q(offset_b[27]) );
  DFQD1BWP12T offset_b_reg_28_ ( .D(n612), .CP(clk), .Q(offset_b[28]) );
  DFQD1BWP12T offset_b_reg_29_ ( .D(n611), .CP(clk), .Q(offset_b[29]) );
  DFQD1BWP12T offset_b_reg_30_ ( .D(n610), .CP(clk), .Q(offset_b[30]) );
  DFQD1BWP12T offset_b_reg_31_ ( .D(n609), .CP(clk), .Q(offset_b[31]) );
  TIEHBWP12T U3 ( .Z(n2) );
  INVD1BWP12T U4 ( .I(n2), .ZN(offset_a[0]) );
  INVD1BWP12T U5 ( .I(n2), .ZN(offset_a[1]) );
  INVD1BWP12T U6 ( .I(n2), .ZN(offset_a[2]) );
  INVD1BWP12T U7 ( .I(n2), .ZN(offset_a[3]) );
  INVD1BWP12T U8 ( .I(n2), .ZN(offset_a[4]) );
  INVD1BWP12T U9 ( .I(n2), .ZN(offset_a[5]) );
  INVD1BWP12T U10 ( .I(n2), .ZN(offset_a[6]) );
  INVD1BWP12T U11 ( .I(n2), .ZN(offset_a[7]) );
  INVD1BWP12T U12 ( .I(n2), .ZN(offset_a[8]) );
  INVD1BWP12T U13 ( .I(n2), .ZN(offset_a[9]) );
  INVD1BWP12T U14 ( .I(n2), .ZN(offset_a[10]) );
  INVD1BWP12T U15 ( .I(n2), .ZN(offset_a[11]) );
  INVD1BWP12T U16 ( .I(n2), .ZN(offset_a[12]) );
  INVD1BWP12T U17 ( .I(n2), .ZN(offset_a[13]) );
  INVD1BWP12T U18 ( .I(n2), .ZN(offset_a[14]) );
  INVD1BWP12T U19 ( .I(n2), .ZN(offset_a[15]) );
  INVD1BWP12T U20 ( .I(n2), .ZN(offset_a[16]) );
  INVD1BWP12T U21 ( .I(n2), .ZN(offset_a[17]) );
  INVD1BWP12T U22 ( .I(n2), .ZN(offset_a[18]) );
  INVD1BWP12T U23 ( .I(n2), .ZN(offset_a[19]) );
  INVD1BWP12T U24 ( .I(n2), .ZN(offset_a[20]) );
  INVD1BWP12T U25 ( .I(n2), .ZN(offset_a[21]) );
  INVD1BWP12T U26 ( .I(n2), .ZN(offset_a[22]) );
  INVD1BWP12T U27 ( .I(n2), .ZN(offset_a[23]) );
  INVD1BWP12T U28 ( .I(n2), .ZN(offset_a[24]) );
  INVD1BWP12T U29 ( .I(n2), .ZN(offset_a[25]) );
  INVD1BWP12T U30 ( .I(n2), .ZN(offset_a[26]) );
  INVD1BWP12T U31 ( .I(n2), .ZN(offset_a[27]) );
  INVD1BWP12T U32 ( .I(n2), .ZN(offset_a[28]) );
  INVD1BWP12T U33 ( .I(n2), .ZN(offset_a[29]) );
  INVD1BWP12T U34 ( .I(n2), .ZN(offset_a[30]) );
  INVD1BWP12T U35 ( .I(n2), .ZN(offset_a[31]) );
  NR2D1BWP12T U36 ( .A1(instruction[8]), .A2(N539), .ZN(n85) );
  INR2D1BWP12T U37 ( .A1(n151), .B1(N704), .ZN(n77) );
  INR2D1BWP12T U38 ( .A1(instruction[15]), .B1(instruction[13]), .ZN(n100) );
  NR2D1BWP12T U39 ( .A1(n74), .A2(n149), .ZN(n166) );
  NR2D1BWP12T U40 ( .A1(instruction[12]), .A2(instruction[11]), .ZN(n502) );
  INVD1BWP12T U41 ( .I(instruction[12]), .ZN(n451) );
  NR2D1BWP12T U42 ( .A1(n356), .A2(N544), .ZN(n80) );
  ND2D1BWP12T U43 ( .A1(n85), .A2(n79), .ZN(n81) );
  ND2D1BWP12T U44 ( .A1(n78), .A2(n447), .ZN(n74) );
  NR4D0BWP12T U45 ( .A1(N705), .A2(N701), .A3(N702), .A4(N703), .ZN(n78) );
  ND2D1BWP12T U46 ( .A1(n80), .A2(N543), .ZN(n177) );
  INVD1BWP12T U47 ( .I(N544), .ZN(n139) );
  INR3D0BWP12T U48 ( .A1(n80), .B1(N543), .B2(N542), .ZN(n84) );
  NR2D1BWP12T U49 ( .A1(N701), .A2(n163), .ZN(n75) );
  ND2D1BWP12T U50 ( .A1(N541), .A2(n84), .ZN(n138) );
  IND2D1BWP12T U51 ( .A1(N705), .B1(n77), .ZN(n70) );
  INVD1BWP12T U52 ( .I(n148), .ZN(n150) );
  ND2D1BWP12T U53 ( .A1(n83), .A2(n139), .ZN(n89) );
  NR2D1BWP12T U54 ( .A1(n89), .A2(n141), .ZN(n174) );
  NR2D1BWP12T U55 ( .A1(n74), .A2(n153), .ZN(n219) );
  NR2D1BWP12T U56 ( .A1(n461), .A2(n493), .ZN(n110) );
  ND2D1BWP12T U57 ( .A1(n79), .A2(n84), .ZN(n90) );
  INVD1BWP12T U58 ( .I(n498), .ZN(n229) );
  NR3D1BWP12T U59 ( .A1(next_step[0]), .A2(N907), .A3(n308), .ZN(n403) );
  INR4D0BWP12T U60 ( .A1(N701), .B1(N703), .B2(N702), .B3(n70), .ZN(n205) );
  NR2D1BWP12T U61 ( .A1(n465), .A2(n376), .ZN(n200) );
  NR2D1BWP12T U62 ( .A1(n81), .A2(n137), .ZN(n202) );
  INVD1BWP12T U63 ( .I(n177), .ZN(n182) );
  NR2D1BWP12T U64 ( .A1(n256), .A2(n259), .ZN(n241) );
  AOI31D1BWP12T U65 ( .A1(n77), .A2(N705), .A3(n71), .B(n166), .ZN(n154) );
  INVD1BWP12T U66 ( .I(n205), .ZN(n152) );
  INVD1BWP12T U67 ( .I(flag_z), .ZN(n56) );
  ND2D1BWP12T U68 ( .A1(flag_c), .A2(n56), .ZN(n58) );
  INVD1BWP12T U69 ( .I(n502), .ZN(n94) );
  INVD1BWP12T U70 ( .I(n303), .ZN(n169) );
  NR2D1BWP12T U71 ( .A1(itstate[6]), .A2(itstate[7]), .ZN(n57) );
  INVD1BWP12T U72 ( .I(itstate[4]), .ZN(n65) );
  ND2D1BWP12T U73 ( .A1(n100), .A2(instruction[14]), .ZN(n93) );
  NR3D1BWP12T U74 ( .A1(n483), .A2(n96), .A3(instruction[9]), .ZN(n462) );
  ND2D1BWP12T U75 ( .A1(n88), .A2(n142), .ZN(n141) );
  ND2D1BWP12T U76 ( .A1(n73), .A2(n150), .ZN(n153) );
  INVD1BWP12T U77 ( .I(n70), .ZN(n73) );
  NR2D1BWP12T U78 ( .A1(n137), .A2(n141), .ZN(n376) );
  INVD1BWP12T U79 ( .I(n174), .ZN(n222) );
  INVD1BWP12T U80 ( .I(n465), .ZN(n173) );
  INR2D1BWP12T U81 ( .A1(N912), .B1(N906), .ZN(n105) );
  OAI22D1BWP12T U82 ( .A1(memory_read_finished), .A2(n157), .B1(
        memory_write_finished), .B2(memory_store_request_BAR), .ZN(n68) );
  NR3D1BWP12T U83 ( .A1(n219), .A2(n190), .A3(n204), .ZN(n358) );
  INVD1BWP12T U84 ( .I(n341), .ZN(n322) );
  ND2D1BWP12T U85 ( .A1(n110), .A2(n490), .ZN(n405) );
  ND2D1BWP12T U86 ( .A1(n312), .A2(n506), .ZN(n511) );
  INVD1BWP12T U87 ( .I(n128), .ZN(n491) );
  NR2D1BWP12T U88 ( .A1(n312), .A2(n404), .ZN(n498) );
  INVD1BWP12T U89 ( .I(n505), .ZN(n499) );
  INVD1BWP12T U90 ( .I(memory_load_request), .ZN(n157) );
  NR2D1BWP12T U91 ( .A1(n451), .A2(n95), .ZN(n492) );
  AOI31D1BWP12T U92 ( .A1(n142), .A2(n200), .A3(n424), .B(n422), .ZN(n187) );
  NR3D1BWP12T U93 ( .A1(N539), .A2(n407), .A3(n90), .ZN(n465) );
  OAI22D1BWP12T U94 ( .A1(n121), .A2(n419), .B1(n231), .B2(n291), .ZN(n394) );
  OAI21D1BWP12T U95 ( .A1(n222), .A2(n390), .B(n278), .ZN(n235) );
  NR2D1BWP12T U96 ( .A1(n403), .A2(n229), .ZN(n126) );
  NR2D1BWP12T U97 ( .A1(n448), .A2(n405), .ZN(n127) );
  NR2D1BWP12T U98 ( .A1(n478), .A2(n419), .ZN(n501) );
  NR2D1BWP12T U99 ( .A1(n478), .A2(n333), .ZN(n416) );
  INVD1BWP12T U100 ( .I(n126), .ZN(n441) );
  INVD1BWP12T U101 ( .I(n127), .ZN(n442) );
  INVD1BWP12T U102 ( .I(n420), .ZN(n506) );
  NR2D1BWP12T U103 ( .A1(n121), .A2(n98), .ZN(n493) );
  NR2D1BWP12T U104 ( .A1(n303), .A2(n348), .ZN(n473) );
  NR2D1BWP12T U105 ( .A1(n471), .A2(n196), .ZN(n220) );
  NR2D1BWP12T U106 ( .A1(n485), .A2(n422), .ZN(n381) );
  NR2D1BWP12T U107 ( .A1(n381), .A2(n459), .ZN(n249) );
  NR2D1BWP12T U108 ( .A1(n451), .A2(n98), .ZN(n256) );
  ND2D1BWP12T U109 ( .A1(n412), .A2(n411), .ZN(n259) );
  NR2D1BWP12T U110 ( .A1(n94), .A2(n98), .ZN(n505) );
  INVD1BWP12T U111 ( .I(n370), .ZN(n485) );
  INVD1BWP12T U112 ( .I(n486), .ZN(n278) );
  ND2D1BWP12T U113 ( .A1(n154), .A2(n155), .ZN(n190) );
  OAI21D1BWP12T U114 ( .A1(instruction[7]), .A2(n152), .B(n160), .ZN(n204) );
  NR2D1BWP12T U115 ( .A1(n169), .A2(n348), .ZN(n471) );
  INVD1BWP12T U116 ( .I(memory_store_request), .ZN(memory_store_request_BAR)
         );
  INVD1BWP12T U117 ( .I(n285), .ZN(n351) );
  MOAI22D0BWP12T U118 ( .A1(flag_n), .A2(flag_v), .B1(flag_n), .B2(flag_v), 
        .ZN(n299) );
  ND2D1BWP12T U119 ( .A1(n299), .A2(n56), .ZN(n292) );
  INVD1BWP12T U120 ( .I(n292), .ZN(n294) );
  INVD1BWP12T U121 ( .I(n58), .ZN(n298) );
  NR2D1BWP12T U122 ( .A1(n95), .A2(n94), .ZN(n404) );
  NR2D1BWP12T U123 ( .A1(n451), .A2(n93), .ZN(n312) );
  NR3D1BWP12T U124 ( .A1(n96), .A2(n169), .A3(n282), .ZN(n448) );
  INVD1BWP12T U125 ( .I(n492), .ZN(n308) );
  INVD1BWP12T U126 ( .I(n231), .ZN(n432) );
  INVD1BWP12T U127 ( .I(instruction[10]), .ZN(n483) );
  INVD1BWP12T U128 ( .I(instruction[9]), .ZN(n488) );
  INVD1BWP12T U129 ( .I(instruction[11]), .ZN(n470) );
  INVD1BWP12T U130 ( .I(n295), .ZN(n282) );
  NR2D1BWP12T U131 ( .A1(instruction[10]), .A2(n499), .ZN(n449) );
  NR2D1BWP12T U132 ( .A1(instruction[13]), .A2(n143), .ZN(n450) );
  INVD1BWP12T U133 ( .I(instruction[8]), .ZN(n407) );
  ND2D1BWP12T U134 ( .A1(n508), .A2(instruction[7]), .ZN(n420) );
  INVD1BWP12T U135 ( .I(n449), .ZN(n280) );
  NR2D1BWP12T U136 ( .A1(n170), .A2(n485), .ZN(n508) );
  ND2D1BWP12T U137 ( .A1(n350), .A2(n328), .ZN(n335) );
  INVD1BWP12T U138 ( .I(instruction[6]), .ZN(n333) );
  INVD1BWP12T U139 ( .I(itstate[5]), .ZN(n329) );
  NR2D1BWP12T U140 ( .A1(instruction[12]), .A2(n93), .ZN(n428) );
  INVD1BWP12T U141 ( .I(n462), .ZN(n422) );
  INR2D1BWP12T U142 ( .A1(n433), .B1(n105), .ZN(n426) );
  INVD1BWP12T U143 ( .I(n508), .ZN(n478) );
  OR2XD1BWP12T U144 ( .A1(n141), .A2(n140), .Z(n198) );
  ND2D1BWP12T U145 ( .A1(N703), .A2(n73), .ZN(n382) );
  ND3D1BWP12T U146 ( .A1(n142), .A2(n222), .A3(n173), .ZN(n355) );
  INVD1BWP12T U147 ( .I(n88), .ZN(n356) );
  INVD1BWP12T U148 ( .I(N546), .ZN(n178) );
  NR2D1BWP12T U149 ( .A1(n105), .A2(n308), .ZN(n144) );
  INVD1BWP12T U150 ( .I(n379), .ZN(n387) );
  INVD1BWP12T U151 ( .I(n274), .ZN(n512) );
  INVD1BWP12T U152 ( .I(n381), .ZN(n390) );
  OAI22D1BWP12T U153 ( .A1(n337), .A2(n336), .B1(n447), .B2(n335), .ZN(n684)
         );
  OAI22D1BWP12T U154 ( .A1(n337), .A2(n334), .B1(n333), .B2(n335), .ZN(n685)
         );
  MOAI22D0BWP12T U155 ( .A1(n337), .A2(n329), .B1(instruction[5]), .B2(n330), 
        .ZN(n686) );
  INVD1BWP12T U156 ( .I(N910), .ZN(next_step[0]) );
  INVD1BWP12T U157 ( .I(next_step[1]), .ZN(N907) );
  AOI21D1BWP12T U158 ( .A1(n512), .A2(step[0]), .B(n106), .ZN(N910) );
  CKND0BWP12T U159 ( .I(N545), .ZN(n34) );
  AOI221D0BWP12T U160 ( .A1(N546), .A2(N545), .B1(n178), .B2(n34), .C(n89), 
        .ZN(n35) );
  NR4D0BWP12T U161 ( .A1(n175), .A2(n202), .A3(n464), .A4(n35), .ZN(n142) );
  AOI21D1BWP12T U162 ( .A1(n51), .A2(n50), .B(n329), .ZN(n64) );
  NR2D1BWP12T U163 ( .A1(n351), .A2(n66), .ZN(n170) );
  NR3D1BWP12T U164 ( .A1(reset), .A2(n67), .A3(n68), .ZN(n370) );
  CKND0BWP12T U165 ( .I(n159), .ZN(n36) );
  AOI211D0BWP12T U166 ( .A1(N707), .A2(N706), .B(n74), .C(N704), .ZN(n37) );
  OAI32D0BWP12T U167 ( .A1(n206), .A2(N706), .A3(n36), .B1(n37), .B2(n206), 
        .ZN(n76) );
  NR4D0BWP12T U168 ( .A1(itstate[3]), .A2(itstate[0]), .A3(itstate[2]), .A4(
        itstate[1]), .ZN(n38) );
  ND4D0BWP12T U169 ( .A1(n329), .A2(n57), .A3(n38), .A4(n65), .ZN(n285) );
  CKND2D0BWP12T U170 ( .A1(alu_opcode[4]), .A2(n512), .ZN(n39) );
  NR4D0BWP12T U171 ( .A1(n448), .A2(n144), .A3(n187), .A4(n395), .ZN(n40) );
  AOI32D0BWP12T U172 ( .A1(n455), .A2(n39), .A3(n40), .B1(n478), .B2(n39), 
        .ZN(n670) );
  AOI211D0BWP12T U173 ( .A1(step[7]), .A2(n512), .B(n387), .C(n365), .ZN(n41)
         );
  AOI32D0BWP12T U174 ( .A1(n198), .A2(n41), .A3(n391), .B1(n390), .B2(n41), 
        .ZN(next_step[7]) );
  AOI31D0BWP12T U175 ( .A1(n188), .A2(n155), .A3(n469), .B(n468), .ZN(n42) );
  NR2D0BWP12T U176 ( .A1(n191), .A2(n42), .ZN(n221) );
  AO31D0BWP12T U177 ( .A1(n176), .A2(n177), .A3(n139), .B(n141), .Z(n43) );
  CKND2D0BWP12T U178 ( .A1(n198), .A2(n43), .ZN(n463) );
  IND4D0BWP12T U179 ( .A1(n295), .B1(instruction[6]), .B2(n447), .B3(n324), 
        .ZN(n44) );
  NR2D0BWP12T U180 ( .A1(n44), .A2(n280), .ZN(n45) );
  OA21D0BWP12T U181 ( .A1(n45), .A2(n395), .B(n508), .Z(n46) );
  AOI31D0BWP12T U182 ( .A1(n293), .A2(n398), .A3(n333), .B(n46), .ZN(n47) );
  AOI32D0BWP12T U183 ( .A1(n286), .A2(n287), .A3(n47), .B1(n285), .B2(n287), 
        .ZN(next_update_flag_v) );
  AOI22D0BWP12T U184 ( .A1(step[1]), .A2(n512), .B1(n144), .B2(n370), .ZN(n48)
         );
  AOI21D0BWP12T U185 ( .A1(N707), .A2(n387), .B(n106), .ZN(n49) );
  OAI211D0BWP12T U186 ( .A1(n178), .A2(n390), .B(n48), .C(n49), .ZN(
        next_step[1]) );
  CKND2D1BWP12T U187 ( .A1(instruction[12]), .A2(instruction[11]), .ZN(n392)
         );
  NR2D1BWP12T U188 ( .A1(instruction[15]), .A2(instruction[14]), .ZN(n352) );
  INVD1BWP12T U189 ( .I(n352), .ZN(n143) );
  TPOAI21D0BWP12T U190 ( .A1(instruction[10]), .A2(n392), .B(n450), .ZN(n343)
         );
  AOI22D0BWP12T U191 ( .A1(itstate[6]), .A2(flag_v), .B1(flag_c), .B2(n57), 
        .ZN(n51) );
  TPOAI21D0BWP12T U192 ( .A1(itstate[6]), .A2(n299), .B(itstate[7]), .ZN(n50)
         );
  CKND2D0BWP12T U193 ( .A1(itstate[6]), .A2(n292), .ZN(n54) );
  INVD1BWP12T U194 ( .I(itstate[6]), .ZN(n334) );
  TPND2D0BWP12T U195 ( .A1(n334), .A2(n58), .ZN(n53) );
  OR2D0BWP12T U196 ( .A1(flag_n), .A2(n334), .Z(n52) );
  INVD1BWP12T U197 ( .I(itstate[7]), .ZN(n336) );
  AOI32D1BWP12T U198 ( .A1(n54), .A2(itstate[7]), .A3(n53), .B1(n52), .B2(n336), .ZN(n55) );
  AOI211XD0BWP12T U199 ( .A1(n57), .A2(n56), .B(itstate[5]), .C(n55), .ZN(n63)
         );
  AOI22D0BWP12T U200 ( .A1(itstate[6]), .A2(flag_n), .B1(flag_z), .B2(n334), 
        .ZN(n60) );
  AOI32D0BWP12T U201 ( .A1(n298), .A2(n334), .A3(n329), .B1(itstate[6]), .B2(
        n294), .ZN(n59) );
  OAI32D0BWP12T U202 ( .A1(itstate[7]), .A2(itstate[5]), .A3(n60), .B1(n59), 
        .B2(n336), .ZN(n61) );
  NR2D1BWP12T U203 ( .A1(n64), .A2(n61), .ZN(n62) );
  OAI32D1BWP12T U204 ( .A1(n65), .A2(n64), .A3(n63), .B1(n62), .B2(itstate[4]), 
        .ZN(n66) );
  AOI21D1BWP12T U205 ( .A1(split_instruction), .A2(stall_to_instructionfetch), 
        .B(instruction_valid), .ZN(n67) );
  IND2D1BWP12T U206 ( .A1(reset), .B1(n68), .ZN(n274) );
  CKND2D1BWP12T U207 ( .A1(instruction[13]), .A2(n352), .ZN(n419) );
  AOI22D0BWP12T U208 ( .A1(n512), .A2(offset_b[1]), .B1(n501), .B2(
        instruction[1]), .ZN(n109) );
  ND3D1BWP12T U209 ( .A1(instruction[13]), .A2(instruction[15]), .A3(
        instruction[14]), .ZN(n95) );
  NR2D1BWP12T U210 ( .A1(n470), .A2(n308), .ZN(n433) );
  INVD1BWP12T U211 ( .I(n428), .ZN(n468) );
  INVD1BWP12T U212 ( .I(instruction[14]), .ZN(n92) );
  ND3D1BWP12T U213 ( .A1(instruction[15]), .A2(instruction[13]), .A3(n92), 
        .ZN(n325) );
  IND2XD1BWP12T U214 ( .A1(n325), .B1(instruction[12]), .ZN(n96) );
  CKND2D0BWP12T U215 ( .A1(n468), .A2(n422), .ZN(n431) );
  INVD1BWP12T U216 ( .I(instruction[7]), .ZN(n447) );
  NR2D2BWP12T U217 ( .A1(N706), .A2(N707), .ZN(n151) );
  TPNR2D0BWP12T U218 ( .A1(N703), .A2(n70), .ZN(n69) );
  ND2D1BWP12T U219 ( .A1(N702), .A2(n69), .ZN(n163) );
  TPNR2D0BWP12T U220 ( .A1(n75), .A2(n205), .ZN(n72) );
  NR4D0BWP12T U221 ( .A1(instruction[7]), .A2(N701), .A3(N702), .A4(N703), 
        .ZN(n71) );
  ND2D1BWP12T U222 ( .A1(N704), .A2(n151), .ZN(n149) );
  NR4D0BWP12T U223 ( .A1(instruction[7]), .A2(N701), .A3(N702), .A4(n382), 
        .ZN(n206) );
  INVD1BWP12T U224 ( .I(N707), .ZN(n159) );
  OAI211D1BWP12T U225 ( .A1(instruction[7]), .A2(n72), .B(n154), .C(n76), .ZN(
        n148) );
  INR2D0BWP12T U226 ( .A1(n75), .B1(instruction[7]), .ZN(n162) );
  INR2D1BWP12T U227 ( .A1(n76), .B1(n162), .ZN(n155) );
  TPND3D0BWP12T U228 ( .A1(instruction[7]), .A2(n78), .A3(n77), .ZN(n160) );
  CKND2D1BWP12T U229 ( .A1(n370), .A2(n428), .ZN(n379) );
  TPNR2D1BWP12T U230 ( .A1(N541), .A2(N540), .ZN(n79) );
  NR3D1BWP12T U231 ( .A1(N543), .A2(N542), .A3(n81), .ZN(n83) );
  NR2D2BWP12T U232 ( .A1(N545), .A2(N546), .ZN(n88) );
  NR4D0BWP12T U233 ( .A1(instruction[8]), .A2(N539), .A3(N540), .A4(n138), 
        .ZN(n175) );
  IND3D1BWP12T U234 ( .A1(N543), .B1(n80), .B2(N542), .ZN(n137) );
  IND2D1BWP12T U235 ( .A1(n90), .B1(N539), .ZN(n176) );
  NR3D1BWP12T U236 ( .A1(N542), .A2(n177), .A3(n81), .ZN(n82) );
  TPAOI31D0BWP12T U237 ( .A1(n88), .A2(N544), .A3(n83), .B(n82), .ZN(n87) );
  IND3D1BWP12T U238 ( .A1(N541), .B1(N540), .B2(n84), .ZN(n140) );
  INR2D1BWP12T U239 ( .A1(n85), .B1(n140), .ZN(n203) );
  INVD1BWP12T U240 ( .I(n203), .ZN(n86) );
  OAI211D1BWP12T U241 ( .A1(instruction[8]), .A2(n176), .B(n87), .C(n86), .ZN(
        n464) );
  NR2D1BWP12T U242 ( .A1(n370), .A2(n512), .ZN(n486) );
  TPNR2D0BWP12T U243 ( .A1(instruction[12]), .A2(n325), .ZN(n120) );
  OAI32D0BWP12T U244 ( .A1(instruction[9]), .A2(instruction[11]), .A3(
        instruction[8]), .B1(n483), .B2(instruction[9]), .ZN(n91) );
  CKND2D1BWP12T U245 ( .A1(instruction[11]), .A2(n451), .ZN(n121) );
  OAI22D0BWP12T U246 ( .A1(n91), .A2(n96), .B1(n95), .B2(n121), .ZN(n129) );
  NR2D1BWP12T U247 ( .A1(n92), .A2(instruction[15]), .ZN(n99) );
  IND2D1BWP12T U248 ( .A1(instruction[13]), .B1(n99), .ZN(n98) );
  CKND2D1BWP12T U249 ( .A1(n143), .A2(n499), .ZN(n243) );
  NR2D1BWP12T U250 ( .A1(instruction[11]), .A2(instruction[10]), .ZN(n303) );
  NR2D1BWP12T U251 ( .A1(instruction[8]), .A2(instruction[9]), .ZN(n295) );
  INVD1BWP12T U252 ( .I(n448), .ZN(n122) );
  TPND2D0BWP12T U253 ( .A1(n498), .A2(n122), .ZN(n269) );
  NR4D0BWP12T U254 ( .A1(n120), .A2(n129), .A3(n243), .A4(n269), .ZN(n184) );
  CKND2D0BWP12T U255 ( .A1(n100), .A2(instruction[12]), .ZN(n97) );
  TPNR2D0BWP12T U256 ( .A1(instruction[14]), .A2(n97), .ZN(n461) );
  CKND2D1BWP12T U257 ( .A1(instruction[13]), .A2(n99), .ZN(n412) );
  INR2D0BWP12T U258 ( .A1(n100), .B1(instruction[14]), .ZN(n101) );
  ND2D1BWP12T U259 ( .A1(n101), .A2(n451), .ZN(n411) );
  CKND2D1BWP12T U260 ( .A1(n110), .A2(n241), .ZN(n270) );
  TPNR2D0BWP12T U261 ( .A1(n170), .A2(n270), .ZN(n186) );
  OAI21D0BWP12T U262 ( .A1(N911), .A2(n470), .B(n492), .ZN(n102) );
  TPAOI31D0BWP12T U263 ( .A1(n184), .A2(n186), .A3(n102), .B(n485), .ZN(n103)
         );
  RCAOI211D0BWP12T U264 ( .A1(n381), .A2(n355), .B(n486), .C(n103), .ZN(n104)
         );
  OAI21D1BWP12T U265 ( .A1(n358), .A2(n379), .B(n104), .ZN(n106) );
  INVD1BWP12T U266 ( .I(instruction[0]), .ZN(n437) );
  OAI22D0BWP12T U267 ( .A1(n126), .A2(n437), .B1(n411), .B2(n333), .ZN(n107)
         );
  TPOAI31D0BWP12T U268 ( .A1(n426), .A2(n431), .A3(n107), .B(n508), .ZN(n108)
         );
  OAI211D0BWP12T U269 ( .A1(n343), .A2(n420), .B(n109), .C(n108), .ZN(n672) );
  AOI22D0BWP12T U270 ( .A1(n512), .A2(offset_b[3]), .B1(n501), .B2(
        instruction[3]), .ZN(n114) );
  INVD1BWP12T U271 ( .I(n120), .ZN(n490) );
  INVD1BWP12T U272 ( .I(instruction[1]), .ZN(n500) );
  OAI22D0BWP12T U273 ( .A1(n127), .A2(n500), .B1(n407), .B2(n411), .ZN(n112)
         );
  INVD0BWP12T U274 ( .I(instruction[2]), .ZN(n342) );
  CKND2D1BWP12T U275 ( .A1(n450), .A2(n392), .ZN(n445) );
  OAI22D0BWP12T U276 ( .A1(n126), .A2(n342), .B1(n488), .B2(n445), .ZN(n111)
         );
  OAI21D0BWP12T U277 ( .A1(n112), .A2(n111), .B(n508), .ZN(n113) );
  OAI211D0BWP12T U278 ( .A1(n420), .A2(n412), .B(n114), .C(n113), .ZN(n674) );
  AOI22D0BWP12T U279 ( .A1(n512), .A2(offset_b[2]), .B1(n501), .B2(
        instruction[2]), .ZN(n118) );
  OAI22D0BWP12T U280 ( .A1(n127), .A2(n437), .B1(n412), .B2(n333), .ZN(n116)
         );
  TPOAI22D0BWP12T U281 ( .A1(n126), .A2(n500), .B1(n343), .B2(n407), .ZN(n115)
         );
  OAI21D0BWP12T U282 ( .A1(n116), .A2(n115), .B(n508), .ZN(n117) );
  OAI211D0BWP12T U283 ( .A1(n420), .A2(n411), .B(n118), .C(n117), .ZN(n673) );
  AO222D1BWP12T U284 ( .A1(n442), .A2(n416), .B1(n441), .B2(n506), .C1(
        offset_b[8]), .C2(n512), .Z(n679) );
  AOI211D0BWP12T U285 ( .A1(n512), .A2(alu_write_to_reg[0]), .B(n381), .C(n486), .ZN(n125) );
  CKND2D1BWP12T U286 ( .A1(instruction[10]), .A2(n505), .ZN(n231) );
  AOI211D0BWP12T U287 ( .A1(n447), .A2(instruction[6]), .B(n488), .C(
        instruction[8]), .ZN(n119) );
  IAO21D0BWP12T U288 ( .A1(n280), .A2(n119), .B(n450), .ZN(n314) );
  OAI21D0BWP12T U289 ( .A1(instruction[8]), .A2(n231), .B(n314), .ZN(n481) );
  CKND2D1BWP12T U290 ( .A1(instruction[8]), .A2(n488), .ZN(n291) );
  AOI21D1BWP12T U291 ( .A1(n119), .A2(n449), .B(n394), .ZN(n354) );
  IND3D1BWP12T U292 ( .A1(n129), .B1(n186), .B2(n354), .ZN(n145) );
  INVD0BWP12T U293 ( .I(n419), .ZN(n260) );
  AOI211XD0BWP12T U294 ( .A1(n260), .A2(n121), .B(n428), .C(n120), .ZN(n484)
         );
  TPND2D0BWP12T U295 ( .A1(instruction[9]), .A2(n432), .ZN(n128) );
  AOI32D0BWP12T U296 ( .A1(n484), .A2(n122), .A3(n128), .B1(n407), .B2(n122), 
        .ZN(n123) );
  AOI211D0BWP12T U297 ( .A1(instruction[0]), .A2(n481), .B(n145), .C(n123), 
        .ZN(n124) );
  AOI32D0BWP12T U298 ( .A1(n126), .A2(n125), .A3(n124), .B1(n485), .B2(n125), 
        .ZN(n641) );
  INVD1BWP12T U299 ( .I(n450), .ZN(n397) );
  CKND2D1BWP12T U300 ( .A1(n241), .A2(n397), .ZN(n496) );
  CKND2D0BWP12T U301 ( .A1(n498), .A2(n127), .ZN(n132) );
  TPNR2D0BWP12T U302 ( .A1(n428), .A2(n260), .ZN(n489) );
  OR2XD1BWP12T U303 ( .A1(n129), .A2(n170), .Z(n268) );
  AOI211D1BWP12T U304 ( .A1(n260), .A2(n502), .B(n491), .C(n268), .ZN(n253) );
  NR2XD0BWP12T U305 ( .A1(instruction[11]), .A2(n308), .ZN(n289) );
  AOI211D0BWP12T U306 ( .A1(n505), .A2(instruction[0]), .B(n289), .C(n144), 
        .ZN(n130) );
  OAI211D1BWP12T U307 ( .A1(n489), .A2(n407), .B(n253), .C(n130), .ZN(n131) );
  RCAOI211D0BWP12T U308 ( .A1(instruction[3]), .A2(n496), .B(n132), .C(n131), 
        .ZN(n134) );
  AOI211D0BWP12T U309 ( .A1(n512), .A2(operand_a[0]), .B(n381), .C(n486), .ZN(
        n133) );
  OAI21D0BWP12T U310 ( .A1(n134), .A2(n485), .B(n133), .ZN(n635) );
  IND3D0BWP12T U311 ( .A1(n405), .B1(n498), .B2(n241), .ZN(n430) );
  CKND2D0BWP12T U312 ( .A1(instruction[12]), .A2(n260), .ZN(n135) );
  AOI32D0BWP12T U313 ( .A1(n308), .A2(n468), .A3(n135), .B1(instruction[11]), 
        .B2(n468), .ZN(n136) );
  AOI211XD0BWP12T U314 ( .A1(n295), .A2(n432), .B(n430), .C(n136), .ZN(n455)
         );
  NR2D1BWP12T U315 ( .A1(n138), .A2(n141), .ZN(n183) );
  RCAOI211D0BWP12T U316 ( .A1(n142), .A2(n356), .B(n183), .C(n463), .ZN(n424)
         );
  NR2D0BWP12T U317 ( .A1(n143), .A2(n392), .ZN(n395) );
  INVD1BWP12T U318 ( .I(alu_write_to_reg[4]), .ZN(n147) );
  OAI21D0BWP12T U319 ( .A1(n426), .A2(n145), .B(n370), .ZN(n146) );
  OAI211D0BWP12T U320 ( .A1(n274), .A2(n147), .B(n146), .C(n278), .ZN(n640) );
  CKND2D1BWP12T U321 ( .A1(instruction[9]), .A2(n256), .ZN(n348) );
  OAI21D1BWP12T U322 ( .A1(N706), .A2(N707), .B(n150), .ZN(n357) );
  OAI22D1BWP12T U323 ( .A1(n382), .A2(n148), .B1(n163), .B2(n153), .ZN(n386)
         );
  INR2XD0BWP12T U324 ( .A1(n357), .B1(n386), .ZN(n188) );
  OR3D1BWP12T U325 ( .A1(N705), .A2(n149), .A3(n148), .Z(n378) );
  ND3D1BWP12T U326 ( .A1(N705), .A2(n151), .A3(n150), .ZN(n362) );
  OAI211D0BWP12T U327 ( .A1(n153), .A2(n152), .B(n378), .C(n362), .ZN(n189) );
  INR3XD0BWP12T U328 ( .A1(n154), .B1(n204), .B2(n189), .ZN(n469) );
  AOI21D1BWP12T U329 ( .A1(n256), .A2(n488), .B(n259), .ZN(n460) );
  INVD1BWP12T U330 ( .I(n461), .ZN(n239) );
  CKND2D1BWP12T U331 ( .A1(n460), .A2(n239), .ZN(n191) );
  CKND2D1BWP12T U332 ( .A1(instruction[11]), .A2(n187), .ZN(n453) );
  OAI21D1BWP12T U333 ( .A1(n221), .A2(n470), .B(n453), .ZN(n156) );
  TPOAI31D0BWP12T U334 ( .A1(n493), .A2(n473), .A3(n156), .B(n508), .ZN(n158)
         );
  OAI21D0BWP12T U335 ( .A1(n274), .A2(n157), .B(n158), .ZN(n683) );
  IOA21D1BWP12T U336 ( .A1(n512), .A2(memory_write_to_reg_enable), .B(n158), 
        .ZN(n650) );
  NR2D0BWP12T U337 ( .A1(n460), .A2(n485), .ZN(n211) );
  CKND2D0BWP12T U338 ( .A1(N706), .A2(n159), .ZN(n161) );
  ND3D0BWP12T U339 ( .A1(n161), .A2(n378), .A3(n160), .ZN(n165) );
  TPNR2D0BWP12T U340 ( .A1(n219), .A2(n162), .ZN(n209) );
  CKND2D0BWP12T U341 ( .A1(n209), .A2(n163), .ZN(n164) );
  TPOAI31D0BWP12T U342 ( .A1(n166), .A2(n165), .A3(n164), .B(n387), .ZN(n167)
         );
  OAI31D0BWP12T U343 ( .A1(n407), .A2(n485), .A3(n239), .B(n167), .ZN(n168) );
  AOI211D0BWP12T U344 ( .A1(instruction[0]), .A2(n211), .B(n486), .C(n168), 
        .ZN(n375) );
  IND3D1BWP12T U345 ( .A1(n170), .B1(n184), .B2(n308), .ZN(n196) );
  OA21XD0BWP12T U346 ( .A1(n428), .A2(n191), .B(n370), .Z(n368) );
  AOI22D0BWP12T U347 ( .A1(memory_write_to_reg[0]), .A2(n512), .B1(n470), .B2(
        n368), .ZN(n172) );
  AOI22D0BWP12T U348 ( .A1(instruction[8]), .A2(n493), .B1(instruction[0]), 
        .B2(n473), .ZN(n171) );
  AOI32D0BWP12T U349 ( .A1(n220), .A2(n172), .A3(n171), .B1(n485), .B2(n172), 
        .ZN(n180) );
  CKND2D0BWP12T U350 ( .A1(instruction[11]), .A2(n173), .ZN(n224) );
  INR4D0BWP12T U351 ( .A1(n176), .B1(n175), .B2(n174), .B3(n183), .ZN(n199) );
  AOI21D0BWP12T U352 ( .A1(n178), .A2(N545), .B(n182), .ZN(n179) );
  CKND2D1BWP12T U353 ( .A1(n199), .A2(n179), .ZN(n371) );
  OAI32D0BWP12T U354 ( .A1(n180), .A2(n224), .A3(n371), .B1(n381), .B2(n180), 
        .ZN(n181) );
  CKND2D1BWP12T U355 ( .A1(n375), .A2(n181), .ZN(n649) );
  NR3XD0BWP12T U356 ( .A1(n355), .A2(N544), .A3(n356), .ZN(n367) );
  IND2D1BWP12T U357 ( .A1(n182), .B1(n367), .ZN(n380) );
  NR3XD0BWP12T U358 ( .A1(n376), .A2(n183), .A3(n380), .ZN(n391) );
  INR2D0BWP12T U359 ( .A1(n184), .B1(n492), .ZN(n185) );
  AOI32D1BWP12T U360 ( .A1(n186), .A2(n278), .A3(n185), .B1(n485), .B2(n278), 
        .ZN(n365) );
  TPND3D0BWP12T U361 ( .A1(n508), .A2(n187), .A3(n470), .ZN(n400) );
  IND2XD1BWP12T U362 ( .A1(n189), .B1(n188), .ZN(n427) );
  AOI211D0BWP12T U363 ( .A1(n470), .A2(n190), .B(n204), .C(n427), .ZN(n192) );
  MOAI22D0BWP12T U364 ( .A1(n192), .A2(n468), .B1(n470), .B2(n191), .ZN(n193)
         );
  OAI21D0BWP12T U365 ( .A1(n471), .A2(n193), .B(n508), .ZN(n194) );
  OAI211D0BWP12T U366 ( .A1(n274), .A2(memory_store_request_BAR), .B(n400), 
        .C(n194), .ZN(n665) );
  NR2D0BWP12T U367 ( .A1(n303), .A2(n239), .ZN(n197) );
  NR2XD0BWP12T U368 ( .A1(n493), .A2(n196), .ZN(n240) );
  IND2D1BWP12T U369 ( .A1(n473), .B1(n240), .ZN(n369) );
  AOI211D0BWP12T U370 ( .A1(n471), .A2(instruction[2]), .B(n197), .C(n369), 
        .ZN(n213) );
  ND3XD0BWP12T U371 ( .A1(n200), .A2(n199), .A3(n198), .ZN(n201) );
  TPOAI31D0BWP12T U372 ( .A1(n203), .A2(n202), .A3(n201), .B(n381), .ZN(n208)
         );
  NR4D0BWP12T U373 ( .A1(n206), .A2(n205), .A3(n204), .A4(n386), .ZN(n207) );
  AOI32D0BWP12T U374 ( .A1(n209), .A2(n208), .A3(n207), .B1(n379), .B2(n208), 
        .ZN(n210) );
  AOI211XD0BWP12T U375 ( .A1(instruction[2]), .A2(n211), .B(n486), .C(n210), 
        .ZN(n217) );
  IND3D0BWP12T U376 ( .A1(n211), .B1(n379), .B2(n390), .ZN(n215) );
  AOI22D0BWP12T U377 ( .A1(instruction[11]), .A2(n215), .B1(n512), .B2(
        memory_store_data_reg[2]), .ZN(n212) );
  OAI211D0BWP12T U378 ( .A1(n213), .A2(n485), .B(n217), .C(n212), .ZN(n653) );
  TPNR2D0BWP12T U379 ( .A1(instruction[10]), .A2(n470), .ZN(n331) );
  AOI22D0BWP12T U380 ( .A1(instruction[10]), .A2(n493), .B1(instruction[2]), 
        .B2(n473), .ZN(n214) );
  OA211D1BWP12T U381 ( .A1(n331), .A2(n239), .B(n220), .C(n214), .Z(n218) );
  AOI22D0BWP12T U382 ( .A1(memory_write_to_reg[2]), .A2(n512), .B1(n470), .B2(
        n215), .ZN(n216) );
  OAI211D0BWP12T U383 ( .A1(n218), .A2(n485), .B(n217), .C(n216), .ZN(n647) );
  TPND2D0BWP12T U384 ( .A1(n428), .A2(n219), .ZN(n232) );
  OAI211D0BWP12T U385 ( .A1(instruction[11]), .A2(n221), .B(n220), .C(n232), 
        .ZN(n223) );
  AOI21D0BWP12T U386 ( .A1(n370), .A2(n223), .B(n235), .ZN(n227) );
  AOI22D0BWP12T U387 ( .A1(n512), .A2(memory_write_to_reg[3]), .B1(n381), .B2(
        n224), .ZN(n225) );
  CKND2D1BWP12T U388 ( .A1(n227), .A2(n225), .ZN(n646) );
  AOI22D0BWP12T U389 ( .A1(memory_write_to_reg[4]), .A2(n512), .B1(n381), .B2(
        n470), .ZN(n226) );
  CKND2D1BWP12T U390 ( .A1(n227), .A2(n226), .ZN(n645) );
  CKND0BWP12T U391 ( .I(memory_address_source_is_reg), .ZN(n228) );
  CKND2D0BWP12T U392 ( .A1(n508), .A2(n428), .ZN(n458) );
  OAI211D0BWP12T U393 ( .A1(n274), .A2(n228), .B(n458), .C(n400), .ZN(n661) );
  NR4D0BWP12T U394 ( .A1(n462), .A2(n492), .A3(n229), .A4(n442), .ZN(n252) );
  IND4D1BWP12T U395 ( .A1(n259), .B1(n343), .B2(n252), .B3(n489), .ZN(n504) );
  OAI32D0BWP12T U396 ( .A1(n486), .A2(n268), .A3(n504), .B1(n370), .B2(n486), 
        .ZN(n266) );
  INVD1BWP12T U397 ( .I(n266), .ZN(n510) );
  AOI21D0BWP12T U398 ( .A1(n512), .A2(operand_b[3]), .B(n510), .ZN(n230) );
  OAI31D0BWP12T U399 ( .A1(n485), .A2(n333), .A3(n231), .B(n230), .ZN(n630) );
  ND2D0BWP12T U400 ( .A1(n470), .A2(n232), .ZN(n233) );
  OAI32D0BWP12T U401 ( .A1(n235), .A2(n369), .A3(n233), .B1(n370), .B2(n235), 
        .ZN(n238) );
  AOI22D0BWP12T U402 ( .A1(n512), .A2(memory_store_data_reg[3]), .B1(n465), 
        .B2(n381), .ZN(n234) );
  TPND2D0BWP12T U403 ( .A1(n238), .A2(n234), .ZN(n652) );
  CKND2D1BWP12T U404 ( .A1(n433), .A2(N911), .ZN(n346) );
  CKND2D1BWP12T U405 ( .A1(n253), .A2(n346), .ZN(n250) );
  AOI211D0BWP12T U406 ( .A1(instruction[9]), .A2(n449), .B(n394), .C(n250), 
        .ZN(n237) );
  AOI21D0BWP12T U407 ( .A1(n512), .A2(alu_opcode[3]), .B(n235), .ZN(n236) );
  OAI21D0BWP12T U408 ( .A1(n237), .A2(n485), .B(n236), .ZN(n669) );
  IOA21D1BWP12T U409 ( .A1(n512), .A2(memory_store_data_reg[4]), .B(n238), 
        .ZN(n651) );
  AO31D0BWP12T U410 ( .A1(n241), .A2(n240), .A3(n239), .B(n485), .Z(n242) );
  CKND2D1BWP12T U411 ( .A1(n278), .A2(n242), .ZN(n459) );
  IOA21D1BWP12T U412 ( .A1(n512), .A2(memory_store_address_reg[3]), .B(n249), 
        .ZN(n657) );
  INR3XD0BWP12T U413 ( .A1(n252), .B1(n428), .B2(n268), .ZN(n262) );
  AOI31D0BWP12T U414 ( .A1(n256), .A2(n483), .A3(n488), .B(n243), .ZN(n244) );
  OAI211D0BWP12T U415 ( .A1(instruction[12]), .A2(n412), .B(n262), .C(n244), 
        .ZN(n245) );
  AOI22D0BWP12T U416 ( .A1(n370), .A2(n245), .B1(n512), .B2(
        load_store_width[1]), .ZN(n246) );
  CKND2D1BWP12T U417 ( .A1(n246), .A2(n278), .ZN(n662) );
  AOI22D0BWP12T U418 ( .A1(n512), .A2(memory_store_address_reg[2]), .B1(n387), 
        .B2(instruction[10]), .ZN(n247) );
  CKND2D1BWP12T U419 ( .A1(n249), .A2(n247), .ZN(n658) );
  AOI22D0BWP12T U420 ( .A1(n512), .A2(memory_store_address_reg[0]), .B1(n387), 
        .B2(instruction[8]), .ZN(n248) );
  CKND2D1BWP12T U421 ( .A1(n249), .A2(n248), .ZN(n660) );
  AOI22D0BWP12T U422 ( .A1(n370), .A2(n250), .B1(n512), .B2(operand_a[4]), 
        .ZN(n251) );
  ND2D0BWP12T U423 ( .A1(n251), .A2(n278), .ZN(n634) );
  INVD1BWP12T U424 ( .I(operand_a[3]), .ZN(n255) );
  CKND2D1BWP12T U425 ( .A1(n253), .A2(n252), .ZN(n276) );
  AOI32D0BWP12T U426 ( .A1(instruction[7]), .A2(n370), .A3(n432), .B1(n276), 
        .B2(n370), .ZN(n254) );
  OAI211D0BWP12T U427 ( .A1(n274), .A2(n255), .B(n254), .C(n278), .ZN(n636) );
  IND2XD1BWP12T U428 ( .A1(n256), .B1(n397), .ZN(n507) );
  AOI22D0BWP12T U429 ( .A1(instruction[5]), .A2(n505), .B1(instruction[8]), 
        .B2(n507), .ZN(n258) );
  CKND2D0BWP12T U430 ( .A1(n512), .A2(operand_b[2]), .ZN(n257) );
  OAI211D0BWP12T U431 ( .A1(n258), .A2(n485), .B(n266), .C(n257), .ZN(n631) );
  AOI211D0BWP12T U432 ( .A1(n260), .A2(n470), .B(instruction[12]), .C(n259), 
        .ZN(n263) );
  AOI22D0BWP12T U433 ( .A1(instruction[8]), .A2(n449), .B1(n432), .B2(n291), 
        .ZN(n261) );
  AOI31D0BWP12T U434 ( .A1(n263), .A2(n262), .A3(n261), .B(n485), .ZN(n264) );
  AO211D0BWP12T U435 ( .A1(n512), .A2(alu_opcode[2]), .B(n264), .C(n486), .Z(
        n668) );
  AOI22D0BWP12T U436 ( .A1(n505), .A2(instruction[3]), .B1(instruction[6]), 
        .B2(n507), .ZN(n267) );
  CKND2D0BWP12T U437 ( .A1(n512), .A2(operand_b[0]), .ZN(n265) );
  OAI211D0BWP12T U438 ( .A1(n267), .A2(n485), .B(n266), .C(n265), .ZN(n633) );
  INVD1BWP12T U439 ( .I(alu_write_to_reg[3]), .ZN(n273) );
  AOI21D0BWP12T U440 ( .A1(instruction[8]), .A2(n491), .B(n492), .ZN(n476) );
  NR4D0BWP12T U441 ( .A1(n462), .A2(n270), .A3(n269), .A4(n268), .ZN(n271) );
  ND3D1BWP12T U442 ( .A1(n354), .A2(n476), .A3(n271), .ZN(n480) );
  AOI32D0BWP12T U443 ( .A1(instruction[7]), .A2(n370), .A3(n432), .B1(n480), 
        .B2(n370), .ZN(n272) );
  OAI211D0BWP12T U444 ( .A1(n274), .A2(n273), .B(n272), .C(n278), .ZN(n642) );
  OAI22D0BWP12T U445 ( .A1(n489), .A2(n483), .B1(n499), .B2(n342), .ZN(n275)
         );
  AOI211D0BWP12T U446 ( .A1(instruction[5]), .A2(n496), .B(n276), .C(n275), 
        .ZN(n279) );
  CKND2D0BWP12T U447 ( .A1(n512), .A2(operand_a[2]), .ZN(n277) );
  OAI211D0BWP12T U448 ( .A1(n279), .A2(n485), .B(n278), .C(n277), .ZN(n637) );
  CKND0BWP12T U449 ( .I(n291), .ZN(n293) );
  TPNR2D0BWP12T U450 ( .A1(n420), .A2(n280), .ZN(n398) );
  ND2XD0BWP12T U451 ( .A1(instruction[8]), .A2(instruction[9]), .ZN(n324) );
  TPNR2D0BWP12T U452 ( .A1(instruction[8]), .A2(n488), .ZN(n281) );
  AOI22D0BWP12T U453 ( .A1(n508), .A2(n394), .B1(n281), .B2(n398), .ZN(n287)
         );
  CKND2D0BWP12T U454 ( .A1(instruction[12]), .A2(n501), .ZN(n286) );
  AOI21D0BWP12T U455 ( .A1(n407), .A2(instruction[6]), .B(n293), .ZN(n283) );
  OAI22D0BWP12T U456 ( .A1(n283), .A2(n478), .B1(n282), .B2(n420), .ZN(n284)
         );
  AOI22D0BWP12T U457 ( .A1(n508), .A2(n450), .B1(n449), .B2(n284), .ZN(n288)
         );
  AOI32D0BWP12T U458 ( .A1(n288), .A2(n287), .A3(n286), .B1(n285), .B2(n287), 
        .ZN(next_update_flag_c) );
  TPND2D0BWP12T U459 ( .A1(n508), .A2(n289), .ZN(n341) );
  AOI22D0BWP12T U460 ( .A1(n512), .A2(offset_b[18]), .B1(instruction[6]), .B2(
        n322), .ZN(n290) );
  ND2D0BWP12T U461 ( .A1(n290), .A2(n511), .ZN(n622) );
  AOI211D0BWP12T U462 ( .A1(n432), .A2(n291), .B(n404), .C(n448), .ZN(n315) );
  AOI221D0BWP12T U463 ( .A1(n295), .A2(n294), .B1(n293), .B2(n292), .C(n470), 
        .ZN(n307) );
  AOI22D0BWP12T U464 ( .A1(instruction[9]), .A2(flag_v), .B1(flag_n), .B2(n488), .ZN(n297) );
  NR2D0BWP12T U465 ( .A1(instruction[8]), .A2(n297), .ZN(n296) );
  AOI211D0BWP12T U466 ( .A1(instruction[8]), .A2(n297), .B(instruction[11]), 
        .C(n296), .ZN(n306) );
  AOI22D0BWP12T U467 ( .A1(instruction[9]), .A2(n299), .B1(n298), .B2(n488), 
        .ZN(n300) );
  MAOI22D0BWP12T U468 ( .A1(n300), .A2(n407), .B1(n300), .B2(n407), .ZN(n304)
         );
  AOI22D0BWP12T U469 ( .A1(instruction[9]), .A2(flag_c), .B1(flag_z), .B2(n488), .ZN(n301) );
  MAOI22D0BWP12T U470 ( .A1(n301), .A2(n407), .B1(n301), .B2(n407), .ZN(n302)
         );
  AOI22D0BWP12T U471 ( .A1(n331), .A2(n304), .B1(n303), .B2(n302), .ZN(n305)
         );
  OAI31D0BWP12T U472 ( .A1(n307), .A2(n306), .A3(n483), .B(n305), .ZN(n311) );
  CKND0BWP12T U473 ( .I(n484), .ZN(n310) );
  CKND2D0BWP12T U474 ( .A1(n308), .A2(n422), .ZN(n309) );
  AOI211D0BWP12T U475 ( .A1(n312), .A2(n311), .B(n310), .C(n309), .ZN(n313) );
  AOI31D0BWP12T U476 ( .A1(n315), .A2(n314), .A3(n313), .B(n478), .ZN(
        next_alu_write_to_reg_enable) );
  AOI22D0BWP12T U477 ( .A1(n512), .A2(offset_b[20]), .B1(instruction[8]), .B2(
        n322), .ZN(n316) );
  ND2D0BWP12T U478 ( .A1(n316), .A2(n511), .ZN(n620) );
  AOI22D0BWP12T U479 ( .A1(n512), .A2(offset_b[22]), .B1(instruction[10]), 
        .B2(n322), .ZN(n317) );
  ND2D0BWP12T U480 ( .A1(n317), .A2(n511), .ZN(n618) );
  AOI22D0BWP12T U481 ( .A1(n512), .A2(offset_b[21]), .B1(instruction[9]), .B2(
        n322), .ZN(n318) );
  ND2D0BWP12T U482 ( .A1(n318), .A2(n511), .ZN(n619) );
  AOI22D0BWP12T U483 ( .A1(n512), .A2(offset_b[16]), .B1(instruction[4]), .B2(
        n322), .ZN(n319) );
  ND2D0BWP12T U484 ( .A1(n319), .A2(n511), .ZN(n624) );
  AOI22D0BWP12T U485 ( .A1(instruction[5]), .A2(n322), .B1(n512), .B2(
        offset_b[17]), .ZN(n320) );
  ND2D0BWP12T U486 ( .A1(n320), .A2(n511), .ZN(n623) );
  AOI22D0BWP12T U487 ( .A1(n512), .A2(offset_b[15]), .B1(instruction[3]), .B2(
        n322), .ZN(n321) );
  ND2D0BWP12T U488 ( .A1(n321), .A2(n511), .ZN(n625) );
  AOI22D0BWP12T U489 ( .A1(n512), .A2(offset_b[19]), .B1(instruction[7]), .B2(
        n322), .ZN(n323) );
  ND2D0BWP12T U490 ( .A1(n323), .A2(n511), .ZN(n621) );
  NR3D0BWP12T U491 ( .A1(itstate[2]), .A2(itstate[1]), .A3(itstate[0]), .ZN(
        n326) );
  NR4D0BWP12T U492 ( .A1(n483), .A2(n325), .A3(n392), .A4(n324), .ZN(n327) );
  AOI211XD0BWP12T U493 ( .A1(itstate[3]), .A2(n326), .B(n327), .C(n485), .ZN(
        n349) );
  TPND2D0BWP12T U494 ( .A1(n370), .A2(n327), .ZN(n436) );
  OR4D1BWP12T U495 ( .A1(instruction[3]), .A2(instruction[2]), .A3(
        instruction[1]), .A4(instruction[0]), .Z(n328) );
  OAI22D0BWP12T U496 ( .A1(reset), .A2(n370), .B1(n436), .B2(n328), .ZN(n435)
         );
  NR2D1BWP12T U497 ( .A1(n349), .A2(n435), .ZN(n337) );
  INVD1BWP12T U498 ( .I(n436), .ZN(n350) );
  INVD1BWP12T U499 ( .I(n335), .ZN(n330) );
  AO222D0BWP12T U500 ( .A1(n435), .A2(itstate[4]), .B1(instruction[4]), .B2(
        n330), .C1(itstate[3]), .C2(n349), .Z(n687) );
  OAI32D0BWP12T U501 ( .A1(n478), .A2(n331), .A3(n348), .B1(n411), .B2(n478), 
        .ZN(n332) );
  AO21D0BWP12T U502 ( .A1(n512), .A2(load_store_width[0]), .B(n332), .Z(n663)
         );
  TPND2D0BWP12T U503 ( .A1(n512), .A2(offset_b[12]), .ZN(n338) );
  OAI211D0BWP12T U504 ( .A1(n437), .A2(n341), .B(n338), .C(n511), .ZN(n628) );
  TPND2D0BWP12T U505 ( .A1(n512), .A2(offset_b[13]), .ZN(n339) );
  OAI211D0BWP12T U506 ( .A1(n500), .A2(n341), .B(n511), .C(n339), .ZN(n627) );
  TPND2D0BWP12T U507 ( .A1(n512), .A2(offset_b[14]), .ZN(n340) );
  OAI211D0BWP12T U508 ( .A1(n342), .A2(n341), .B(n511), .C(n340), .ZN(n626) );
  AOI22D0BWP12T U509 ( .A1(n512), .A2(offset_b[0]), .B1(n501), .B2(
        instruction[0]), .ZN(n345) );
  IND2XD0BWP12T U510 ( .A1(n343), .B1(n416), .ZN(n344) );
  OAI211D0BWP12T U511 ( .A1(n346), .A2(n478), .B(n345), .C(n344), .ZN(n671) );
  TPND2D0BWP12T U512 ( .A1(n512), .A2(memorycontroller_sign_extend), .ZN(n347)
         );
  TPOAI31D0BWP12T U513 ( .A1(n470), .A2(n478), .A3(n348), .B(n347), .ZN(n664)
         );
  AO222D0BWP12T U514 ( .A1(n435), .A2(itstate[2]), .B1(instruction[2]), .B2(
        n350), .C1(itstate[1]), .C2(n349), .Z(n689) );
  AO222D0BWP12T U515 ( .A1(n435), .A2(itstate[1]), .B1(instruction[1]), .B2(
        n350), .C1(itstate[0]), .C2(n349), .Z(n690) );
  AO222D0BWP12T U516 ( .A1(n435), .A2(itstate[3]), .B1(instruction[3]), .B2(
        n350), .C1(itstate[2]), .C2(n349), .Z(n688) );
  OAI211D0BWP12T U517 ( .A1(n352), .A2(n449), .B(n370), .C(n351), .ZN(n353) );
  OAI21D1BWP12T U518 ( .A1(n354), .A2(n478), .B(n353), .ZN(next_update_flag_n)
         );
  NR2D0BWP12T U519 ( .A1(n356), .A2(n355), .ZN(n361) );
  INVD0BWP12T U520 ( .I(n365), .ZN(n360) );
  TPND2D0BWP12T U521 ( .A1(n358), .A2(n357), .ZN(n363) );
  AOI22D0BWP12T U522 ( .A1(n512), .A2(step[2]), .B1(n387), .B2(n363), .ZN(n359) );
  OAI211D1BWP12T U523 ( .A1(n361), .A2(n390), .B(n360), .C(n359), .ZN(
        next_step[2]) );
  INVD1BWP12T U524 ( .I(n362), .ZN(n364) );
  OAI32D1BWP12T U525 ( .A1(n365), .A2(n364), .A3(n363), .B1(n387), .B2(n365), 
        .ZN(n377) );
  CKND2D0BWP12T U526 ( .A1(n512), .A2(step[3]), .ZN(n366) );
  OAI211D1BWP12T U527 ( .A1(n367), .A2(n390), .B(n377), .C(n366), .ZN(
        next_step[3]) );
  AOI22D0BWP12T U528 ( .A1(instruction[11]), .A2(n368), .B1(n512), .B2(
        memory_store_data_reg[0]), .ZN(n374) );
  AOI32D0BWP12T U529 ( .A1(instruction[0]), .A2(n370), .A3(n471), .B1(n369), 
        .B2(n370), .ZN(n373) );
  OAI21D0BWP12T U530 ( .A1(instruction[11]), .A2(n371), .B(n381), .ZN(n372) );
  ND4D1BWP12T U531 ( .A1(n375), .A2(n374), .A3(n373), .A4(n372), .ZN(n655) );
  INVD1BWP12T U532 ( .I(n376), .ZN(n423) );
  OAI21D1BWP12T U533 ( .A1(n379), .A2(n378), .B(n377), .ZN(n385) );
  TPAOI21D0BWP12T U534 ( .A1(n381), .A2(n380), .B(n385), .ZN(n421) );
  INVD1BWP12T U535 ( .I(n382), .ZN(n383) );
  AOI22D0BWP12T U536 ( .A1(n512), .A2(step[5]), .B1(n387), .B2(n383), .ZN(n384) );
  OAI211D1BWP12T U537 ( .A1(n390), .A2(n423), .B(n421), .C(n384), .ZN(
        next_step[5]) );
  INVD0BWP12T U538 ( .I(n385), .ZN(n389) );
  AOI22D0BWP12T U539 ( .A1(n512), .A2(step[6]), .B1(n387), .B2(n386), .ZN(n388) );
  OAI211D1BWP12T U540 ( .A1(n391), .A2(n390), .B(n389), .C(n388), .ZN(
        next_step[6]) );
  CKND0BWP12T U541 ( .I(n392), .ZN(n393) );
  AOI22D0BWP12T U542 ( .A1(n448), .A2(n506), .B1(n501), .B2(n393), .ZN(n402)
         );
  RCAOI211D0BWP12T U543 ( .A1(instruction[9]), .A2(n395), .B(n426), .C(n394), 
        .ZN(n396) );
  OAI32D0BWP12T U544 ( .A1(n478), .A2(instruction[12]), .A3(n397), .B1(n396), 
        .B2(n478), .ZN(n399) );
  AOI211XD0BWP12T U545 ( .A1(n512), .A2(alu_opcode[1]), .B(n399), .C(n398), 
        .ZN(n401) );
  ND3D1BWP12T U546 ( .A1(n402), .A2(n401), .A3(n400), .ZN(n667) );
  OAI21D1BWP12T U547 ( .A1(n404), .A2(n403), .B(n508), .ZN(n410) );
  AOI22D0BWP12T U548 ( .A1(n512), .A2(offset_b[9]), .B1(n506), .B2(n405), .ZN(
        n406) );
  OAI211D1BWP12T U549 ( .A1(n407), .A2(n410), .B(n406), .C(n511), .ZN(n680) );
  TPND2D0BWP12T U550 ( .A1(n512), .A2(offset_b[11]), .ZN(n408) );
  OAI211D1BWP12T U551 ( .A1(n483), .A2(n410), .B(n511), .C(n408), .ZN(n682) );
  TPND2D0BWP12T U552 ( .A1(n512), .A2(offset_b[10]), .ZN(n409) );
  OAI211D1BWP12T U553 ( .A1(n488), .A2(n410), .B(n511), .C(n409), .ZN(n681) );
  INVD1BWP12T U554 ( .I(n411), .ZN(n439) );
  AOI22D0BWP12T U555 ( .A1(instruction[10]), .A2(n439), .B1(instruction[4]), 
        .B2(n441), .ZN(n415) );
  AOI22D1BWP12T U556 ( .A1(instruction[5]), .A2(n501), .B1(n512), .B2(
        offset_b[5]), .ZN(n414) );
  INVD1BWP12T U557 ( .I(n412), .ZN(n440) );
  AOI22D0BWP12T U558 ( .A1(instruction[9]), .A2(n440), .B1(instruction[3]), 
        .B2(n442), .ZN(n413) );
  AOI32D1BWP12T U559 ( .A1(n415), .A2(n414), .A3(n413), .B1(n478), .B2(n414), 
        .ZN(n676) );
  AOI22D1BWP12T U560 ( .A1(n512), .A2(offset_b[7]), .B1(n416), .B2(n441), .ZN(
        n418) );
  ND3D0BWP12T U561 ( .A1(instruction[5]), .A2(n508), .A3(n442), .ZN(n417) );
  OAI211D1BWP12T U562 ( .A1(n420), .A2(n419), .B(n418), .C(n417), .ZN(n678) );
  IOA21D1BWP12T U563 ( .A1(n512), .A2(step[4]), .B(n421), .ZN(next_step[4]) );
  AOI21D0BWP12T U564 ( .A1(n424), .A2(n423), .B(n422), .ZN(n425) );
  AOI211XD0BWP12T U565 ( .A1(n428), .A2(n427), .B(n426), .C(n425), .ZN(n429)
         );
  MOAI22D0BWP12T U566 ( .A1(n429), .A2(n478), .B1(split_instruction), .B2(n512), .ZN(n693) );
  NR4D0BWP12T U567 ( .A1(n433), .A2(n432), .A3(n431), .A4(n430), .ZN(n434) );
  MOAI22D0BWP12T U568 ( .A1(n434), .A2(n478), .B1(stall_to_instructionfetch), 
        .B2(n512), .ZN(n692) );
  MOAI22D0BWP12T U569 ( .A1(n437), .A2(n436), .B1(itstate[0]), .B2(n435), .ZN(
        n691) );
  AO222D1BWP12T U570 ( .A1(n440), .A2(instruction[10]), .B1(instruction[4]), 
        .B2(n442), .C1(instruction[5]), .C2(n441), .Z(n438) );
  AO222D0BWP12T U571 ( .A1(n438), .A2(n508), .B1(instruction[6]), .B2(n501), 
        .C1(n512), .C2(offset_b[6]), .Z(n677) );
  AOI22D0BWP12T U572 ( .A1(instruction[8]), .A2(n440), .B1(instruction[9]), 
        .B2(n439), .ZN(n444) );
  AOI22D1BWP12T U573 ( .A1(instruction[2]), .A2(n442), .B1(instruction[3]), 
        .B2(n441), .ZN(n443) );
  OAI211D1BWP12T U574 ( .A1(n483), .A2(n445), .B(n444), .C(n443), .ZN(n446) );
  AO222D0BWP12T U575 ( .A1(n446), .A2(n508), .B1(instruction[4]), .B2(n501), 
        .C1(n512), .C2(offset_b[4]), .Z(n675) );
  AOI22D0BWP12T U576 ( .A1(n449), .A2(instruction[6]), .B1(n448), .B2(n447), 
        .ZN(n454) );
  OAI211D0BWP12T U577 ( .A1(n451), .A2(n488), .B(instruction[11]), .C(n450), 
        .ZN(n452) );
  ND4D1BWP12T U578 ( .A1(n455), .A2(n454), .A3(n453), .A4(n452), .ZN(n456) );
  AOI31D0BWP12T U579 ( .A1(n492), .A2(N910), .A3(next_step[1]), .B(n456), .ZN(
        n457) );
  MOAI22D0BWP12T U580 ( .A1(n457), .A2(n478), .B1(n512), .B2(alu_opcode[0]), 
        .ZN(n666) );
  MOAI22D0BWP12T U581 ( .A1(n488), .A2(n458), .B1(n512), .B2(
        memory_store_address_reg[1]), .ZN(n659) );
  AO21D0BWP12T U582 ( .A1(n512), .A2(memory_store_address_reg[4]), .B(n459), 
        .Z(n656) );
  MAOI22D0BWP12T U583 ( .A1(instruction[9]), .A2(n461), .B1(n460), .B2(n500), 
        .ZN(n467) );
  OAI31D0BWP12T U584 ( .A1(n465), .A2(n464), .A3(n463), .B(n462), .ZN(n466) );
  OAI211D1BWP12T U585 ( .A1(n469), .A2(n468), .B(n467), .C(n466), .ZN(n474) );
  AOI22D0BWP12T U586 ( .A1(n471), .A2(instruction[1]), .B1(n470), .B2(n474), 
        .ZN(n472) );
  MOAI22D0BWP12T U587 ( .A1(n472), .A2(n478), .B1(n512), .B2(
        memory_store_data_reg[1]), .ZN(n654) );
  AOI222D0BWP12T U588 ( .A1(n474), .A2(instruction[11]), .B1(instruction[1]), 
        .B2(n473), .C1(instruction[9]), .C2(n493), .ZN(n475) );
  MOAI22D0BWP12T U589 ( .A1(n475), .A2(n478), .B1(n512), .B2(
        memory_write_to_reg[1]), .ZN(n648) );
  OAI211D0BWP12T U590 ( .A1(n484), .A2(n488), .B(n498), .C(n476), .ZN(n477) );
  AOI21D0BWP12T U591 ( .A1(instruction[1]), .A2(n481), .B(n477), .ZN(n479) );
  MOAI22D0BWP12T U592 ( .A1(n479), .A2(n478), .B1(n512), .B2(
        alu_write_to_reg[1]), .ZN(n644) );
  AOI21D0BWP12T U593 ( .A1(instruction[2]), .A2(n481), .B(n480), .ZN(n482) );
  OAI32D0BWP12T U594 ( .A1(n485), .A2(n484), .A3(n483), .B1(n482), .B2(n485), 
        .ZN(n487) );
  AO211D0BWP12T U595 ( .A1(n512), .A2(alu_write_to_reg[2]), .B(n487), .C(n486), 
        .Z(n643) );
  OAI22D0BWP12T U596 ( .A1(instruction[11]), .A2(n490), .B1(n489), .B2(n488), 
        .ZN(n495) );
  OR3XD0BWP12T U597 ( .A1(n493), .A2(n492), .A3(n491), .Z(n494) );
  AOI211D0BWP12T U598 ( .A1(instruction[4]), .A2(n496), .B(n495), .C(n494), 
        .ZN(n497) );
  OAI211D0BWP12T U599 ( .A1(n500), .A2(n499), .B(n498), .C(n497), .ZN(n503) );
  AO222D0BWP12T U600 ( .A1(n503), .A2(n508), .B1(n512), .B2(operand_a[1]), 
        .C1(n502), .C2(n501), .Z(n638) );
  AO21D0BWP12T U601 ( .A1(n505), .A2(instruction[4]), .B(n504), .Z(n509) );
  AO222D0BWP12T U602 ( .A1(n509), .A2(n508), .B1(n507), .B2(n506), .C1(
        operand_b[1]), .C2(n512), .Z(n632) );
  AO21D0BWP12T U603 ( .A1(n512), .A2(operand_b[4]), .B(n510), .Z(n629) );
  IOA21D0BWP12T U604 ( .A1(n512), .A2(offset_b[23]), .B(n511), .ZN(n617) );
  IOA21D0BWP12T U605 ( .A1(n512), .A2(offset_b[24]), .B(n511), .ZN(n616) );
  IOA21D0BWP12T U606 ( .A1(n512), .A2(offset_b[25]), .B(n511), .ZN(n615) );
  IOA21D0BWP12T U607 ( .A1(n512), .A2(offset_b[26]), .B(n511), .ZN(n614) );
  IOA21D0BWP12T U608 ( .A1(n512), .A2(offset_b[27]), .B(n511), .ZN(n613) );
  IOA21D0BWP12T U609 ( .A1(n512), .A2(offset_b[28]), .B(n511), .ZN(n612) );
  IOA21D0BWP12T U610 ( .A1(n512), .A2(offset_b[29]), .B(n511), .ZN(n611) );
  IOA21D0BWP12T U611 ( .A1(n512), .A2(offset_b[30]), .B(n511), .ZN(n610) );
  IOA21D0BWP12T U612 ( .A1(n512), .A2(offset_b[31]), .B(n511), .ZN(n609) );
endmodule


module ALU_VARIABLE ( a, b, op, c_in, result, c_out, z, n, v );
  input [31:0] a;
  input [31:0] b;
  input [3:0] op;
  output [31:0] result;
  input c_in;
  output c_out, z, n, v;
  wire   n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168;
  tri   [31:0] a;
  tri   [31:0] b;
  tri   [31:0] result;

  OAI21D1BWP12T U3 ( .A1(b[0]), .A2(n4636), .B(n4128), .ZN(n3211) );
  OAI32D1BWP12T U4 ( .A1(n4313), .A2(n4671), .A3(n4670), .B1(n4343), .B2(n4313), .ZN(n4346) );
  OAI21D1BWP12T U5 ( .A1(a[6]), .A2(a[5]), .B(n5424), .ZN(n3286) );
  ND2D1BWP12T U6 ( .A1(b[1]), .A2(n5951), .ZN(n4009) );
  ND2D1BWP12T U7 ( .A1(n3211), .A2(n3212), .ZN(n4538) );
  ND2D1BWP12T U8 ( .A1(b[0]), .A2(a[16]), .ZN(n3488) );
  NR2D1BWP12T U9 ( .A1(n5964), .A2(b[0]), .ZN(n3483) );
  NR2D1BWP12T U10 ( .A1(b[0]), .A2(a[20]), .ZN(n4971) );
  ND2D1BWP12T U11 ( .A1(a[9]), .A2(n4344), .ZN(n4667) );
  OAI32D1BWP12T U12 ( .A1(n4694), .A2(a[28]), .A3(n5901), .B1(n5892), .B2(
        n4694), .ZN(n4695) );
  NR2D1BWP12T U13 ( .A1(a[11]), .A2(n5423), .ZN(n4640) );
  ND2D1BWP12T U14 ( .A1(a[11]), .A2(n4131), .ZN(n4636) );
  NR2D1BWP12T U15 ( .A1(a[5]), .A2(n5419), .ZN(n4645) );
  INVD1BWP12T U16 ( .I(n3301), .ZN(n4641) );
  INVD1BWP12T U17 ( .I(n3302), .ZN(n4642) );
  ND2D1BWP12T U18 ( .A1(b[0]), .A2(a[9]), .ZN(n3573) );
  OAI21D1BWP12T U19 ( .A1(a[4]), .A2(a[3]), .B(n5419), .ZN(n3307) );
  INVD1BWP12T U20 ( .I(n5380), .ZN(n4453) );
  INVD1BWP12T U21 ( .I(n5444), .ZN(n3358) );
  NR2D1BWP12T U22 ( .A1(a[3]), .A2(n3320), .ZN(n4661) );
  ND2D1BWP12T U23 ( .A1(b[0]), .A2(a[14]), .ZN(n3487) );
  FA1D0BWP12T U24 ( .A(n3293), .B(n3292), .CI(n3291), .CO(n3330), .S(n3294) );
  INVD1BWP12T U25 ( .I(n3450), .ZN(n5453) );
  RCIAO21D0BWP12T U26 ( .A1(n4631), .A2(b[0]), .B(n4634), .ZN(n3282) );
  FA1D0BWP12T U27 ( .A(n3274), .B(n3273), .CI(n3272), .CO(n3259), .S(n3327) );
  NR2D1BWP12T U28 ( .A1(n4699), .A2(a[8]), .ZN(n3450) );
  INVD1BWP12T U29 ( .I(n5442), .ZN(n3359) );
  FA1D0BWP12T U30 ( .A(n3276), .B(n3275), .CI(n3278), .CO(n3268), .S(n3326) );
  FA1D0BWP12T U31 ( .A(n3264), .B(n3263), .CI(n3262), .CO(n3243), .S(n3266) );
  INVD1BWP12T U32 ( .I(b[9]), .ZN(n4482) );
  ND2D1BWP12T U33 ( .A1(b[9]), .A2(n3509), .ZN(n5454) );
  FA1D0BWP12T U34 ( .A(n3261), .B(n3260), .CI(n3259), .CO(n3335), .S(n3267) );
  INVD1BWP12T U35 ( .I(n3424), .ZN(n3361) );
  FA1D0BWP12T U36 ( .A(n3249), .B(n3244), .CI(n3243), .CO(n3332), .S(n3337) );
  INVD1BWP12T U37 ( .I(n5395), .ZN(n3364) );
  FA1D0BWP12T U38 ( .A(n4539), .B(n4538), .CI(n4537), .CO(n4543), .S(n4547) );
  MAOI22D0BWP12T U39 ( .A1(b[1]), .A2(n3593), .B1(n3481), .B2(b[1]), .ZN(n3537) );
  ND2D1BWP12T U40 ( .A1(b[3]), .A2(b[2]), .ZN(n3627) );
  INVD1BWP12T U41 ( .I(a[8]), .ZN(n3360) );
  MOAI22D0BWP12T U42 ( .A1(n3572), .A2(n5256), .B1(n3493), .B2(n3492), .ZN(
        n5241) );
  ND2D1BWP12T U43 ( .A1(b[0]), .A2(a[26]), .ZN(n3761) );
  NR2D1BWP12T U44 ( .A1(b[0]), .A2(a[24]), .ZN(n3400) );
  NR2D1BWP12T U45 ( .A1(b[2]), .A2(n5237), .ZN(n3497) );
  NR2D1BWP12T U46 ( .A1(b[1]), .A2(n5593), .ZN(n4603) );
  ND2D1BWP12T U47 ( .A1(b[2]), .A2(a[31]), .ZN(n4599) );
  INVD1BWP12T U48 ( .I(n3430), .ZN(n3482) );
  ND2D1BWP12T U49 ( .A1(b[0]), .A2(a[20]), .ZN(n4956) );
  ND2D1BWP12T U50 ( .A1(b[0]), .A2(a[29]), .ZN(n3817) );
  INVD1BWP12T U51 ( .I(b[1]), .ZN(n4419) );
  INVD1BWP12T U52 ( .I(n3455), .ZN(n5122) );
  INVD1BWP12T U53 ( .I(n5191), .ZN(n5123) );
  INVD1BWP12T U54 ( .I(n3567), .ZN(n3565) );
  INVD1BWP12T U55 ( .I(a[30]), .ZN(n4738) );
  INVD1BWP12T U56 ( .I(n5086), .ZN(n3572) );
  NR2D1BWP12T U57 ( .A1(n3430), .A2(n3485), .ZN(n5086) );
  INVD1BWP12T U58 ( .I(n4974), .ZN(n5181) );
  INVD1BWP12T U59 ( .I(n5085), .ZN(n5178) );
  INVD1BWP12T U60 ( .I(n3382), .ZN(n5250) );
  INVD1BWP12T U61 ( .I(n3536), .ZN(n5177) );
  INVD1BWP12T U62 ( .I(b[17]), .ZN(n4838) );
  ND2D1BWP12T U63 ( .A1(a[6]), .A2(a[5]), .ZN(n5424) );
  ND2D1BWP12T U64 ( .A1(a[4]), .A2(a[3]), .ZN(n5419) );
  NR2D1BWP12T U65 ( .A1(b[2]), .A2(n5421), .ZN(n5439) );
  NR2D1BWP12T U66 ( .A1(b[6]), .A2(n3577), .ZN(n5438) );
  NR2D1BWP12T U67 ( .A1(n4555), .A2(a[6]), .ZN(n5458) );
  ND2D1BWP12T U68 ( .A1(n5379), .A2(a[0]), .ZN(n5436) );
  NR2D1BWP12T U69 ( .A1(b[0]), .A2(b[1]), .ZN(n3430) );
  INVD1BWP12T U70 ( .I(n5246), .ZN(n5099) );
  OAI21D1BWP12T U71 ( .A1(n4759), .A2(n5799), .B(n5436), .ZN(n4758) );
  INVD1BWP12T U72 ( .I(b[0]), .ZN(n5379) );
  NR2D1BWP12T U73 ( .A1(n5471), .A2(n5439), .ZN(n3632) );
  IND2D1BWP12T U74 ( .A1(n5467), .B1(n3321), .ZN(n3639) );
  AOI211D1BWP12T U75 ( .A1(n3630), .A2(n5240), .B(n3629), .C(n3628), .ZN(n5495) );
  INVD1BWP12T U76 ( .I(n3632), .ZN(n3640) );
  NR2D1BWP12T U77 ( .A1(n3645), .A2(b[4]), .ZN(n3653) );
  INVD1BWP12T U78 ( .I(n3723), .ZN(n3691) );
  NR2D1BWP12T U79 ( .A1(a[2]), .A2(a[1]), .ZN(n3341) );
  NR2D1BWP12T U80 ( .A1(n5472), .A2(n5440), .ZN(n3723) );
  INVD1BWP12T U81 ( .I(a[3]), .ZN(n3363) );
  OAI211D1BWP12T U82 ( .A1(b[3]), .A2(n3718), .B(n3717), .C(n3716), .ZN(n3721)
         );
  AOI21D1BWP12T U83 ( .A1(n5238), .A2(n3713), .B(b[4]), .ZN(n3717) );
  IND2D1BWP12T U84 ( .A1(n5094), .B1(n3710), .ZN(n3712) );
  ND2D1BWP12T U85 ( .A1(n3324), .A2(n3323), .ZN(n3670) );
  INVD1BWP12T U86 ( .I(n3674), .ZN(n3675) );
  INVD1BWP12T U87 ( .I(n3682), .ZN(n3685) );
  AOI211D1BWP12T U88 ( .A1(n3430), .A2(a[12]), .B(n5211), .C(n3206), .ZN(n3664) );
  ND2D1BWP12T U89 ( .A1(b[0]), .A2(a[15]), .ZN(n3205) );
  AOI21D1BWP12T U90 ( .A1(n3709), .A2(b[4]), .B(n3358), .ZN(n3682) );
  ND2D1BWP12T U91 ( .A1(n5638), .A2(n5052), .ZN(n3346) );
  INVD1BWP12T U92 ( .I(a[5]), .ZN(n3300) );
  INVD1BWP12T U93 ( .I(b[5]), .ZN(n4490) );
  NR2D1BWP12T U94 ( .A1(n5459), .A2(n5447), .ZN(n3622) );
  OAI211D1BWP12T U95 ( .A1(n3707), .A2(n3599), .B(n3598), .C(n3597), .ZN(n3615) );
  INVD1BWP12T U96 ( .I(n5100), .ZN(n3599) );
  AOI21D1BWP12T U97 ( .A1(n5240), .A2(n5099), .B(b[4]), .ZN(n3598) );
  INVD1BWP12T U98 ( .I(n3622), .ZN(n3620) );
  INVD1BWP12T U99 ( .I(n3535), .ZN(n3608) );
  INVD1BWP12T U100 ( .I(n3534), .ZN(n3609) );
  FA1D0BWP12T U101 ( .A(n3312), .B(n3311), .CI(n3310), .CO(n3306), .S(n3313)
         );
  OA21D1BWP12T U102 ( .A1(n3299), .A2(n3298), .B(n3297), .Z(n3312) );
  NR2D1BWP12T U103 ( .A1(n3482), .A2(b[2]), .ZN(n3569) );
  AN2D1BWP12T U104 ( .A1(n3592), .A2(n3607), .Z(n3588) );
  INVD1BWP12T U105 ( .I(n4493), .ZN(n3589) );
  OAI22D1BWP12T U106 ( .A1(n5394), .A2(n3588), .B1(a[6]), .B2(b[6]), .ZN(n3548) );
  INVD1BWP12T U107 ( .I(b[7]), .ZN(n4450) );
  INVD1BWP12T U108 ( .I(n3521), .ZN(n3522) );
  INVD1BWP12T U109 ( .I(n4495), .ZN(n3549) );
  AOI22D1BWP12T U110 ( .A1(b[0]), .A2(a[2]), .B1(a[3]), .B2(n5379), .ZN(n3610)
         );
  ND2D1BWP12T U111 ( .A1(n5210), .A2(b[1]), .ZN(n5128) );
  INVD1BWP12T U112 ( .I(b[8]), .ZN(n4699) );
  NR2D1BWP12T U113 ( .A1(n3548), .A2(n3533), .ZN(n3449) );
  ND2D1BWP12T U114 ( .A1(n5452), .A2(n3522), .ZN(n3472) );
  ND2D1BWP12T U115 ( .A1(n5453), .A2(n3466), .ZN(n3473) );
  OAI211D1BWP12T U116 ( .A1(n3664), .A2(n3707), .B(n3454), .C(n3453), .ZN(
        n5513) );
  AOI21D1BWP12T U117 ( .A1(n5240), .A2(n5106), .B(b[4]), .ZN(n3454) );
  FA1D0BWP12T U118 ( .A(n3328), .B(n3327), .CI(n3326), .CO(n3277), .S(n3329)
         );
  RCIAO21D0BWP12T U119 ( .A1(n5393), .A2(n3449), .B(n3457), .ZN(n3478) );
  INVD1BWP12T U120 ( .I(n3498), .ZN(n5500) );
  INVD1BWP12T U121 ( .I(n5816), .ZN(n5010) );
  OAI211D1BWP12T U122 ( .A1(n3594), .A2(n3627), .B(n3495), .C(n3494), .ZN(
        n3498) );
  AOI21D1BWP12T U123 ( .A1(n5242), .A2(n5099), .B(b[4]), .ZN(n3495) );
  AOI22D1BWP12T U124 ( .A1(n3360), .A2(b[8]), .B1(n3472), .B2(n3359), .ZN(
        n3518) );
  ND2D1BWP12T U125 ( .A1(n3435), .A2(n5454), .ZN(n4343) );
  FA1D0BWP12T U126 ( .A(n3268), .B(n3267), .CI(n3266), .CO(n3265), .S(n3269)
         );
  INVD1BWP12T U127 ( .I(b[10]), .ZN(n4646) );
  ND2D1BWP12T U128 ( .A1(n4482), .A2(a[9]), .ZN(n3435) );
  AOI211D1BWP12T U129 ( .A1(n3430), .A2(a[14]), .B(n5144), .C(n3406), .ZN(
        n5118) );
  INVD1BWP12T U130 ( .I(n3443), .ZN(n3444) );
  ND2D1BWP12T U131 ( .A1(n3424), .A2(n5455), .ZN(n3446) );
  INVD1BWP12T U132 ( .I(n5521), .ZN(n3496) );
  FA1D0BWP12T U133 ( .A(n3337), .B(n3336), .CI(n3335), .CO(n3376), .S(n3254)
         );
  ND2D1BWP12T U134 ( .A1(n3420), .A2(n3444), .ZN(n3394) );
  NR2D1BWP12T U135 ( .A1(b[3]), .A2(n5030), .ZN(n5015) );
  FA1D0BWP12T U136 ( .A(n3334), .B(n3333), .CI(n3332), .CO(n4551), .S(n3377)
         );
  INVD1BWP12T U137 ( .I(a[12]), .ZN(n4791) );
  AOI21D1BWP12T U138 ( .A1(n3364), .A2(n3368), .B(n3378), .ZN(n4836) );
  NR2D1BWP12T U139 ( .A1(n3749), .A2(b[11]), .ZN(n3357) );
  INVD1BWP12T U140 ( .I(n3393), .ZN(n4148) );
  MOAI22D0BWP12T U141 ( .A1(b[11]), .A2(a[11]), .B1(n3394), .B2(n3364), .ZN(
        n4790) );
  OAI211D1BWP12T U142 ( .A1(n5122), .A2(n5286), .B(n3348), .C(n3347), .ZN(
        n5206) );
  ND2D1BWP12T U143 ( .A1(n4744), .A2(n4742), .ZN(n3365) );
  INVD1BWP12T U144 ( .I(n4745), .ZN(n3392) );
  NR2D1BWP12T U145 ( .A1(n3357), .A2(n3191), .ZN(n3393) );
  NR2D1BWP12T U146 ( .A1(a[11]), .A2(n4741), .ZN(n3191) );
  FA1D0BWP12T U147 ( .A(n4548), .B(n4547), .CI(n4546), .CO(n5360), .S(n4550)
         );
  ND2D1BWP12T U148 ( .A1(n5541), .A2(b[4]), .ZN(n5521) );
  INVD1BWP12T U149 ( .I(b[14]), .ZN(n5390) );
  MAOI22D0BWP12T U150 ( .A1(b[2]), .A2(n3537), .B1(n3708), .B2(b[2]), .ZN(
        n5078) );
  ND2D1BWP12T U151 ( .A1(n5570), .A2(n5770), .ZN(n5070) );
  OAI22D1BWP12T U152 ( .A1(n4419), .A2(n3398), .B1(n3401), .B2(b[1]), .ZN(
        n5105) );
  INVD1BWP12T U153 ( .I(n3627), .ZN(n5238) );
  ND2D1BWP12T U154 ( .A1(n4983), .A2(b[3]), .ZN(n5171) );
  NR2D1BWP12T U155 ( .A1(n3572), .A2(n5159), .ZN(n5211) );
  INVD1BWP12T U156 ( .I(n3564), .ZN(n3566) );
  AOI22D1BWP12T U157 ( .A1(b[0]), .A2(a[1]), .B1(a[2]), .B2(n5379), .ZN(n3563)
         );
  ND2D1BWP12T U158 ( .A1(n3414), .A2(n3413), .ZN(n5026) );
  MOAI22D0BWP12T U159 ( .A1(n5131), .A2(n3563), .B1(a[0]), .B2(n5098), .ZN(
        n5028) );
  ND2D1BWP12T U160 ( .A1(n3418), .A2(n3417), .ZN(n5202) );
  INVD1BWP12T U161 ( .I(n3538), .ZN(n3706) );
  AOI32D1BWP12T U162 ( .A1(n5220), .A2(n3761), .A3(n4008), .B1(n3480), .B2(
        n5220), .ZN(n3708) );
  AOI211D1BWP12T U163 ( .A1(n5254), .A2(n5178), .B(n3370), .C(n3369), .ZN(
        n5173) );
  INVD1BWP12T U164 ( .I(n3663), .ZN(n5240) );
  AOI21D1BWP12T U165 ( .A1(n5240), .A2(n5117), .B(n5273), .ZN(n5538) );
  INVD1BWP12T U166 ( .I(n5705), .ZN(n5201) );
  ND2D1BWP12T U167 ( .A1(n5632), .A2(b[4]), .ZN(n5204) );
  INVD1BWP12T U168 ( .I(n3707), .ZN(n5242) );
  ND2D1BWP12T U169 ( .A1(n5638), .A2(n5057), .ZN(n5062) );
  ND2D1BWP12T U170 ( .A1(a[0]), .A2(b[3]), .ZN(n5198) );
  ND2D1BWP12T U171 ( .A1(n4419), .A2(b[2]), .ZN(n5047) );
  INVD1BWP12T U172 ( .I(n5150), .ZN(n5256) );
  NR2D1BWP12T U173 ( .A1(b[2]), .A2(n3571), .ZN(n3431) );
  AOI22D1BWP12T U174 ( .A1(b[0]), .A2(n4603), .B1(a[30]), .B2(n3430), .ZN(
        n5277) );
  ND2D1BWP12T U175 ( .A1(b[3]), .A2(a[31]), .ZN(n5541) );
  INVD1BWP12T U176 ( .I(n5284), .ZN(n5255) );
  ND2D1BWP12T U177 ( .A1(n4599), .A2(n3383), .ZN(n3705) );
  ND2D1BWP12T U178 ( .A1(n3482), .A2(b[2]), .ZN(n5143) );
  INVD1BWP12T U179 ( .I(b[3]), .ZN(n5136) );
  INVD1BWP12T U180 ( .I(n5286), .ZN(n5192) );
  NR2D1BWP12T U181 ( .A1(n3572), .A2(n5143), .ZN(n5254) );
  NR2D1BWP12T U182 ( .A1(n5703), .A2(n5705), .ZN(n5258) );
  INVD1BWP12T U183 ( .I(n5204), .ZN(n5168) );
  ND2D1BWP12T U184 ( .A1(b[2]), .A2(b[1]), .ZN(n5045) );
  ND2D1BWP12T U185 ( .A1(n3201), .A2(n3200), .ZN(n4997) );
  INVD1BWP12T U186 ( .I(n5262), .ZN(n5288) );
  NR2D1BWP12T U187 ( .A1(n4995), .A2(n3569), .ZN(n5290) );
  INVD1BWP12T U188 ( .I(n5131), .ZN(n5057) );
  NR2D1BWP12T U189 ( .A1(b[3]), .A2(b[2]), .ZN(n5525) );
  AOI222D1BWP12T U190 ( .A1(n3646), .A2(n3568), .B1(n5262), .B2(n3567), .C1(
        n3566), .C2(n5254), .ZN(n5146) );
  ND2D1BWP12T U191 ( .A1(a[31]), .A2(n5826), .ZN(n5669) );
  ND2D1BWP12T U192 ( .A1(n3572), .A2(n3568), .ZN(n5286) );
  NR2D1BWP12T U193 ( .A1(n5086), .A2(n3568), .ZN(n5262) );
  INVD1BWP12T U194 ( .I(n5254), .ZN(n5282) );
  INVD1BWP12T U195 ( .I(n5258), .ZN(n5280) );
  INVD1BWP12T U196 ( .I(n5290), .ZN(n5263) );
  NR2D1BWP12T U197 ( .A1(n5136), .A2(b[4]), .ZN(n5079) );
  INVD1BWP12T U198 ( .I(n5045), .ZN(n5051) );
  INVD1BWP12T U199 ( .I(n5047), .ZN(n5052) );
  INVD1BWP12T U200 ( .I(n5128), .ZN(n5095) );
  INVD1BWP12T U201 ( .I(n5145), .ZN(n4995) );
  ND4D1BWP12T U202 ( .A1(n3199), .A2(n3198), .A3(n3197), .A4(n3196), .ZN(n5528) );
  NR4D0BWP12T U203 ( .A1(b[27]), .A2(b[26]), .A3(b[16]), .A4(b[31]), .ZN(n3199) );
  NR4D0BWP12T U204 ( .A1(b[30]), .A2(b[20]), .A3(b[19]), .A4(b[11]), .ZN(n3198) );
  NR4D0BWP12T U205 ( .A1(b[22]), .A2(b[21]), .A3(b[18]), .A4(b[15]), .ZN(n3197) );
  NR4D0BWP12T U206 ( .A1(b[28]), .A2(b[25]), .A3(b[23]), .A4(b[13]), .ZN(n3193) );
  NR4D0BWP12T U207 ( .A1(b[10]), .A2(b[9]), .A3(b[6]), .A4(b[5]), .ZN(n3192)
         );
  OR2XD1BWP12T U208 ( .A1(op[0]), .A2(n5622), .Z(n3356) );
  ND2D1BWP12T U209 ( .A1(op[0]), .A2(n5622), .ZN(n3343) );
  ND2D1BWP12T U210 ( .A1(n3202), .A2(op[2]), .ZN(n3355) );
  ND2D1BWP12T U211 ( .A1(op[0]), .A2(op[1]), .ZN(n3362) );
  INVD1BWP12T U212 ( .I(n5528), .ZN(n5570) );
  ND2D1BWP12T U213 ( .A1(n3430), .A2(n5525), .ZN(n5632) );
  INVD1BWP12T U214 ( .I(n5492), .ZN(n5634) );
  ND2D1BWP12T U215 ( .A1(op[3]), .A2(n5594), .ZN(n5623) );
  INVD1BWP12T U216 ( .I(a[0]), .ZN(n5633) );
  NR2D1BWP12T U217 ( .A1(b[1]), .A2(a[1]), .ZN(n5807) );
  NR2D1BWP12T U218 ( .A1(n5383), .A2(n5807), .ZN(n5797) );
  ND2D1BWP12T U219 ( .A1(b[1]), .A2(a[1]), .ZN(n5806) );
  NR2D1BWP12T U220 ( .A1(n5805), .A2(b[1]), .ZN(n5804) );
  NR2D1BWP12T U221 ( .A1(n5379), .A2(a[0]), .ZN(n5799) );
  INVD1BWP12T U222 ( .I(n5797), .ZN(n5798) );
  INVD1BWP12T U223 ( .I(a[1]), .ZN(n5805) );
  INVD1BWP12T U224 ( .I(n3429), .ZN(n5830) );
  NR2D1BWP12T U225 ( .A1(n5210), .A2(a[2]), .ZN(n5471) );
  INVD1BWP12T U226 ( .I(n5495), .ZN(n3645) );
  NR2D1BWP12T U227 ( .A1(n3653), .A2(n6009), .ZN(n5494) );
  NR2D1BWP12T U228 ( .A1(n5421), .A2(n5210), .ZN(n5384) );
  NR2D1BWP12T U229 ( .A1(n5528), .A2(b[4]), .ZN(n5670) );
  OAI21D1BWP12T U230 ( .A1(n3634), .A2(n3633), .B(n3699), .ZN(n5410) );
  INVD1BWP12T U231 ( .I(a[2]), .ZN(n5421) );
  INVD1BWP12T U232 ( .I(b[2]), .ZN(n5210) );
  NR2D1BWP12T U233 ( .A1(n5136), .A2(a[3]), .ZN(n5472) );
  NR2D1BWP12T U234 ( .A1(b[3]), .A2(n3363), .ZN(n5440) );
  ND2D1BWP12T U235 ( .A1(n3341), .A2(n5633), .ZN(n3698) );
  OAI22D1BWP12T U236 ( .A1(n3609), .A2(n5128), .B1(n3610), .B2(n5131), .ZN(
        n5032) );
  OAI22D1BWP12T U237 ( .A1(n3610), .A2(n5288), .B1(n3609), .B2(n5282), .ZN(
        n5172) );
  AOI211D1BWP12T U238 ( .A1(b[4]), .A2(n5996), .B(n3719), .C(n5528), .ZN(n5549) );
  NR2D1BWP12T U239 ( .A1(n3363), .A2(n5136), .ZN(n5385) );
  OAI21D1BWP12T U240 ( .A1(n5110), .A2(n5703), .B(n3721), .ZN(n5082) );
  FA1D0BWP12T U241 ( .A(n3670), .B(n3669), .CI(n3668), .CO(n3602), .S(n5310)
         );
  ND2D1BWP12T U242 ( .A1(n5703), .A2(a[4]), .ZN(n5444) );
  NR2D1BWP12T U243 ( .A1(a[3]), .A2(n3698), .ZN(n3697) );
  INVD1BWP12T U244 ( .I(n5536), .ZN(n3666) );
  ND2D1BWP12T U245 ( .A1(b[4]), .A2(a[4]), .ZN(n5386) );
  INVD1BWP12T U246 ( .I(a[4]), .ZN(n3709) );
  ND2D1BWP12T U247 ( .A1(n3300), .A2(n4490), .ZN(n3607) );
  NR2D1BWP12T U248 ( .A1(b[5]), .A2(n3300), .ZN(n5447) );
  MAOI22D0BWP12T U249 ( .A1(n3622), .A2(n3621), .B1(n3622), .B2(n3621), .ZN(
        n4867) );
  NR2D1BWP12T U250 ( .A1(n3300), .A2(n4490), .ZN(n3600) );
  OAI21D1BWP12T U251 ( .A1(n5971), .A2(n5703), .B(n3615), .ZN(n5271) );
  OA21D1BWP12T U252 ( .A1(n5703), .A2(n5972), .B(n3615), .Z(n5551) );
  OAI222D1BWP12T U253 ( .A1(n3608), .A2(n5288), .B1(n3609), .B2(n5286), .C1(
        n3610), .C2(n5282), .ZN(n5281) );
  OAI222D1BWP12T U254 ( .A1(n5128), .A2(n3610), .B1(n5047), .B2(n3609), .C1(
        n5131), .C2(n3608), .ZN(n5036) );
  NR2D1BWP12T U255 ( .A1(n3569), .A2(n5541), .ZN(n5539) );
  INVD1BWP12T U256 ( .I(n5116), .ZN(n3583) );
  ND2D1BWP12T U257 ( .A1(b[4]), .A2(n5538), .ZN(n3584) );
  ND2D1BWP12T U258 ( .A1(n3584), .A2(n3583), .ZN(n5511) );
  INVD1BWP12T U259 ( .I(n5067), .ZN(n5008) );
  INVD1BWP12T U260 ( .I(b[6]), .ZN(n4555) );
  INVD1BWP12T U261 ( .I(a[6]), .ZN(n3577) );
  NR2D1BWP12T U262 ( .A1(a[7]), .A2(b[7]), .ZN(n3533) );
  ND2D1BWP12T U263 ( .A1(n3528), .A2(b[7]), .ZN(n5452) );
  MAOI22D0BWP12T U264 ( .A1(n3550), .A2(n3549), .B1(n3550), .B2(n3549), .ZN(
        n4866) );
  NR2D1BWP12T U265 ( .A1(n3528), .A2(n4450), .ZN(n3526) );
  ND2D1BWP12T U266 ( .A1(a[7]), .A2(n4450), .ZN(n3525) );
  INVD1BWP12T U267 ( .I(a[7]), .ZN(n3528) );
  INVD1BWP12T U268 ( .I(b[4]), .ZN(n5703) );
  NR2D1BWP12T U269 ( .A1(n5070), .A2(n6138), .ZN(n5817) );
  NR2D1BWP12T U270 ( .A1(a[8]), .A2(b[8]), .ZN(n3457) );
  ND2D1BWP12T U271 ( .A1(a[8]), .A2(n4699), .ZN(n3466) );
  MAOI22D0BWP12T U272 ( .A1(n3475), .A2(n3474), .B1(n3475), .B2(n3474), .ZN(
        n4872) );
  ND2D1BWP12T U273 ( .A1(a[8]), .A2(b[8]), .ZN(n3458) );
  INVD1BWP12T U274 ( .I(n5513), .ZN(n3469) );
  OAI222D1BWP12T U275 ( .A1(n5062), .A2(n4995), .B1(n3469), .B2(n5925), .C1(
        n5263), .C2(n5706), .ZN(n5219) );
  INVD1BWP12T U276 ( .I(n3435), .ZN(n3503) );
  MOAI22D0BWP12T U277 ( .A1(n4211), .A2(n3517), .B1(n4211), .B2(n3517), .ZN(
        n4871) );
  MAOI22D0BWP12T U278 ( .A1(n3479), .A2(n4343), .B1(n3479), .B2(n4343), .ZN(
        n4924) );
  OAI22D1BWP12T U279 ( .A1(n5136), .A2(n5010), .B1(n5066), .B2(b[3]), .ZN(
        n5021) );
  OAI21D1BWP12T U280 ( .A1(n5845), .A2(n5703), .B(n3498), .ZN(n3499) );
  ND2D1BWP12T U281 ( .A1(b[9]), .A2(a[9]), .ZN(n5387) );
  MAOI22D0BWP12T U282 ( .A1(n3518), .A2(n4343), .B1(n3518), .B2(n4343), .ZN(
        n4770) );
  NR2D1BWP12T U283 ( .A1(n3576), .A2(n3342), .ZN(n3510) );
  INVD1BWP12T U284 ( .I(n4343), .ZN(n4211) );
  INVD1BWP12T U285 ( .I(a[9]), .ZN(n3509) );
  ND2D1BWP12T U286 ( .A1(n4646), .A2(n3421), .ZN(n3420) );
  ND2D1BWP12T U287 ( .A1(n4646), .A2(a[10]), .ZN(n3424) );
  ND2D1BWP12T U288 ( .A1(b[10]), .A2(a[10]), .ZN(n3423) );
  MAOI22D0BWP12T U289 ( .A1(n3446), .A2(n3445), .B1(n3446), .B2(n3445), .ZN(
        n4874) );
  OAI21D1BWP12T U290 ( .A1(n5136), .A2(n3650), .B(n3412), .ZN(n5113) );
  MOAI22D0BWP12T U291 ( .A1(n5705), .A2(n5200), .B1(n5202), .B2(n5705), .ZN(
        n5084) );
  ND2D1BWP12T U292 ( .A1(n5769), .A2(n5136), .ZN(n5498) );
  AOI21D1BWP12T U293 ( .A1(b[4]), .A2(n5498), .B(n3432), .ZN(n5507) );
  AOI32D1BWP12T U294 ( .A1(n3496), .A2(n3433), .A3(n5540), .B1(n3432), .B2(
        n3433), .ZN(n5557) );
  ND2D1BWP12T U295 ( .A1(n6092), .A2(n6096), .ZN(n3693) );
  INVD1BWP12T U296 ( .I(a[10]), .ZN(n3421) );
  ND2D1BWP12T U297 ( .A1(n3510), .A2(n3509), .ZN(n3508) );
  NR2D1BWP12T U298 ( .A1(n3343), .A2(n3504), .ZN(n5374) );
  NR2D1BWP12T U299 ( .A1(b[4]), .A2(n6115), .ZN(n5815) );
  NR2D1BWP12T U300 ( .A1(n3362), .A2(n3344), .ZN(n3429) );
  INVD1BWP12T U301 ( .I(n4058), .ZN(n3378) );
  ND2D1BWP12T U302 ( .A1(b[11]), .A2(a[11]), .ZN(n4057) );
  INVD1BWP12T U303 ( .I(n3357), .ZN(n4743) );
  AOI21D1BWP12T U304 ( .A1(b[3]), .A2(n5032), .B(n5015), .ZN(n4980) );
  AOI22D1BWP12T U305 ( .A1(n5201), .A2(n5172), .B1(n5173), .B2(n5705), .ZN(
        n5147) );
  IOA21D1BWP12T U306 ( .A1(n5757), .A2(b[4]), .B(n3384), .ZN(n5083) );
  NR2D1BWP12T U307 ( .A1(a[10]), .A2(n3508), .ZN(n3410) );
  NR2D1BWP12T U308 ( .A1(n3355), .A2(n5592), .ZN(n5826) );
  INVD1BWP12T U309 ( .I(b[11]), .ZN(n4741) );
  INVD1BWP12T U310 ( .I(a[11]), .ZN(n3749) );
  NR2D1BWP12T U311 ( .A1(n6145), .A2(n5870), .ZN(n5600) );
  FA1D0BWP12T U312 ( .A(n4551), .B(n4550), .CI(n4549), .CO(n5359), .S(n5368)
         );
  ND2D1BWP12T U313 ( .A1(a[12]), .A2(n4792), .ZN(n4742) );
  ND2D1BWP12T U314 ( .A1(b[12]), .A2(n4791), .ZN(n4744) );
  MAOI22D0BWP12T U315 ( .A1(n3365), .A2(n4836), .B1(n3365), .B2(n4836), .ZN(
        n4875) );
  AO21D1BWP12T U316 ( .A1(n5723), .A2(b[4]), .B(n3349), .Z(n5272) );
  AOI31D1BWP12T U317 ( .A1(b[4]), .A2(n5723), .A3(n5532), .B(n3349), .ZN(n5516) );
  MAOI22D0BWP12T U318 ( .A1(n3365), .A2(n4790), .B1(n3365), .B2(n4790), .ZN(
        n4826) );
  AOI22D1BWP12T U319 ( .A1(n5258), .A2(n5227), .B1(n5290), .B2(n5206), .ZN(
        n5092) );
  MAOI22D0BWP12T U320 ( .A1(n4982), .A2(n5014), .B1(n5070), .B2(n4997), .ZN(
        n4999) );
  INVD1BWP12T U321 ( .I(b[12]), .ZN(n4792) );
  ND2D1BWP12T U322 ( .A1(n3410), .A2(n3749), .ZN(n3727) );
  NR2D1BWP12T U323 ( .A1(n5528), .A2(n5866), .ZN(n5621) );
  INVD1BWP12T U324 ( .I(n5859), .ZN(n5635) );
  INVD1BWP12T U325 ( .I(n5600), .ZN(n5620) );
  NR2D1BWP12T U326 ( .A1(n5570), .A2(n5669), .ZN(n5859) );
  INVD1BWP12T U327 ( .I(n5826), .ZN(n5866) );
  INVD1BWP12T U328 ( .I(a[13]), .ZN(n5872) );
  NR2D1BWP12T U329 ( .A1(n5889), .A2(n6135), .ZN(n6048) );
  ND2D1BWP12T U330 ( .A1(n5632), .A2(n5171), .ZN(n5705) );
  NR2D1BWP12T U331 ( .A1(n5263), .A2(n6115), .ZN(n5698) );
  INVD1BWP12T U332 ( .I(a[17]), .ZN(n5679) );
  OAI21D1BWP12T U333 ( .A1(n5769), .A2(n5136), .B(n3651), .ZN(n6009) );
  MAOI22D0BWP12T U334 ( .A1(n5240), .A2(n5278), .B1(b[3]), .B2(n3658), .ZN(
        n6071) );
  NR2D1BWP12T U335 ( .A1(n3362), .A2(n3504), .ZN(n6074) );
  OAI21D1BWP12T U336 ( .A1(n5274), .A2(n3663), .B(n3614), .ZN(n5971) );
  INVD1BWP12T U337 ( .I(a[21]), .ZN(n5964) );
  OAI21D1BWP12T U338 ( .A1(n4983), .A2(n5541), .B(n3541), .ZN(n5937) );
  INVD1BWP12T U339 ( .I(a[23]), .ZN(n5951) );
  INVD1BWP12T U340 ( .I(a[22]), .ZN(n6155) );
  AOI22D1BWP12T U341 ( .A1(n5525), .A2(n5104), .B1(n5242), .B2(n5278), .ZN(
        n5925) );
  INVD1BWP12T U342 ( .I(a[24]), .ZN(n5912) );
  NR2D1BWP12T U343 ( .A1(b[3]), .A2(n5138), .ZN(n5845) );
  NR2D1BWP12T U344 ( .A1(n3356), .A2(n3344), .ZN(n6052) );
  INVD1BWP12T U345 ( .I(a[25]), .ZN(n5833) );
  INVD1BWP12T U346 ( .I(n6048), .ZN(n6133) );
  AOI21D1BWP12T U347 ( .A1(n5277), .A2(b[2]), .B(n3431), .ZN(n5769) );
  NR2D1BWP12T U348 ( .A1(b[4]), .A2(b[3]), .ZN(n5770) );
  NR2D1BWP12T U349 ( .A1(n5528), .A2(n5830), .ZN(n5870) );
  INVD1BWP12T U350 ( .I(a[26]), .ZN(n5787) );
  INVD1BWP12T U351 ( .I(a[27]), .ZN(n5758) );
  NR2D1BWP12T U352 ( .A1(n3343), .A2(n3344), .ZN(n6135) );
  NR2D1BWP12T U353 ( .A1(n3504), .A2(n5592), .ZN(n6150) );
  INVD1BWP12T U354 ( .I(a[29]), .ZN(n5901) );
  INVD1BWP12T U355 ( .I(n5146), .ZN(n6111) );
  NR2D1BWP12T U356 ( .A1(n5623), .A2(n3343), .ZN(n6151) );
  INVD1BWP12T U357 ( .I(n6045), .ZN(n6128) );
  INVD1BWP12T U358 ( .I(n6150), .ZN(n6092) );
  INVD1BWP12T U359 ( .I(n6145), .ZN(n6115) );
  INVD1BWP12T U360 ( .I(n6160), .ZN(n6113) );
  NR2D1BWP12T U361 ( .A1(n3356), .A2(n3355), .ZN(n6122) );
  INVD1BWP12T U362 ( .I(n6164), .ZN(n6120) );
  INVD1BWP12T U363 ( .I(n6162), .ZN(n6126) );
  OR2XD1BWP12T U364 ( .A1(op[0]), .A2(op[1]), .Z(n5592) );
  INVD1BWP12T U365 ( .I(a[31]), .ZN(n5593) );
  INVD1BWP12T U366 ( .I(n6135), .ZN(n6096) );
  NR2D1BWP12T U367 ( .A1(n3362), .A2(n3355), .ZN(n6145) );
  INVD1BWP12T U368 ( .I(n5090), .ZN(n5608) );
  INVD1BWP12T U369 ( .I(op[1]), .ZN(n5622) );
  INVD1BWP12T U370 ( .I(n5374), .ZN(n6130) );
  INVD1BWP12T U371 ( .I(n6074), .ZN(n6156) );
  INVD1BWP12T U372 ( .I(n6151), .ZN(n6034) );
  INVD1BWP12T U373 ( .I(n6052), .ZN(n6138) );
  NR2D1BWP12T U374 ( .A1(n5623), .A2(n3356), .ZN(n6160) );
  NR2D1BWP12T U375 ( .A1(n3355), .A2(n3343), .ZN(n6164) );
  NR2D1BWP12T U376 ( .A1(n5623), .A2(n3362), .ZN(n6162) );
  INVD1BWP12T U377 ( .I(n6122), .ZN(n6167) );
  OAI32D1BWP12T U378 ( .A1(n5613), .A2(b[31]), .A3(a[31]), .B1(n5587), .B2(
        n5613), .ZN(n5589) );
  ND2D1BWP12T U379 ( .A1(a[2]), .A2(n5808), .ZN(n3642) );
  AOI211D1BWP12T U380 ( .A1(n5698), .A2(n5172), .B(n3704), .C(n3703), .ZN(
        n3726) );
  OAI22D1BWP12T U381 ( .A1(n5600), .A2(n5082), .B1(n4761), .B2(n6167), .ZN(
        n3724) );
  ND2D1BWP12T U382 ( .A1(n5817), .A2(n5014), .ZN(n3678) );
  MOAI22D0BWP12T U383 ( .A1(n5600), .A2(n5271), .B1(n6160), .B2(n4922), .ZN(
        n3617) );
  AOI22D1BWP12T U384 ( .A1(n5698), .A2(n5281), .B1(n5817), .B2(n5036), .ZN(
        n3611) );
  NR2D1BWP12T U385 ( .A1(n3586), .A2(n3585), .ZN(n3591) );
  MAOI22D0BWP12T U386 ( .A1(n4767), .A2(n6122), .B1(n4816), .B2(n6120), .ZN(
        n3590) );
  OAI22D1BWP12T U387 ( .A1(n4926), .A2(n6113), .B1(n5600), .B2(n5511), .ZN(
        n3585) );
  OAI22D1BWP12T U388 ( .A1(n5372), .A2(n6130), .B1(n6048), .B2(n3525), .ZN(
        n3547) );
  MAOI22D0BWP12T U389 ( .A1(n6074), .A2(n3528), .B1(n6096), .B2(n5452), .ZN(
        n3531) );
  FA1D0BWP12T U390 ( .A(n3247), .B(n3246), .CI(n3245), .CO(n3241), .S(n3336)
         );
  AOI21D0BWP12T U391 ( .A1(n4211), .A2(n3518), .B(n3503), .ZN(n3397) );
  AOI22D0BWP12T U392 ( .A1(n3608), .A2(n5192), .B1(n5262), .B2(n5178), .ZN(
        n3123) );
  AOI22D0BWP12T U393 ( .A1(n5177), .A2(n5254), .B1(n5255), .B2(n3610), .ZN(
        n3124) );
  CKND2D0BWP12T U394 ( .A1(n3123), .A2(n3124), .ZN(n5259) );
  CKND2D0BWP12T U395 ( .A1(n3563), .A2(n3562), .ZN(n3125) );
  AOI22D0BWP12T U396 ( .A1(n5095), .A2(n3564), .B1(n5051), .B2(n5436), .ZN(
        n3126) );
  CKND2D0BWP12T U397 ( .A1(n5057), .A2(n3565), .ZN(n3127) );
  OAI211D0BWP12T U398 ( .A1(n5210), .A2(n3125), .B(n3126), .C(n3127), .ZN(
        n5067) );
  CKND2D0BWP12T U399 ( .A1(n3423), .A2(n3368), .ZN(n3128) );
  MAOI22D0BWP12T U400 ( .A1(n3393), .A2(n3128), .B1(n3393), .B2(n3128), .ZN(
        n4876) );
  MAOI22D0BWP12T U401 ( .A1(n6122), .A2(n4766), .B1(n4872), .B2(n6126), .ZN(
        n3476) );
  INR2D0BWP12T U402 ( .A1(n5143), .B1(n3569), .ZN(n3568) );
  IAO21D0BWP12T U403 ( .A1(n5798), .A2(n5634), .B(n5383), .ZN(n3631) );
  IAO21D0BWP12T U404 ( .A1(n3640), .A2(n3639), .B(n5471), .ZN(n3692) );
  INVD1BWP12T U405 ( .I(n3294), .ZN(n3295) );
  FA1D0BWP12T U406 ( .A(n3297), .B(n3296), .CI(n3295), .CO(n3524), .S(n3556)
         );
  IAO21D0BWP12T U407 ( .A1(n3619), .A2(n3620), .B(n5447), .ZN(n3587) );
  AOI21D1BWP12T U408 ( .A1(n5238), .A2(n3708), .B(b[4]), .ZN(n3375) );
  OAI211D1BWP12T U409 ( .A1(n3663), .A2(n3538), .B(n3375), .C(n3374), .ZN(
        n3384) );
  IND2D0BWP12T U410 ( .A1(n5642), .B1(n5645), .ZN(n4917) );
  NR2D0BWP12T U411 ( .A1(n3400), .A2(n3728), .ZN(n3129) );
  MAOI22D0BWP12T U412 ( .A1(n5086), .A2(n5229), .B1(n3129), .B2(n3204), .ZN(
        n5104) );
  CKND0BWP12T U413 ( .I(n5128), .ZN(n3130) );
  AOI21D0BWP12T U414 ( .A1(n5210), .A2(n3566), .B(n3130), .ZN(n3131) );
  AOI22D0BWP12T U415 ( .A1(n5095), .A2(n3563), .B1(n3346), .B2(n3131), .ZN(
        n5014) );
  CKND0BWP12T U416 ( .I(n3419), .ZN(n3132) );
  MAOI222D0BWP12T U417 ( .A(n3254), .B(n3265), .C(n3132), .ZN(n3331) );
  MAOI22D0BWP12T U418 ( .A1(n3265), .A2(n3254), .B1(n3265), .B2(n3254), .ZN(
        n3133) );
  MAOI22D0BWP12T U419 ( .A1(n3419), .A2(n3133), .B1(n3419), .B2(n3133), .ZN(
        n5341) );
  CKND2D0BWP12T U420 ( .A1(n3423), .A2(n3394), .ZN(n3134) );
  MAOI22D0BWP12T U421 ( .A1(n4148), .A2(n3134), .B1(n4148), .B2(n3134), .ZN(
        n4823) );
  INVD1BWP12T U422 ( .I(n5021), .ZN(n3513) );
  MAOI22D0BWP12T U423 ( .A1(n5826), .A2(n5548), .B1(n3499), .B2(n5646), .ZN(
        n3516) );
  AOI32D1BWP12T U424 ( .A1(n4419), .A2(n4330), .A3(n3488), .B1(n3373), .B2(
        b[1]), .ZN(n3713) );
  AOI21D0BWP12T U425 ( .A1(n5798), .A2(n4758), .B(n5804), .ZN(n3638) );
  IAO21D0BWP12T U426 ( .A1(n3632), .A2(n3631), .B(n5384), .ZN(n3690) );
  IND2D1BWP12T U427 ( .A1(n3307), .B1(b[0]), .ZN(n3318) );
  FA1D0BWP12T U428 ( .A(n3318), .B(n3317), .CI(n3316), .CO(n3603), .S(n3669)
         );
  IOA21D0BWP12T U429 ( .A1(n3682), .A2(n3683), .B(n5444), .ZN(n3616) );
  OAI21D0BWP12T U430 ( .A1(n3279), .A2(n3280), .B(n3278), .ZN(n3135) );
  MAOI22D0BWP12T U431 ( .A1(n3284), .A2(n3135), .B1(n3284), .B2(n3135), .ZN(
        n3136) );
  MAOI22D0BWP12T U432 ( .A1(n3330), .A2(n3136), .B1(n3330), .B2(n3136), .ZN(
        n3288) );
  CKND0BWP12T U433 ( .I(n3330), .ZN(n3137) );
  MAOI222D0BWP12T U434 ( .A(n3284), .B(n3137), .C(n3135), .ZN(n3456) );
  AOI21D0BWP12T U435 ( .A1(n4837), .A2(n4862), .B(n5642), .ZN(n4860) );
  IAO21D0BWP12T U436 ( .A1(n4891), .A2(n4931), .B(n5696), .ZN(n4911) );
  AOI21D0BWP12T U437 ( .A1(n4941), .A2(n4754), .B(n6012), .ZN(n4753) );
  IAO21D0BWP12T U438 ( .A1(n4936), .A2(n4894), .B(n5437), .ZN(n4938) );
  IAO21D0BWP12T U439 ( .A1(n4908), .A2(n4783), .B(n6132), .ZN(n4751) );
  IOA21D0BWP12T U440 ( .A1(n5917), .A2(n4904), .B(n5916), .ZN(n4905) );
  OA21D0BWP12T U441 ( .A1(n5752), .A2(n4750), .B(n5431), .Z(n4788) );
  IOA21D0BWP12T U442 ( .A1(n5887), .A2(n4902), .B(n4901), .ZN(n4950) );
  OAI22D0BWP12T U443 ( .A1(n3610), .A2(n5286), .B1(n5288), .B2(n5177), .ZN(
        n3138) );
  OAI22D0BWP12T U444 ( .A1(n5282), .A2(n3608), .B1(n3609), .B2(n5284), .ZN(
        n3139) );
  NR2D0BWP12T U445 ( .A1(n3138), .A2(n3139), .ZN(n5090) );
  NR2D0BWP12T U446 ( .A1(n3588), .A2(n3600), .ZN(n3140) );
  MAOI22D0BWP12T U447 ( .A1(n3140), .A2(n3589), .B1(n3140), .B2(n3589), .ZN(
        n4816) );
  IAO21D0BWP12T U448 ( .A1(n4148), .A2(n4889), .B(n3357), .ZN(n3141) );
  MAOI22D0BWP12T U449 ( .A1(n3365), .A2(n3141), .B1(n3365), .B2(n3141), .ZN(
        n4930) );
  AOI22D0BWP12T U450 ( .A1(n5052), .A2(n5230), .B1(n5057), .B2(n5231), .ZN(
        n3142) );
  OAI22D0BWP12T U451 ( .A1(n4995), .A2(n5014), .B1(n5054), .B2(n4996), .ZN(
        n3143) );
  AOI211D0BWP12T U452 ( .A1(n5056), .A2(n4997), .B(n5528), .C(n3143), .ZN(
        n3144) );
  AOI22D0BWP12T U453 ( .A1(n5229), .A2(n5095), .B1(n5051), .B2(n5228), .ZN(
        n3145) );
  AOI32D0BWP12T U454 ( .A1(n3142), .A2(n3144), .A3(n3145), .B1(n5081), .B2(
        n3144), .ZN(n5732) );
  INVD1BWP12T U455 ( .I(n5011), .ZN(n3439) );
  AOI211D1BWP12T U456 ( .A1(n5815), .A2(n5113), .B(n3441), .C(n3440), .ZN(
        n3448) );
  OAI32D1BWP12T U457 ( .A1(n4419), .A2(n3400), .A3(n3399), .B1(b[1]), .B2(
        n3398), .ZN(n3570) );
  FA1D0BWP12T U458 ( .A(n3234), .B(n3233), .CI(n3232), .CO(n4528), .S(n3333)
         );
  OA21D0BWP12T U459 ( .A1(n3211), .A2(n3212), .B(n4538), .Z(n3146) );
  CKND0BWP12T U460 ( .I(n3242), .ZN(n3147) );
  CKND0BWP12T U461 ( .I(n3241), .ZN(n3148) );
  MAOI222D0BWP12T U462 ( .A(n3146), .B(n3147), .C(n3148), .ZN(n4546) );
  MAOI22D0BWP12T U463 ( .A1(n3146), .A2(n3147), .B1(n3146), .B2(n3147), .ZN(
        n3149) );
  MAOI22D0BWP12T U464 ( .A1(n3241), .A2(n3149), .B1(n3241), .B2(n3149), .ZN(
        n3334) );
  IAO21D0BWP12T U465 ( .A1(n3638), .A2(n3640), .B(n5439), .ZN(n3722) );
  IAO21D0BWP12T U466 ( .A1(n3723), .A2(n3690), .B(n5385), .ZN(n3674) );
  IAO21D0BWP12T U467 ( .A1(n3620), .A2(n3616), .B(n5459), .ZN(n3582) );
  IAO21D0BWP12T U468 ( .A1(n3587), .A2(n3589), .B(n5438), .ZN(n3521) );
  OAI32D1BWP12T U469 ( .A1(n4419), .A2(n3404), .A3(n3403), .B1(n3451), .B2(
        b[1]), .ZN(n3630) );
  IAO21D0BWP12T U470 ( .A1(n4809), .A2(n4917), .B(n5642), .ZN(n4808) );
  AOI21D0BWP12T U471 ( .A1(n5858), .A2(n4915), .B(n5478), .ZN(n4913) );
  IOA21D0BWP12T U472 ( .A1(n4857), .A2(n4756), .B(n5469), .ZN(n4754) );
  IAO21D0BWP12T U473 ( .A1(n4909), .A2(n4910), .B(n5994), .ZN(n4936) );
  IOA21D0BWP12T U474 ( .A1(n4939), .A2(n4755), .B(n5965), .ZN(n4783) );
  AO21D0BWP12T U475 ( .A1(n4896), .A2(n4947), .B(n5943), .Z(n4904) );
  AOI21D0BWP12T U476 ( .A1(n4419), .A2(n3593), .B(n5210), .ZN(n3150) );
  OAI22D0BWP12T U477 ( .A1(n4419), .A2(n4599), .B1(n3150), .B2(n3497), .ZN(
        n5531) );
  IAO21D0BWP12T U478 ( .A1(n4847), .A2(n4782), .B(n5838), .ZN(n4787) );
  AOI32D1BWP12T U479 ( .A1(n3405), .A2(n3203), .A3(n3817), .B1(n4600), .B2(
        n3203), .ZN(n5278) );
  IOA21D0BWP12T U480 ( .A1(n4898), .A2(n4944), .B(n5431), .ZN(n4900) );
  IOA21D0BWP12T U481 ( .A1(n5887), .A2(n4748), .B(n4901), .ZN(n4749) );
  MOAI22D0BWP12T U482 ( .A1(n3603), .A2(n3313), .B1(n3603), .B2(n3313), .ZN(
        n3151) );
  MAOI22D0BWP12T U483 ( .A1(n3602), .A2(n3151), .B1(n3602), .B2(n3151), .ZN(
        n5348) );
  MAOI222D0BWP12T U484 ( .A(n3313), .B(n3152), .C(n3153), .ZN(n3555) );
  CKND0BWP12T U485 ( .I(n3602), .ZN(n3152) );
  CKND0BWP12T U486 ( .I(n3603), .ZN(n3153) );
  AOI22D0BWP12T U487 ( .A1(n5525), .A2(n3715), .B1(n5242), .B2(n3714), .ZN(
        n3154) );
  OAI211D0BWP12T U488 ( .A1(n5136), .A2(n5080), .B(n5703), .C(n3154), .ZN(
        n5109) );
  MAOI22D0BWP12T U489 ( .A1(n3325), .A2(n3329), .B1(n3325), .B2(n3329), .ZN(
        n3155) );
  MAOI22D0BWP12T U490 ( .A1(n3456), .A2(n3155), .B1(n3456), .B2(n3155), .ZN(
        n5338) );
  CKND0BWP12T U491 ( .I(n3456), .ZN(n3156) );
  MAOI222D0BWP12T U492 ( .A(n3325), .B(n3329), .C(n3156), .ZN(n3502) );
  NR2D0BWP12T U493 ( .A1(n3449), .A2(n3526), .ZN(n3157) );
  MAOI22D0BWP12T U494 ( .A1(n3157), .A2(n3473), .B1(n3157), .B2(n3473), .ZN(
        n4817) );
  OA22D0BWP12T U495 ( .A1(n5263), .A2(n5259), .B1(n5280), .B2(n5269), .Z(n3158) );
  CKND2D0BWP12T U496 ( .A1(n3499), .A2(n3158), .ZN(n5140) );
  AOI22D0BWP12T U497 ( .A1(n5095), .A2(n5283), .B1(n5057), .B2(n5289), .ZN(
        n3159) );
  OAI22D0BWP12T U498 ( .A1(n4995), .A2(n5036), .B1(n5054), .B2(n5033), .ZN(
        n3160) );
  AOI211D0BWP12T U499 ( .A1(n5056), .A2(n5034), .B(n5528), .C(n3160), .ZN(
        n3161) );
  AOI22D0BWP12T U500 ( .A1(n5052), .A2(n5287), .B1(n5051), .B2(n5285), .ZN(
        n3162) );
  AOI32D0BWP12T U501 ( .A1(n3159), .A2(n3161), .A3(n3162), .B1(n5081), .B2(
        n3161), .ZN(n5898) );
  NR2D1BWP12T U502 ( .A1(n3410), .A2(n3749), .ZN(n3387) );
  OAI22D1BWP12T U503 ( .A1(n6048), .A2(n4743), .B1(n4057), .B2(n6128), .ZN(
        n3379) );
  OAI22D1BWP12T U504 ( .A1(n3387), .A2(n3386), .B1(n4933), .B2(n6113), .ZN(
        n3388) );
  OAI22D1BWP12T U505 ( .A1(n4980), .A2(n5631), .B1(n5600), .B2(n5083), .ZN(
        n3389) );
  NR4D0BWP12T U506 ( .A1(n3391), .A2(n3390), .A3(n3389), .A4(n3388), .ZN(n3396) );
  FA1D0BWP12T U507 ( .A(n4530), .B(n4529), .CI(n4528), .CO(n4534), .S(n4548)
         );
  CKND0BWP12T U508 ( .I(n3488), .ZN(n3163) );
  OAI32D0BWP12T U509 ( .A1(n5253), .A2(n4378), .A3(n3163), .B1(n3493), .B2(
        n5253), .ZN(n5246) );
  OAI32D1BWP12T U510 ( .A1(b[1]), .A2(n3402), .A3(n4970), .B1(n3401), .B2(
        n4419), .ZN(n5121) );
  ND2D1BWP12T U511 ( .A1(n4266), .A2(n4956), .ZN(n3371) );
  OAI32D1BWP12T U512 ( .A1(n4419), .A2(n3483), .A3(n3484), .B1(b[1]), .B2(
        n3371), .ZN(n3538) );
  ND2D1BWP12T U513 ( .A1(a[0]), .A2(b[2]), .ZN(n3319) );
  AOI32D1BWP12T U514 ( .A1(n3321), .A2(n5809), .A3(n3319), .B1(b[2]), .B2(
        n4455), .ZN(n3634) );
  AO21D0BWP12T U515 ( .A1(n3640), .A2(n3637), .B(n5384), .Z(n3696) );
  IAO21D0BWP12T U516 ( .A1(n3722), .A2(n3691), .B(n5440), .ZN(n3681) );
  IAO21D0BWP12T U517 ( .A1(n3582), .A2(n3589), .B(n5458), .ZN(n3540) );
  IAO21D0BWP12T U518 ( .A1(n3397), .A2(n3446), .B(n3361), .ZN(n4745) );
  OA21D0BWP12T U519 ( .A1(n4912), .A2(n4911), .B(n5434), .Z(n4940) );
  IAO21D0BWP12T U520 ( .A1(n4784), .A2(n4894), .B(n5437), .ZN(n4755) );
  IOA21D0BWP12T U521 ( .A1(n5917), .A2(n4752), .B(n5460), .ZN(n4782) );
  IOA21D0BWP12T U522 ( .A1(n4897), .A2(n4945), .B(n5430), .ZN(n4944) );
  IAO21D0BWP12T U523 ( .A1(n4788), .A2(n5727), .B(n5432), .ZN(n4748) );
  IAO21D0BWP12T U524 ( .A1(n4951), .A2(n4950), .B(n5433), .ZN(n5580) );
  CKND0BWP12T U525 ( .I(n3653), .ZN(n3164) );
  AOI32D0BWP12T U526 ( .A1(n3646), .A2(n3164), .A3(n3720), .B1(n5703), .B2(
        n3164), .ZN(n5091) );
  AOI211D1BWP12T U527 ( .A1(n5238), .A2(n5106), .B(b[4]), .C(n3665), .ZN(n5112) );
  MOAI22D0BWP12T U528 ( .A1(n3556), .A2(n3306), .B1(n3556), .B2(n3306), .ZN(
        n3165) );
  MAOI22D0BWP12T U529 ( .A1(n3555), .A2(n3165), .B1(n3555), .B2(n3165), .ZN(
        n5311) );
  MAOI222D0BWP12T U530 ( .A(n3306), .B(n3166), .C(n3167), .ZN(n3523) );
  CKND0BWP12T U531 ( .I(n3555), .ZN(n3166) );
  CKND0BWP12T U532 ( .I(n3556), .ZN(n3167) );
  NR2D0BWP12T U533 ( .A1(n5128), .A2(n3535), .ZN(n3168) );
  OAI22D0BWP12T U534 ( .A1(n3534), .A2(n5045), .B1(n3536), .B2(n5131), .ZN(
        n3169) );
  AOI211D0BWP12T U535 ( .A1(n5052), .A2(n3610), .B(n3168), .C(n3169), .ZN(
        n5024) );
  CKND2D0BWP12T U536 ( .A1(n3472), .A2(n3525), .ZN(n3170) );
  MOAI22D0BWP12T U537 ( .A1(n3473), .A2(n3170), .B1(n3473), .B2(n3170), .ZN(
        n4766) );
  CKND0BWP12T U538 ( .I(n3502), .ZN(n3171) );
  MAOI222D0BWP12T U539 ( .A(n3269), .B(n3277), .C(n3171), .ZN(n3419) );
  MAOI22D0BWP12T U540 ( .A1(n3277), .A2(n3269), .B1(n3277), .B2(n3269), .ZN(
        n3172) );
  MAOI22D0BWP12T U541 ( .A1(n3502), .A2(n3172), .B1(n3502), .B2(n3172), .ZN(
        n5339) );
  MOAI22D0BWP12T U542 ( .A1(n5858), .A2(n4808), .B1(n5858), .B2(n4808), .ZN(
        n5880) );
  OAI22D1BWP12T U543 ( .A1(n3209), .A2(n4792), .B1(n4744), .B2(n6096), .ZN(
        n3339) );
  FA1D0BWP12T U544 ( .A(n4524), .B(n4523), .CI(n4522), .CO(n4536), .S(n4529)
         );
  FA1D0BWP12T U545 ( .A(n4518), .B(n4517), .CI(n4516), .CO(n4531), .S(n4539)
         );
  MAOI222D0BWP12T U546 ( .A(n4273), .B(n4261), .C(n4252), .ZN(n4274) );
  MOAI22D0BWP12T U547 ( .A1(n4261), .A2(n4252), .B1(n4261), .B2(n4252), .ZN(
        n3173) );
  MAOI22D0BWP12T U548 ( .A1(n4273), .A2(n3173), .B1(n4273), .B2(n3173), .ZN(
        n4338) );
  AOI22D1BWP12T U549 ( .A1(n3480), .A2(n5758), .B1(n3409), .B2(n3408), .ZN(
        n3571) );
  MOAI22D0BWP12T U550 ( .A1(b[0]), .A2(a[26]), .B1(n3817), .B2(b[1]), .ZN(
        n3409) );
  CKND0BWP12T U551 ( .I(n5797), .ZN(n3174) );
  OAI21D0BWP12T U552 ( .A1(n4810), .A2(n3174), .B(n5806), .ZN(n3637) );
  IAO21D0BWP12T U553 ( .A1(n3692), .A2(n3691), .B(n5472), .ZN(n3683) );
  ND2D1BWP12T U554 ( .A1(b[0]), .A2(a[7]), .ZN(n3661) );
  IAO21D0BWP12T U555 ( .A1(n3681), .A2(n3685), .B(n3358), .ZN(n3619) );
  AOI32D1BWP12T U556 ( .A1(n3487), .A2(b[1]), .A3(n3372), .B1(n3489), .B2(
        n4419), .ZN(n3714) );
  AOI21D0BWP12T U557 ( .A1(n4495), .A2(n3550), .B(n3533), .ZN(n3475) );
  IAO21D0BWP12T U558 ( .A1(n4858), .A2(n4806), .B(n6046), .ZN(n4824) );
  IAO21D0BWP12T U559 ( .A1(n4891), .A2(n4776), .B(n5696), .ZN(n4756) );
  IAO21D0BWP12T U560 ( .A1(n4940), .A2(n4892), .B(n6017), .ZN(n4909) );
  AOI22D0BWP12T U561 ( .A1(n5052), .A2(n5177), .B1(n5178), .B2(n5095), .ZN(
        n3175) );
  AOI22D0BWP12T U562 ( .A1(n5051), .A2(n3608), .B1(n5250), .B2(n5057), .ZN(
        n3176) );
  CKND2D0BWP12T U563 ( .A1(n3175), .A2(n3176), .ZN(n5030) );
  AOI21D0BWP12T U564 ( .A1(n4893), .A2(n4753), .B(n5994), .ZN(n4784) );
  OA21D0BWP12T U565 ( .A1(n4895), .A2(n4938), .B(n5961), .Z(n4907) );
  IAO21D0BWP12T U566 ( .A1(n4751), .A2(n4946), .B(n5943), .ZN(n4752) );
  ND2D1BWP12T U567 ( .A1(n4266), .A2(n3491), .ZN(n5150) );
  IOA21D0BWP12T U568 ( .A1(n4906), .A2(n4905), .B(n5429), .ZN(n4945) );
  IAO21D0BWP12T U569 ( .A1(n4787), .A2(n5772), .B(n5773), .ZN(n4750) );
  AOI21D0BWP12T U570 ( .A1(n4899), .A2(n4900), .B(n5432), .ZN(n4902) );
  IAO21D0BWP12T U571 ( .A1(n4951), .A2(n4749), .B(n5433), .ZN(n5579) );
  OA21D0BWP12T U572 ( .A1(n3324), .A2(n3323), .B(n3670), .Z(n3177) );
  OAI21D0BWP12T U573 ( .A1(n3322), .A2(n3710), .B(n4657), .ZN(n3178) );
  CKND0BWP12T U574 ( .I(n3699), .ZN(n3179) );
  MAOI222D0BWP12T U575 ( .A(n3177), .B(n3178), .C(n3179), .ZN(n3668) );
  MAOI22D0BWP12T U576 ( .A1(n3177), .A2(n3178), .B1(n3177), .B2(n3178), .ZN(
        n3180) );
  MAOI22D0BWP12T U577 ( .A1(n3699), .A2(n3180), .B1(n3699), .B2(n3180), .ZN(
        n5373) );
  CKND0BWP12T U578 ( .I(n3524), .ZN(n3181) );
  CKND0BWP12T U579 ( .I(n3523), .ZN(n3182) );
  MAOI222D0BWP12T U580 ( .A(n3288), .B(n3181), .C(n3182), .ZN(n3325) );
  MAOI22D0BWP12T U581 ( .A1(n3288), .A2(n3181), .B1(n3288), .B2(n3181), .ZN(
        n3183) );
  MAOI22D0BWP12T U582 ( .A1(n3523), .A2(n3183), .B1(n3523), .B2(n3183), .ZN(
        n5372) );
  CKND2D0BWP12T U583 ( .A1(n3467), .A2(n3525), .ZN(n3184) );
  MAOI22D0BWP12T U584 ( .A1(n3473), .A2(n3184), .B1(n3473), .B2(n3184), .ZN(
        n4927) );
  AOI211D1BWP12T U585 ( .A1(n5525), .A2(n3630), .B(b[4]), .C(n3407), .ZN(n3412) );
  CKND0BWP12T U586 ( .I(n3377), .ZN(n3185) );
  CKND0BWP12T U587 ( .I(n3376), .ZN(n3186) );
  MAOI222D0BWP12T U588 ( .A(n3331), .B(n3185), .C(n3186), .ZN(n4549) );
  MAOI22D0BWP12T U589 ( .A1(n3331), .A2(n3185), .B1(n3331), .B2(n3185), .ZN(
        n3187) );
  MAOI22D0BWP12T U590 ( .A1(n3376), .A2(n3187), .B1(n3376), .B2(n3187), .ZN(
        n5358) );
  IOA21D0BWP12T U591 ( .A1(n3392), .A2(n3393), .B(n4743), .ZN(n3188) );
  MOAI22D0BWP12T U592 ( .A1(n3365), .A2(n3188), .B1(n3365), .B2(n3188), .ZN(
        n4774) );
  AOI22D0BWP12T U593 ( .A1(n5262), .A2(n3455), .B1(n5254), .B2(n3567), .ZN(
        n3189) );
  OAI21D0BWP12T U594 ( .A1(n5284), .A2(n3563), .B(n3189), .ZN(n3190) );
  AOI21D0BWP12T U595 ( .A1(n5192), .A2(n3566), .B(n3190), .ZN(n5706) );
  OAI32D1BWP12T U596 ( .A1(n5858), .A2(b[14]), .A3(n6093), .B1(n6096), .B2(
        n5858), .ZN(n5860) );
  INVD1BWP12T U597 ( .I(n4455), .ZN(n5809) );
  IND2XD1BWP12T U598 ( .A1(n3526), .B1(n3458), .ZN(n5393) );
  NR2XD0BWP12T U599 ( .A1(n3577), .A2(n4555), .ZN(n3558) );
  OR2D1BWP12T U600 ( .A1(n3558), .A2(n3600), .Z(n5394) );
  MAOI222D1BWP12T U601 ( .A(a[0]), .B(b[0]), .C(c_in), .ZN(n4810) );
  CKND1BWP12T U602 ( .I(n5806), .ZN(n5383) );
  MAOI222D1BWP12T U603 ( .A(b[3]), .B(a[3]), .C(n3696), .ZN(n3684) );
  MAOI222D1BWP12T U604 ( .A(n5703), .B(n3709), .C(n3684), .ZN(n3592) );
  MAOI222D1BWP12T U605 ( .A(b[9]), .B(a[9]), .C(n3478), .ZN(n3443) );
  CKND2D0BWP12T U606 ( .A1(n3423), .A2(n4057), .ZN(n5395) );
  INVD1BWP12T U607 ( .I(op[3]), .ZN(n3202) );
  INVD1BWP12T U608 ( .I(op[2]), .ZN(n5594) );
  NR2D0BWP12T U609 ( .A1(n3361), .A2(n3503), .ZN(n5446) );
  CKND2D1BWP12T U610 ( .A1(n3466), .A2(n3525), .ZN(n5442) );
  NR2XD0BWP12T U611 ( .A1(n4490), .A2(a[5]), .ZN(n5459) );
  AOI22D0BWP12T U612 ( .A1(n5633), .A2(b[0]), .B1(n5805), .B2(b[1]), .ZN(n5467) );
  CKND0BWP12T U613 ( .I(n5804), .ZN(n3321) );
  NR2D1BWP12T U614 ( .A1(n5458), .A2(n5438), .ZN(n4493) );
  CKND2D0BWP12T U615 ( .A1(n3540), .A2(n5452), .ZN(n3467) );
  AOI21D0BWP12T U616 ( .A1(n3359), .A2(n3467), .B(n3450), .ZN(n3479) );
  CKND2D0BWP12T U617 ( .A1(n3479), .A2(n5454), .ZN(n3434) );
  AOI22D0BWP12T U618 ( .A1(b[10]), .A2(n3421), .B1(n5446), .B2(n3434), .ZN(
        n3385) );
  INVD1BWP12T U619 ( .I(n3385), .ZN(n4889) );
  ND4D0BWP12T U620 ( .A1(n3192), .A2(n4838), .A3(n4699), .A4(n4450), .ZN(n3195) );
  ND3D0BWP12T U621 ( .A1(n3193), .A2(n5390), .A3(n4792), .ZN(n3194) );
  NR4D0BWP12T U622 ( .A1(b[29]), .A2(b[24]), .A3(n3195), .A4(n3194), .ZN(n3196) );
  CKND2D0BWP12T U623 ( .A1(n5570), .A2(n5079), .ZN(n5068) );
  INVD1BWP12T U624 ( .I(n5068), .ZN(n4982) );
  CKND0BWP12T U625 ( .I(n5436), .ZN(n5638) );
  OAI22D1BWP12T U626 ( .A1(n5379), .A2(a[3]), .B1(a[4]), .B2(b[0]), .ZN(n3564)
         );
  OAI22D1BWP12T U627 ( .A1(n5379), .A2(n3509), .B1(n3421), .B2(b[0]), .ZN(
        n5191) );
  OAI22D1BWP12T U628 ( .A1(n5379), .A2(n3528), .B1(n3360), .B2(b[0]), .ZN(
        n3455) );
  AOI22D0BWP12T U629 ( .A1(n5095), .A2(n5123), .B1(n5122), .B2(n5052), .ZN(
        n3201) );
  CKND2D1BWP12T U630 ( .A1(n5210), .A2(n4419), .ZN(n5131) );
  OAI22D1BWP12T U631 ( .A1(n5379), .A2(n3749), .B1(n4791), .B2(b[0]), .ZN(
        n5193) );
  CKND0BWP12T U632 ( .I(n5193), .ZN(n5158) );
  OAI22D1BWP12T U633 ( .A1(n5379), .A2(n3300), .B1(n3577), .B2(b[0]), .ZN(
        n3567) );
  AOI22D0BWP12T U634 ( .A1(n5057), .A2(n5158), .B1(n5051), .B2(n3565), .ZN(
        n3200) );
  ND2D1BWP12T U635 ( .A1(n5594), .A2(n3202), .ZN(n3344) );
  NR2D1BWP12T U636 ( .A1(n5379), .A2(n4419), .ZN(n3485) );
  INVD0BWP12T U637 ( .I(n3485), .ZN(n3405) );
  CKND2D1BWP12T U638 ( .A1(n5379), .A2(b[1]), .ZN(n3562) );
  CKND0BWP12T U639 ( .I(n3562), .ZN(n3204) );
  AOI22D0BWP12T U640 ( .A1(a[30]), .A2(n3204), .B1(a[28]), .B2(n3430), .ZN(
        n3203) );
  NR2XD0BWP12T U641 ( .A1(a[31]), .A2(n4419), .ZN(n4600) );
  CKND2D1BWP12T U642 ( .A1(n5278), .A2(n5525), .ZN(n5723) );
  CKND0BWP12T U643 ( .I(n5525), .ZN(n5245) );
  CKND2D1BWP12T U644 ( .A1(n5245), .A2(a[31]), .ZN(n5532) );
  AOI22D1BWP12T U645 ( .A1(b[0]), .A2(a[25]), .B1(a[26]), .B2(n5379), .ZN(
        n5229) );
  NR2D0BWP12T U646 ( .A1(a[27]), .A2(n4419), .ZN(n3728) );
  OAI22D0BWP12T U647 ( .A1(n5379), .A2(a[23]), .B1(a[22]), .B2(b[0]), .ZN(
        n3398) );
  NR2D0BWP12T U648 ( .A1(a[21]), .A2(n5379), .ZN(n4172) );
  OR2D1BWP12T U649 ( .A1(n4971), .A2(n4172), .Z(n3401) );
  OAI22D0BWP12T U650 ( .A1(n5210), .A2(n5104), .B1(n5105), .B2(b[2]), .ZN(
        n3658) );
  AOI22D1BWP12T U651 ( .A1(b[0]), .A2(a[13]), .B1(a[14]), .B2(n5379), .ZN(
        n5159) );
  TPNR2D0BWP12T U652 ( .A1(n4419), .A2(n3205), .ZN(n3206) );
  CKND0BWP12T U653 ( .I(n3664), .ZN(n5134) );
  CKND2D1BWP12T U654 ( .A1(n5136), .A2(b[2]), .ZN(n3707) );
  OAI22D1BWP12T U655 ( .A1(n5379), .A2(a[17]), .B1(a[18]), .B2(b[0]), .ZN(
        n5188) );
  TPNR2D0BWP12T U656 ( .A1(n3572), .A2(n5188), .ZN(n5212) );
  AOI22D0BWP12T U657 ( .A1(a[19]), .A2(n3485), .B1(a[16]), .B2(n3430), .ZN(
        n3207) );
  IND2XD1BWP12T U658 ( .A1(n5212), .B1(n3207), .ZN(n5106) );
  AOI22D0BWP12T U659 ( .A1(n5525), .A2(n5134), .B1(n5242), .B2(n5106), .ZN(
        n3208) );
  OA211D0BWP12T U660 ( .A1(n3658), .A2(n5136), .B(n3208), .C(n5703), .Z(n3349)
         );
  NR2D1BWP12T U661 ( .A1(n5592), .A2(op[2]), .ZN(n6045) );
  CKND2D1BWP12T U662 ( .A1(op[2]), .A2(op[3]), .ZN(n3504) );
  AOI21D0BWP12T U663 ( .A1(a[12]), .A2(n6045), .B(n6150), .ZN(n3209) );
  CKND2D1BWP12T U664 ( .A1(a[0]), .A2(n5805), .ZN(n4470) );
  NR2D1BWP12T U665 ( .A1(n5805), .A2(a[0]), .ZN(n5380) );
  NR2D1BWP12T U666 ( .A1(n5633), .A2(n5805), .ZN(n4455) );
  AOI22D0BWP12T U667 ( .A1(n5380), .A2(n4646), .B1(n4455), .B2(n4741), .ZN(
        n3210) );
  OAI21D0BWP12T U668 ( .A1(n4741), .A2(n4470), .B(n3210), .ZN(n3212) );
  CKND2D0BWP12T U669 ( .A1(a[10]), .A2(a[9]), .ZN(n5423) );
  OA21D0BWP12T U670 ( .A1(a[10]), .A2(a[9]), .B(n5423), .Z(n4131) );
  TPND3D0BWP12T U671 ( .A1(n3421), .A2(n3509), .A3(a[11]), .ZN(n4128) );
  NR2D0BWP12T U672 ( .A1(n5421), .A2(n5805), .ZN(n3322) );
  OR2XD1BWP12T U673 ( .A1(n3341), .A2(n3322), .Z(n3320) );
  NR2D1BWP12T U674 ( .A1(n3363), .A2(n3320), .ZN(n4660) );
  CKND2D1BWP12T U675 ( .A1(n3322), .A2(n3363), .ZN(n4658) );
  CKND2D1BWP12T U676 ( .A1(a[3]), .A2(n3341), .ZN(n4657) );
  AOI22D0BWP12T U677 ( .A1(b[8]), .A2(n4658), .B1(n4657), .B2(n4699), .ZN(
        n3213) );
  AOI221D0BWP12T U678 ( .A1(n4661), .A2(b[9]), .B1(n4660), .B2(n4482), .C(
        n3213), .ZN(n3240) );
  OAI22D1BWP12T U679 ( .A1(n5379), .A2(n3421), .B1(n3749), .B2(b[0]), .ZN(
        n3382) );
  CKND0BWP12T U680 ( .I(n4640), .ZN(n4129) );
  CKND2D0BWP12T U681 ( .A1(n4129), .A2(n4128), .ZN(n4210) );
  CKND2D1BWP12T U682 ( .A1(n4131), .A2(n3749), .ZN(n4637) );
  AOI22D0BWP12T U683 ( .A1(b[1]), .A2(n4637), .B1(n4636), .B2(n4419), .ZN(
        n3214) );
  AOI21D0BWP12T U684 ( .A1(n3382), .A2(n4210), .B(n3214), .ZN(n3239) );
  NR2D1BWP12T U685 ( .A1(a[7]), .A2(n5424), .ZN(n4635) );
  NR3D1BWP12T U686 ( .A1(a[6]), .A2(a[5]), .A3(n3528), .ZN(n4634) );
  CKND0BWP12T U687 ( .I(n3286), .ZN(n4494) );
  CKND2D1BWP12T U688 ( .A1(n4494), .A2(n3528), .ZN(n4632) );
  ND2D1BWP12T U689 ( .A1(a[7]), .A2(n4494), .ZN(n4631) );
  AOI22D0BWP12T U690 ( .A1(b[5]), .A2(n4632), .B1(n4631), .B2(n4490), .ZN(
        n3215) );
  AOI221D0BWP12T U691 ( .A1(n4635), .A2(b[4]), .B1(n4634), .B2(n5703), .C(
        n3215), .ZN(n3238) );
  AOI22D0BWP12T U692 ( .A1(b[4]), .A2(n4632), .B1(n4631), .B2(n5703), .ZN(
        n3216) );
  AOI221D0BWP12T U693 ( .A1(n4635), .A2(b[3]), .B1(n4634), .B2(n5136), .C(
        n3216), .ZN(n3247) );
  NR2XD0BWP12T U694 ( .A1(n3307), .A2(a[5]), .ZN(n3302) );
  NR3D1BWP12T U695 ( .A1(a[4]), .A2(a[3]), .A3(n3300), .ZN(n4644) );
  NR2D1BWP12T U696 ( .A1(n4645), .A2(n4644), .ZN(n3304) );
  TPNR2D0BWP12T U697 ( .A1(n3300), .A2(n3307), .ZN(n3301) );
  OAI22D0BWP12T U698 ( .A1(n3622), .A2(n3304), .B1(b[6]), .B2(n4641), .ZN(
        n3217) );
  AOI21D0BWP12T U699 ( .A1(b[6]), .A2(n3302), .B(n3217), .ZN(n3246) );
  AOI22D0BWP12T U700 ( .A1(b[7]), .A2(n4658), .B1(n4657), .B2(n4450), .ZN(
        n3218) );
  AOI221D0BWP12T U701 ( .A1(n4661), .A2(b[8]), .B1(n4660), .B2(n4699), .C(
        n3218), .ZN(n3245) );
  AOI22D0BWP12T U702 ( .A1(b[7]), .A2(n4642), .B1(n4641), .B2(n4450), .ZN(
        n3219) );
  AOI221D0BWP12T U703 ( .A1(n4645), .A2(b[6]), .B1(n4644), .B2(n4555), .C(
        n3219), .ZN(n3234) );
  TPNR2D0BWP12T U704 ( .A1(n3360), .A2(n3528), .ZN(n5414) );
  CKND2D0BWP12T U705 ( .A1(n3509), .A2(n5414), .ZN(n4341) );
  CKND1BWP12T U706 ( .I(n4341), .ZN(n4671) );
  CKND2D0BWP12T U707 ( .A1(n3360), .A2(n3528), .ZN(n3342) );
  NR2D1BWP12T U708 ( .A1(n3509), .A2(n3342), .ZN(n4670) );
  INR2XD0BWP12T U709 ( .A1(n3342), .B1(n5414), .ZN(n4344) );
  CKND2D1BWP12T U710 ( .A1(n4344), .A2(n3509), .ZN(n4668) );
  AOI22D0BWP12T U711 ( .A1(b[3]), .A2(n4668), .B1(n4667), .B2(n5136), .ZN(
        n3220) );
  AOI221D0BWP12T U712 ( .A1(n4671), .A2(b[2]), .B1(n4670), .B2(n5210), .C(
        n3220), .ZN(n3233) );
  OAI22D0BWP12T U713 ( .A1(b[9]), .A2(n4453), .B1(n4646), .B2(n4470), .ZN(
        n3221) );
  AOI21D0BWP12T U714 ( .A1(n4455), .A2(n4646), .B(n3221), .ZN(n3226) );
  AOI22D0BWP12T U715 ( .A1(b[2]), .A2(n4668), .B1(n4667), .B2(n5210), .ZN(
        n3222) );
  AOI221D0BWP12T U716 ( .A1(n4671), .A2(b[1]), .B1(n4670), .B2(n4419), .C(
        n3222), .ZN(n3225) );
  ND2D0BWP12T U717 ( .A1(b[0]), .A2(n4131), .ZN(n3224) );
  OAI22D0BWP12T U718 ( .A1(n3622), .A2(n3307), .B1(n3304), .B2(n3685), .ZN(
        n3250) );
  AOI22D0BWP12T U719 ( .A1(n5380), .A2(n4699), .B1(n4455), .B2(n4482), .ZN(
        n3223) );
  OAI21D0BWP12T U720 ( .A1(n4482), .A2(n4470), .B(n3223), .ZN(n3251) );
  TPND2D0BWP12T U721 ( .A1(n3250), .A2(n3251), .ZN(n3249) );
  FA1D0BWP12T U722 ( .A(n3226), .B(n3225), .CI(n3224), .CO(n3232), .S(n3244)
         );
  AOI22D0BWP12T U723 ( .A1(b[1]), .A2(n4668), .B1(n4667), .B2(n4419), .ZN(
        n3227) );
  OAI22D1BWP12T U724 ( .A1(n5379), .A2(n3360), .B1(n3509), .B2(b[0]), .ZN(
        n5085) );
  OAI32D0BWP12T U725 ( .A1(n3227), .A2(n4671), .A3(n4670), .B1(n5085), .B2(
        n3227), .ZN(n3264) );
  AOI22D0BWP12T U726 ( .A1(b[6]), .A2(n4658), .B1(n4657), .B2(n4555), .ZN(
        n3228) );
  AOI221D1BWP12T U727 ( .A1(n4661), .A2(b[7]), .B1(n4660), .B2(n4450), .C(
        n3228), .ZN(n3263) );
  CKND2D0BWP12T U728 ( .A1(a[9]), .A2(n5379), .ZN(n3490) );
  IAO21D0BWP12T U729 ( .A1(n5414), .A2(n3490), .B(n4670), .ZN(n3262) );
  AOI22D0BWP12T U730 ( .A1(b[8]), .A2(n4642), .B1(n4641), .B2(n4699), .ZN(
        n3229) );
  AOI221D0BWP12T U731 ( .A1(n4645), .A2(b[7]), .B1(n4644), .B2(n4450), .C(
        n3229), .ZN(n4530) );
  AOI22D1BWP12T U732 ( .A1(a[12]), .A2(n3749), .B1(a[11]), .B2(n4791), .ZN(
        n4488) );
  OR2XD0BWP12T U733 ( .A1(n4488), .A2(n5379), .Z(n4524) );
  AOI22D0BWP12T U734 ( .A1(b[9]), .A2(n4658), .B1(n4657), .B2(n4482), .ZN(
        n3230) );
  AOI221D1BWP12T U735 ( .A1(n4661), .A2(b[10]), .B1(n4660), .B2(n4646), .C(
        n3230), .ZN(n4523) );
  OAI22D0BWP12T U736 ( .A1(b[11]), .A2(n4453), .B1(n4792), .B2(n4470), .ZN(
        n3231) );
  AOI21D0BWP12T U737 ( .A1(n4455), .A2(n4792), .B(n3231), .ZN(n4522) );
  CKND1BWP12T U738 ( .I(n4128), .ZN(n4639) );
  AOI22D0BWP12T U739 ( .A1(b[2]), .A2(n4637), .B1(n4636), .B2(n5210), .ZN(
        n3235) );
  AOI221D0BWP12T U740 ( .A1(n4640), .A2(b[1]), .B1(n4639), .B2(n4419), .C(
        n3235), .ZN(n4518) );
  AOI22D0BWP12T U741 ( .A1(b[4]), .A2(n4668), .B1(n4667), .B2(n5703), .ZN(
        n3236) );
  AOI221D0BWP12T U742 ( .A1(n4671), .A2(b[3]), .B1(n4670), .B2(n5136), .C(
        n3236), .ZN(n4517) );
  AOI22D0BWP12T U743 ( .A1(b[6]), .A2(n4632), .B1(n4631), .B2(n4555), .ZN(
        n3237) );
  AOI221D0BWP12T U744 ( .A1(n4635), .A2(b[5]), .B1(n4634), .B2(n4490), .C(
        n3237), .ZN(n4516) );
  FA1D0BWP12T U745 ( .A(n3240), .B(n3239), .CI(n3238), .CO(n4537), .S(n3242)
         );
  AOI22D0BWP12T U746 ( .A1(b[3]), .A2(n4632), .B1(n4631), .B2(n5136), .ZN(
        n3248) );
  AOI221D0BWP12T U747 ( .A1(n4635), .A2(b[2]), .B1(n4634), .B2(n5210), .C(
        n3248), .ZN(n3261) );
  RCOAI21D0BWP12T U748 ( .A1(n3251), .A2(n3250), .B(n3249), .ZN(n3260) );
  ND2D0BWP12T U749 ( .A1(b[0]), .A2(n4344), .ZN(n3274) );
  OAI22D0BWP12T U750 ( .A1(b[7]), .A2(n4453), .B1(n4699), .B2(n4470), .ZN(
        n3252) );
  AOI21D0BWP12T U751 ( .A1(n4455), .A2(n4699), .B(n3252), .ZN(n3273) );
  AOI22D0BWP12T U752 ( .A1(b[5]), .A2(n4658), .B1(n4657), .B2(n4490), .ZN(
        n3253) );
  AOI221D0BWP12T U753 ( .A1(n4661), .A2(b[6]), .B1(n4660), .B2(n4555), .C(
        n3253), .ZN(n3272) );
  OAI22D0BWP12T U754 ( .A1(b[4]), .A2(n4641), .B1(n3304), .B2(n3691), .ZN(
        n3255) );
  RCAOI21D0BWP12T U755 ( .A1(b[4]), .A2(n3302), .B(n3255), .ZN(n3276) );
  AOI22D0BWP12T U756 ( .A1(b[2]), .A2(n4632), .B1(n4631), .B2(n5210), .ZN(
        n3256) );
  AOI221D1BWP12T U757 ( .A1(n4635), .A2(b[1]), .B1(n4634), .B2(n4419), .C(
        n3256), .ZN(n3275) );
  AOI22D0BWP12T U758 ( .A1(n5380), .A2(n4555), .B1(n4455), .B2(n4450), .ZN(
        n3257) );
  OAI21D0BWP12T U759 ( .A1(n4450), .A2(n4470), .B(n3257), .ZN(n3279) );
  AOI22D0BWP12T U760 ( .A1(b[2]), .A2(n4645), .B1(n4644), .B2(n5210), .ZN(
        n3258) );
  OAI221D0BWP12T U761 ( .A1(b[3]), .A2(n4641), .B1(n5136), .B2(n4642), .C(
        n3258), .ZN(n3280) );
  ND2D1BWP12T U762 ( .A1(n3279), .A2(n3280), .ZN(n3278) );
  OAI22D1BWP12T U763 ( .A1(n5379), .A2(n3577), .B1(n3528), .B2(b[0]), .ZN(
        n3536) );
  OR2D0BWP12T U764 ( .A1(n4635), .A2(n4634), .Z(n4492) );
  AOI22D0BWP12T U765 ( .A1(b[1]), .A2(n4632), .B1(n4631), .B2(n4419), .ZN(
        n3270) );
  AOI21D0BWP12T U766 ( .A1(n3536), .A2(n4492), .B(n3270), .ZN(n3283) );
  AOI22D0BWP12T U767 ( .A1(b[4]), .A2(n4658), .B1(n4657), .B2(n5703), .ZN(
        n3271) );
  AOI221D0BWP12T U768 ( .A1(n4661), .A2(b[5]), .B1(n4660), .B2(n4490), .C(
        n3271), .ZN(n3281) );
  FA1D0BWP12T U769 ( .A(n3283), .B(n3282), .CI(n3281), .CO(n3328), .S(n3284)
         );
  AOI22D0BWP12T U770 ( .A1(n5380), .A2(n4490), .B1(n4455), .B2(n4555), .ZN(
        n3285) );
  OAI21D0BWP12T U771 ( .A1(n4555), .A2(n4470), .B(n3285), .ZN(n3293) );
  TPNR2D0BWP12T U772 ( .A1(n5379), .A2(n3286), .ZN(n3292) );
  AOI22D0BWP12T U773 ( .A1(b[1]), .A2(n4645), .B1(n4644), .B2(n4419), .ZN(
        n3287) );
  OAI221D0BWP12T U774 ( .A1(b[2]), .A2(n4641), .B1(n5210), .B2(n4642), .C(
        n3287), .ZN(n3291) );
  AO21D0BWP12T U775 ( .A1(n5379), .A2(n3301), .B(n4644), .Z(n3298) );
  AOI22D0BWP12T U776 ( .A1(n5380), .A2(n5703), .B1(n4455), .B2(n4490), .ZN(
        n3289) );
  OAI21D0BWP12T U777 ( .A1(n4490), .A2(n4470), .B(n3289), .ZN(n3299) );
  ND2D0BWP12T U778 ( .A1(n3298), .A2(n3299), .ZN(n3297) );
  AOI21D0BWP12T U779 ( .A1(n4658), .A2(n4657), .B(n3723), .ZN(n3290) );
  AOI221D1BWP12T U780 ( .A1(n4661), .A2(b[4]), .B1(n4660), .B2(n5703), .C(
        n3290), .ZN(n3296) );
  OAI22D1BWP12T U781 ( .A1(n5379), .A2(n3709), .B1(n3300), .B2(b[0]), .ZN(
        n3535) );
  AOI22D0BWP12T U782 ( .A1(b[1]), .A2(n3302), .B1(n3301), .B2(n4419), .ZN(
        n3303) );
  OAI21D0BWP12T U783 ( .A1(n3608), .A2(n3304), .B(n3303), .ZN(n3311) );
  OA22XD1BWP12T U784 ( .A1(n4657), .A2(b[2]), .B1(n5210), .B2(n4658), .Z(n3305) );
  OAI21D0BWP12T U785 ( .A1(n3723), .A2(n3320), .B(n3305), .ZN(n3310) );
  AOI22D0BWP12T U786 ( .A1(b[1]), .A2(n4658), .B1(n4657), .B2(n4419), .ZN(
        n3308) );
  AOI221D1BWP12T U787 ( .A1(n4661), .A2(b[2]), .B1(n4660), .B2(n5210), .C(
        n3308), .ZN(n3317) );
  OAI22D0BWP12T U788 ( .A1(b[3]), .A2(n4453), .B1(n5703), .B2(n4470), .ZN(
        n3309) );
  AOI21D0BWP12T U789 ( .A1(n4455), .A2(n5703), .B(n3309), .ZN(n3316) );
  OAI211D0BWP12T U790 ( .A1(n5210), .A2(a[0]), .B(n5198), .C(a[1]), .ZN(n3314)
         );
  OAI21D1BWP12T U791 ( .A1(a[1]), .A2(n5198), .B(n3314), .ZN(n3324) );
  TPAOI22D0BWP12T U792 ( .A1(b[1]), .A2(n4661), .B1(n4660), .B2(n4419), .ZN(
        n3315) );
  AOI32D0BWP12T U793 ( .A1(n4658), .A2(n3315), .A3(n4657), .B1(n3610), .B2(
        n3315), .ZN(n3323) );
  AOI32D1BWP12T U794 ( .A1(n3321), .A2(n5379), .A3(n4453), .B1(b[0]), .B2(
        n3320), .ZN(n3633) );
  CKND2D1BWP12T U795 ( .A1(n3634), .A2(n3633), .ZN(n3699) );
  CKND2D0BWP12T U796 ( .A1(a[3]), .A2(n5379), .ZN(n3710) );
  NR2D1BWP12T U797 ( .A1(n3356), .A2(n3504), .ZN(n5889) );
  OAI22D1BWP12T U798 ( .A1(n5368), .A2(n6130), .B1(n6048), .B2(n4742), .ZN(
        n3338) );
  RCAOI211D0BWP12T U799 ( .A1(n5621), .A2(n5516), .B(n3339), .C(n3338), .ZN(
        n3340) );
  OAI211D1BWP12T U800 ( .A1(n4999), .A2(n6138), .B(n3340), .C(n5635), .ZN(
        n3354) );
  CKND2D1BWP12T U801 ( .A1(n3697), .A2(n3709), .ZN(n3676) );
  NR2XD0BWP12T U802 ( .A1(a[5]), .A2(n3676), .ZN(n3601) );
  CKND2D1BWP12T U803 ( .A1(n3601), .A2(n3577), .ZN(n3576) );
  OAI21D1BWP12T U804 ( .A1(n3727), .A2(n6034), .B(n6092), .ZN(n3351) );
  INVD0BWP12T U805 ( .I(n3569), .ZN(n4983) );
  CKND2D0BWP12T U806 ( .A1(n3566), .A2(n5262), .ZN(n3345) );
  OAI211D1BWP12T U807 ( .A1(n3563), .A2(n5282), .B(n3346), .C(n3345), .ZN(
        n5227) );
  TPNR2D0BWP12T U808 ( .A1(n5703), .A2(n5136), .ZN(n5145) );
  CKND2D1BWP12T U809 ( .A1(n5143), .A2(n5086), .ZN(n5284) );
  TPAOI22D0BWP12T U810 ( .A1(n5254), .A2(n5191), .B1(n5255), .B2(n3567), .ZN(
        n3348) );
  CKND2D0BWP12T U811 ( .A1(n5193), .A2(n5262), .ZN(n3347) );
  OAI21D1BWP12T U812 ( .A1(n5092), .A2(n6115), .B(n5272), .ZN(n3350) );
  AOI22D1BWP12T U813 ( .A1(a[12]), .A2(n3351), .B1(n5620), .B2(n3350), .ZN(
        n3352) );
  CKND2D1BWP12T U814 ( .A1(n6151), .A2(n3727), .ZN(n3386) );
  AOI32D1BWP12T U815 ( .A1(n6156), .A2(n3352), .A3(n3386), .B1(a[12]), .B2(
        n3352), .ZN(n3353) );
  AOI211D1BWP12T U816 ( .A1(n6160), .A2(n4930), .B(n3354), .C(n3353), .ZN(
        n3367) );
  INVD1BWP12T U817 ( .I(c_in), .ZN(n4759) );
  CKND2D1BWP12T U818 ( .A1(b[10]), .A2(n3421), .ZN(n5455) );
  NR2D1BWP12T U819 ( .A1(n5633), .A2(n5379), .ZN(n5492) );
  MAOI222D1BWP12T U820 ( .A(n3675), .B(a[4]), .C(b[4]), .ZN(n3621) );
  INR2XD0BWP12T U821 ( .A1(n3607), .B1(n3621), .ZN(n3553) );
  OAI22D0BWP12T U822 ( .A1(n5394), .A2(n3553), .B1(a[6]), .B2(b[6]), .ZN(n3550) );
  NR2XD0BWP12T U823 ( .A1(n3533), .A2(n3526), .ZN(n4495) );
  MAOI222D1BWP12T U824 ( .A(a[8]), .B(b[8]), .C(n3475), .ZN(n3517) );
  MAOI222D1BWP12T U825 ( .A(n4482), .B(n3509), .C(n3517), .ZN(n3445) );
  CKND2D0BWP12T U826 ( .A1(n3445), .A2(n3420), .ZN(n3368) );
  ND2XD0BWP12T U827 ( .A1(n4741), .A2(n3749), .ZN(n4058) );
  AOI22D1BWP12T U828 ( .A1(n6122), .A2(n4774), .B1(n6162), .B2(n4875), .ZN(
        n3366) );
  OAI211D1BWP12T U829 ( .A1(n4826), .A2(n6120), .B(n3367), .C(n3366), .ZN(
        result[12]) );
  OAI21D0BWP12T U830 ( .A1(n5805), .A2(b[0]), .B(n5634), .ZN(n3534) );
  NR2XD0BWP12T U831 ( .A1(n3536), .A2(n5286), .ZN(n3370) );
  OAI22D0BWP12T U832 ( .A1(n3535), .A2(n5284), .B1(n3382), .B2(n5288), .ZN(
        n3369) );
  CKND2D1BWP12T U833 ( .A1(n5168), .A2(n6145), .ZN(n3427) );
  AOI22D1BWP12T U834 ( .A1(b[0]), .A2(n4738), .B1(n5901), .B2(n5379), .ZN(
        n3593) );
  OAI22D0BWP12T U835 ( .A1(n5379), .A2(a[28]), .B1(a[27]), .B2(b[0]), .ZN(
        n3481) );
  OR2D1BWP12T U836 ( .A1(n3537), .A2(b[2]), .Z(n3383) );
  NR2D0BWP12T U837 ( .A1(b[3]), .A2(n3383), .ZN(n5542) );
  CKND0BWP12T U838 ( .I(n5532), .ZN(n5523) );
  IAO21D0BWP12T U839 ( .A1(n5542), .A2(n5523), .B(n5528), .ZN(n5750) );
  CKND2D1BWP12T U840 ( .A1(n5210), .A2(b[3]), .ZN(n3663) );
  TPNR2D0BWP12T U841 ( .A1(n5379), .A2(n6155), .ZN(n3484) );
  CKND2D1BWP12T U842 ( .A1(a[19]), .A2(n5379), .ZN(n4266) );
  OAI22D1BWP12T U843 ( .A1(n5379), .A2(n5912), .B1(n5833), .B2(b[0]), .ZN(
        n5018) );
  CKND2D0BWP12T U844 ( .A1(n5018), .A2(n5086), .ZN(n5220) );
  CKND2D0BWP12T U845 ( .A1(n4419), .A2(a[23]), .ZN(n4008) );
  TPNR2D0BWP12T U846 ( .A1(n5379), .A2(b[1]), .ZN(n3480) );
  CKND2D0BWP12T U847 ( .A1(a[13]), .A2(n5379), .ZN(n3372) );
  AOI22D0BWP12T U848 ( .A1(b[0]), .A2(a[12]), .B1(a[11]), .B2(n5379), .ZN(
        n3489) );
  CKND2D1BWP12T U849 ( .A1(a[15]), .A2(n5379), .ZN(n4330) );
  OAI22D0BWP12T U850 ( .A1(n5379), .A2(a[18]), .B1(a[17]), .B2(b[0]), .ZN(
        n3373) );
  AOI22D0BWP12T U851 ( .A1(n5525), .A2(n3714), .B1(n5242), .B2(n3713), .ZN(
        n3374) );
  OA21XD0BWP12T U852 ( .A1(n5670), .A2(n5750), .B(n3384), .Z(n5558) );
  MOAI22D0BWP12T U853 ( .A1(n5147), .A2(n3427), .B1(n5826), .B2(n5558), .ZN(
        n3391) );
  OAI32D1BWP12T U854 ( .A1(a[11]), .A2(n4741), .A3(n6096), .B1(n6156), .B2(
        a[11]), .ZN(n3381) );
  OAI22D1BWP12T U855 ( .A1(n5358), .A2(n6130), .B1(n3378), .B2(n6092), .ZN(
        n3380) );
  OR4D1BWP12T U856 ( .A1(n5859), .A2(n3381), .A3(n3380), .A4(n3379), .Z(n3390)
         );
  ND2D1BWP12T U857 ( .A1(n5670), .A2(n6052), .ZN(n5631) );
  ND3D0BWP12T U858 ( .A1(n5136), .A2(n5143), .A3(n3705), .ZN(n5757) );
  AOI22D0BWP12T U859 ( .A1(n3393), .A2(n4889), .B1(n4148), .B2(n3385), .ZN(
        n4933) );
  AOI22D1BWP12T U860 ( .A1(n3393), .A2(n3392), .B1(n4148), .B2(n4745), .ZN(
        n4775) );
  AOI22D1BWP12T U861 ( .A1(n4775), .A2(n6122), .B1(n4823), .B2(n6164), .ZN(
        n3395) );
  OAI211D1BWP12T U862 ( .A1(n4876), .A2(n6126), .B(n3396), .C(n3395), .ZN(
        result[11]) );
  INVD1BWP12T U863 ( .I(n3446), .ZN(n3442) );
  MAOI22D0BWP12T U864 ( .A1(n3442), .A2(n3397), .B1(n3442), .B2(n3397), .ZN(
        n4771) );
  NR2D0BWP12T U865 ( .A1(a[25]), .A2(n5379), .ZN(n3399) );
  NR2XD0BWP12T U866 ( .A1(b[0]), .A2(a[18]), .ZN(n3402) );
  TPNR2D0BWP12T U867 ( .A1(a[19]), .A2(n5379), .ZN(n4970) );
  AOI22D1BWP12T U868 ( .A1(b[2]), .A2(n3570), .B1(n5121), .B2(n5210), .ZN(
        n3650) );
  NR2D0BWP12T U869 ( .A1(a[13]), .A2(n5379), .ZN(n3404) );
  NR2XD0BWP12T U870 ( .A1(b[0]), .A2(a[12]), .ZN(n3403) );
  AOI22D0BWP12T U871 ( .A1(b[0]), .A2(a[11]), .B1(a[10]), .B2(n5379), .ZN(
        n3451) );
  OAI22D1BWP12T U872 ( .A1(n5379), .A2(a[15]), .B1(a[16]), .B2(b[0]), .ZN(
        n5208) );
  NR2XD0BWP12T U873 ( .A1(n5208), .A2(n3572), .ZN(n5144) );
  NR2XD0BWP12T U874 ( .A1(n5679), .A2(n3405), .ZN(n3406) );
  NR2XD0BWP12T U875 ( .A1(n5118), .A2(n3707), .ZN(n3407) );
  ND3D0BWP12T U876 ( .A1(a[28]), .A2(b[1]), .A3(n5379), .ZN(n3408) );
  AO211D1BWP12T U877 ( .A1(a[10]), .A2(n3508), .B(n3410), .C(n6034), .Z(n3411)
         );
  OAI31D1BWP12T U878 ( .A1(n3412), .A2(n5498), .A3(n6115), .B(n3411), .ZN(
        n3441) );
  NR2D0BWP12T U879 ( .A1(b[0]), .A2(n5128), .ZN(n5098) );
  INVD1BWP12T U880 ( .I(n5028), .ZN(n3415) );
  AOI22D0BWP12T U881 ( .A1(n5095), .A2(n5122), .B1(n5051), .B2(n3564), .ZN(
        n3414) );
  TPAOI22D0BWP12T U882 ( .A1(n5057), .A2(n5123), .B1(n5052), .B2(n3565), .ZN(
        n3413) );
  AOI22D1BWP12T U883 ( .A1(b[3]), .A2(n3415), .B1(n5026), .B2(n5136), .ZN(
        n5011) );
  CKND2D0BWP12T U884 ( .A1(n5570), .A2(n5113), .ZN(n3432) );
  OAI22D1BWP12T U885 ( .A1(n5086), .A2(n3563), .B1(n3562), .B2(n5633), .ZN(
        n3646) );
  INR2D1BWP12T U886 ( .A1(n3646), .B1(n3568), .ZN(n5200) );
  NR2D0BWP12T U887 ( .A1(n3572), .A2(n3455), .ZN(n3416) );
  AOI22D0BWP12T U888 ( .A1(b[2]), .A2(n3416), .B1(n5255), .B2(n3564), .ZN(
        n3418) );
  AOI22D0BWP12T U889 ( .A1(n3565), .A2(n5192), .B1(n5123), .B2(n5262), .ZN(
        n3417) );
  OA211D1BWP12T U890 ( .A1(n3421), .A2(n6150), .B(n3420), .C(n3693), .Z(n3422)
         );
  RCAOI21D0BWP12T U891 ( .A1(n5374), .A2(n5341), .B(n3422), .ZN(n3426) );
  OAI222D1BWP12T U892 ( .A1(n6133), .A2(n3424), .B1(a[10]), .B2(n6074), .C1(
        n3423), .C2(n6045), .ZN(n3425) );
  OAI211D1BWP12T U893 ( .A1(n5084), .A2(n3427), .B(n3426), .C(n3425), .ZN(
        n3428) );
  AOI21D1BWP12T U894 ( .A1(n5507), .A2(n3429), .B(n3428), .ZN(n3438) );
  CKND2D0BWP12T U895 ( .A1(a[31]), .A2(n5528), .ZN(n3433) );
  OAI22D0BWP12T U896 ( .A1(n3482), .A2(n4738), .B1(n5593), .B2(n3430), .ZN(
        n5524) );
  IAO21D1BWP12T U897 ( .A1(n5210), .A2(n5524), .B(n3431), .ZN(n3652) );
  CKND2D0BWP12T U898 ( .A1(n3652), .A2(n5136), .ZN(n5540) );
  CKND2D0BWP12T U899 ( .A1(n3435), .A2(n3434), .ZN(n3436) );
  MAOI22D0BWP12T U900 ( .A1(n3442), .A2(n3436), .B1(n3442), .B2(n3436), .ZN(
        n4929) );
  TPAOI22D0BWP12T U901 ( .A1(n5826), .A2(n5557), .B1(n6160), .B2(n4929), .ZN(
        n3437) );
  OAI211D1BWP12T U902 ( .A1(n3439), .A2(n5631), .B(n3438), .C(n3437), .ZN(
        n3440) );
  AOI22D1BWP12T U903 ( .A1(n3444), .A2(n3446), .B1(n3443), .B2(n3442), .ZN(
        n4822) );
  RCAOI22D0BWP12T U904 ( .A1(n6164), .A2(n4822), .B1(n6162), .B2(n4874), .ZN(
        n3447) );
  OAI211D1BWP12T U905 ( .A1(n4771), .A2(n6167), .B(n3448), .C(n3447), .ZN(
        result[10]) );
  CKND2D0BWP12T U906 ( .A1(a[8]), .A2(n5379), .ZN(n3452) );
  AOI32D1BWP12T U907 ( .A1(n3573), .A2(n4419), .A3(n3452), .B1(n3451), .B2(
        b[1]), .ZN(n5135) );
  AOI22D1BWP12T U908 ( .A1(n5525), .A2(n5135), .B1(n5238), .B2(n5105), .ZN(
        n3453) );
  INVD1BWP12T U909 ( .I(n5889), .ZN(n6093) );
  OAI22D1BWP12T U910 ( .A1(n3457), .A2(n6092), .B1(a[8]), .B2(n6156), .ZN(
        n3460) );
  INVD0BWP12T U911 ( .I(n3473), .ZN(n3474) );
  OAI22D1BWP12T U912 ( .A1(n3458), .A2(n6128), .B1(n3474), .B2(n6096), .ZN(
        n3459) );
  RCAOI211D0BWP12T U913 ( .A1(n5338), .A2(n5374), .B(n3460), .C(n3459), .ZN(
        n3465) );
  AOI22D0BWP12T U914 ( .A1(n5057), .A2(n5122), .B1(n5095), .B2(n3565), .ZN(
        n3462) );
  AOI22D0BWP12T U915 ( .A1(n5052), .A2(n3564), .B1(n5051), .B2(n3563), .ZN(
        n3461) );
  CKND2D1BWP12T U916 ( .A1(n3462), .A2(n3461), .ZN(n5055) );
  RCOAI22D0BWP12T U917 ( .A1(n5055), .A2(n5070), .B1(n5062), .B2(n5068), .ZN(
        n5044) );
  CKND1BWP12T U918 ( .I(n3576), .ZN(n3529) );
  ND2XD0BWP12T U919 ( .A1(n3529), .A2(n3528), .ZN(n3527) );
  AOI211D1BWP12T U920 ( .A1(a[8]), .A2(n3527), .B(n3510), .C(n6034), .ZN(n3463) );
  RCAOI211D0BWP12T U921 ( .A1(n6052), .A2(n5044), .B(n3463), .C(n5859), .ZN(
        n3464) );
  OAI211D1BWP12T U922 ( .A1(n3466), .A2(n6093), .B(n3465), .C(n3464), .ZN(
        n3471) );
  AOI21D0BWP12T U923 ( .A1(b[4]), .A2(n5925), .B(n5528), .ZN(n5512) );
  ND2D0BWP12T U924 ( .A1(n5830), .A2(n5866), .ZN(n3636) );
  NR2D0BWP12T U925 ( .A1(n5136), .A2(n5669), .ZN(n5837) );
  AOI211D1BWP12T U926 ( .A1(n5512), .A2(n3636), .B(n5815), .C(n5837), .ZN(
        n3468) );
  OAI22D1BWP12T U927 ( .A1(n3469), .A2(n3468), .B1(n4927), .B2(n6113), .ZN(
        n3470) );
  AOI211XD0BWP12T U928 ( .A1(n6145), .A2(n5219), .B(n3471), .C(n3470), .ZN(
        n3477) );
  OAI211D1BWP12T U929 ( .A1(n4817), .A2(n6120), .B(n3477), .C(n3476), .ZN(
        result[8]) );
  MAOI22D0BWP12T U930 ( .A1(n4343), .A2(n3478), .B1(n4343), .B2(n3478), .ZN(
        n4821) );
  CKND0BWP12T U931 ( .I(n3480), .ZN(n3493) );
  OAI222D1BWP12T U932 ( .A1(n3482), .A2(n5833), .B1(n4419), .B2(n3481), .C1(
        n5787), .C2(n3493), .ZN(n5237) );
  TPND2D0BWP12T U933 ( .A1(n5136), .A2(n5531), .ZN(n5848) );
  CKND0BWP12T U934 ( .I(n3483), .ZN(n4957) );
  CKND2D0BWP12T U935 ( .A1(n3562), .A2(n4957), .ZN(n3486) );
  AOI222D1BWP12T U936 ( .A1(n4009), .A2(n3486), .B1(a[24]), .B2(n3485), .C1(
        n4419), .C2(n3484), .ZN(n3594) );
  NR2XD0BWP12T U937 ( .A1(n5872), .A2(b[1]), .ZN(n4378) );
  CKND2D0BWP12T U938 ( .A1(n4330), .A2(n3487), .ZN(n4974) );
  NR2D0BWP12T U939 ( .A1(n3572), .A2(n5181), .ZN(n5253) );
  CKND2D1BWP12T U940 ( .A1(b[0]), .A2(a[10]), .ZN(n3539) );
  AOI32D1BWP12T U941 ( .A1(n3490), .A2(n4419), .A3(n3539), .B1(n3489), .B2(
        b[1]), .ZN(n5100) );
  CKND2D1BWP12T U942 ( .A1(b[0]), .A2(a[18]), .ZN(n3491) );
  CKND2D0BWP12T U943 ( .A1(a[17]), .A2(n4419), .ZN(n4328) );
  CKND2D0BWP12T U944 ( .A1(n4328), .A2(n4956), .ZN(n3492) );
  AOI22D0BWP12T U945 ( .A1(n5525), .A2(n5100), .B1(n5240), .B2(n5241), .ZN(
        n3494) );
  AOI211XD0BWP12T U946 ( .A1(n3496), .A2(n5848), .B(n5500), .C(n5528), .ZN(
        n5548) );
  AOI32D1BWP12T U947 ( .A1(a[31]), .A2(b[1]), .A3(n5379), .B1(n3593), .B2(
        n4419), .ZN(n5274) );
  AO21D0BWP12T U948 ( .A1(b[2]), .A2(n5274), .B(n3497), .Z(n5138) );
  INVD1BWP12T U949 ( .I(n5870), .ZN(n5646) );
  CKND2D0BWP12T U950 ( .A1(n5262), .A2(n3534), .ZN(n5269) );
  NR2D0BWP12T U951 ( .A1(n5131), .A2(n3609), .ZN(n5816) );
  NR2D0BWP12T U952 ( .A1(n5131), .A2(n5085), .ZN(n3501) );
  OAI22D0BWP12T U953 ( .A1(n5128), .A2(n3536), .B1(n5047), .B2(n3535), .ZN(
        n3500) );
  AO211D0BWP12T U954 ( .A1(n3610), .A2(n5051), .B(n3501), .C(n3500), .Z(n5066)
         );
  OAI22D1BWP12T U955 ( .A1(n4211), .A2(n6096), .B1(a[9]), .B2(n6156), .ZN(
        n3507) );
  AOI21D0BWP12T U956 ( .A1(b[9]), .A2(n5622), .B(n3503), .ZN(n3505) );
  OR2XD0BWP12T U957 ( .A1(op[0]), .A2(n3504), .Z(n5671) );
  OAI22D1BWP12T U958 ( .A1(n3505), .A2(n5671), .B1(n5387), .B2(n6128), .ZN(
        n3506) );
  RCAOI211D0BWP12T U959 ( .A1(n5339), .A2(n5374), .B(n3507), .C(n3506), .ZN(
        n3512) );
  OAI211D1BWP12T U960 ( .A1(n3510), .A2(n3509), .B(n6151), .C(n3508), .ZN(
        n3511) );
  OAI211D1BWP12T U961 ( .A1(n3513), .A2(n5631), .B(n3512), .C(n3511), .ZN(
        n3514) );
  RCAOI211D0BWP12T U962 ( .A1(n6145), .A2(n5140), .B(n5859), .C(n3514), .ZN(
        n3515) );
  OAI211D1BWP12T U963 ( .A1(n4924), .A2(n6113), .B(n3516), .C(n3515), .ZN(
        n3520) );
  OAI22D1BWP12T U964 ( .A1(n4871), .A2(n6126), .B1(n6167), .B2(n4770), .ZN(
        n3519) );
  AO211D1BWP12T U965 ( .A1(n6164), .A2(n4821), .B(n3520), .C(n3519), .Z(
        result[9]) );
  AOI22D0BWP12T U966 ( .A1(n4495), .A2(n3522), .B1(n3549), .B2(n3521), .ZN(
        n4763) );
  AOI21D0BWP12T U967 ( .A1(n3526), .A2(n6045), .B(n6150), .ZN(n3532) );
  OAI211D0BWP12T U968 ( .A1(n3529), .A2(n3528), .B(n6151), .C(n3527), .ZN(
        n3530) );
  OAI211D1BWP12T U969 ( .A1(n3533), .A2(n3532), .B(n3531), .C(n3530), .ZN(
        n3546) );
  AOI22D1BWP12T U970 ( .A1(n5024), .A2(n5817), .B1(n5698), .B2(n5608), .ZN(
        n3544) );
  TPND2D0BWP12T U971 ( .A1(n5136), .A2(n5078), .ZN(n3541) );
  CKND0BWP12T U972 ( .I(n3541), .ZN(n5533) );
  OAI22D0BWP12T U973 ( .A1(n5210), .A2(n3706), .B1(n3713), .B2(b[2]), .ZN(
        n5080) );
  CKND2D0BWP12T U974 ( .A1(a[7]), .A2(n5379), .ZN(n3595) );
  AOI32D1BWP12T U975 ( .A1(n3595), .A2(n3572), .A3(n3539), .B1(n5086), .B2(
        n5178), .ZN(n3715) );
  OA21XD1BWP12T U976 ( .A1(n5521), .A2(n5533), .B(n5109), .Z(n5518) );
  MAOI22D0BWP12T U977 ( .A1(n3540), .A2(n3549), .B1(n3540), .B2(n3549), .ZN(
        n4921) );
  AOI22D0BWP12T U978 ( .A1(n5621), .A2(n5518), .B1(n6160), .B2(n4921), .ZN(
        n3543) );
  OAI211D1BWP12T U979 ( .A1(n5703), .A2(n5937), .B(n5109), .C(n5620), .ZN(
        n3542) );
  ND3D1BWP12T U980 ( .A1(n3544), .A2(n3543), .A3(n3542), .ZN(n3545) );
  NR4D0BWP12T U981 ( .A1(n5859), .A2(n3547), .A3(n3546), .A4(n3545), .ZN(n3552) );
  MAOI22D0BWP12T U982 ( .A1(n3549), .A2(n3548), .B1(n3549), .B2(n3548), .ZN(
        n4815) );
  RCAOI22D0BWP12T U983 ( .A1(n6164), .A2(n4815), .B1(n6162), .B2(n4866), .ZN(
        n3551) );
  OAI211D1BWP12T U984 ( .A1(n4763), .A2(n6167), .B(n3552), .C(n3551), .ZN(
        result[7]) );
  NR2D0BWP12T U985 ( .A1(n3553), .A2(n3600), .ZN(n3554) );
  MAOI22D0BWP12T U986 ( .A1(n3554), .A2(n3589), .B1(n3554), .B2(n3589), .ZN(
        n4869) );
  AOI22D0BWP12T U987 ( .A1(n6045), .A2(n3558), .B1(n6074), .B2(n3577), .ZN(
        n3557) );
  OAI211D1BWP12T U988 ( .A1(n5311), .A2(n6130), .B(n3557), .C(n5635), .ZN(
        n3561) );
  OAI22D0BWP12T U989 ( .A1(n3558), .A2(n6096), .B1(b[6]), .B2(n6093), .ZN(
        n3560) );
  TPND2D0BWP12T U990 ( .A1(n3577), .A2(n4555), .ZN(n3559) );
  OAI32D0BWP12T U991 ( .A1(n3561), .A2(n6150), .A3(n3560), .B1(n3559), .B2(
        n3561), .ZN(n3581) );
  AOI22D1BWP12T U992 ( .A1(n5008), .A2(n5817), .B1(n5698), .B2(n6111), .ZN(
        n3580) );
  CKND0BWP12T U993 ( .I(n5277), .ZN(n5117) );
  AOI22D0BWP12T U994 ( .A1(b[2]), .A2(n3571), .B1(n3570), .B2(n5210), .ZN(
        n5119) );
  NR2XD0BWP12T U995 ( .A1(b[3]), .A2(n5119), .ZN(n5273) );
  CKND2D0BWP12T U996 ( .A1(a[6]), .A2(n5379), .ZN(n3660) );
  AOI32D1BWP12T U997 ( .A1(n3573), .A2(n3572), .A3(n3660), .B1(n5122), .B2(
        n5086), .ZN(n3625) );
  AOI22D0BWP12T U998 ( .A1(n5242), .A2(n3630), .B1(n5238), .B2(n5121), .ZN(
        n3574) );
  TPOAI21D0BWP12T U999 ( .A1(n5118), .A2(n3663), .B(n3574), .ZN(n3575) );
  RCAOI211D0BWP12T U1000 ( .A1(n5525), .A2(n3625), .B(b[4]), .C(n3575), .ZN(
        n5116) );
  OAI211D1BWP12T U1001 ( .A1(n5539), .A2(n3584), .B(n5621), .C(n3583), .ZN(
        n3579) );
  OAI211D0BWP12T U1002 ( .A1(n3601), .A2(n3577), .B(n6151), .C(n3576), .ZN(
        n3578) );
  ND4D1BWP12T U1003 ( .A1(n3581), .A2(n3580), .A3(n3579), .A4(n3578), .ZN(
        n3586) );
  MAOI22D0BWP12T U1004 ( .A1(n3582), .A2(n3589), .B1(n3582), .B2(n3589), .ZN(
        n4926) );
  MAOI22D0BWP12T U1005 ( .A1(n3589), .A2(n3587), .B1(n3589), .B2(n3587), .ZN(
        n4767) );
  OAI211D1BWP12T U1006 ( .A1(n4869), .A2(n6126), .B(n3591), .C(n3590), .ZN(
        result[6]) );
  MAOI22D0BWP12T U1007 ( .A1(n3622), .A2(n3592), .B1(n3622), .B2(n3592), .ZN(
        n4819) );
  OAI22D0BWP12T U1008 ( .A1(n5131), .A2(n3593), .B1(a[31]), .B2(n5057), .ZN(
        n5519) );
  CKND0BWP12T U1009 ( .I(n3594), .ZN(n5239) );
  AOI22D1BWP12T U1010 ( .A1(n5525), .A2(n5239), .B1(n5242), .B2(n5237), .ZN(
        n3614) );
  OAI21D0BWP12T U1011 ( .A1(n5519), .A2(n5136), .B(n3614), .ZN(n5972) );
  CKND2D1BWP12T U1012 ( .A1(b[0]), .A2(a[8]), .ZN(n3596) );
  OAI22D0BWP12T U1013 ( .A1(n5379), .A2(a[6]), .B1(a[5]), .B2(b[0]), .ZN(n3711) );
  AOI32D1BWP12T U1014 ( .A1(n3596), .A2(b[1]), .A3(n3595), .B1(n3711), .B2(
        n4419), .ZN(n5096) );
  TPAOI22D0BWP12T U1015 ( .A1(n5525), .A2(n5096), .B1(n5238), .B2(n5241), .ZN(
        n3597) );
  AOI22D0BWP12T U1016 ( .A1(n3600), .A2(n6045), .B1(n5447), .B2(n6133), .ZN(
        n3613) );
  OAI21D0BWP12T U1017 ( .A1(a[5]), .A2(n6096), .B(n6092), .ZN(n3606) );
  RCAOI211D0BWP12T U1018 ( .A1(a[5]), .A2(n3676), .B(n3601), .C(n6034), .ZN(
        n3605) );
  OAI22D0BWP12T U1019 ( .A1(n5348), .A2(n6130), .B1(a[5]), .B2(n6156), .ZN(
        n3604) );
  RCAOI211D0BWP12T U1020 ( .A1(n3607), .A2(n3606), .B(n3605), .C(n3604), .ZN(
        n3612) );
  ND4D1BWP12T U1021 ( .A1(n3613), .A2(n3612), .A3(n3611), .A4(n5635), .ZN(
        n3618) );
  MAOI22D0BWP12T U1022 ( .A1(n3622), .A2(n3616), .B1(n3622), .B2(n3616), .ZN(
        n4922) );
  AOI211XD0BWP12T U1023 ( .A1(n5551), .A2(n5621), .B(n3618), .C(n3617), .ZN(
        n3624) );
  MAOI22D0BWP12T U1024 ( .A1(n3620), .A2(n3619), .B1(n3620), .B2(n3619), .ZN(
        n4768) );
  AOI22D0BWP12T U1025 ( .A1(n6122), .A2(n4768), .B1(n6162), .B2(n4867), .ZN(
        n3623) );
  OAI211D1BWP12T U1026 ( .A1(n4819), .A2(n6120), .B(n3624), .C(n3623), .ZN(
        result[5]) );
  AOI22D0BWP12T U1027 ( .A1(b[0]), .A2(a[3]), .B1(a[2]), .B2(n5379), .ZN(n5127) );
  OAI22D0BWP12T U1028 ( .A1(n5379), .A2(a[5]), .B1(a[4]), .B2(b[0]), .ZN(n3659) );
  MOAI22D0BWP12T U1029 ( .A1(n3625), .A2(n5210), .B1(n3659), .B2(n5095), .ZN(
        n3626) );
  RCAOI211D0BWP12T U1030 ( .A1(n5057), .A2(n5127), .B(b[3]), .C(n3626), .ZN(
        n3629) );
  NR2XD0BWP12T U1031 ( .A1(n5118), .A2(n3627), .ZN(n3628) );
  MOAI22D0BWP12T U1032 ( .A1(n3632), .A2(n3631), .B1(n3632), .B2(n3631), .ZN(
        n4863) );
  OAI22D1BWP12T U1033 ( .A1(n4863), .A2(n6126), .B1(n5410), .B2(n6130), .ZN(
        n3635) );
  AOI31D1BWP12T U1034 ( .A1(n5670), .A2(n3645), .A3(n3636), .B(n3635), .ZN(
        n3657) );
  MAOI22D0BWP12T U1035 ( .A1(n3640), .A2(n3637), .B1(n3640), .B2(n3637), .ZN(
        n4814) );
  IND2XD0BWP12T U1036 ( .A1(n5070), .B1(n5028), .ZN(n5009) );
  MAOI22D0BWP12T U1037 ( .A1(n4814), .A2(n6164), .B1(n6138), .B2(n5009), .ZN(
        n3656) );
  MAOI22D0BWP12T U1038 ( .A1(n3640), .A2(n3638), .B1(n3640), .B2(n3638), .ZN(
        n4760) );
  MAOI22D0BWP12T U1039 ( .A1(n3640), .A2(n3639), .B1(n3640), .B2(n3639), .ZN(
        n4919) );
  TPAOI22D0BWP12T U1040 ( .A1(n6045), .A2(n5384), .B1(n6074), .B2(n5421), .ZN(
        n3644) );
  CKND2D0BWP12T U1041 ( .A1(n5633), .A2(n5805), .ZN(n5808) );
  MOAI22D0BWP12T U1042 ( .A1(n5210), .A2(n6092), .B1(n5471), .B2(n6135), .ZN(
        n3641) );
  AOI31D0BWP12T U1043 ( .A1(n6151), .A2(n3698), .A3(n3642), .B(n3641), .ZN(
        n3643) );
  OAI211D1BWP12T U1044 ( .A1(n4919), .A2(n6113), .B(n3644), .C(n3643), .ZN(
        n3649) );
  TPNR2D0BWP12T U1045 ( .A1(n5136), .A2(n5143), .ZN(n3720) );
  AOI32D1BWP12T U1046 ( .A1(n6133), .A2(a[2]), .A3(n5210), .B1(n6150), .B2(
        a[2]), .ZN(n3647) );
  OAI211D1BWP12T U1047 ( .A1(n6115), .A2(n5091), .B(n5635), .C(n3647), .ZN(
        n3648) );
  RCAOI211D0BWP12T U1048 ( .A1(n4760), .A2(n6122), .B(n3649), .C(n3648), .ZN(
        n3655) );
  CKND2D0BWP12T U1049 ( .A1(n5136), .A2(n3650), .ZN(n3651) );
  OAI21D1BWP12T U1050 ( .A1(n3652), .A2(n5136), .B(n3651), .ZN(n6008) );
  NR2XD0BWP12T U1051 ( .A1(n3653), .A2(n6008), .ZN(n5517) );
  AOI22D1BWP12T U1052 ( .A1(n5494), .A2(n5620), .B1(n5517), .B2(n5621), .ZN(
        n3654) );
  ND4D1BWP12T U1053 ( .A1(n3657), .A2(n3656), .A3(n3655), .A4(n3654), .ZN(
        result[2]) );
  OAI21D0BWP12T U1054 ( .A1(n5136), .A2(n4599), .B(n6071), .ZN(n5536) );
  AOI32D0BWP12T U1055 ( .A1(n3661), .A2(b[1]), .A3(n3660), .B1(n3659), .B2(
        n4419), .ZN(n5129) );
  AOI22D0BWP12T U1056 ( .A1(n5525), .A2(n5129), .B1(n5242), .B2(n5135), .ZN(
        n3662) );
  OAI21D1BWP12T U1057 ( .A1(n3664), .A2(n3663), .B(n3662), .ZN(n3665) );
  AOI211XD0BWP12T U1058 ( .A1(b[4]), .A2(n3666), .B(n5112), .C(n5528), .ZN(
        n5550) );
  NR2XD0BWP12T U1059 ( .A1(b[4]), .A2(a[4]), .ZN(n3667) );
  INVD1BWP12T U1060 ( .I(n3693), .ZN(n5939) );
  RCAOI211D0BWP12T U1061 ( .A1(a[4]), .A2(n6092), .B(n3667), .C(n5939), .ZN(
        n3673) );
  TPOAI22D0BWP12T U1062 ( .A1(a[4]), .A2(n6156), .B1(n6048), .B2(n5444), .ZN(
        n3672) );
  OAI22D1BWP12T U1063 ( .A1(n5310), .A2(n6130), .B1(n5386), .B2(n6128), .ZN(
        n3671) );
  NR4D0BWP12T U1064 ( .A1(n5859), .A2(n3673), .A3(n3672), .A4(n3671), .ZN(
        n3680) );
  AOI22D0BWP12T U1065 ( .A1(n3675), .A2(n3685), .B1(n3674), .B2(n3682), .ZN(
        n4868) );
  INVD1BWP12T U1066 ( .I(n5227), .ZN(n5213) );
  NR2XD0BWP12T U1067 ( .A1(n5213), .A2(n5263), .ZN(n5157) );
  AOI22D0BWP12T U1068 ( .A1(n4868), .A2(n6162), .B1(n5157), .B2(n6145), .ZN(
        n3679) );
  OAI211D1BWP12T U1069 ( .A1(n3697), .A2(n3709), .B(n6151), .C(n3676), .ZN(
        n3677) );
  ND4D1BWP12T U1070 ( .A1(n3680), .A2(n3679), .A3(n3678), .A4(n3677), .ZN(
        n3689) );
  MAOI22D0BWP12T U1071 ( .A1(n3682), .A2(n3681), .B1(n3682), .B2(n3681), .ZN(
        n4762) );
  MOAI22D0BWP12T U1072 ( .A1(n3683), .A2(n3685), .B1(n3683), .B2(n3685), .ZN(
        n4923) );
  MOAI22D0BWP12T U1073 ( .A1(n3685), .A2(n3684), .B1(n3685), .B2(n3684), .ZN(
        n4813) );
  AOI22D0BWP12T U1074 ( .A1(n4923), .A2(n6160), .B1(n6164), .B2(n4813), .ZN(
        n3687) );
  AO211D1BWP12T U1075 ( .A1(n6071), .A2(b[4]), .B(n5112), .C(n5600), .Z(n3686)
         );
  OAI211D1BWP12T U1076 ( .A1(n6167), .A2(n4762), .B(n3687), .C(n3686), .ZN(
        n3688) );
  AO211D1BWP12T U1077 ( .A1(n5550), .A2(n5826), .B(n3689), .C(n3688), .Z(
        result[4]) );
  MAOI22D0BWP12T U1078 ( .A1(n3691), .A2(n3690), .B1(n3691), .B2(n3690), .ZN(
        n4864) );
  MAOI22D0BWP12T U1079 ( .A1(n3692), .A2(n3691), .B1(n3692), .B2(n3691), .ZN(
        n4918) );
  AOI22D1BWP12T U1080 ( .A1(n5385), .A2(n6045), .B1(n5440), .B2(n6133), .ZN(
        n3695) );
  AOI22D1BWP12T U1081 ( .A1(n6150), .A2(a[3]), .B1(n3693), .B2(n5472), .ZN(
        n3694) );
  OAI211D1BWP12T U1082 ( .A1(n4918), .A2(n6113), .B(n3695), .C(n3694), .ZN(
        n3704) );
  MAOI22D0BWP12T U1083 ( .A1(n3723), .A2(n3696), .B1(n3723), .B2(n3696), .ZN(
        n4811) );
  RCAOI211D0BWP12T U1084 ( .A1(a[3]), .A2(n3698), .B(n3697), .C(n6034), .ZN(
        n3701) );
  OAI22D1BWP12T U1085 ( .A1(a[3]), .A2(n6156), .B1(n5373), .B2(n6130), .ZN(
        n3700) );
  AOI211D1BWP12T U1086 ( .A1(n5817), .A2(n5032), .B(n3701), .C(n3700), .ZN(
        n3702) );
  OAI211D1BWP12T U1087 ( .A1(n6120), .A2(n4811), .B(n3702), .C(n5635), .ZN(
        n3703) );
  OAI222D1BWP12T U1088 ( .A1(n3708), .A2(n3707), .B1(n5245), .B2(n3706), .C1(
        n5136), .C2(n3705), .ZN(n5996) );
  TPNR2D0BWP12T U1089 ( .A1(n5379), .A2(n3709), .ZN(n5094) );
  MAOI22D0BWP12T U1090 ( .A1(n5057), .A2(n3712), .B1(n5128), .B2(n3711), .ZN(
        n3718) );
  AOI22D1BWP12T U1091 ( .A1(n5242), .A2(n3715), .B1(n5240), .B2(n3714), .ZN(
        n3716) );
  CKND1BWP12T U1092 ( .I(n3721), .ZN(n3719) );
  NR2D1BWP12T U1093 ( .A1(n3720), .A2(n5996), .ZN(n5110) );
  MAOI22D0BWP12T U1094 ( .A1(n3723), .A2(n3722), .B1(n3723), .B2(n3722), .ZN(
        n4761) );
  AOI21D1BWP12T U1095 ( .A1(n5549), .A2(n5826), .B(n3724), .ZN(n3725) );
  OAI211D1BWP12T U1096 ( .A1(n4864), .A2(n6126), .B(n3726), .C(n3725), .ZN(
        result[3]) );
  INVD1BWP12T U1097 ( .I(b[31]), .ZN(n5595) );
  OAI22D1BWP12T U1098 ( .A1(n5595), .A2(a[31]), .B1(n5593), .B2(b[31]), .ZN(
        n5457) );
  ND2D1BWP12T U1099 ( .A1(n6113), .A2(n6167), .ZN(n5582) );
  NR2D1BWP12T U1100 ( .A1(a[12]), .A2(n3727), .ZN(n5873) );
  NR2D1BWP12T U1101 ( .A1(a[14]), .A2(a[13]), .ZN(n3747) );
  ND2D1BWP12T U1102 ( .A1(n5873), .A2(n3747), .ZN(n6036) );
  NR2D1BWP12T U1103 ( .A1(a[15]), .A2(n6036), .ZN(n6035) );
  INVD1BWP12T U1104 ( .I(a[16]), .ZN(n5710) );
  ND2D1BWP12T U1105 ( .A1(n6035), .A2(n5710), .ZN(n5709) );
  INVD1BWP12T U1106 ( .I(a[18]), .ZN(n6024) );
  ND2D1BWP12T U1107 ( .A1(n6024), .A2(n5679), .ZN(n4267) );
  NR2D1BWP12T U1108 ( .A1(n5709), .A2(n4267), .ZN(n5984) );
  INVD1BWP12T U1109 ( .I(a[20]), .ZN(n6082) );
  INVD1BWP12T U1110 ( .I(a[19]), .ZN(n5988) );
  ND2D1BWP12T U1111 ( .A1(n6082), .A2(n5988), .ZN(n4173) );
  INVD1BWP12T U1112 ( .I(n4173), .ZN(n3729) );
  ND2D1BWP12T U1113 ( .A1(n5984), .A2(n3729), .ZN(n6081) );
  NR2D1BWP12T U1114 ( .A1(a[21]), .A2(n6081), .ZN(n6152) );
  NR2D1BWP12T U1115 ( .A1(a[23]), .A2(a[22]), .ZN(n3751) );
  ND2D1BWP12T U1116 ( .A1(n6152), .A2(n3751), .ZN(n5734) );
  INVD1BWP12T U1117 ( .I(n5734), .ZN(n5950) );
  ND4D1BWP12T U1118 ( .A1(n5901), .A2(n5833), .A3(n5912), .A4(n5950), .ZN(
        n5564) );
  NR2D1BWP12T U1119 ( .A1(a[27]), .A2(a[26]), .ZN(n5733) );
  INVD1BWP12T U1120 ( .I(n5733), .ZN(n5736) );
  NR2D1BWP12T U1121 ( .A1(a[28]), .A2(n5736), .ZN(n5900) );
  IND2D1BWP12T U1122 ( .A1(n5564), .B1(n5900), .ZN(n5493) );
  NR2D1BWP12T U1123 ( .A1(a[30]), .A2(n5493), .ZN(n5581) );
  ND2D1BWP12T U1124 ( .A1(a[31]), .A2(n5581), .ZN(n5611) );
  NR2D1BWP12T U1125 ( .A1(n5611), .A2(n6034), .ZN(n4736) );
  OAI22D1BWP12T U1126 ( .A1(n5787), .A2(a[25]), .B1(n5833), .B2(a[26]), .ZN(
        n4557) );
  AOI22D1BWP12T U1127 ( .A1(a[27]), .A2(b[2]), .B1(n5210), .B2(n5758), .ZN(
        n3746) );
  ND2D1BWP12T U1128 ( .A1(a[27]), .A2(a[26]), .ZN(n5415) );
  IND2D1BWP12T U1129 ( .A1(n4557), .B1(n5415), .ZN(n3777) );
  NR2D1BWP12T U1130 ( .A1(n5733), .A2(n3777), .ZN(n4558) );
  AO21D1BWP12T U1131 ( .A1(a[27]), .A2(n4419), .B(n3728), .Z(n3778) );
  AOI22D1BWP12T U1132 ( .A1(n4557), .A2(n3746), .B1(n4558), .B2(n3778), .ZN(
        n3874) );
  OAI22D1BWP12T U1133 ( .A1(n5912), .A2(a[23]), .B1(n5951), .B2(a[24]), .ZN(
        n3973) );
  AOI22D1BWP12T U1134 ( .A1(a[25]), .A2(b[4]), .B1(n5703), .B2(n5833), .ZN(
        n3741) );
  INVD1BWP12T U1135 ( .I(n3973), .ZN(n4701) );
  ND2D1BWP12T U1136 ( .A1(a[25]), .A2(a[24]), .ZN(n5416) );
  OAI211D1BWP12T U1137 ( .A1(a[25]), .A2(a[24]), .B(n4701), .C(n5416), .ZN(
        n4702) );
  INVD1BWP12T U1138 ( .I(n4702), .ZN(n3966) );
  AOI22D1BWP12T U1139 ( .A1(a[25]), .A2(b[3]), .B1(n5136), .B2(n5833), .ZN(
        n3891) );
  AOI22D1BWP12T U1140 ( .A1(n3973), .A2(n3741), .B1(n3966), .B2(n3891), .ZN(
        n3873) );
  NR2D1BWP12T U1141 ( .A1(n6082), .A2(n5988), .ZN(n5413) );
  AN2D1BWP12T U1142 ( .A1(n5413), .A2(n5964), .Z(n4676) );
  NR2D1BWP12T U1143 ( .A1(n5964), .A2(n4173), .ZN(n4675) );
  NR2D1BWP12T U1144 ( .A1(n3729), .A2(n5413), .ZN(n4236) );
  ND2D1BWP12T U1145 ( .A1(n4236), .A2(n5964), .ZN(n4673) );
  ND2D1BWP12T U1146 ( .A1(a[21]), .A2(n4236), .ZN(n4672) );
  AOI22D1BWP12T U1147 ( .A1(b[8]), .A2(n4673), .B1(n4672), .B2(n4699), .ZN(
        n3730) );
  AOI221D1BWP12T U1148 ( .A1(n4676), .A2(b[7]), .B1(n4675), .B2(n4450), .C(
        n3730), .ZN(n3872) );
  INVD1BWP12T U1149 ( .I(a[28]), .ZN(n5737) );
  AOI22D1BWP12T U1150 ( .A1(a[28]), .A2(a[27]), .B1(n5758), .B2(n5737), .ZN(
        n4694) );
  ND2D1BWP12T U1151 ( .A1(b[0]), .A2(n4694), .ZN(n3889) );
  OA211D1BWP12T U1152 ( .A1(n5737), .A2(n5758), .B(a[29]), .C(n3889), .Z(n3733) );
  INVD1BWP12T U1153 ( .I(b[29]), .ZN(n4841) );
  INVD1BWP12T U1154 ( .I(b[28]), .ZN(n5722) );
  AOI22D1BWP12T U1155 ( .A1(n5380), .A2(n5722), .B1(n4455), .B2(n4841), .ZN(
        n3731) );
  OAI21D1BWP12T U1156 ( .A1(n4841), .A2(n4470), .B(n3731), .ZN(n3732) );
  ND2D1BWP12T U1157 ( .A1(n3733), .A2(n3732), .ZN(n3814) );
  OAI21D1BWP12T U1158 ( .A1(n3733), .A2(n3732), .B(n3814), .ZN(n3757) );
  INVD1BWP12T U1159 ( .I(b[20]), .ZN(n6067) );
  INVD1BWP12T U1160 ( .I(b[21]), .ZN(n4740) );
  AOI22D1BWP12T U1161 ( .A1(b[21]), .A2(n4668), .B1(n4667), .B2(n4740), .ZN(
        n3734) );
  AOI221D1BWP12T U1162 ( .A1(n4671), .A2(b[20]), .B1(n4670), .B2(n6067), .C(
        n3734), .ZN(n3788) );
  INVD1BWP12T U1163 ( .I(a[15]), .ZN(n6042) );
  NR3D1BWP12T U1164 ( .A1(a[17]), .A2(n5710), .A3(n6042), .ZN(n4329) );
  ND3D1BWP12T U1165 ( .A1(n5710), .A2(n6042), .A3(a[17]), .ZN(n4324) );
  INVD1BWP12T U1166 ( .I(n4324), .ZN(n4331) );
  AOI22D1BWP12T U1167 ( .A1(a[16]), .A2(a[15]), .B1(n6042), .B2(n5710), .ZN(
        n4359) );
  ND2D1BWP12T U1168 ( .A1(n4359), .A2(n5679), .ZN(n4553) );
  ND2D1BWP12T U1169 ( .A1(a[17]), .A2(n4359), .ZN(n4554) );
  INVD1BWP12T U1170 ( .I(b[13]), .ZN(n5476) );
  AOI22D1BWP12T U1171 ( .A1(b[13]), .A2(n4553), .B1(n4554), .B2(n5476), .ZN(
        n3735) );
  AOI221D1BWP12T U1172 ( .A1(n4329), .A2(b[12]), .B1(n4331), .B2(n4792), .C(
        n3735), .ZN(n3787) );
  INVD1BWP12T U1173 ( .I(b[22]), .ZN(n4839) );
  INVD1BWP12T U1174 ( .I(b[23]), .ZN(n5940) );
  AOI22D1BWP12T U1175 ( .A1(b[23]), .A2(n4632), .B1(n4631), .B2(n5940), .ZN(
        n3736) );
  AOI221D1BWP12T U1176 ( .A1(n4635), .A2(b[22]), .B1(n4634), .B2(n4839), .C(
        n3736), .ZN(n3786) );
  INVD1BWP12T U1177 ( .I(b[24]), .ZN(n5918) );
  INVD1BWP12T U1178 ( .I(b[25]), .ZN(n4739) );
  AOI22D1BWP12T U1179 ( .A1(b[25]), .A2(n4642), .B1(n4641), .B2(n4739), .ZN(
        n3737) );
  AOI221D1BWP12T U1180 ( .A1(n4645), .A2(b[24]), .B1(n4644), .B2(n5918), .C(
        n3737), .ZN(n3772) );
  AOI22D1BWP12T U1181 ( .A1(b[22]), .A2(n4632), .B1(n4631), .B2(n4839), .ZN(
        n3738) );
  AOI221D1BWP12T U1182 ( .A1(n4635), .A2(b[21]), .B1(n4634), .B2(n4740), .C(
        n3738), .ZN(n3769) );
  AOI22D1BWP12T U1183 ( .A1(b[12]), .A2(n4553), .B1(n4554), .B2(n4792), .ZN(
        n3739) );
  AOI221D1BWP12T U1184 ( .A1(n4329), .A2(b[11]), .B1(n4331), .B2(n4741), .C(
        n3739), .ZN(n3768) );
  INVD1BWP12T U1185 ( .I(b[19]), .ZN(n5989) );
  AOI22D1BWP12T U1186 ( .A1(b[20]), .A2(n4668), .B1(n4667), .B2(n6067), .ZN(
        n3740) );
  AOI221D1BWP12T U1187 ( .A1(n4671), .A2(b[19]), .B1(n4670), .B2(n5989), .C(
        n3740), .ZN(n3767) );
  AOI22D1BWP12T U1188 ( .A1(a[25]), .A2(b[5]), .B1(n4490), .B2(n5833), .ZN(
        n3785) );
  AOI22D1BWP12T U1189 ( .A1(n3973), .A2(n3785), .B1(n3966), .B2(n3741), .ZN(
        n3808) );
  INVD1BWP12T U1190 ( .I(b[18]), .ZN(n6010) );
  AOI22D1BWP12T U1191 ( .A1(b[19]), .A2(n4637), .B1(n4636), .B2(n5989), .ZN(
        n3742) );
  AOI221D1BWP12T U1192 ( .A1(n4640), .A2(b[18]), .B1(n4639), .B2(n6010), .C(
        n3742), .ZN(n3807) );
  AOI22D1BWP12T U1193 ( .A1(b[9]), .A2(n4673), .B1(n4672), .B2(n4482), .ZN(
        n3743) );
  AOI221D1BWP12T U1194 ( .A1(n4676), .A2(b[8]), .B1(n4675), .B2(n4699), .C(
        n3743), .ZN(n3806) );
  NR2D1BWP12T U1195 ( .A1(n6024), .A2(n5679), .ZN(n4268) );
  INVD1BWP12T U1196 ( .I(n4268), .ZN(n3744) );
  NR2D1BWP12T U1197 ( .A1(a[19]), .A2(n3744), .ZN(n4692) );
  NR2D1BWP12T U1198 ( .A1(n5988), .A2(n4267), .ZN(n4691) );
  INR2D1BWP12T U1199 ( .A1(n4267), .B1(n4268), .ZN(n4270) );
  ND2D1BWP12T U1200 ( .A1(n4270), .A2(n5988), .ZN(n4689) );
  ND2D1BWP12T U1201 ( .A1(a[19]), .A2(n4270), .ZN(n4688) );
  AOI22D1BWP12T U1202 ( .A1(b[11]), .A2(n4689), .B1(n4688), .B2(n4741), .ZN(
        n3745) );
  AOI221D1BWP12T U1203 ( .A1(n4692), .A2(b[10]), .B1(n4691), .B2(n4646), .C(
        n3745), .ZN(n3795) );
  AOI22D1BWP12T U1204 ( .A1(a[27]), .A2(b[3]), .B1(n5136), .B2(n5758), .ZN(
        n3801) );
  AOI22D1BWP12T U1205 ( .A1(n4557), .A2(n3801), .B1(n4558), .B2(n3746), .ZN(
        n3794) );
  INVD1BWP12T U1206 ( .I(b[15]), .ZN(n4890) );
  ND2D1BWP12T U1207 ( .A1(n4890), .A2(n6042), .ZN(n6043) );
  ND2D1BWP12T U1208 ( .A1(b[15]), .A2(a[15]), .ZN(n5392) );
  ND2D1BWP12T U1209 ( .A1(n6043), .A2(n5392), .ZN(n4858) );
  INVD1BWP12T U1210 ( .I(n4858), .ZN(n4914) );
  INVD1BWP12T U1211 ( .I(a[14]), .ZN(n5874) );
  NR2D1BWP12T U1212 ( .A1(n5874), .A2(n5872), .ZN(n5412) );
  NR2D1BWP12T U1213 ( .A1(n3747), .A2(n5412), .ZN(n4452) );
  ND2D1BWP12T U1214 ( .A1(n6042), .A2(n5412), .ZN(n3779) );
  ND2D1BWP12T U1215 ( .A1(a[15]), .A2(n3747), .ZN(n4422) );
  AOI22D1BWP12T U1216 ( .A1(b[14]), .A2(n3779), .B1(n4422), .B2(n5390), .ZN(
        n3748) );
  AOI21D1BWP12T U1217 ( .A1(n4914), .A2(n4452), .B(n3748), .ZN(n3793) );
  NR2D1BWP12T U1218 ( .A1(a[13]), .A2(n4488), .ZN(n4666) );
  NR2D1BWP12T U1219 ( .A1(n4488), .A2(n5872), .ZN(n4665) );
  NR3D1BWP12T U1220 ( .A1(n4791), .A2(n3749), .A3(a[13]), .ZN(n4007) );
  INVD1BWP12T U1221 ( .I(n4007), .ZN(n4663) );
  NR3D1BWP12T U1222 ( .A1(n5872), .A2(a[12]), .A3(a[11]), .ZN(n4476) );
  INVD1BWP12T U1223 ( .I(n4476), .ZN(n4662) );
  INVD1BWP12T U1224 ( .I(b[16]), .ZN(n4793) );
  AOI22D1BWP12T U1225 ( .A1(b[16]), .A2(n4663), .B1(n4662), .B2(n4793), .ZN(
        n3750) );
  AOI221D1BWP12T U1226 ( .A1(n4666), .A2(b[17]), .B1(n4665), .B2(n4838), .C(
        n3750), .ZN(n3869) );
  OAI22D1BWP12T U1227 ( .A1(n6155), .A2(a[21]), .B1(n5964), .B2(a[22]), .ZN(
        n4648) );
  AOI22D1BWP12T U1228 ( .A1(a[23]), .A2(b[6]), .B1(n4555), .B2(n5951), .ZN(
        n3759) );
  ND2D1BWP12T U1229 ( .A1(a[23]), .A2(a[22]), .ZN(n5418) );
  IND2D1BWP12T U1230 ( .A1(n4648), .B1(n5418), .ZN(n4060) );
  NR2D1BWP12T U1231 ( .A1(n3751), .A2(n4060), .ZN(n4649) );
  AOI22D1BWP12T U1232 ( .A1(a[23]), .A2(b[5]), .B1(n4490), .B2(n5951), .ZN(
        n3875) );
  AOI22D1BWP12T U1233 ( .A1(n4648), .A2(n3759), .B1(n4649), .B2(n3875), .ZN(
        n3776) );
  NR2D1BWP12T U1234 ( .A1(b[13]), .A2(a[13]), .ZN(n5642) );
  ND2D1BWP12T U1235 ( .A1(b[13]), .A2(a[13]), .ZN(n5645) );
  ND2D1BWP12T U1236 ( .A1(n3779), .A2(n4422), .ZN(n4421) );
  ND2D1BWP12T U1237 ( .A1(n4452), .A2(n6042), .ZN(n4684) );
  ND2D1BWP12T U1238 ( .A1(a[15]), .A2(n4452), .ZN(n4683) );
  AOI22D1BWP12T U1239 ( .A1(b[14]), .A2(n4684), .B1(n4683), .B2(n5390), .ZN(
        n3752) );
  AOI21D1BWP12T U1240 ( .A1(n4917), .A2(n4421), .B(n3752), .ZN(n3775) );
  AOI22D1BWP12T U1241 ( .A1(b[10]), .A2(n4689), .B1(n4688), .B2(n4646), .ZN(
        n3753) );
  AOI221D1BWP12T U1242 ( .A1(n4692), .A2(b[9]), .B1(n4691), .B2(n4482), .C(
        n3753), .ZN(n3774) );
  OAI22D1BWP12T U1243 ( .A1(b[27]), .A2(n4453), .B1(n5722), .B2(n4470), .ZN(
        n3754) );
  AOI21D1BWP12T U1244 ( .A1(n4455), .A2(n5722), .B(n3754), .ZN(n3888) );
  INVD1BWP12T U1245 ( .I(b[26]), .ZN(n5784) );
  AOI22D1BWP12T U1246 ( .A1(b[25]), .A2(n4658), .B1(n4657), .B2(n4739), .ZN(
        n3755) );
  AOI221D1BWP12T U1247 ( .A1(n4661), .A2(b[26]), .B1(n4660), .B2(n5784), .C(
        n3755), .ZN(n3887) );
  FA1D0BWP12T U1248 ( .A(n3758), .B(n3757), .CI(n3756), .CO(n3858), .S(n3866)
         );
  AOI22D1BWP12T U1249 ( .A1(a[23]), .A2(b[7]), .B1(n4450), .B2(n5951), .ZN(
        n3784) );
  AOI22D1BWP12T U1250 ( .A1(n4648), .A2(n3784), .B1(n4649), .B2(n3759), .ZN(
        n3798) );
  AOI22D1BWP12T U1251 ( .A1(a[29]), .A2(b[1]), .B1(n4419), .B2(n5901), .ZN(
        n3804) );
  ND2D1BWP12T U1252 ( .A1(a[28]), .A2(n5901), .ZN(n5892) );
  OAI22D1BWP12T U1253 ( .A1(n5379), .A2(n5737), .B1(n5901), .B2(b[0]), .ZN(
        n4960) );
  AOI22D1BWP12T U1254 ( .A1(n3804), .A2(n4694), .B1(n4695), .B2(n4960), .ZN(
        n3797) );
  INVD1BWP12T U1255 ( .I(b[27]), .ZN(n5751) );
  AOI22D1BWP12T U1256 ( .A1(b[26]), .A2(n4658), .B1(n4657), .B2(n5784), .ZN(
        n3760) );
  AOI221D1BWP12T U1257 ( .A1(n4661), .A2(b[27]), .B1(n4660), .B2(n5751), .C(
        n3760), .ZN(n3796) );
  NR2D1BWP12T U1258 ( .A1(b[0]), .A2(a[26]), .ZN(n3762) );
  OAI211D1BWP12T U1259 ( .A1(n3762), .A2(n5833), .B(a[27]), .C(n3761), .ZN(
        n3906) );
  AOI22D1BWP12T U1260 ( .A1(b[7]), .A2(n4673), .B1(n4672), .B2(n4450), .ZN(
        n3763) );
  AOI221D1BWP12T U1261 ( .A1(n4676), .A2(b[6]), .B1(n4675), .B2(n4555), .C(
        n3763), .ZN(n3905) );
  AOI22D1BWP12T U1262 ( .A1(b[23]), .A2(n4642), .B1(n4641), .B2(n5940), .ZN(
        n3764) );
  AOI221D1BWP12T U1263 ( .A1(n4645), .A2(b[22]), .B1(n4644), .B2(n4839), .C(
        n3764), .ZN(n3904) );
  AOI22D1BWP12T U1264 ( .A1(b[10]), .A2(n4329), .B1(n4331), .B2(n4646), .ZN(
        n3765) );
  OAI221D1BWP12T U1265 ( .A1(b[11]), .A2(n4554), .B1(n4741), .B2(n4553), .C(
        n3765), .ZN(n3911) );
  AOI22D1BWP12T U1266 ( .A1(n5380), .A2(n5784), .B1(n4455), .B2(n5751), .ZN(
        n3766) );
  OAI21D1BWP12T U1267 ( .A1(n5751), .A2(n4470), .B(n3766), .ZN(n3912) );
  ND2D1BWP12T U1268 ( .A1(n3911), .A2(n3912), .ZN(n3910) );
  FA1D0BWP12T U1269 ( .A(n3769), .B(n3768), .CI(n3767), .CO(n3771), .S(n3884)
         );
  FA1D0BWP12T U1270 ( .A(n3772), .B(n3771), .CI(n3770), .CO(n3857), .S(n3882)
         );
  AOI22D1BWP12T U1271 ( .A1(b[15]), .A2(n4663), .B1(n4662), .B2(n4890), .ZN(
        n3773) );
  AOI221D1BWP12T U1272 ( .A1(n4666), .A2(b[16]), .B1(n4665), .B2(n4793), .C(
        n3773), .ZN(n3896) );
  FA1D0BWP12T U1273 ( .A(n3776), .B(n3775), .CI(n3774), .CO(n3868), .S(n3895)
         );
  AOI22D1BWP12T U1274 ( .A1(b[0]), .A2(a[26]), .B1(a[27]), .B2(n5379), .ZN(
        n5283) );
  MAOI22D0BWP12T U1275 ( .A1(n4557), .A2(n3778), .B1(n5283), .B2(n3777), .ZN(
        n3937) );
  INVD1BWP12T U1276 ( .I(n3779), .ZN(n4687) );
  INVD1BWP12T U1277 ( .I(n4422), .ZN(n4686) );
  AOI22D1BWP12T U1278 ( .A1(b[13]), .A2(n4684), .B1(n4683), .B2(n5476), .ZN(
        n3780) );
  AOI221D1BWP12T U1279 ( .A1(n4687), .A2(b[12]), .B1(n4686), .B2(n4792), .C(
        n3780), .ZN(n3936) );
  AOI22D1BWP12T U1280 ( .A1(b[14]), .A2(n4663), .B1(n4662), .B2(n5390), .ZN(
        n3781) );
  AOI221D1BWP12T U1281 ( .A1(n4666), .A2(b[15]), .B1(n4665), .B2(n4890), .C(
        n3781), .ZN(n3935) );
  AOI22D1BWP12T U1282 ( .A1(b[10]), .A2(n4673), .B1(n4672), .B2(n4646), .ZN(
        n3782) );
  AOI221D1BWP12T U1283 ( .A1(n4676), .A2(b[9]), .B1(n4675), .B2(n4482), .C(
        n3782), .ZN(n3831) );
  AOI22D1BWP12T U1284 ( .A1(b[20]), .A2(n4637), .B1(n4636), .B2(n6067), .ZN(
        n3783) );
  AOI221D1BWP12T U1285 ( .A1(n4640), .A2(b[19]), .B1(n4639), .B2(n5989), .C(
        n3783), .ZN(n3825) );
  AOI22D1BWP12T U1286 ( .A1(a[23]), .A2(b[8]), .B1(n4699), .B2(n5951), .ZN(
        n3848) );
  AOI22D1BWP12T U1287 ( .A1(n4648), .A2(n3848), .B1(n4649), .B2(n3784), .ZN(
        n3824) );
  AOI22D1BWP12T U1288 ( .A1(a[25]), .A2(b[6]), .B1(n4555), .B2(n5833), .ZN(
        n3846) );
  AOI22D1BWP12T U1289 ( .A1(n3973), .A2(n3846), .B1(n3966), .B2(n3785), .ZN(
        n3823) );
  FA1D0BWP12T U1290 ( .A(n3788), .B(n3787), .CI(n3786), .CO(n3829), .S(n3756)
         );
  AOI22D1BWP12T U1291 ( .A1(b[16]), .A2(n4684), .B1(n4683), .B2(n4793), .ZN(
        n3789) );
  AOI21D1BWP12T U1292 ( .A1(n4914), .A2(n4421), .B(n3789), .ZN(n3828) );
  AOI22D1BWP12T U1293 ( .A1(b[26]), .A2(n4642), .B1(n4641), .B2(n5784), .ZN(
        n3790) );
  AOI221D1BWP12T U1294 ( .A1(n4645), .A2(b[25]), .B1(n4644), .B2(n4739), .C(
        n3790), .ZN(n3845) );
  AOI22D1BWP12T U1295 ( .A1(b[14]), .A2(n4553), .B1(n4554), .B2(n5390), .ZN(
        n3791) );
  AOI221D1BWP12T U1296 ( .A1(n4329), .A2(b[13]), .B1(n4331), .B2(n5476), .C(
        n3791), .ZN(n3844) );
  AOI22D1BWP12T U1297 ( .A1(b[12]), .A2(n4689), .B1(n4688), .B2(n4792), .ZN(
        n3792) );
  AOI221D1BWP12T U1298 ( .A1(n4692), .A2(b[11]), .B1(n4691), .B2(n4741), .C(
        n3792), .ZN(n3843) );
  FA1D0BWP12T U1299 ( .A(n3795), .B(n3794), .CI(n3793), .CO(n3826), .S(n3870)
         );
  FA1D0BWP12T U1300 ( .A(n3798), .B(n3797), .CI(n3796), .CO(n3813), .S(n3865)
         );
  INVD1BWP12T U1301 ( .I(b[30]), .ZN(n4737) );
  OAI22D1BWP12T U1302 ( .A1(b[29]), .A2(n4453), .B1(n4737), .B2(n4470), .ZN(
        n3799) );
  AOI21D1BWP12T U1303 ( .A1(n4455), .A2(n4737), .B(n3799), .ZN(n3852) );
  AOI22D1BWP12T U1304 ( .A1(b[27]), .A2(n4658), .B1(n4657), .B2(n5751), .ZN(
        n3800) );
  AOI221D1BWP12T U1305 ( .A1(n4661), .A2(b[28]), .B1(n4660), .B2(n5722), .C(
        n3800), .ZN(n3851) );
  ND2D1BWP12T U1306 ( .A1(a[30]), .A2(a[29]), .ZN(n5417) );
  NR2D1BWP12T U1307 ( .A1(a[30]), .A2(a[29]), .ZN(n4604) );
  INR2D1BWP12T U1308 ( .A1(n5417), .B1(n4604), .ZN(n4598) );
  ND2D1BWP12T U1309 ( .A1(b[0]), .A2(n4598), .ZN(n3850) );
  AOI22D1BWP12T U1310 ( .A1(a[27]), .A2(b[4]), .B1(n5703), .B2(n5758), .ZN(
        n3847) );
  AOI22D1BWP12T U1311 ( .A1(n4557), .A2(n3847), .B1(n4558), .B2(n3801), .ZN(
        n3810) );
  AOI22D1BWP12T U1312 ( .A1(b[24]), .A2(n4632), .B1(n4631), .B2(n5918), .ZN(
        n3802) );
  AOI221D1BWP12T U1313 ( .A1(n4635), .A2(b[23]), .B1(n4634), .B2(n5940), .C(
        n3802), .ZN(n3855) );
  AOI22D1BWP12T U1314 ( .A1(b[17]), .A2(n4663), .B1(n4662), .B2(n4838), .ZN(
        n3803) );
  AOI221D1BWP12T U1315 ( .A1(n4666), .A2(b[18]), .B1(n4665), .B2(n6010), .C(
        n3803), .ZN(n3834) );
  AOI22D1BWP12T U1316 ( .A1(a[29]), .A2(b[2]), .B1(n5210), .B2(n5901), .ZN(
        n3841) );
  AOI22D1BWP12T U1317 ( .A1(n4694), .A2(n3841), .B1(n4695), .B2(n3804), .ZN(
        n3833) );
  AOI22D1BWP12T U1318 ( .A1(b[22]), .A2(n4668), .B1(n4667), .B2(n4839), .ZN(
        n3805) );
  AOI221D1BWP12T U1319 ( .A1(n4671), .A2(b[21]), .B1(n4670), .B2(n4740), .C(
        n3805), .ZN(n3832) );
  FA1D0BWP12T U1320 ( .A(n3808), .B(n3807), .CI(n3806), .CO(n3853), .S(n3770)
         );
  FA1D0BWP12T U1321 ( .A(n3811), .B(n3810), .CI(n3809), .CO(n4570), .S(n3862)
         );
  FA1D0BWP12T U1322 ( .A(n3814), .B(n3813), .CI(n3812), .CO(n4616), .S(n3811)
         );
  AOI22D1BWP12T U1323 ( .A1(b[23]), .A2(n4668), .B1(n4667), .B2(n5940), .ZN(
        n3815) );
  AOI221D1BWP12T U1324 ( .A1(n4671), .A2(b[22]), .B1(n4670), .B2(n4839), .C(
        n3815), .ZN(n4562) );
  ND2D1BWP12T U1325 ( .A1(n4604), .A2(n5379), .ZN(n3816) );
  OAI32D1BWP12T U1326 ( .A1(a[31]), .A2(n4738), .A3(n3817), .B1(n3816), .B2(
        n5593), .ZN(n3818) );
  OAI32D1BWP12T U1327 ( .A1(n3818), .A2(n4600), .A3(n4603), .B1(n4598), .B2(
        n3818), .ZN(n4561) );
  AOI22D1BWP12T U1328 ( .A1(b[28]), .A2(n4658), .B1(n4657), .B2(n5722), .ZN(
        n3819) );
  AOI221D1BWP12T U1329 ( .A1(n4661), .A2(b[29]), .B1(n4660), .B2(n4841), .C(
        n3819), .ZN(n4560) );
  AOI22D1BWP12T U1330 ( .A1(a[1]), .A2(b[31]), .B1(n5595), .B2(n5805), .ZN(
        n3820) );
  AOI22D1BWP12T U1331 ( .A1(a[0]), .A2(n3820), .B1(n5380), .B2(n4737), .ZN(
        n3822) );
  ND3D1BWP12T U1332 ( .A1(a[31]), .A2(n5417), .A3(n3850), .ZN(n3821) );
  NR2D1BWP12T U1333 ( .A1(n3822), .A2(n3821), .ZN(n4698) );
  AO21D1BWP12T U1334 ( .A1(n3822), .A2(n3821), .B(n4698), .Z(n4708) );
  FA1D0BWP12T U1335 ( .A(n3825), .B(n3824), .CI(n3823), .CO(n4707), .S(n3830)
         );
  FA1D0BWP12T U1336 ( .A(n3828), .B(n3827), .CI(n3826), .CO(n4614), .S(n3863)
         );
  FA1D0BWP12T U1337 ( .A(n3831), .B(n3830), .CI(n3829), .CO(n4568), .S(n3864)
         );
  FA1D0BWP12T U1338 ( .A(n3834), .B(n3833), .CI(n3832), .CO(n4586), .S(n3854)
         );
  AOI22D1BWP12T U1339 ( .A1(b[13]), .A2(n4689), .B1(n4688), .B2(n5476), .ZN(
        n3835) );
  AOI221D1BWP12T U1340 ( .A1(n4692), .A2(b[12]), .B1(n4691), .B2(n4792), .C(
        n3835), .ZN(n4585) );
  AOI22D1BWP12T U1341 ( .A1(b[11]), .A2(n4673), .B1(n4672), .B2(n4741), .ZN(
        n3836) );
  AOI221D1BWP12T U1342 ( .A1(n4676), .A2(b[10]), .B1(n4675), .B2(n4646), .C(
        n3836), .ZN(n4712) );
  AOI22D1BWP12T U1343 ( .A1(b[15]), .A2(n4553), .B1(n4554), .B2(n4890), .ZN(
        n3837) );
  AOI221D1BWP12T U1344 ( .A1(n4329), .A2(b[14]), .B1(n4331), .B2(n5390), .C(
        n3837), .ZN(n4711) );
  AOI22D1BWP12T U1345 ( .A1(b[27]), .A2(n4642), .B1(n4641), .B2(n5751), .ZN(
        n3838) );
  AOI221D1BWP12T U1346 ( .A1(n4645), .A2(b[26]), .B1(n4644), .B2(n5784), .C(
        n3838), .ZN(n4710) );
  AOI22D1BWP12T U1347 ( .A1(b[25]), .A2(n4632), .B1(n4631), .B2(n4739), .ZN(
        n3839) );
  AOI221D1BWP12T U1348 ( .A1(n4635), .A2(b[24]), .B1(n4634), .B2(n5918), .C(
        n3839), .ZN(n4613) );
  AOI22D1BWP12T U1349 ( .A1(b[17]), .A2(n4684), .B1(n4683), .B2(n4838), .ZN(
        n3840) );
  AOI221D1BWP12T U1350 ( .A1(n4687), .A2(b[16]), .B1(n4686), .B2(n4793), .C(
        n3840), .ZN(n4565) );
  AOI22D1BWP12T U1351 ( .A1(a[29]), .A2(b[3]), .B1(n5136), .B2(n5901), .ZN(
        n4696) );
  AOI22D1BWP12T U1352 ( .A1(n4696), .A2(n4694), .B1(n4695), .B2(n3841), .ZN(
        n4564) );
  AOI22D1BWP12T U1353 ( .A1(b[18]), .A2(n4663), .B1(n4662), .B2(n6010), .ZN(
        n3842) );
  AOI221D1BWP12T U1354 ( .A1(n4666), .A2(b[19]), .B1(n4665), .B2(n5989), .C(
        n3842), .ZN(n4563) );
  FA1D0BWP12T U1355 ( .A(n3845), .B(n3844), .CI(n3843), .CO(n4611), .S(n3827)
         );
  AOI22D1BWP12T U1356 ( .A1(a[25]), .A2(n4450), .B1(b[7]), .B2(n5833), .ZN(
        n4703) );
  MAOI22D0BWP12T U1357 ( .A1(n3966), .A2(n3846), .B1(n4703), .B2(n4701), .ZN(
        n4607) );
  AOI22D1BWP12T U1358 ( .A1(a[27]), .A2(b[5]), .B1(n4490), .B2(n5758), .ZN(
        n4559) );
  AOI22D1BWP12T U1359 ( .A1(n4559), .A2(n4557), .B1(n4558), .B2(n3847), .ZN(
        n4578) );
  AOI22D1BWP12T U1360 ( .A1(a[23]), .A2(b[9]), .B1(n4482), .B2(n5951), .ZN(
        n4650) );
  AOI22D1BWP12T U1361 ( .A1(n4650), .A2(n4648), .B1(n4649), .B2(n3848), .ZN(
        n4577) );
  AOI22D1BWP12T U1362 ( .A1(b[21]), .A2(n4637), .B1(n4636), .B2(n4740), .ZN(
        n3849) );
  AOI221D1BWP12T U1363 ( .A1(n4640), .A2(b[20]), .B1(n4639), .B2(n6067), .C(
        n3849), .ZN(n4576) );
  FA1D0BWP12T U1364 ( .A(n3852), .B(n3851), .CI(n3850), .CO(n4605), .S(n3812)
         );
  FA1D0BWP12T U1365 ( .A(n3855), .B(n3854), .CI(n3853), .CO(n4572), .S(n3809)
         );
  FA1D0BWP12T U1366 ( .A(n3858), .B(n3857), .CI(n3856), .CO(n4571), .S(n3861)
         );
  FA1D0BWP12T U1367 ( .A(n3861), .B(n3860), .CI(n3859), .CO(n4610), .S(n3921)
         );
  FA1D0BWP12T U1368 ( .A(n3864), .B(n3863), .CI(n3862), .CO(n4581), .S(n3920)
         );
  FA1D0BWP12T U1369 ( .A(n3867), .B(n3866), .CI(n3865), .CO(n3860), .S(n3880)
         );
  FA1D0BWP12T U1370 ( .A(n3870), .B(n3869), .CI(n3868), .CO(n3856), .S(n3879)
         );
  AOI22D1BWP12T U1371 ( .A1(b[24]), .A2(n4642), .B1(n4641), .B2(n5918), .ZN(
        n3871) );
  AOI221D1BWP12T U1372 ( .A1(n4645), .A2(b[23]), .B1(n4644), .B2(n5940), .C(
        n3871), .ZN(n3902) );
  FA1D0BWP12T U1373 ( .A(n3874), .B(n3873), .CI(n3872), .CO(n3758), .S(n3901)
         );
  AOI22D1BWP12T U1374 ( .A1(a[23]), .A2(b[4]), .B1(n5703), .B2(n5951), .ZN(
        n3938) );
  AOI22D1BWP12T U1375 ( .A1(n4648), .A2(n3875), .B1(n4649), .B2(n3938), .ZN(
        n3915) );
  AOI22D1BWP12T U1376 ( .A1(b[21]), .A2(n4632), .B1(n4631), .B2(n4740), .ZN(
        n3876) );
  AOI221D1BWP12T U1377 ( .A1(n4635), .A2(b[20]), .B1(n4634), .B2(n6067), .C(
        n3876), .ZN(n3914) );
  AOI22D1BWP12T U1378 ( .A1(b[24]), .A2(n4658), .B1(n4657), .B2(n5918), .ZN(
        n3877) );
  AOI221D1BWP12T U1379 ( .A1(n4661), .A2(b[25]), .B1(n4660), .B2(n4739), .C(
        n3877), .ZN(n3913) );
  FA1D0BWP12T U1380 ( .A(n3880), .B(n3879), .CI(n3878), .CO(n3919), .S(n3927)
         );
  FA1D0BWP12T U1381 ( .A(n3883), .B(n3882), .CI(n3881), .CO(n3859), .S(n3924)
         );
  FA1D0BWP12T U1382 ( .A(n3885), .B(n3910), .CI(n3884), .CO(n3883), .S(n3930)
         );
  AOI22D1BWP12T U1383 ( .A1(b[18]), .A2(n4637), .B1(n4636), .B2(n6010), .ZN(
        n3886) );
  AOI221D1BWP12T U1384 ( .A1(n4640), .A2(b[17]), .B1(n4639), .B2(n4838), .C(
        n3886), .ZN(n3899) );
  FA1D0BWP12T U1385 ( .A(n3889), .B(n3888), .CI(n3887), .CO(n3867), .S(n3898)
         );
  AOI22D1BWP12T U1386 ( .A1(b[17]), .A2(n4637), .B1(n4636), .B2(n4838), .ZN(
        n3890) );
  AOI221D1BWP12T U1387 ( .A1(n4640), .A2(b[16]), .B1(n4639), .B2(n4793), .C(
        n3890), .ZN(n3949) );
  AOI22D1BWP12T U1388 ( .A1(a[25]), .A2(b[2]), .B1(n5210), .B2(n5833), .ZN(
        n3918) );
  AOI22D1BWP12T U1389 ( .A1(n3973), .A2(n3891), .B1(n3966), .B2(n3918), .ZN(
        n3948) );
  ND2D1BWP12T U1390 ( .A1(b[0]), .A2(n4557), .ZN(n3954) );
  AOI22D1BWP12T U1391 ( .A1(b[23]), .A2(n4658), .B1(n4657), .B2(n5940), .ZN(
        n3892) );
  AOI221D1BWP12T U1392 ( .A1(n4661), .A2(b[24]), .B1(n4660), .B2(n5918), .C(
        n3892), .ZN(n3953) );
  OAI22D1BWP12T U1393 ( .A1(b[25]), .A2(n4453), .B1(n5784), .B2(n4470), .ZN(
        n3893) );
  AOI21D1BWP12T U1394 ( .A1(n4455), .A2(n5784), .B(n3893), .ZN(n3952) );
  FA1D0BWP12T U1395 ( .A(n3896), .B(n3895), .CI(n3894), .CO(n3881), .S(n3928)
         );
  FA1D0BWP12T U1396 ( .A(n3899), .B(n3898), .CI(n3897), .CO(n3922), .S(n3929)
         );
  FA1D0BWP12T U1397 ( .A(n3902), .B(n3901), .CI(n3900), .CO(n3878), .S(n3933)
         );
  AOI22D1BWP12T U1398 ( .A1(b[9]), .A2(n4689), .B1(n4688), .B2(n4482), .ZN(
        n3903) );
  AOI221D1BWP12T U1399 ( .A1(n4692), .A2(b[8]), .B1(n4691), .B2(n4699), .C(
        n3903), .ZN(n3960) );
  FA1D0BWP12T U1400 ( .A(n3906), .B(n3905), .CI(n3904), .CO(n3885), .S(n3959)
         );
  AOI22D1BWP12T U1401 ( .A1(b[10]), .A2(n4553), .B1(n4554), .B2(n4646), .ZN(
        n3907) );
  AOI221D1BWP12T U1402 ( .A1(n4329), .A2(b[9]), .B1(n4331), .B2(n4482), .C(
        n3907), .ZN(n3964) );
  AOI22D1BWP12T U1403 ( .A1(b[18]), .A2(n4668), .B1(n4667), .B2(n6010), .ZN(
        n3908) );
  AOI221D1BWP12T U1404 ( .A1(n4671), .A2(b[17]), .B1(n4670), .B2(n4838), .C(
        n3908), .ZN(n3963) );
  NR2D1BWP12T U1405 ( .A1(n4007), .A2(n4476), .ZN(n4489) );
  NR2D1BWP12T U1406 ( .A1(n4489), .A2(n4917), .ZN(n3909) );
  AOI221D1BWP12T U1407 ( .A1(n4666), .A2(b[14]), .B1(n4665), .B2(n5390), .C(
        n3909), .ZN(n3962) );
  OAI21D1BWP12T U1408 ( .A1(n3912), .A2(n3911), .B(n3910), .ZN(n3946) );
  FA1D0BWP12T U1409 ( .A(n3915), .B(n3914), .CI(n3913), .CO(n3900), .S(n3945)
         );
  AOI22D1BWP12T U1410 ( .A1(b[6]), .A2(n4673), .B1(n4672), .B2(n4555), .ZN(
        n3916) );
  AOI221D1BWP12T U1411 ( .A1(n4676), .A2(b[5]), .B1(n4675), .B2(n4490), .C(
        n3916), .ZN(n3993) );
  AOI22D1BWP12T U1412 ( .A1(b[16]), .A2(n4637), .B1(n4636), .B2(n4793), .ZN(
        n3917) );
  AOI221D1BWP12T U1413 ( .A1(n4640), .A2(b[15]), .B1(n4639), .B2(n4890), .C(
        n3917), .ZN(n3992) );
  AOI22D1BWP12T U1414 ( .A1(a[25]), .A2(b[1]), .B1(n4419), .B2(n5833), .ZN(
        n3967) );
  AOI22D1BWP12T U1415 ( .A1(n3973), .A2(n3918), .B1(n3966), .B2(n3967), .ZN(
        n3991) );
  FA1D0BWP12T U1416 ( .A(n3921), .B(n3920), .CI(n3919), .CO(n4608), .S(n3977)
         );
  FA1D0BWP12T U1417 ( .A(n3924), .B(n3923), .CI(n3922), .CO(n3976), .S(n3926)
         );
  FA1D0BWP12T U1418 ( .A(n3927), .B(n3926), .CI(n3925), .CO(n3978), .S(n3981)
         );
  FA1D0BWP12T U1419 ( .A(n3930), .B(n3929), .CI(n3928), .CO(n3923), .S(n3943)
         );
  FA1D0BWP12T U1420 ( .A(n3933), .B(n3932), .CI(n3931), .CO(n3925), .S(n3942)
         );
  AOI22D1BWP12T U1421 ( .A1(b[19]), .A2(n4668), .B1(n4667), .B2(n5989), .ZN(
        n3934) );
  AOI221D1BWP12T U1422 ( .A1(n4671), .A2(b[18]), .B1(n4670), .B2(n6010), .C(
        n3934), .ZN(n4024) );
  FA1D0BWP12T U1423 ( .A(n3937), .B(n3936), .CI(n3935), .CO(n3894), .S(n4023)
         );
  AOI22D1BWP12T U1424 ( .A1(a[23]), .A2(b[3]), .B1(n5136), .B2(n5951), .ZN(
        n3956) );
  AOI22D1BWP12T U1425 ( .A1(n4648), .A2(n3938), .B1(n4649), .B2(n3956), .ZN(
        n3972) );
  AOI22D1BWP12T U1426 ( .A1(b[8]), .A2(n4689), .B1(n4688), .B2(n4699), .ZN(
        n3939) );
  AOI221D1BWP12T U1427 ( .A1(n4692), .A2(b[7]), .B1(n4691), .B2(n4450), .C(
        n3939), .ZN(n3971) );
  AOI22D1BWP12T U1428 ( .A1(b[22]), .A2(n4642), .B1(n4641), .B2(n4839), .ZN(
        n3940) );
  AOI221D1BWP12T U1429 ( .A1(n4645), .A2(b[21]), .B1(n4644), .B2(n4740), .C(
        n3940), .ZN(n3970) );
  FA1D0BWP12T U1430 ( .A(n3943), .B(n3942), .CI(n3941), .CO(n3980), .S(n3984)
         );
  FA1D0BWP12T U1431 ( .A(n3946), .B(n3945), .CI(n3944), .CO(n3931), .S(n3987)
         );
  FA1D0BWP12T U1432 ( .A(n3949), .B(n3948), .CI(n3947), .CO(n3897), .S(n3986)
         );
  AOI22D1BWP12T U1433 ( .A1(n5380), .A2(n5918), .B1(n4455), .B2(n4739), .ZN(
        n3950) );
  OAI21D1BWP12T U1434 ( .A1(n4739), .A2(n4470), .B(n3950), .ZN(n4014) );
  AOI22D1BWP12T U1435 ( .A1(b[8]), .A2(n4329), .B1(n4331), .B2(n4699), .ZN(
        n3951) );
  OAI221D1BWP12T U1436 ( .A1(b[9]), .A2(n4554), .B1(n4482), .B2(n4553), .C(
        n3951), .ZN(n4015) );
  ND2D1BWP12T U1437 ( .A1(n4014), .A2(n4015), .ZN(n4013) );
  FA1D0BWP12T U1438 ( .A(n3954), .B(n3953), .CI(n3952), .CO(n3947), .S(n3995)
         );
  AOI22D1BWP12T U1439 ( .A1(b[22]), .A2(n4658), .B1(n4657), .B2(n4839), .ZN(
        n3955) );
  AOI221D1BWP12T U1440 ( .A1(n4661), .A2(b[23]), .B1(n4660), .B2(n5940), .C(
        n3955), .ZN(n4069) );
  AOI22D1BWP12T U1441 ( .A1(a[23]), .A2(b[2]), .B1(n5210), .B2(n5951), .ZN(
        n4010) );
  AOI22D1BWP12T U1442 ( .A1(n4648), .A2(n3956), .B1(n4649), .B2(n4010), .ZN(
        n4068) );
  AOI22D1BWP12T U1443 ( .A1(b[15]), .A2(n4637), .B1(n4636), .B2(n4890), .ZN(
        n3957) );
  AOI221D1BWP12T U1444 ( .A1(n4640), .A2(b[14]), .B1(n4639), .B2(n5390), .C(
        n3957), .ZN(n4067) );
  FA1D0BWP12T U1445 ( .A(n3960), .B(n3959), .CI(n3958), .CO(n3932), .S(n3990)
         );
  AOI22D1BWP12T U1446 ( .A1(b[20]), .A2(n4632), .B1(n4631), .B2(n6067), .ZN(
        n3961) );
  AOI221D1BWP12T U1447 ( .A1(n4635), .A2(b[19]), .B1(n4634), .B2(n5989), .C(
        n3961), .ZN(n4002) );
  FA1D0BWP12T U1448 ( .A(n3964), .B(n3963), .CI(n3962), .CO(n3958), .S(n4001)
         );
  AOI22D1BWP12T U1449 ( .A1(b[19]), .A2(n4632), .B1(n4631), .B2(n5989), .ZN(
        n3965) );
  AOI221D1BWP12T U1450 ( .A1(n4635), .A2(b[18]), .B1(n4634), .B2(n6010), .C(
        n3965), .ZN(n4018) );
  AOI22D1BWP12T U1451 ( .A1(n3967), .A2(n3973), .B1(n3966), .B2(n5018), .ZN(
        n4017) );
  AOI22D1BWP12T U1452 ( .A1(b[17]), .A2(n4668), .B1(n4667), .B2(n4838), .ZN(
        n3968) );
  AOI221D1BWP12T U1453 ( .A1(n4671), .A2(b[16]), .B1(n4670), .B2(n4793), .C(
        n3968), .ZN(n4016) );
  AOI22D1BWP12T U1454 ( .A1(b[12]), .A2(n4684), .B1(n4683), .B2(n4792), .ZN(
        n3969) );
  AOI221D1BWP12T U1455 ( .A1(n4687), .A2(b[11]), .B1(n4686), .B2(n4741), .C(
        n3969), .ZN(n4036) );
  FA1D0BWP12T U1456 ( .A(n3972), .B(n3971), .CI(n3970), .CO(n4022), .S(n4035)
         );
  ND2D1BWP12T U1457 ( .A1(b[0]), .A2(n3973), .ZN(n4053) );
  OAI211D1BWP12T U1458 ( .A1(n5912), .A2(n5951), .B(a[25]), .C(n4053), .ZN(
        n4005) );
  AOI22D1BWP12T U1459 ( .A1(b[11]), .A2(n4684), .B1(n4683), .B2(n4741), .ZN(
        n3974) );
  AOI221D1BWP12T U1460 ( .A1(n4687), .A2(b[10]), .B1(n4686), .B2(n4646), .C(
        n3974), .ZN(n4004) );
  AOI22D1BWP12T U1461 ( .A1(b[7]), .A2(n4689), .B1(n4688), .B2(n4450), .ZN(
        n3975) );
  AOI221D1BWP12T U1462 ( .A1(n4692), .A2(b[6]), .B1(n4691), .B2(n4555), .C(
        n3975), .ZN(n4003) );
  FA1D0BWP12T U1463 ( .A(n3978), .B(n3977), .CI(n3976), .CO(n4705), .S(n5319)
         );
  FA1D0BWP12T U1464 ( .A(n3981), .B(n3980), .CI(n3979), .CO(n5320), .S(n5344)
         );
  FA1D0BWP12T U1465 ( .A(n3984), .B(n3983), .CI(n3982), .CO(n3979), .S(n4030)
         );
  FA1D0BWP12T U1466 ( .A(n3987), .B(n3986), .CI(n3985), .CO(n3983), .S(n4033)
         );
  FA1D0BWP12T U1467 ( .A(n3990), .B(n3989), .CI(n3988), .CO(n3982), .S(n4027)
         );
  FA1D0BWP12T U1468 ( .A(n3993), .B(n3992), .CI(n3991), .CO(n3944), .S(n4039)
         );
  FA1D0BWP12T U1469 ( .A(n4013), .B(n3995), .CI(n3994), .CO(n3985), .S(n4038)
         );
  AOI22D1BWP12T U1470 ( .A1(b[5]), .A2(n4673), .B1(n4672), .B2(n4490), .ZN(
        n3996) );
  AOI221D1BWP12T U1471 ( .A1(n4676), .A2(b[4]), .B1(n4675), .B2(n5703), .C(
        n3996), .ZN(n4066) );
  AOI22D1BWP12T U1472 ( .A1(b[21]), .A2(n4642), .B1(n4641), .B2(n4740), .ZN(
        n3997) );
  AOI221D1BWP12T U1473 ( .A1(n4645), .A2(b[20]), .B1(n4644), .B2(n6067), .C(
        n3997), .ZN(n4065) );
  OAI22D1BWP12T U1474 ( .A1(b[23]), .A2(n4453), .B1(n5918), .B2(n4470), .ZN(
        n3998) );
  AOI21D1BWP12T U1475 ( .A1(n4455), .A2(n5918), .B(n3998), .ZN(n4052) );
  AOI22D1BWP12T U1476 ( .A1(b[21]), .A2(n4658), .B1(n4657), .B2(n4740), .ZN(
        n3999) );
  AOI221D1BWP12T U1477 ( .A1(n4661), .A2(b[22]), .B1(n4660), .B2(n4839), .C(
        n3999), .ZN(n4051) );
  FA1D0BWP12T U1478 ( .A(n4002), .B(n4001), .CI(n4000), .CO(n3989), .S(n4042)
         );
  FA1D0BWP12T U1479 ( .A(n4005), .B(n4004), .CI(n4003), .CO(n4034), .S(n4045)
         );
  OAI22D1BWP12T U1480 ( .A1(b[12]), .A2(n4662), .B1(n4488), .B2(n4917), .ZN(
        n4006) );
  AOI21D1BWP12T U1481 ( .A1(b[12]), .A2(n4007), .B(n4006), .ZN(n4044) );
  ND2D1BWP12T U1482 ( .A1(n4009), .A2(n4008), .ZN(n4061) );
  AOI22D1BWP12T U1483 ( .A1(n4648), .A2(n4010), .B1(n4649), .B2(n4061), .ZN(
        n4056) );
  AOI22D1BWP12T U1484 ( .A1(b[10]), .A2(n4684), .B1(n4683), .B2(n4646), .ZN(
        n4011) );
  AOI221D1BWP12T U1485 ( .A1(n4687), .A2(b[9]), .B1(n4686), .B2(n4482), .C(
        n4011), .ZN(n4055) );
  AOI22D1BWP12T U1486 ( .A1(b[6]), .A2(n4689), .B1(n4688), .B2(n4555), .ZN(
        n4012) );
  AOI221D1BWP12T U1487 ( .A1(n4692), .A2(b[5]), .B1(n4691), .B2(n4490), .C(
        n4012), .ZN(n4054) );
  OAI21D1BWP12T U1488 ( .A1(n4015), .A2(n4014), .B(n4013), .ZN(n4105) );
  FA1D0BWP12T U1489 ( .A(n4018), .B(n4017), .CI(n4016), .CO(n4000), .S(n4104)
         );
  AOI22D1BWP12T U1490 ( .A1(b[14]), .A2(n4637), .B1(n4636), .B2(n5390), .ZN(
        n4019) );
  AOI221D1BWP12T U1491 ( .A1(n4640), .A2(b[13]), .B1(n4639), .B2(n5476), .C(
        n4019), .ZN(n4050) );
  AOI22D1BWP12T U1492 ( .A1(b[20]), .A2(n4642), .B1(n4641), .B2(n6067), .ZN(
        n4020) );
  AOI221D1BWP12T U1493 ( .A1(n4645), .A2(b[19]), .B1(n4644), .B2(n5989), .C(
        n4020), .ZN(n4049) );
  AOI22D1BWP12T U1494 ( .A1(b[4]), .A2(n4673), .B1(n4672), .B2(n5703), .ZN(
        n4021) );
  AOI221D1BWP12T U1495 ( .A1(n4676), .A2(b[3]), .B1(n4675), .B2(n5136), .C(
        n4021), .ZN(n4048) );
  FA1D0BWP12T U1496 ( .A(n4024), .B(n4023), .CI(n4022), .CO(n3941), .S(n4031)
         );
  FA1D0BWP12T U1497 ( .A(n4027), .B(n4026), .CI(n4025), .CO(n4028), .S(n4032)
         );
  FA1D0BWP12T U1498 ( .A(n4030), .B(n4029), .CI(n4028), .CO(n5343), .S(n5317)
         );
  FA1D0BWP12T U1499 ( .A(n4033), .B(n4032), .CI(n4031), .CO(n4029), .S(n4116)
         );
  FA1D0BWP12T U1500 ( .A(n4036), .B(n4035), .CI(n4034), .CO(n3988), .S(n4110)
         );
  FA1D0BWP12T U1501 ( .A(n4039), .B(n4038), .CI(n4037), .CO(n4026), .S(n4075)
         );
  FA1D0BWP12T U1502 ( .A(n4042), .B(n4041), .CI(n4040), .CO(n4025), .S(n4074)
         );
  FA1D0BWP12T U1503 ( .A(n4045), .B(n4044), .CI(n4043), .CO(n4041), .S(n4078)
         );
  ND2D1BWP12T U1504 ( .A1(b[0]), .A2(n4648), .ZN(n4125) );
  OAI211D1BWP12T U1505 ( .A1(n6155), .A2(n5964), .B(a[23]), .C(n4125), .ZN(
        n4155) );
  AOI22D1BWP12T U1506 ( .A1(b[17]), .A2(n4632), .B1(n4631), .B2(n4838), .ZN(
        n4046) );
  AOI221D1BWP12T U1507 ( .A1(n4635), .A2(b[16]), .B1(n4634), .B2(n4793), .C(
        n4046), .ZN(n4154) );
  AOI22D1BWP12T U1508 ( .A1(b[20]), .A2(n4658), .B1(n4657), .B2(n6067), .ZN(
        n4047) );
  AOI221D1BWP12T U1509 ( .A1(n4661), .A2(b[21]), .B1(n4660), .B2(n4740), .C(
        n4047), .ZN(n4153) );
  FA1D0BWP12T U1510 ( .A(n4050), .B(n4049), .CI(n4048), .CO(n4103), .S(n4121)
         );
  FA1D0BWP12T U1511 ( .A(n4053), .B(n4052), .CI(n4051), .CO(n4064), .S(n4120)
         );
  FA1D0BWP12T U1512 ( .A(n4056), .B(n4055), .CI(n4054), .CO(n4043), .S(n4158)
         );
  OAI33D1BWP12T U1513 ( .A1(a[12]), .A2(n4058), .A3(n5872), .B1(n4791), .B2(
        n4057), .B3(a[13]), .ZN(n4059) );
  AOI221D1BWP12T U1514 ( .A1(n4666), .A2(b[12]), .B1(n4665), .B2(n4792), .C(
        n4059), .ZN(n4157) );
  AOI22D1BWP12T U1515 ( .A1(b[0]), .A2(a[22]), .B1(a[23]), .B2(n5379), .ZN(
        n5285) );
  MAOI22D0BWP12T U1516 ( .A1(n4648), .A2(n4061), .B1(n5285), .B2(n4060), .ZN(
        n4096) );
  AOI22D1BWP12T U1517 ( .A1(b[10]), .A2(n4663), .B1(n4662), .B2(n4646), .ZN(
        n4062) );
  AOI221D1BWP12T U1518 ( .A1(n4666), .A2(b[11]), .B1(n4665), .B2(n4741), .C(
        n4062), .ZN(n4095) );
  AOI22D1BWP12T U1519 ( .A1(b[9]), .A2(n4684), .B1(n4683), .B2(n4482), .ZN(
        n4063) );
  AOI221D1BWP12T U1520 ( .A1(n4687), .A2(b[8]), .B1(n4686), .B2(n4699), .C(
        n4063), .ZN(n4094) );
  FA1D0BWP12T U1521 ( .A(n4066), .B(n4065), .CI(n4064), .CO(n4037), .S(n4081)
         );
  FA1D0BWP12T U1522 ( .A(n4069), .B(n4068), .CI(n4067), .CO(n3994), .S(n4080)
         );
  AOI22D1BWP12T U1523 ( .A1(b[16]), .A2(n4668), .B1(n4667), .B2(n4793), .ZN(
        n4070) );
  AOI221D1BWP12T U1524 ( .A1(n4671), .A2(b[15]), .B1(n4670), .B2(n4890), .C(
        n4070), .ZN(n4086) );
  AOI22D1BWP12T U1525 ( .A1(b[8]), .A2(n4553), .B1(n4554), .B2(n4699), .ZN(
        n4071) );
  AOI221D1BWP12T U1526 ( .A1(n4329), .A2(b[7]), .B1(n4331), .B2(n4450), .C(
        n4071), .ZN(n4085) );
  AOI22D1BWP12T U1527 ( .A1(b[18]), .A2(n4632), .B1(n4631), .B2(n6010), .ZN(
        n4072) );
  AOI221D1BWP12T U1528 ( .A1(n4635), .A2(b[17]), .B1(n4634), .B2(n4838), .C(
        n4072), .ZN(n4084) );
  FA1D0BWP12T U1529 ( .A(n4075), .B(n4074), .CI(n4073), .CO(n4114), .S(n4109)
         );
  FA1D0BWP12T U1530 ( .A(n4078), .B(n4077), .CI(n4076), .CO(n4073), .S(n4113)
         );
  FA1D0BWP12T U1531 ( .A(n4081), .B(n4080), .CI(n4079), .CO(n4108), .S(n4112)
         );
  AOI22D1BWP12T U1532 ( .A1(n5380), .A2(n4839), .B1(n4455), .B2(n5940), .ZN(
        n4082) );
  OAI21D1BWP12T U1533 ( .A1(n5940), .A2(n4470), .B(n4082), .ZN(n4151) );
  AOI22D1BWP12T U1534 ( .A1(b[6]), .A2(n4329), .B1(n4331), .B2(n4555), .ZN(
        n4083) );
  OAI221D1BWP12T U1535 ( .A1(b[7]), .A2(n4554), .B1(n4450), .B2(n4553), .C(
        n4083), .ZN(n4152) );
  ND2D1BWP12T U1536 ( .A1(n4151), .A2(n4152), .ZN(n4150) );
  FA1D0BWP12T U1537 ( .A(n4086), .B(n4085), .CI(n4084), .CO(n4079), .S(n4107)
         );
  AOI22D1BWP12T U1538 ( .A1(b[13]), .A2(n4637), .B1(n4636), .B2(n5476), .ZN(
        n4087) );
  AOI221D1BWP12T U1539 ( .A1(n4640), .A2(b[12]), .B1(n4639), .B2(n4792), .C(
        n4087), .ZN(n4100) );
  AOI22D1BWP12T U1540 ( .A1(b[3]), .A2(n4673), .B1(n4672), .B2(n5136), .ZN(
        n4088) );
  AOI221D1BWP12T U1541 ( .A1(n4676), .A2(b[2]), .B1(n4675), .B2(n5210), .C(
        n4088), .ZN(n4099) );
  AOI22D1BWP12T U1542 ( .A1(b[19]), .A2(n4642), .B1(n4641), .B2(n5989), .ZN(
        n4089) );
  AOI221D1BWP12T U1543 ( .A1(n4645), .A2(b[18]), .B1(n4644), .B2(n6010), .C(
        n4089), .ZN(n4098) );
  AOI22D1BWP12T U1544 ( .A1(b[15]), .A2(n4668), .B1(n4667), .B2(n4890), .ZN(
        n4090) );
  AOI221D1BWP12T U1545 ( .A1(n4671), .A2(b[14]), .B1(n4670), .B2(n5390), .C(
        n4090), .ZN(n4135) );
  AOI22D1BWP12T U1546 ( .A1(b[16]), .A2(n4632), .B1(n4631), .B2(n4793), .ZN(
        n4091) );
  AOI221D1BWP12T U1547 ( .A1(n4635), .A2(b[15]), .B1(n4634), .B2(n4890), .C(
        n4091), .ZN(n4139) );
  AOI22D1BWP12T U1548 ( .A1(b[6]), .A2(n4553), .B1(n4554), .B2(n4555), .ZN(
        n4092) );
  AOI221D1BWP12T U1549 ( .A1(n4329), .A2(b[5]), .B1(n4331), .B2(n4490), .C(
        n4092), .ZN(n4138) );
  AOI22D1BWP12T U1550 ( .A1(b[9]), .A2(n4663), .B1(n4662), .B2(n4482), .ZN(
        n4093) );
  AOI221D1BWP12T U1551 ( .A1(n4666), .A2(b[10]), .B1(n4665), .B2(n4646), .C(
        n4093), .ZN(n4137) );
  FA1D0BWP12T U1552 ( .A(n4096), .B(n4095), .CI(n4094), .CO(n4156), .S(n4133)
         );
  AOI22D1BWP12T U1553 ( .A1(b[5]), .A2(n4689), .B1(n4688), .B2(n4490), .ZN(
        n4097) );
  AOI221D1BWP12T U1554 ( .A1(n4692), .A2(b[4]), .B1(n4691), .B2(n5703), .C(
        n4097), .ZN(n4196) );
  FA1D0BWP12T U1555 ( .A(n4100), .B(n4099), .CI(n4098), .CO(n4106), .S(n4195)
         );
  AOI22D1BWP12T U1556 ( .A1(b[14]), .A2(n4668), .B1(n4667), .B2(n5390), .ZN(
        n4101) );
  AOI221D1BWP12T U1557 ( .A1(n4671), .A2(b[13]), .B1(n4670), .B2(n5476), .C(
        n4101), .ZN(n4127) );
  OAI22D1BWP12T U1558 ( .A1(b[21]), .A2(n4453), .B1(n4839), .B2(n4470), .ZN(
        n4102) );
  AOI21D1BWP12T U1559 ( .A1(n4455), .A2(n4839), .B(n4102), .ZN(n4126) );
  FA1D0BWP12T U1560 ( .A(n4105), .B(n4104), .CI(n4103), .CO(n4040), .S(n4144)
         );
  FA1D0BWP12T U1561 ( .A(n4150), .B(n4107), .CI(n4106), .CO(n4143), .S(n4119)
         );
  FA1D0BWP12T U1562 ( .A(n4110), .B(n4109), .CI(n4108), .CO(n4115), .S(n4180)
         );
  FA1D0BWP12T U1563 ( .A(n4113), .B(n4112), .CI(n4111), .CO(n4179), .S(n4145)
         );
  FA1D0BWP12T U1564 ( .A(n4116), .B(n4115), .CI(n4114), .CO(n5316), .S(n5346)
         );
  FA1D0BWP12T U1565 ( .A(n4119), .B(n4118), .CI(n4117), .CO(n4111), .S(n4187)
         );
  FA1D0BWP12T U1566 ( .A(n4122), .B(n4121), .CI(n4120), .CO(n4077), .S(n4186)
         );
  AOI22D1BWP12T U1567 ( .A1(n5380), .A2(n6067), .B1(n4455), .B2(n4740), .ZN(
        n4123) );
  OAI21D1BWP12T U1568 ( .A1(n4740), .A2(n4470), .B(n4123), .ZN(n4204) );
  AOI22D1BWP12T U1569 ( .A1(b[4]), .A2(n4329), .B1(n4331), .B2(n5703), .ZN(
        n4124) );
  OAI221D1BWP12T U1570 ( .A1(b[5]), .A2(n4554), .B1(n4490), .B2(n4553), .C(
        n4124), .ZN(n4205) );
  ND2D1BWP12T U1571 ( .A1(n4204), .A2(n4205), .ZN(n4203) );
  FA1D0BWP12T U1572 ( .A(n4127), .B(n4126), .CI(n4125), .CO(n4194), .S(n4164)
         );
  AOI22D1BWP12T U1573 ( .A1(b[10]), .A2(n4129), .B1(n4128), .B2(n4646), .ZN(
        n4130) );
  AOI21D1BWP12T U1574 ( .A1(n4131), .A2(n4148), .B(n4130), .ZN(n4235) );
  INVD1BWP12T U1575 ( .I(n4672), .ZN(n4175) );
  AOI21D1BWP12T U1576 ( .A1(n4175), .A2(n5379), .B(n4675), .ZN(n4234) );
  AOI22D1BWP12T U1577 ( .A1(b[18]), .A2(n4658), .B1(n4657), .B2(n6010), .ZN(
        n4132) );
  AOI221D1BWP12T U1578 ( .A1(n4661), .A2(b[19]), .B1(n4660), .B2(n5989), .C(
        n4132), .ZN(n4233) );
  FA1D0BWP12T U1579 ( .A(n4135), .B(n4134), .CI(n4133), .CO(n4118), .S(n4160)
         );
  AOI22D1BWP12T U1580 ( .A1(b[19]), .A2(n4658), .B1(n4657), .B2(n5989), .ZN(
        n4136) );
  AOI221D1BWP12T U1581 ( .A1(n4661), .A2(b[20]), .B1(n4660), .B2(n6067), .C(
        n4136), .ZN(n4167) );
  FA1D0BWP12T U1582 ( .A(n4139), .B(n4138), .CI(n4137), .CO(n4134), .S(n4166)
         );
  AOI22D1BWP12T U1583 ( .A1(b[17]), .A2(n4642), .B1(n4641), .B2(n4838), .ZN(
        n4140) );
  AOI221D1BWP12T U1584 ( .A1(n4645), .A2(b[16]), .B1(n4644), .B2(n4793), .C(
        n4140), .ZN(n4229) );
  AOI22D1BWP12T U1585 ( .A1(b[3]), .A2(n4689), .B1(n4688), .B2(n5136), .ZN(
        n4141) );
  AOI221D1BWP12T U1586 ( .A1(n4692), .A2(b[2]), .B1(n4691), .B2(n5210), .C(
        n4141), .ZN(n4228) );
  AOI22D1BWP12T U1587 ( .A1(b[7]), .A2(n4684), .B1(n4683), .B2(n4450), .ZN(
        n4142) );
  AOI221D1BWP12T U1588 ( .A1(n4687), .A2(b[6]), .B1(n4686), .B2(n4555), .C(
        n4142), .ZN(n4227) );
  FA1D0BWP12T U1589 ( .A(n4145), .B(n4144), .CI(n4143), .CO(n4181), .S(n4183)
         );
  AOI22D1BWP12T U1590 ( .A1(b[18]), .A2(n4642), .B1(n4641), .B2(n6010), .ZN(
        n4146) );
  AOI221D1BWP12T U1591 ( .A1(n4645), .A2(b[17]), .B1(n4644), .B2(n4838), .C(
        n4146), .ZN(n4171) );
  AOI22D1BWP12T U1592 ( .A1(b[12]), .A2(n4637), .B1(n4636), .B2(n4792), .ZN(
        n4147) );
  AOI21D1BWP12T U1593 ( .A1(n4148), .A2(n4210), .B(n4147), .ZN(n4170) );
  AOI22D1BWP12T U1594 ( .A1(b[4]), .A2(n4689), .B1(n4688), .B2(n5703), .ZN(
        n4149) );
  AOI221D1BWP12T U1595 ( .A1(n4692), .A2(b[3]), .B1(n4691), .B2(n5136), .C(
        n4149), .ZN(n4169) );
  OAI21D1BWP12T U1596 ( .A1(n4152), .A2(n4151), .B(n4150), .ZN(n4192) );
  FA1D0BWP12T U1597 ( .A(n4155), .B(n4154), .CI(n4153), .CO(n4122), .S(n4191)
         );
  FA1D0BWP12T U1598 ( .A(n4158), .B(n4157), .CI(n4156), .CO(n4076), .S(n4189)
         );
  FA1D0BWP12T U1599 ( .A(n4161), .B(n4160), .CI(n4159), .CO(n4185), .S(n4216)
         );
  AOI22D1BWP12T U1600 ( .A1(b[2]), .A2(n4673), .B1(n4672), .B2(n5210), .ZN(
        n4162) );
  AOI221D1BWP12T U1601 ( .A1(n4676), .A2(b[1]), .B1(n4675), .B2(n4419), .C(
        n4162), .ZN(n4202) );
  FA1D0BWP12T U1602 ( .A(n4203), .B(n4164), .CI(n4163), .CO(n4161), .S(n4201)
         );
  FA1D0BWP12T U1603 ( .A(n4167), .B(n4166), .CI(n4165), .CO(n4159), .S(n4200)
         );
  AOI22D1BWP12T U1604 ( .A1(b[8]), .A2(n4684), .B1(n4683), .B2(n4699), .ZN(
        n4168) );
  AOI221D1BWP12T U1605 ( .A1(n4687), .A2(b[7]), .B1(n4686), .B2(n4450), .C(
        n4168), .ZN(n4199) );
  FA1D0BWP12T U1606 ( .A(n4171), .B(n4170), .CI(n4169), .CO(n4193), .S(n4198)
         );
  INVD1BWP12T U1607 ( .I(n4673), .ZN(n4176) );
  MOAI22D0BWP12T U1608 ( .A1(n4173), .A2(n4957), .B1(n4172), .B2(n5413), .ZN(
        n4174) );
  AOI221D1BWP12T U1609 ( .A1(n4176), .A2(b[1]), .B1(n4175), .B2(n4419), .C(
        n4174), .ZN(n4208) );
  AOI22D1BWP12T U1610 ( .A1(b[13]), .A2(n4668), .B1(n4667), .B2(n5476), .ZN(
        n4177) );
  AOI221D1BWP12T U1611 ( .A1(n4671), .A2(b[12]), .B1(n4670), .B2(n4792), .C(
        n4177), .ZN(n4207) );
  AOI22D1BWP12T U1612 ( .A1(b[15]), .A2(n4632), .B1(n4631), .B2(n4890), .ZN(
        n4178) );
  AOI221D1BWP12T U1613 ( .A1(n4635), .A2(b[14]), .B1(n4634), .B2(n5390), .C(
        n4178), .ZN(n4206) );
  FA1D0BWP12T U1614 ( .A(n4181), .B(n4180), .CI(n4179), .CO(n5347), .S(n5366)
         );
  FA1D0BWP12T U1615 ( .A(n4184), .B(n4183), .CI(n4182), .CO(n5367), .S(n5364)
         );
  FA1D0BWP12T U1616 ( .A(n4187), .B(n4186), .CI(n4185), .CO(n4184), .S(n4241)
         );
  FA1D0BWP12T U1617 ( .A(n4190), .B(n4189), .CI(n4188), .CO(n4182), .S(n4240)
         );
  FA1D0BWP12T U1618 ( .A(n4193), .B(n4192), .CI(n4191), .CO(n4190), .S(n4219)
         );
  FA1D0BWP12T U1619 ( .A(n4196), .B(n4195), .CI(n4194), .CO(n4117), .S(n4218)
         );
  FA1D0BWP12T U1620 ( .A(n4199), .B(n4198), .CI(n4197), .CO(n4214), .S(n4222)
         );
  FA1D0BWP12T U1621 ( .A(n4202), .B(n4201), .CI(n4200), .CO(n4215), .S(n4221)
         );
  OAI21D1BWP12T U1622 ( .A1(n4205), .A2(n4204), .B(n4203), .ZN(n4232) );
  FA1D0BWP12T U1623 ( .A(n4208), .B(n4207), .CI(n4206), .CO(n4197), .S(n4231)
         );
  AOI22D1BWP12T U1624 ( .A1(b[10]), .A2(n4637), .B1(n4636), .B2(n4646), .ZN(
        n4209) );
  AOI21D1BWP12T U1625 ( .A1(n4211), .A2(n4210), .B(n4209), .ZN(n4251) );
  AOI22D1BWP12T U1626 ( .A1(b[2]), .A2(n4689), .B1(n4688), .B2(n5210), .ZN(
        n4212) );
  AOI221D1BWP12T U1627 ( .A1(n4692), .A2(b[1]), .B1(n4691), .B2(n4419), .C(
        n4212), .ZN(n4250) );
  AOI22D1BWP12T U1628 ( .A1(b[6]), .A2(n4684), .B1(n4683), .B2(n4555), .ZN(
        n4213) );
  AOI221D1BWP12T U1629 ( .A1(n4687), .A2(b[5]), .B1(n4686), .B2(n4490), .C(
        n4213), .ZN(n4249) );
  FA1D0BWP12T U1630 ( .A(n4216), .B(n4215), .CI(n4214), .CO(n4188), .S(n4291)
         );
  FA1D0BWP12T U1631 ( .A(n4219), .B(n4218), .CI(n4217), .CO(n4239), .S(n4290)
         );
  FA1D0BWP12T U1632 ( .A(n4222), .B(n4221), .CI(n4220), .CO(n4217), .S(n4244)
         );
  AOI22D1BWP12T U1633 ( .A1(b[8]), .A2(n4663), .B1(n4662), .B2(n4699), .ZN(
        n4223) );
  AOI221D1BWP12T U1634 ( .A1(n4666), .A2(b[9]), .B1(n4665), .B2(n4482), .C(
        n4223), .ZN(n4282) );
  AOI22D1BWP12T U1635 ( .A1(b[4]), .A2(n4553), .B1(n4554), .B2(n5703), .ZN(
        n4224) );
  AOI221D1BWP12T U1636 ( .A1(n4329), .A2(b[3]), .B1(n4331), .B2(n5136), .C(
        n4224), .ZN(n4255) );
  AOI22D1BWP12T U1637 ( .A1(b[12]), .A2(n4668), .B1(n4667), .B2(n4792), .ZN(
        n4225) );
  AOI221D1BWP12T U1638 ( .A1(n4671), .A2(b[11]), .B1(n4670), .B2(n4741), .C(
        n4225), .ZN(n4254) );
  AOI22D1BWP12T U1639 ( .A1(b[14]), .A2(n4632), .B1(n4631), .B2(n5390), .ZN(
        n4226) );
  AOI221D1BWP12T U1640 ( .A1(n4635), .A2(b[13]), .B1(n4634), .B2(n5476), .C(
        n4226), .ZN(n4253) );
  FA1D0BWP12T U1641 ( .A(n4229), .B(n4228), .CI(n4227), .CO(n4165), .S(n4280)
         );
  FA1D0BWP12T U1642 ( .A(n4232), .B(n4231), .CI(n4230), .CO(n4220), .S(n4285)
         );
  FA1D0BWP12T U1643 ( .A(n4235), .B(n4234), .CI(n4233), .CO(n4163), .S(n4284)
         );
  ND2D1BWP12T U1644 ( .A1(b[0]), .A2(n4236), .ZN(n4265) );
  OAI22D1BWP12T U1645 ( .A1(b[19]), .A2(n4453), .B1(n6067), .B2(n4470), .ZN(
        n4237) );
  AOI21D1BWP12T U1646 ( .A1(n4455), .A2(n6067), .B(n4237), .ZN(n4264) );
  AOI22D1BWP12T U1647 ( .A1(b[17]), .A2(n4658), .B1(n4657), .B2(n4838), .ZN(
        n4238) );
  AOI221D1BWP12T U1648 ( .A1(n4661), .A2(b[18]), .B1(n4660), .B2(n6010), .C(
        n4238), .ZN(n4263) );
  FA1D0BWP12T U1649 ( .A(n4241), .B(n4240), .CI(n4239), .CO(n5363), .S(n5334)
         );
  FA1D0BWP12T U1650 ( .A(n4244), .B(n4243), .CI(n4242), .CO(n4289), .S(n4294)
         );
  AOI22D1BWP12T U1651 ( .A1(b[9]), .A2(n4637), .B1(n4636), .B2(n4482), .ZN(
        n4245) );
  AOI221D1BWP12T U1652 ( .A1(n4640), .A2(b[8]), .B1(n4639), .B2(n4699), .C(
        n4245), .ZN(n4309) );
  AOI22D1BWP12T U1653 ( .A1(b[13]), .A2(n4632), .B1(n4631), .B2(n5476), .ZN(
        n4246) );
  AOI221D1BWP12T U1654 ( .A1(n4635), .A2(b[12]), .B1(n4634), .B2(n4792), .C(
        n4246), .ZN(n4308) );
  AOI22D1BWP12T U1655 ( .A1(b[16]), .A2(n4658), .B1(n4657), .B2(n4793), .ZN(
        n4247) );
  AOI221D1BWP12T U1656 ( .A1(n4661), .A2(b[17]), .B1(n4660), .B2(n4838), .C(
        n4247), .ZN(n4307) );
  AOI22D1BWP12T U1657 ( .A1(b[7]), .A2(n4663), .B1(n4662), .B2(n4450), .ZN(
        n4248) );
  AOI221D1BWP12T U1658 ( .A1(n4666), .A2(b[8]), .B1(n4665), .B2(n4699), .C(
        n4248), .ZN(n4276) );
  FA1D0BWP12T U1659 ( .A(n4251), .B(n4250), .CI(n4249), .CO(n4230), .S(n4275)
         );
  FA1D0BWP12T U1660 ( .A(n4255), .B(n4254), .CI(n4253), .CO(n4281), .S(n4279)
         );
  AOI22D1BWP12T U1661 ( .A1(n5380), .A2(n6010), .B1(n4455), .B2(n5989), .ZN(
        n4256) );
  OAI21D1BWP12T U1662 ( .A1(n5989), .A2(n4470), .B(n4256), .ZN(n4305) );
  AOI22D1BWP12T U1663 ( .A1(b[2]), .A2(n4329), .B1(n4331), .B2(n5210), .ZN(
        n4257) );
  OAI221D1BWP12T U1664 ( .A1(b[3]), .A2(n4554), .B1(n5136), .B2(n4553), .C(
        n4257), .ZN(n4306) );
  ND2D1BWP12T U1665 ( .A1(n4305), .A2(n4306), .ZN(n4304) );
  AOI22D1BWP12T U1666 ( .A1(b[15]), .A2(n4642), .B1(n4641), .B2(n4890), .ZN(
        n4258) );
  AOI221D1BWP12T U1667 ( .A1(n4645), .A2(b[14]), .B1(n4644), .B2(n5390), .C(
        n4258), .ZN(n4316) );
  AOI22D1BWP12T U1668 ( .A1(b[5]), .A2(n4684), .B1(n4683), .B2(n4490), .ZN(
        n4259) );
  AOI221D1BWP12T U1669 ( .A1(n4687), .A2(b[4]), .B1(n4686), .B2(n5703), .C(
        n4259), .ZN(n4315) );
  AOI22D1BWP12T U1670 ( .A1(b[6]), .A2(n4663), .B1(n4662), .B2(n4555), .ZN(
        n4260) );
  AOI221D1BWP12T U1671 ( .A1(n4666), .A2(b[7]), .B1(n4665), .B2(n4450), .C(
        n4260), .ZN(n4314) );
  AOI22D1BWP12T U1672 ( .A1(b[16]), .A2(n4642), .B1(n4641), .B2(n4793), .ZN(
        n4262) );
  AOI221D1BWP12T U1673 ( .A1(n4645), .A2(b[15]), .B1(n4644), .B2(n4890), .C(
        n4262), .ZN(n4288) );
  FA1D0BWP12T U1674 ( .A(n4265), .B(n4264), .CI(n4263), .CO(n4283), .S(n4287)
         );
  RCIAO21D0BWP12T U1675 ( .A1(n4266), .A2(n4268), .B(n4691), .ZN(n4322) );
  MAOI22D0BWP12T U1676 ( .A1(n4970), .A2(n4268), .B1(n4267), .B2(n4266), .ZN(
        n4269) );
  OA221D1BWP12T U1677 ( .A1(n4689), .A2(n4419), .B1(n4688), .B2(b[1]), .C(
        n4269), .Z(n4321) );
  ND2D1BWP12T U1678 ( .A1(b[0]), .A2(n4270), .ZN(n4327) );
  OAI22D1BWP12T U1679 ( .A1(b[17]), .A2(n4453), .B1(n6010), .B2(n4470), .ZN(
        n4271) );
  AOI21D1BWP12T U1680 ( .A1(n4455), .A2(n6010), .B(n4271), .ZN(n4326) );
  AOI22D1BWP12T U1681 ( .A1(b[15]), .A2(n4658), .B1(n4657), .B2(n4890), .ZN(
        n4272) );
  AOI221D1BWP12T U1682 ( .A1(n4661), .A2(b[16]), .B1(n4660), .B2(n4793), .C(
        n4272), .ZN(n4325) );
  INVD1BWP12T U1683 ( .I(n4274), .ZN(n4297) );
  FA1D0BWP12T U1684 ( .A(n4277), .B(n4276), .CI(n4275), .CO(n4296), .S(n4252)
         );
  FA1D0BWP12T U1685 ( .A(n4279), .B(n4304), .CI(n4278), .CO(n4295), .S(n4261)
         );
  FA1D0BWP12T U1686 ( .A(n4282), .B(n4281), .CI(n4280), .CO(n4243), .S(n4300)
         );
  FA1D0BWP12T U1687 ( .A(n4285), .B(n4284), .CI(n4283), .CO(n4242), .S(n4299)
         );
  FA1D0BWP12T U1688 ( .A(n4288), .B(n4287), .CI(n4286), .CO(n4298), .S(n4273)
         );
  FA1D0BWP12T U1689 ( .A(n4291), .B(n4290), .CI(n4289), .CO(n5335), .S(n5331)
         );
  FA1D0BWP12T U1690 ( .A(n4294), .B(n4293), .CI(n4292), .CO(n5332), .S(n5314)
         );
  FA1D0BWP12T U1691 ( .A(n4297), .B(n4296), .CI(n4295), .CO(n4293), .S(n4364)
         );
  FA1D0BWP12T U1692 ( .A(n4300), .B(n4299), .CI(n4298), .CO(n4292), .S(n4363)
         );
  AOI22D1BWP12T U1693 ( .A1(b[8]), .A2(n4637), .B1(n4636), .B2(n4699), .ZN(
        n4301) );
  AOI221D1BWP12T U1694 ( .A1(n4640), .A2(b[7]), .B1(n4639), .B2(n4450), .C(
        n4301), .ZN(n4356) );
  AOI22D1BWP12T U1695 ( .A1(b[14]), .A2(n4642), .B1(n4641), .B2(n5390), .ZN(
        n4302) );
  AOI221D1BWP12T U1696 ( .A1(n4645), .A2(b[13]), .B1(n4644), .B2(n5476), .C(
        n4302), .ZN(n4355) );
  AOI22D1BWP12T U1697 ( .A1(b[4]), .A2(n4684), .B1(n4683), .B2(n5703), .ZN(
        n4303) );
  AOI221D1BWP12T U1698 ( .A1(n4687), .A2(b[3]), .B1(n4686), .B2(n5136), .C(
        n4303), .ZN(n4354) );
  OAI21D1BWP12T U1699 ( .A1(n4306), .A2(n4305), .B(n4304), .ZN(n4318) );
  FA1D0BWP12T U1700 ( .A(n4309), .B(n4308), .CI(n4307), .CO(n4277), .S(n4317)
         );
  AOI22D1BWP12T U1701 ( .A1(b[11]), .A2(n4668), .B1(n4667), .B2(n4741), .ZN(
        n4310) );
  AOI221D1BWP12T U1702 ( .A1(n4671), .A2(b[10]), .B1(n4670), .B2(n4646), .C(
        n4310), .ZN(n4351) );
  AOI22D1BWP12T U1703 ( .A1(b[2]), .A2(n4553), .B1(n4554), .B2(n5210), .ZN(
        n4311) );
  AOI221D1BWP12T U1704 ( .A1(n4329), .A2(b[1]), .B1(n4331), .B2(n4419), .C(
        n4311), .ZN(n4348) );
  AOI22D1BWP12T U1705 ( .A1(b[5]), .A2(n4663), .B1(n4662), .B2(n4490), .ZN(
        n4312) );
  AOI221D1BWP12T U1706 ( .A1(n4666), .A2(b[6]), .B1(n4665), .B2(n4555), .C(
        n4312), .ZN(n4347) );
  AOI22D1BWP12T U1707 ( .A1(b[10]), .A2(n4668), .B1(n4667), .B2(n4646), .ZN(
        n4313) );
  FA1D0BWP12T U1708 ( .A(n4316), .B(n4315), .CI(n4314), .CO(n4278), .S(n4349)
         );
  FA1D0BWP12T U1709 ( .A(n4319), .B(n4318), .CI(n4317), .CO(n4337), .S(n4373)
         );
  FA1D0BWP12T U1710 ( .A(n4322), .B(n4321), .CI(n4320), .CO(n4286), .S(n4372)
         );
  AOI22D1BWP12T U1711 ( .A1(n5380), .A2(n4793), .B1(n4455), .B2(n4838), .ZN(
        n4323) );
  OAI21D1BWP12T U1712 ( .A1(n4838), .A2(n4470), .B(n4323), .ZN(n4375) );
  OAI21D1BWP12T U1713 ( .A1(b[0]), .A2(n4554), .B(n4324), .ZN(n4376) );
  ND2D1BWP12T U1714 ( .A1(n4375), .A2(n4376), .ZN(n4374) );
  FA1D0BWP12T U1715 ( .A(n4327), .B(n4326), .CI(n4325), .CO(n4320), .S(n4353)
         );
  OAI21D1BWP12T U1716 ( .A1(a[17]), .A2(n4419), .B(n4328), .ZN(n4332) );
  AOI222D1BWP12T U1717 ( .A1(n4332), .A2(n4359), .B1(n5379), .B2(n4331), .C1(
        n4330), .C2(n4329), .ZN(n4392) );
  AOI22D1BWP12T U1718 ( .A1(b[7]), .A2(n4637), .B1(n4636), .B2(n4450), .ZN(
        n4333) );
  AOI221D1BWP12T U1719 ( .A1(n4640), .A2(b[6]), .B1(n4639), .B2(n4555), .C(
        n4333), .ZN(n4391) );
  AOI22D1BWP12T U1720 ( .A1(b[14]), .A2(n4658), .B1(n4657), .B2(n5390), .ZN(
        n4334) );
  AOI221D1BWP12T U1721 ( .A1(n4661), .A2(b[15]), .B1(n4660), .B2(n4890), .C(
        n4334), .ZN(n4390) );
  FA1D0BWP12T U1722 ( .A(n4337), .B(n4336), .CI(n4335), .CO(n4362), .S(n4367)
         );
  INVD1BWP12T U1723 ( .I(n4338), .ZN(n4366) );
  AOI22D1BWP12T U1724 ( .A1(b[12]), .A2(n4632), .B1(n4631), .B2(n4792), .ZN(
        n4339) );
  AOI221D1BWP12T U1725 ( .A1(n4635), .A2(b[11]), .B1(n4634), .B2(n4741), .C(
        n4339), .ZN(n4386) );
  AOI22D1BWP12T U1726 ( .A1(b[13]), .A2(n4642), .B1(n4641), .B2(n5476), .ZN(
        n4340) );
  AOI221D1BWP12T U1727 ( .A1(n4645), .A2(b[12]), .B1(n4644), .B2(n4792), .C(
        n4340), .ZN(n4383) );
  MAOI22D0BWP12T U1728 ( .A1(b[8]), .A2(n4341), .B1(n4670), .B2(b[8]), .ZN(
        n4342) );
  AOI21D1BWP12T U1729 ( .A1(n4344), .A2(n4343), .B(n4342), .ZN(n4382) );
  AOI22D1BWP12T U1730 ( .A1(b[11]), .A2(n4632), .B1(n4631), .B2(n4741), .ZN(
        n4345) );
  AOI221D1BWP12T U1731 ( .A1(n4635), .A2(b[10]), .B1(n4634), .B2(n4646), .C(
        n4345), .ZN(n4381) );
  FA1D0BWP12T U1732 ( .A(n4348), .B(n4347), .CI(n4346), .CO(n4350), .S(n4384)
         );
  FA1D0BWP12T U1733 ( .A(n4351), .B(n4350), .CI(n4349), .CO(n4336), .S(n4369)
         );
  FA1D0BWP12T U1734 ( .A(n4374), .B(n4353), .CI(n4352), .CO(n4371), .S(n4401)
         );
  FA1D0BWP12T U1735 ( .A(n4356), .B(n4355), .CI(n4354), .CO(n4319), .S(n4400)
         );
  AOI22D1BWP12T U1736 ( .A1(b[3]), .A2(n4684), .B1(n4683), .B2(n5136), .ZN(
        n4357) );
  AOI221D1BWP12T U1737 ( .A1(n4687), .A2(b[2]), .B1(n4686), .B2(n5210), .C(
        n4357), .ZN(n4389) );
  AOI22D1BWP12T U1738 ( .A1(b[4]), .A2(n4663), .B1(n4662), .B2(n5703), .ZN(
        n4358) );
  AOI221D1BWP12T U1739 ( .A1(n4666), .A2(b[5]), .B1(n4665), .B2(n4490), .C(
        n4358), .ZN(n4388) );
  ND2D1BWP12T U1740 ( .A1(b[0]), .A2(n4359), .ZN(n4413) );
  OAI22D1BWP12T U1741 ( .A1(b[15]), .A2(n4453), .B1(n4793), .B2(n4470), .ZN(
        n4360) );
  AOI21D1BWP12T U1742 ( .A1(n4455), .A2(n4793), .B(n4360), .ZN(n4412) );
  AOI22D1BWP12T U1743 ( .A1(b[13]), .A2(n4658), .B1(n4657), .B2(n5476), .ZN(
        n4361) );
  AOI221D1BWP12T U1744 ( .A1(n4661), .A2(b[14]), .B1(n4660), .B2(n5390), .C(
        n4361), .ZN(n4411) );
  FA1D0BWP12T U1745 ( .A(n4364), .B(n4363), .CI(n4362), .CO(n5313), .S(n5328)
         );
  FA1D0BWP12T U1746 ( .A(n4367), .B(n4366), .CI(n4365), .CO(n5329), .S(n5323)
         );
  FA1D0BWP12T U1747 ( .A(n4370), .B(n4369), .CI(n4368), .CO(n4365), .S(n4426)
         );
  FA1D0BWP12T U1748 ( .A(n4373), .B(n4372), .CI(n4371), .CO(n4335), .S(n4425)
         );
  OAI21D1BWP12T U1749 ( .A1(n4376), .A2(n4375), .B(n4374), .ZN(n4404) );
  AOI22D1BWP12T U1750 ( .A1(b[12]), .A2(n4642), .B1(n4641), .B2(n4792), .ZN(
        n4377) );
  AOI221D1BWP12T U1751 ( .A1(n4645), .A2(b[11]), .B1(n4644), .B2(n4741), .C(
        n4377), .ZN(n4407) );
  AOI21D1BWP12T U1752 ( .A1(n5872), .A2(b[1]), .B(n4378), .ZN(n4487) );
  AOI22D1BWP12T U1753 ( .A1(b[2]), .A2(n4684), .B1(n4683), .B2(n5210), .ZN(
        n4379) );
  AOI21D1BWP12T U1754 ( .A1(n4487), .A2(n4421), .B(n4379), .ZN(n4406) );
  AOI22D1BWP12T U1755 ( .A1(b[3]), .A2(n4663), .B1(n4662), .B2(n5136), .ZN(
        n4380) );
  AOI221D1BWP12T U1756 ( .A1(n4666), .A2(b[4]), .B1(n4665), .B2(n5703), .C(
        n4380), .ZN(n4405) );
  FA1D0BWP12T U1757 ( .A(n4383), .B(n4382), .CI(n4381), .CO(n4385), .S(n4402)
         );
  FA1D0BWP12T U1758 ( .A(n4386), .B(n4385), .CI(n4384), .CO(n4370), .S(n4397)
         );
  FA1D0BWP12T U1759 ( .A(n4389), .B(n4388), .CI(n4387), .CO(n4399), .S(n4435)
         );
  FA1D0BWP12T U1760 ( .A(n4392), .B(n4391), .CI(n4390), .CO(n4352), .S(n4434)
         );
  AOI22D1BWP12T U1761 ( .A1(b[6]), .A2(n4637), .B1(n4636), .B2(n4555), .ZN(
        n4393) );
  AOI221D1BWP12T U1762 ( .A1(n4640), .A2(b[5]), .B1(n4639), .B2(n4490), .C(
        n4393), .ZN(n4416) );
  AOI22D1BWP12T U1763 ( .A1(b[8]), .A2(n4668), .B1(n4667), .B2(n4699), .ZN(
        n4394) );
  AOI221D1BWP12T U1764 ( .A1(n4671), .A2(b[7]), .B1(n4670), .B2(n4450), .C(
        n4394), .ZN(n4415) );
  AOI22D1BWP12T U1765 ( .A1(b[10]), .A2(n4632), .B1(n4631), .B2(n4646), .ZN(
        n4395) );
  AOI221D1BWP12T U1766 ( .A1(n4635), .A2(b[9]), .B1(n4634), .B2(n4482), .C(
        n4395), .ZN(n4414) );
  FA1D0BWP12T U1767 ( .A(n4398), .B(n4397), .CI(n4396), .CO(n4424), .S(n4429)
         );
  FA1D0BWP12T U1768 ( .A(n4401), .B(n4400), .CI(n4399), .CO(n4368), .S(n4428)
         );
  FA1D0BWP12T U1769 ( .A(n4404), .B(n4403), .CI(n4402), .CO(n4398), .S(n4432)
         );
  FA1D0BWP12T U1770 ( .A(n4407), .B(n4406), .CI(n4405), .CO(n4403), .S(n4462)
         );
  AOI22D1BWP12T U1771 ( .A1(b[12]), .A2(n4658), .B1(n4657), .B2(n4792), .ZN(
        n4408) );
  AOI221D1BWP12T U1772 ( .A1(n4661), .A2(b[13]), .B1(n4660), .B2(n5476), .C(
        n4408), .ZN(n4446) );
  AOI22D1BWP12T U1773 ( .A1(b[11]), .A2(n4642), .B1(n4641), .B2(n4741), .ZN(
        n4409) );
  AOI221D1BWP12T U1774 ( .A1(n4645), .A2(b[10]), .B1(n4644), .B2(n4646), .C(
        n4409), .ZN(n4445) );
  AOI22D1BWP12T U1775 ( .A1(b[9]), .A2(n4632), .B1(n4631), .B2(n4482), .ZN(
        n4410) );
  AOI221D1BWP12T U1776 ( .A1(n4635), .A2(b[8]), .B1(n4634), .B2(n4699), .C(
        n4410), .ZN(n4444) );
  FA1D0BWP12T U1777 ( .A(n4413), .B(n4412), .CI(n4411), .CO(n4387), .S(n4460)
         );
  FA1D0BWP12T U1778 ( .A(n4416), .B(n4415), .CI(n4414), .CO(n4433), .S(n4437)
         );
  AOI22D1BWP12T U1779 ( .A1(b[4]), .A2(n4640), .B1(n4639), .B2(n5703), .ZN(
        n4417) );
  OAI221D1BWP12T U1780 ( .A1(b[5]), .A2(n4636), .B1(n4490), .B2(n4637), .C(
        n4417), .ZN(n4439) );
  AOI22D1BWP12T U1781 ( .A1(n5380), .A2(n5390), .B1(n4455), .B2(n4890), .ZN(
        n4418) );
  OAI21D1BWP12T U1782 ( .A1(n4890), .A2(n4470), .B(n4418), .ZN(n4440) );
  ND2D1BWP12T U1783 ( .A1(n4439), .A2(n4440), .ZN(n4438) );
  AOI22D1BWP12T U1784 ( .A1(b[1]), .A2(n4684), .B1(n4683), .B2(n4419), .ZN(
        n4420) );
  AOI21D1BWP12T U1785 ( .A1(n4974), .A2(n4421), .B(n4420), .ZN(n4449) );
  OA21D1BWP12T U1786 ( .A1(n4683), .A2(b[0]), .B(n4422), .Z(n4448) );
  AOI22D1BWP12T U1787 ( .A1(b[2]), .A2(n4663), .B1(n4662), .B2(n5210), .ZN(
        n4423) );
  AOI221D1BWP12T U1788 ( .A1(n4666), .A2(b[3]), .B1(n4665), .B2(n5136), .C(
        n4423), .ZN(n4447) );
  FA1D0BWP12T U1789 ( .A(n4426), .B(n4425), .CI(n4424), .CO(n5322), .S(n5325)
         );
  FA1D0BWP12T U1790 ( .A(n4429), .B(n4428), .CI(n4427), .CO(n5326), .S(n5309)
         );
  FA1D0BWP12T U1791 ( .A(n4432), .B(n4431), .CI(n4430), .CO(n4427), .S(n4480)
         );
  FA1D0BWP12T U1792 ( .A(n4435), .B(n4434), .CI(n4433), .CO(n4396), .S(n4479)
         );
  FA1D0BWP12T U1793 ( .A(n4437), .B(n4438), .CI(n4436), .CO(n4430), .S(n4459)
         );
  OAI21D1BWP12T U1794 ( .A1(n4440), .A2(n4439), .B(n4438), .ZN(n4465) );
  AOI22D1BWP12T U1795 ( .A1(b[4]), .A2(n4637), .B1(n4636), .B2(n5703), .ZN(
        n4441) );
  AOI221D1BWP12T U1796 ( .A1(n4640), .A2(b[3]), .B1(n4639), .B2(n5136), .C(
        n4441), .ZN(n4486) );
  NR2D1BWP12T U1797 ( .A1(n4489), .A2(n4487), .ZN(n4442) );
  AOI221D1BWP12T U1798 ( .A1(n4666), .A2(b[2]), .B1(n4665), .B2(n5210), .C(
        n4442), .ZN(n4485) );
  AOI22D1BWP12T U1799 ( .A1(b[6]), .A2(n4668), .B1(n4667), .B2(n4555), .ZN(
        n4443) );
  AOI221D1BWP12T U1800 ( .A1(n4671), .A2(b[5]), .B1(n4670), .B2(n4490), .C(
        n4443), .ZN(n4484) );
  FA1D0BWP12T U1801 ( .A(n4446), .B(n4445), .CI(n4444), .CO(n4461), .S(n4463)
         );
  FA1D0BWP12T U1802 ( .A(n4449), .B(n4448), .CI(n4447), .CO(n4436), .S(n4468)
         );
  AOI22D1BWP12T U1803 ( .A1(b[7]), .A2(n4668), .B1(n4667), .B2(n4450), .ZN(
        n4451) );
  AOI221D1BWP12T U1804 ( .A1(n4671), .A2(b[6]), .B1(n4670), .B2(n4555), .C(
        n4451), .ZN(n4467) );
  ND2D1BWP12T U1805 ( .A1(b[0]), .A2(n4452), .ZN(n4474) );
  OAI22D1BWP12T U1806 ( .A1(b[13]), .A2(n4453), .B1(n5390), .B2(n4470), .ZN(
        n4454) );
  AOI21D1BWP12T U1807 ( .A1(n4455), .A2(n5390), .B(n4454), .ZN(n4473) );
  AOI22D1BWP12T U1808 ( .A1(b[11]), .A2(n4658), .B1(n4657), .B2(n4741), .ZN(
        n4456) );
  AOI221D1BWP12T U1809 ( .A1(n4661), .A2(b[12]), .B1(n4660), .B2(n4792), .C(
        n4456), .ZN(n4472) );
  FA1D0BWP12T U1810 ( .A(n4459), .B(n4458), .CI(n4457), .CO(n4478), .S(n4506)
         );
  FA1D0BWP12T U1811 ( .A(n4462), .B(n4461), .CI(n4460), .CO(n4431), .S(n4505)
         );
  FA1D0BWP12T U1812 ( .A(n4465), .B(n4464), .CI(n4463), .CO(n4458), .S(n4500)
         );
  FA1D0BWP12T U1813 ( .A(n4468), .B(n4467), .CI(n4466), .CO(n4457), .S(n4499)
         );
  AOI22D1BWP12T U1814 ( .A1(n5380), .A2(n4792), .B1(n4455), .B2(n5476), .ZN(
        n4469) );
  OAI21D1BWP12T U1815 ( .A1(n5476), .A2(n4470), .B(n4469), .ZN(n4511) );
  AOI22D1BWP12T U1816 ( .A1(b[2]), .A2(n4640), .B1(n4639), .B2(n5210), .ZN(
        n4471) );
  OAI221D1BWP12T U1817 ( .A1(b[3]), .A2(n4636), .B1(n5136), .B2(n4637), .C(
        n4471), .ZN(n4512) );
  ND2D1BWP12T U1818 ( .A1(n4511), .A2(n4512), .ZN(n4510) );
  FA1D0BWP12T U1819 ( .A(n4474), .B(n4473), .CI(n4472), .CO(n4466), .S(n4497)
         );
  AOI22D1BWP12T U1820 ( .A1(b[9]), .A2(n4642), .B1(n4641), .B2(n4482), .ZN(
        n4475) );
  AOI221D0BWP12T U1821 ( .A1(n4645), .A2(b[8]), .B1(n4644), .B2(n4699), .C(
        n4475), .ZN(n4527) );
  AOI21D1BWP12T U1822 ( .A1(n4665), .A2(n5379), .B(n4476), .ZN(n4526) );
  AOI22D1BWP12T U1823 ( .A1(b[10]), .A2(n4658), .B1(n4657), .B2(n4646), .ZN(
        n4477) );
  AOI221D1BWP12T U1824 ( .A1(n4661), .A2(b[11]), .B1(n4660), .B2(n4741), .C(
        n4477), .ZN(n4525) );
  FA1D0BWP12T U1825 ( .A(n4480), .B(n4479), .CI(n4478), .CO(n5308), .S(n5356)
         );
  AOI22D1BWP12T U1826 ( .A1(b[10]), .A2(n4642), .B1(n4641), .B2(n4646), .ZN(
        n4481) );
  AOI221D1BWP12T U1827 ( .A1(n4645), .A2(b[9]), .B1(n4644), .B2(n4482), .C(
        n4481), .ZN(n4521) );
  AOI22D1BWP12T U1828 ( .A1(b[8]), .A2(n4632), .B1(n4631), .B2(n4699), .ZN(
        n4483) );
  AOI21D1BWP12T U1829 ( .A1(n4495), .A2(n4492), .B(n4483), .ZN(n4503) );
  FA1D0BWP12T U1830 ( .A(n4486), .B(n4485), .CI(n4484), .CO(n4464), .S(n4502)
         );
  AOI22D1BWP12T U1831 ( .A1(b[0]), .A2(a[12]), .B1(a[13]), .B2(n5379), .ZN(
        n5249) );
  OA22D1BWP12T U1832 ( .A1(n5249), .A2(n4489), .B1(n4488), .B2(n4487), .Z(
        n4515) );
  AOI22D1BWP12T U1833 ( .A1(b[5]), .A2(n4668), .B1(n4667), .B2(n4490), .ZN(
        n4491) );
  AOI221D1BWP12T U1834 ( .A1(n4671), .A2(b[4]), .B1(n4670), .B2(n5703), .C(
        n4491), .ZN(n4514) );
  AOI22D1BWP12T U1835 ( .A1(n4495), .A2(n4494), .B1(n4493), .B2(n4492), .ZN(
        n4513) );
  FA1D0BWP12T U1836 ( .A(n4510), .B(n4497), .CI(n4496), .CO(n4498), .S(n4519)
         );
  FA1D0BWP12T U1837 ( .A(n4500), .B(n4499), .CI(n4498), .CO(n4504), .S(n4508)
         );
  FA1D0BWP12T U1838 ( .A(n4503), .B(n4502), .CI(n4501), .CO(n4507), .S(n4520)
         );
  FA1D0BWP12T U1839 ( .A(n4506), .B(n4505), .CI(n4504), .CO(n5357), .S(n5353)
         );
  FA1D0BWP12T U1840 ( .A(n4509), .B(n4508), .CI(n4507), .CO(n5354), .S(n5306)
         );
  OAI21D1BWP12T U1841 ( .A1(n4512), .A2(n4511), .B(n4510), .ZN(n4533) );
  FA1D0BWP12T U1842 ( .A(n4515), .B(n4514), .CI(n4513), .CO(n4501), .S(n4532)
         );
  FA1D0BWP12T U1843 ( .A(n4521), .B(n4520), .CI(n4519), .CO(n4509), .S(n4541)
         );
  FA1D0BWP12T U1844 ( .A(n4527), .B(n4526), .CI(n4525), .CO(n4496), .S(n4535)
         );
  FA1D0BWP12T U1845 ( .A(n4533), .B(n4532), .CI(n4531), .CO(n4542), .S(n4545)
         );
  FA1D0BWP12T U1846 ( .A(n4536), .B(n4535), .CI(n4534), .CO(n4540), .S(n4544)
         );
  FA1D0BWP12T U1847 ( .A(n4542), .B(n4541), .CI(n4540), .CO(n5305), .S(n5350)
         );
  FA1D0BWP12T U1848 ( .A(n4545), .B(n4544), .CI(n4543), .CO(n5351), .S(n5361)
         );
  OA33D1BWP12T U1849 ( .A1(n5710), .A2(n5392), .A3(a[17]), .B1(n5679), .B2(
        n6043), .B3(a[16]), .Z(n4552) );
  OAI221D1BWP12T U1850 ( .A1(b[16]), .A2(n4554), .B1(n4793), .B2(n4553), .C(
        n4552), .ZN(n4630) );
  AOI22D1BWP12T U1851 ( .A1(a[27]), .A2(b[6]), .B1(n4555), .B2(n5758), .ZN(
        n4556) );
  AOI22D1BWP12T U1852 ( .A1(n4559), .A2(n4558), .B1(n4557), .B2(n4556), .ZN(
        n4628) );
  FA1D0BWP12T U1853 ( .A(n4562), .B(n4561), .CI(n4560), .CO(n4567), .S(n4709)
         );
  FA1D0BWP12T U1854 ( .A(n4565), .B(n4564), .CI(n4563), .CO(n4566), .S(n4612)
         );
  MAOI22D0BWP12T U1855 ( .A1(n4567), .A2(n4566), .B1(n4567), .B2(n4566), .ZN(
        n4597) );
  FA1D0BWP12T U1856 ( .A(n4570), .B(n4569), .CI(n4568), .CO(n4575), .S(n4580)
         );
  FA1D0BWP12T U1857 ( .A(n4573), .B(n4572), .CI(n4571), .CO(n4574), .S(n4579)
         );
  MAOI22D0BWP12T U1858 ( .A1(n4575), .A2(n4574), .B1(n4575), .B2(n4574), .ZN(
        n4595) );
  FA1D0BWP12T U1859 ( .A(n4578), .B(n4577), .CI(n4576), .CO(n4583), .S(n4606)
         );
  FA1D0BWP12T U1860 ( .A(n4581), .B(n4580), .CI(n4579), .CO(n4582), .S(n4609)
         );
  MAOI22D0BWP12T U1861 ( .A1(n4583), .A2(n4582), .B1(n4583), .B2(n4582), .ZN(
        n4593) );
  FA1D0BWP12T U1862 ( .A(n4586), .B(n4585), .CI(n4584), .CO(n4591), .S(n4589)
         );
  FA1D0BWP12T U1863 ( .A(n4589), .B(n4588), .CI(n4587), .CO(n4590), .S(n4573)
         );
  MAOI22D0BWP12T U1864 ( .A1(n4591), .A2(n4590), .B1(n4591), .B2(n4590), .ZN(
        n4592) );
  MAOI22D0BWP12T U1865 ( .A1(n4593), .A2(n4592), .B1(n4593), .B2(n4592), .ZN(
        n4594) );
  MAOI22D0BWP12T U1866 ( .A1(n4595), .A2(n4594), .B1(n4595), .B2(n4594), .ZN(
        n4596) );
  MAOI22D0BWP12T U1867 ( .A1(n4597), .A2(n4596), .B1(n4597), .B2(n4596), .ZN(
        n4626) );
  OA211D1BWP12T U1868 ( .A1(b[2]), .A2(a[31]), .B(n4599), .C(n4598), .Z(n4602)
         );
  INR2D1BWP12T U1869 ( .A1(n4600), .B1(n5417), .ZN(n4601) );
  AOI211D1BWP12T U1870 ( .A1(n4604), .A2(n4603), .B(n4602), .C(n4601), .ZN(
        n4624) );
  FA1D0BWP12T U1871 ( .A(n4607), .B(n4606), .CI(n4605), .CO(n4622), .S(n4587)
         );
  FA1D0BWP12T U1872 ( .A(n4610), .B(n4609), .CI(n4608), .CO(n4620), .S(n4706)
         );
  FA1D0BWP12T U1873 ( .A(n4613), .B(n4612), .CI(n4611), .CO(n4618), .S(n4588)
         );
  FA1D0BWP12T U1874 ( .A(n4616), .B(n4615), .CI(n4614), .CO(n4617), .S(n4569)
         );
  MOAI22D0BWP12T U1875 ( .A1(n4618), .A2(n4617), .B1(n4618), .B2(n4617), .ZN(
        n4619) );
  MAOI22D0BWP12T U1876 ( .A1(n4620), .A2(n4619), .B1(n4620), .B2(n4619), .ZN(
        n4621) );
  MAOI22D0BWP12T U1877 ( .A1(n4622), .A2(n4621), .B1(n4622), .B2(n4621), .ZN(
        n4623) );
  MAOI22D0BWP12T U1878 ( .A1(n4624), .A2(n4623), .B1(n4624), .B2(n4623), .ZN(
        n4625) );
  MAOI22D0BWP12T U1879 ( .A1(n4626), .A2(n4625), .B1(n4626), .B2(n4625), .ZN(
        n4627) );
  MAOI22D0BWP12T U1880 ( .A1(n4628), .A2(n4627), .B1(n4628), .B2(n4627), .ZN(
        n4629) );
  MAOI22D0BWP12T U1881 ( .A1(n4630), .A2(n4629), .B1(n4630), .B2(n4629), .ZN(
        n4732) );
  AOI22D1BWP12T U1882 ( .A1(b[26]), .A2(n4632), .B1(n4631), .B2(n5784), .ZN(
        n4633) );
  AOI221D1BWP12T U1883 ( .A1(n4635), .A2(b[25]), .B1(n4634), .B2(n4739), .C(
        n4633), .ZN(n4656) );
  AOI22D1BWP12T U1884 ( .A1(b[22]), .A2(n4637), .B1(n4636), .B2(n4839), .ZN(
        n4638) );
  AOI221D1BWP12T U1885 ( .A1(n4640), .A2(b[21]), .B1(n4639), .B2(n4740), .C(
        n4638), .ZN(n4654) );
  AOI22D1BWP12T U1886 ( .A1(b[28]), .A2(n4642), .B1(n4641), .B2(n5722), .ZN(
        n4643) );
  AOI221D1BWP12T U1887 ( .A1(n4645), .A2(b[27]), .B1(n4644), .B2(n5751), .C(
        n4643), .ZN(n4652) );
  AOI22D1BWP12T U1888 ( .A1(a[23]), .A2(b[10]), .B1(n4646), .B2(n5951), .ZN(
        n4647) );
  AOI22D1BWP12T U1889 ( .A1(n4650), .A2(n4649), .B1(n4648), .B2(n4647), .ZN(
        n4651) );
  MAOI22D0BWP12T U1890 ( .A1(n4652), .A2(n4651), .B1(n4652), .B2(n4651), .ZN(
        n4653) );
  MAOI22D0BWP12T U1891 ( .A1(n4654), .A2(n4653), .B1(n4654), .B2(n4653), .ZN(
        n4655) );
  MAOI22D0BWP12T U1892 ( .A1(n4656), .A2(n4655), .B1(n4656), .B2(n4655), .ZN(
        n4730) );
  AOI22D1BWP12T U1893 ( .A1(b[29]), .A2(n4658), .B1(n4657), .B2(n4841), .ZN(
        n4659) );
  AOI221D1BWP12T U1894 ( .A1(n4661), .A2(b[30]), .B1(n4660), .B2(n4737), .C(
        n4659), .ZN(n4682) );
  AOI22D1BWP12T U1895 ( .A1(b[19]), .A2(n4663), .B1(n4662), .B2(n5989), .ZN(
        n4664) );
  AOI221D1BWP12T U1896 ( .A1(n4666), .A2(b[20]), .B1(n4665), .B2(n6067), .C(
        n4664), .ZN(n4680) );
  AOI22D1BWP12T U1897 ( .A1(b[24]), .A2(n4668), .B1(n4667), .B2(n5918), .ZN(
        n4669) );
  AOI221D1BWP12T U1898 ( .A1(n4671), .A2(b[23]), .B1(n4670), .B2(n5940), .C(
        n4669), .ZN(n4678) );
  AOI22D1BWP12T U1899 ( .A1(b[12]), .A2(n4673), .B1(n4672), .B2(n4792), .ZN(
        n4674) );
  AOI221D1BWP12T U1900 ( .A1(n4676), .A2(b[11]), .B1(n4675), .B2(n4741), .C(
        n4674), .ZN(n4677) );
  MAOI22D0BWP12T U1901 ( .A1(n4678), .A2(n4677), .B1(n4678), .B2(n4677), .ZN(
        n4679) );
  MAOI22D0BWP12T U1902 ( .A1(n4680), .A2(n4679), .B1(n4680), .B2(n4679), .ZN(
        n4681) );
  MAOI22D0BWP12T U1903 ( .A1(n4682), .A2(n4681), .B1(n4682), .B2(n4681), .ZN(
        n4728) );
  AOI22D1BWP12T U1904 ( .A1(b[18]), .A2(n4684), .B1(n4683), .B2(n6010), .ZN(
        n4685) );
  AOI221D1BWP12T U1905 ( .A1(n4687), .A2(b[17]), .B1(n4686), .B2(n4838), .C(
        n4685), .ZN(n4726) );
  AOI22D1BWP12T U1906 ( .A1(b[14]), .A2(n4689), .B1(n4688), .B2(n5390), .ZN(
        n4690) );
  AOI221D1BWP12T U1907 ( .A1(n4692), .A2(b[13]), .B1(n4691), .B2(n5476), .C(
        n4690), .ZN(n4724) );
  AOI22D1BWP12T U1908 ( .A1(a[29]), .A2(b[4]), .B1(n5703), .B2(n5901), .ZN(
        n4693) );
  AOI22D1BWP12T U1909 ( .A1(n4696), .A2(n4695), .B1(n4694), .B2(n4693), .ZN(
        n4697) );
  MAOI22D0BWP12T U1910 ( .A1(n4698), .A2(n4697), .B1(n4698), .B2(n4697), .ZN(
        n4722) );
  OAI32D1BWP12T U1911 ( .A1(a[1]), .A2(n5595), .A3(n5633), .B1(b[31]), .B2(
        n5805), .ZN(n4720) );
  AOI22D1BWP12T U1912 ( .A1(a[25]), .A2(n4699), .B1(b[8]), .B2(n5833), .ZN(
        n4700) );
  OAI22D1BWP12T U1913 ( .A1(n4703), .A2(n4702), .B1(n4701), .B2(n4700), .ZN(
        n4718) );
  FA1D0BWP12T U1914 ( .A(n4706), .B(n4705), .CI(n4704), .CO(n4716), .S(n5597)
         );
  FA1D0BWP12T U1915 ( .A(n4709), .B(n4708), .CI(n4707), .CO(n4714), .S(n4615)
         );
  FA1D0BWP12T U1916 ( .A(n4712), .B(n4711), .CI(n4710), .CO(n4713), .S(n4584)
         );
  MOAI22D0BWP12T U1917 ( .A1(n4714), .A2(n4713), .B1(n4714), .B2(n4713), .ZN(
        n4715) );
  MAOI22D0BWP12T U1918 ( .A1(n4716), .A2(n4715), .B1(n4716), .B2(n4715), .ZN(
        n4717) );
  MAOI22D0BWP12T U1919 ( .A1(n4718), .A2(n4717), .B1(n4718), .B2(n4717), .ZN(
        n4719) );
  MAOI22D0BWP12T U1920 ( .A1(n4720), .A2(n4719), .B1(n4720), .B2(n4719), .ZN(
        n4721) );
  MAOI22D0BWP12T U1921 ( .A1(n4722), .A2(n4721), .B1(n4722), .B2(n4721), .ZN(
        n4723) );
  MAOI22D0BWP12T U1922 ( .A1(n4724), .A2(n4723), .B1(n4724), .B2(n4723), .ZN(
        n4725) );
  MAOI22D0BWP12T U1923 ( .A1(n4726), .A2(n4725), .B1(n4726), .B2(n4725), .ZN(
        n4727) );
  MAOI22D0BWP12T U1924 ( .A1(n4728), .A2(n4727), .B1(n4728), .B2(n4727), .ZN(
        n4729) );
  MAOI22D0BWP12T U1925 ( .A1(n4730), .A2(n4729), .B1(n4730), .B2(n4729), .ZN(
        n4731) );
  MAOI22D0BWP12T U1926 ( .A1(n4732), .A2(n4731), .B1(n4732), .B2(n4731), .ZN(
        n4734) );
  ND2D1BWP12T U1927 ( .A1(n5374), .A2(n4734), .ZN(n5588) );
  INVD1BWP12T U1928 ( .I(n5597), .ZN(n4733) );
  OAI32D1BWP12T U1929 ( .A1(n5597), .A2(n4734), .A3(n6130), .B1(n5588), .B2(
        n4733), .ZN(n4735) );
  AO211D1BWP12T U1930 ( .A1(n5457), .A2(n5582), .B(n4736), .C(n4735), .Z(v) );
  NR2D1BWP12T U1931 ( .A1(n4737), .A2(a[30]), .ZN(n5475) );
  NR2D1BWP12T U1932 ( .A1(n4738), .A2(b[30]), .ZN(n5433) );
  NR2D1BWP12T U1933 ( .A1(n5475), .A2(n5433), .ZN(n6097) );
  INVD1BWP12T U1934 ( .I(n6097), .ZN(n4951) );
  NR2D1BWP12T U1935 ( .A1(n4841), .A2(a[29]), .ZN(n5474) );
  INVD1BWP12T U1936 ( .I(n5474), .ZN(n4901) );
  NR2D1BWP12T U1937 ( .A1(b[29]), .A2(n5901), .ZN(n5890) );
  NR2D1BWP12T U1938 ( .A1(n5474), .A2(n5890), .ZN(n5887) );
  ND2D1BWP12T U1939 ( .A1(n5722), .A2(a[28]), .ZN(n5721) );
  INVD1BWP12T U1940 ( .I(n5721), .ZN(n5432) );
  ND2D1BWP12T U1941 ( .A1(n5751), .A2(a[27]), .ZN(n5431) );
  ND2D1BWP12T U1942 ( .A1(n5784), .A2(a[26]), .ZN(n5430) );
  INVD1BWP12T U1943 ( .I(n5430), .ZN(n5773) );
  ND2D1BWP12T U1944 ( .A1(n4739), .A2(a[25]), .ZN(n5429) );
  INVD1BWP12T U1945 ( .I(n5429), .ZN(n5838) );
  ND2D1BWP12T U1946 ( .A1(b[25]), .A2(n5833), .ZN(n5840) );
  ND2D1BWP12T U1947 ( .A1(n5429), .A2(n5840), .ZN(n4847) );
  ND2D1BWP12T U1948 ( .A1(b[24]), .A2(n5912), .ZN(n5460) );
  ND2D1BWP12T U1949 ( .A1(n5918), .A2(a[24]), .ZN(n5916) );
  ND2D1BWP12T U1950 ( .A1(n5916), .A2(n5460), .ZN(n4800) );
  INVD1BWP12T U1951 ( .I(n4800), .ZN(n5917) );
  NR2D1BWP12T U1952 ( .A1(b[23]), .A2(n5951), .ZN(n5943) );
  ND2D1BWP12T U1953 ( .A1(n4839), .A2(a[22]), .ZN(n5435) );
  INVD1BWP12T U1954 ( .I(n5435), .ZN(n6132) );
  NR2D1BWP12T U1955 ( .A1(n4839), .A2(a[22]), .ZN(n6134) );
  NR2D1BWP12T U1956 ( .A1(n6132), .A2(n6134), .ZN(n4851) );
  INVD1BWP12T U1957 ( .I(n4851), .ZN(n4908) );
  ND2D1BWP12T U1958 ( .A1(b[21]), .A2(n5964), .ZN(n5965) );
  ND2D1BWP12T U1959 ( .A1(n4740), .A2(a[21]), .ZN(n5961) );
  ND2D1BWP12T U1960 ( .A1(n5965), .A2(n5961), .ZN(n4895) );
  INVD1BWP12T U1961 ( .I(n4895), .ZN(n4939) );
  NR2D1BWP12T U1962 ( .A1(b[20]), .A2(n6082), .ZN(n5437) );
  NR2D1BWP12T U1963 ( .A1(b[19]), .A2(n5988), .ZN(n5994) );
  NR2D1BWP12T U1964 ( .A1(n6010), .A2(a[18]), .ZN(n6012) );
  NR2D1BWP12T U1965 ( .A1(b[18]), .A2(n6024), .ZN(n6017) );
  NR2D1BWP12T U1966 ( .A1(n6012), .A2(n6017), .ZN(n4941) );
  ND2D1BWP12T U1967 ( .A1(b[17]), .A2(n5679), .ZN(n5469) );
  ND2D1BWP12T U1968 ( .A1(n4838), .A2(a[17]), .ZN(n5434) );
  ND2D1BWP12T U1969 ( .A1(n5469), .A2(n5434), .ZN(n4912) );
  INVD1BWP12T U1970 ( .I(n4912), .ZN(n4857) );
  NR2D1BWP12T U1971 ( .A1(b[16]), .A2(n5710), .ZN(n5696) );
  NR2D1BWP12T U1972 ( .A1(n4793), .A2(a[16]), .ZN(n5692) );
  NR2D1BWP12T U1973 ( .A1(n5696), .A2(n5692), .ZN(n4932) );
  INVD1BWP12T U1974 ( .I(n4932), .ZN(n4891) );
  OAI21D1BWP12T U1975 ( .A1(a[11]), .A2(n4741), .B(n4744), .ZN(n5461) );
  ND2D1BWP12T U1976 ( .A1(n4743), .A2(n4742), .ZN(n5443) );
  ND2D1BWP12T U1977 ( .A1(n4744), .A2(n5443), .ZN(n4888) );
  OA21D1BWP12T U1978 ( .A1(n4745), .A2(n5461), .B(n4888), .Z(n4769) );
  MAOI222D1BWP12T U1979 ( .A(n5872), .B(b[13]), .C(n4769), .ZN(n4757) );
  ND2D1BWP12T U1980 ( .A1(a[14]), .A2(n5390), .ZN(n4778) );
  NR2D1BWP12T U1981 ( .A1(n5390), .A2(a[14]), .ZN(n5478) );
  INR2D1BWP12T U1982 ( .A1(n4778), .B1(n5478), .ZN(n5858) );
  ND2D1BWP12T U1983 ( .A1(n4757), .A2(n5858), .ZN(n4777) );
  ND2D1BWP12T U1984 ( .A1(a[15]), .A2(n4890), .ZN(n6047) );
  ND2D1BWP12T U1985 ( .A1(n4778), .A2(n6047), .ZN(n5441) );
  INVD1BWP12T U1986 ( .I(n5441), .ZN(n4746) );
  NR2D1BWP12T U1987 ( .A1(n4890), .A2(a[15]), .ZN(n6044) );
  AO21D1BWP12T U1988 ( .A1(n4777), .A2(n4746), .B(n6044), .Z(n4776) );
  NR2D1BWP12T U1989 ( .A1(n5989), .A2(a[19]), .ZN(n5468) );
  NR2D1BWP12T U1990 ( .A1(n5994), .A2(n5468), .ZN(n4893) );
  NR2D1BWP12T U1991 ( .A1(n6067), .A2(a[20]), .ZN(n6068) );
  NR2D1BWP12T U1992 ( .A1(n5437), .A2(n6068), .ZN(n4937) );
  INVD1BWP12T U1993 ( .I(n4937), .ZN(n4894) );
  NR2D1BWP12T U1994 ( .A1(n5940), .A2(a[23]), .ZN(n5473) );
  NR2D1BWP12T U1995 ( .A1(n5943), .A2(n5473), .ZN(n4896) );
  INVD1BWP12T U1996 ( .I(n4896), .ZN(n4946) );
  NR2D1BWP12T U1997 ( .A1(n5784), .A2(a[26]), .ZN(n5463) );
  NR2D1BWP12T U1998 ( .A1(n5773), .A2(n5463), .ZN(n4897) );
  INVD1BWP12T U1999 ( .I(n4897), .ZN(n5772) );
  ND2D1BWP12T U2000 ( .A1(b[27]), .A2(n5758), .ZN(n4747) );
  ND2D1BWP12T U2001 ( .A1(n5431), .A2(n4747), .ZN(n5752) );
  ND2D1BWP12T U2002 ( .A1(b[28]), .A2(n5737), .ZN(n5464) );
  ND2D1BWP12T U2003 ( .A1(n5721), .A2(n5464), .ZN(n5727) );
  MAOI22D0BWP12T U2004 ( .A1(n4951), .A2(n4749), .B1(n4951), .B2(n4749), .ZN(
        n6123) );
  INVD1BWP12T U2005 ( .I(n5887), .ZN(n4903) );
  MAOI22D0BWP12T U2006 ( .A1(n4903), .A2(n4748), .B1(n4903), .B2(n4748), .ZN(
        n5907) );
  INVD1BWP12T U2007 ( .I(n5457), .ZN(n5596) );
  MAOI22D0BWP12T U2008 ( .A1(n5596), .A2(n5579), .B1(n5596), .B2(n5579), .ZN(
        n5619) );
  MAOI22D0BWP12T U2009 ( .A1(n5752), .A2(n4750), .B1(n5752), .B2(n4750), .ZN(
        n5765) );
  MAOI22D0BWP12T U2010 ( .A1(n4946), .A2(n4751), .B1(n4946), .B2(n4751), .ZN(
        n5960) );
  MAOI22D0BWP12T U2011 ( .A1(n4800), .A2(n4752), .B1(n4800), .B2(n4752), .ZN(
        n5932) );
  MAOI22D0BWP12T U2012 ( .A1(n4893), .A2(n4753), .B1(n4893), .B2(n4753), .ZN(
        n6004) );
  INVD1BWP12T U2013 ( .I(n4941), .ZN(n4892) );
  MAOI22D0BWP12T U2014 ( .A1(n4892), .A2(n4754), .B1(n4892), .B2(n4754), .ZN(
        n6033) );
  MAOI22D0BWP12T U2015 ( .A1(n4895), .A2(n4755), .B1(n4895), .B2(n4755), .ZN(
        n5980) );
  MAOI22D0BWP12T U2016 ( .A1(n4857), .A2(n4756), .B1(n4857), .B2(n4756), .ZN(
        n5690) );
  MAOI22D0BWP12T U2017 ( .A1(n4757), .A2(n5858), .B1(n4757), .B2(n5858), .ZN(
        n5881) );
  MAOI22D0BWP12T U2018 ( .A1(n5798), .A2(n4758), .B1(n5798), .B2(n4758), .ZN(
        n5813) );
  INVD1BWP12T U2019 ( .I(n5799), .ZN(n5796) );
  ND2D1BWP12T U2020 ( .A1(n5796), .A2(n5436), .ZN(n5573) );
  INVD1BWP12T U2021 ( .I(n5573), .ZN(n5624) );
  AOI22D0BWP12T U2022 ( .A1(n5624), .A2(c_in), .B1(n5573), .B2(n4759), .ZN(
        n5627) );
  NR4D0BWP12T U2023 ( .A1(n4760), .A2(n5813), .A3(n5627), .A4(n6167), .ZN(
        n4764) );
  ND4D1BWP12T U2024 ( .A1(n4764), .A2(n4763), .A3(n4762), .A4(n4761), .ZN(
        n4765) );
  NR4D0BWP12T U2025 ( .A1(n4768), .A2(n4767), .A3(n4766), .A4(n4765), .ZN(
        n4772) );
  MAOI22D0BWP12T U2026 ( .A1(n4769), .A2(n4917), .B1(n4769), .B2(n4917), .ZN(
        n5659) );
  ND4D1BWP12T U2027 ( .A1(n4772), .A2(n5659), .A3(n4771), .A4(n4770), .ZN(
        n4773) );
  NR4D0BWP12T U2028 ( .A1(n5881), .A2(n4775), .A3(n4774), .A4(n4773), .ZN(
        n4780) );
  MAOI22D0BWP12T U2029 ( .A1(n4932), .A2(n4776), .B1(n4932), .B2(n4776), .ZN(
        n5720) );
  ND2D1BWP12T U2030 ( .A1(n4778), .A2(n4777), .ZN(n4779) );
  MAOI22D0BWP12T U2031 ( .A1(n4914), .A2(n4779), .B1(n4914), .B2(n4779), .ZN(
        n6064) );
  ND4D1BWP12T U2032 ( .A1(n5690), .A2(n4780), .A3(n5720), .A4(n6064), .ZN(
        n4781) );
  NR4D0BWP12T U2033 ( .A1(n6004), .A2(n6033), .A3(n5980), .A4(n4781), .ZN(
        n4785) );
  INVD1BWP12T U2034 ( .I(n4847), .ZN(n4906) );
  MAOI22D0BWP12T U2035 ( .A1(n4782), .A2(n4906), .B1(n4782), .B2(n4906), .ZN(
        n5856) );
  MOAI22D0BWP12T U2036 ( .A1(n4908), .A2(n4783), .B1(n4908), .B2(n4783), .ZN(
        n6168) );
  MAOI22D0BWP12T U2037 ( .A1(n4937), .A2(n4784), .B1(n4937), .B2(n4784), .ZN(
        n6087) );
  ND4D1BWP12T U2038 ( .A1(n4785), .A2(n5856), .A3(n6168), .A4(n6087), .ZN(
        n4786) );
  NR4D0BWP12T U2039 ( .A1(n5765), .A2(n5960), .A3(n5932), .A4(n4786), .ZN(
        n4789) );
  MOAI22D0BWP12T U2040 ( .A1(n5772), .A2(n4787), .B1(n5772), .B2(n4787), .ZN(
        n5791) );
  INVD1BWP12T U2041 ( .I(n5727), .ZN(n4899) );
  MAOI22D0BWP12T U2042 ( .A1(n4899), .A2(n4788), .B1(n4899), .B2(n4788), .ZN(
        n5742) );
  ND4D1BWP12T U2043 ( .A1(n5619), .A2(n4789), .A3(n5791), .A4(n5742), .ZN(
        n5578) );
  NR2D1BWP12T U2044 ( .A1(b[28]), .A2(a[28]), .ZN(n4840) );
  NR2D1BWP12T U2045 ( .A1(b[20]), .A2(a[20]), .ZN(n6075) );
  ND2D1BWP12T U2046 ( .A1(b[17]), .A2(a[17]), .ZN(n5673) );
  INVD1BWP12T U2047 ( .I(n5673), .ZN(n5674) );
  INVD1BWP12T U2048 ( .I(n5392), .ZN(n6046) );
  MAOI222D1BWP12T U2049 ( .A(n4792), .B(n4791), .C(n4790), .ZN(n4809) );
  MAOI222D1BWP12T U2050 ( .A(b[14]), .B(a[14]), .C(n4808), .ZN(n4806) );
  MAOI222D1BWP12T U2051 ( .A(n4824), .B(n5710), .C(n4793), .ZN(n4807) );
  OAI22D1BWP12T U2052 ( .A1(b[17]), .A2(a[17]), .B1(n5674), .B2(n4807), .ZN(
        n4804) );
  MAOI222D1BWP12T U2053 ( .A(n6010), .B(n6024), .C(n4804), .ZN(n4805) );
  MAOI222D1BWP12T U2054 ( .A(b[19]), .B(a[19]), .C(n4805), .ZN(n4801) );
  NR2D1BWP12T U2055 ( .A1(n6075), .A2(n4801), .ZN(n4828) );
  ND2D1BWP12T U2056 ( .A1(b[21]), .A2(a[21]), .ZN(n5962) );
  ND2D1BWP12T U2057 ( .A1(b[20]), .A2(a[20]), .ZN(n6066) );
  ND2D1BWP12T U2058 ( .A1(n5962), .A2(n6066), .ZN(n5396) );
  OAI22D1BWP12T U2059 ( .A1(b[21]), .A2(a[21]), .B1(n4828), .B2(n5396), .ZN(
        n4802) );
  MAOI222D1BWP12T U2060 ( .A(n4839), .B(n6155), .C(n4802), .ZN(n4798) );
  MAOI222D1BWP12T U2061 ( .A(b[23]), .B(a[23]), .C(n4798), .ZN(n4799) );
  MAOI222D1BWP12T U2062 ( .A(n5918), .B(n5912), .C(n4799), .ZN(n4803) );
  MAOI222D1BWP12T U2063 ( .A(b[25]), .B(a[25]), .C(n4803), .ZN(n4795) );
  MAOI222D1BWP12T U2064 ( .A(n5784), .B(n5787), .C(n4795), .ZN(n4794) );
  MAOI222D1BWP12T U2065 ( .A(a[27]), .B(b[27]), .C(n4794), .ZN(n4797) );
  OR2XD1BWP12T U2066 ( .A1(n4840), .A2(n4797), .Z(n4834) );
  ND2D1BWP12T U2067 ( .A1(b[28]), .A2(a[28]), .ZN(n4842) );
  OA21D1BWP12T U2068 ( .A1(n5901), .A2(n4841), .B(n4842), .Z(n5389) );
  AOI22D1BWP12T U2069 ( .A1(n4841), .A2(n5901), .B1(n4834), .B2(n5389), .ZN(
        n4796) );
  MAOI22D0BWP12T U2070 ( .A1(n6097), .A2(n4796), .B1(n6097), .B2(n4796), .ZN(
        n6121) );
  MAOI22D0BWP12T U2071 ( .A1(n5752), .A2(n4794), .B1(n5752), .B2(n4794), .ZN(
        n5764) );
  MAOI22D0BWP12T U2072 ( .A1(n4897), .A2(n4795), .B1(n4897), .B2(n4795), .ZN(
        n5795) );
  MAOI222D1BWP12T U2073 ( .A(b[30]), .B(a[30]), .C(n4796), .ZN(n5586) );
  MAOI22D0BWP12T U2074 ( .A1(n5596), .A2(n5586), .B1(n5596), .B2(n5586), .ZN(
        n5615) );
  MAOI22D0BWP12T U2075 ( .A1(n5727), .A2(n4797), .B1(n5727), .B2(n4797), .ZN(
        n5746) );
  MAOI22D0BWP12T U2076 ( .A1(n4896), .A2(n4798), .B1(n4896), .B2(n4798), .ZN(
        n5957) );
  MAOI22D0BWP12T U2077 ( .A1(n4800), .A2(n4799), .B1(n4800), .B2(n4799), .ZN(
        n5935) );
  MAOI22D0BWP12T U2078 ( .A1(n4937), .A2(n4801), .B1(n4937), .B2(n4801), .ZN(
        n6091) );
  MAOI22D0BWP12T U2079 ( .A1(n4851), .A2(n4802), .B1(n4851), .B2(n4802), .ZN(
        n6163) );
  MAOI22D0BWP12T U2080 ( .A1(n4847), .A2(n4803), .B1(n4847), .B2(n4803), .ZN(
        n5852) );
  MAOI22D0BWP12T U2081 ( .A1(n4892), .A2(n4804), .B1(n4892), .B2(n4804), .ZN(
        n6030) );
  MAOI22D0BWP12T U2082 ( .A1(n4893), .A2(n4805), .B1(n4893), .B2(n4805), .ZN(
        n6007) );
  MOAI22D0BWP12T U2083 ( .A1(n4914), .A2(n4806), .B1(n4914), .B2(n4806), .ZN(
        n6061) );
  MAOI22D0BWP12T U2084 ( .A1(n4912), .A2(n4807), .B1(n4912), .B2(n4807), .ZN(
        n5687) );
  INVD1BWP12T U2085 ( .I(n4917), .ZN(n4837) );
  MOAI22D0BWP12T U2086 ( .A1(n4837), .A2(n4809), .B1(n4837), .B2(n4809), .ZN(
        n5660) );
  MOAI22D0BWP12T U2087 ( .A1(n4810), .A2(n5798), .B1(n4810), .B2(n5798), .ZN(
        n5803) );
  ND4D1BWP12T U2088 ( .A1(n5627), .A2(n6164), .A3(n4811), .A4(n5803), .ZN(
        n4812) );
  NR4D0BWP12T U2089 ( .A1(n4815), .A2(n4814), .A3(n4813), .A4(n4812), .ZN(
        n4818) );
  ND4D1BWP12T U2090 ( .A1(n4819), .A2(n4818), .A3(n4817), .A4(n4816), .ZN(
        n4820) );
  NR4D0BWP12T U2091 ( .A1(n4823), .A2(n4822), .A3(n4821), .A4(n4820), .ZN(
        n4825) );
  MOAI22D0BWP12T U2092 ( .A1(n4932), .A2(n4824), .B1(n4932), .B2(n4824), .ZN(
        n5714) );
  ND4D1BWP12T U2093 ( .A1(n4826), .A2(n5660), .A3(n4825), .A4(n5714), .ZN(
        n4827) );
  NR4D0BWP12T U2094 ( .A1(n6061), .A2(n5687), .A3(n5880), .A4(n4827), .ZN(
        n4830) );
  IND2D1BWP12T U2095 ( .A1(n4828), .B1(n6066), .ZN(n4829) );
  MAOI22D0BWP12T U2096 ( .A1(n4939), .A2(n4829), .B1(n4939), .B2(n4829), .ZN(
        n5979) );
  ND4D1BWP12T U2097 ( .A1(n6030), .A2(n6007), .A3(n4830), .A4(n5979), .ZN(
        n4831) );
  NR4D0BWP12T U2098 ( .A1(n6091), .A2(n6163), .A3(n5852), .A4(n4831), .ZN(
        n4832) );
  ND4D1BWP12T U2099 ( .A1(n5746), .A2(n5957), .A3(n5935), .A4(n4832), .ZN(
        n4833) );
  NR4D0BWP12T U2100 ( .A1(n5764), .A2(n5795), .A3(n5615), .A4(n4833), .ZN(
        n5576) );
  ND2D1BWP12T U2101 ( .A1(n4842), .A2(n4834), .ZN(n4835) );
  MAOI22D0BWP12T U2102 ( .A1(n5887), .A2(n4835), .B1(n5887), .B2(n4835), .ZN(
        n5911) );
  MAOI222D1BWP12T U2103 ( .A(b[12]), .B(a[12]), .C(n4836), .ZN(n4862) );
  MAOI222D1BWP12T U2104 ( .A(b[14]), .B(a[14]), .C(n4860), .ZN(n4859) );
  AOI22D1BWP12T U2105 ( .A1(n5392), .A2(n4859), .B1(n4890), .B2(n6042), .ZN(
        n4861) );
  MAOI222D1BWP12T U2106 ( .A(b[16]), .B(a[16]), .C(n4861), .ZN(n4856) );
  AOI22D1BWP12T U2107 ( .A1(n4838), .A2(n5679), .B1(n5673), .B2(n4856), .ZN(
        n4854) );
  MAOI222D1BWP12T U2108 ( .A(b[18]), .B(a[18]), .C(n4854), .ZN(n4855) );
  MAOI222D1BWP12T U2109 ( .A(n5989), .B(n5988), .C(n4855), .ZN(n4852) );
  INVD1BWP12T U2110 ( .I(n4852), .ZN(n4853) );
  NR2D1BWP12T U2111 ( .A1(n6075), .A2(n4853), .ZN(n4879) );
  OAI22D1BWP12T U2112 ( .A1(b[21]), .A2(a[21]), .B1(n4879), .B2(n5396), .ZN(
        n4850) );
  MAOI222D1BWP12T U2113 ( .A(n4839), .B(n6155), .C(n4850), .ZN(n4885) );
  MAOI222D1BWP12T U2114 ( .A(a[23]), .B(b[23]), .C(n4885), .ZN(n4849) );
  MAOI222D1BWP12T U2115 ( .A(n5918), .B(n5912), .C(n4849), .ZN(n4848) );
  MAOI222D1BWP12T U2116 ( .A(b[25]), .B(a[25]), .C(n4848), .ZN(n4884) );
  MAOI222D1BWP12T U2117 ( .A(n4884), .B(n5784), .C(n5787), .ZN(n4883) );
  MAOI222D1BWP12T U2118 ( .A(b[27]), .B(a[27]), .C(n4883), .ZN(n4846) );
  OR2XD1BWP12T U2119 ( .A1(n4840), .A2(n4846), .Z(n4843) );
  AOI22D1BWP12T U2120 ( .A1(n4843), .A2(n5389), .B1(n4841), .B2(n5901), .ZN(
        n4845) );
  MAOI22D0BWP12T U2121 ( .A1(n6097), .A2(n4845), .B1(n6097), .B2(n4845), .ZN(
        n6127) );
  ND2D1BWP12T U2122 ( .A1(n4843), .A2(n4842), .ZN(n4844) );
  MAOI22D0BWP12T U2123 ( .A1(n4903), .A2(n4844), .B1(n4903), .B2(n4844), .ZN(
        n5908) );
  MAOI222D1BWP12T U2124 ( .A(b[30]), .B(a[30]), .C(n4845), .ZN(n5583) );
  MAOI22D0BWP12T U2125 ( .A1(n5596), .A2(n5583), .B1(n5596), .B2(n5583), .ZN(
        n5616) );
  MAOI22D0BWP12T U2126 ( .A1(n4846), .A2(n4899), .B1(n4846), .B2(n4899), .ZN(
        n5743) );
  MAOI22D0BWP12T U2127 ( .A1(n4848), .A2(n4847), .B1(n4848), .B2(n4847), .ZN(
        n5853) );
  MAOI22D0BWP12T U2128 ( .A1(n5917), .A2(n4849), .B1(n5917), .B2(n4849), .ZN(
        n5931) );
  MAOI22D0BWP12T U2129 ( .A1(n4851), .A2(n4850), .B1(n4851), .B2(n4850), .ZN(
        n6161) );
  AOI22D1BWP12T U2130 ( .A1(n4853), .A2(n4894), .B1(n4852), .B2(n4937), .ZN(
        n6088) );
  MAOI22D0BWP12T U2131 ( .A1(n4854), .A2(n4941), .B1(n4854), .B2(n4941), .ZN(
        n6029) );
  MAOI22D0BWP12T U2132 ( .A1(n4893), .A2(n4855), .B1(n4893), .B2(n4855), .ZN(
        n6003) );
  MAOI22D0BWP12T U2133 ( .A1(n4857), .A2(n4856), .B1(n4857), .B2(n4856), .ZN(
        n5686) );
  MAOI22D0BWP12T U2134 ( .A1(n4859), .A2(n4858), .B1(n4859), .B2(n4858), .ZN(
        n6060) );
  MAOI22D0BWP12T U2135 ( .A1(n4860), .A2(n5858), .B1(n4860), .B2(n5858), .ZN(
        n5884) );
  MAOI22D0BWP12T U2136 ( .A1(n4861), .A2(n4932), .B1(n4861), .B2(n4932), .ZN(
        n5715) );
  MAOI22D0BWP12T U2137 ( .A1(n4862), .A2(n4917), .B1(n4862), .B2(n4917), .ZN(
        n5663) );
  OAI22D1BWP12T U2138 ( .A1(n5798), .A2(n5634), .B1(n5797), .B2(n5492), .ZN(
        n5801) );
  ND4D1BWP12T U2139 ( .A1(n6162), .A2(n4864), .A3(n4863), .A4(n5801), .ZN(
        n4865) );
  NR4D0BWP12T U2140 ( .A1(n4868), .A2(n4867), .A3(n4866), .A4(n4865), .ZN(
        n4870) );
  ND4D1BWP12T U2141 ( .A1(n4872), .A2(n4871), .A3(n4870), .A4(n4869), .ZN(
        n4873) );
  NR4D0BWP12T U2142 ( .A1(n5663), .A2(n4875), .A3(n4874), .A4(n4873), .ZN(
        n4877) );
  ND4D1BWP12T U2143 ( .A1(n5884), .A2(n5715), .A3(n4877), .A4(n4876), .ZN(
        n4878) );
  NR4D0BWP12T U2144 ( .A1(n6003), .A2(n5686), .A3(n6060), .A4(n4878), .ZN(
        n4881) );
  IND2D1BWP12T U2145 ( .A1(n4879), .B1(n6066), .ZN(n4880) );
  MAOI22D0BWP12T U2146 ( .A1(n4939), .A2(n4880), .B1(n4939), .B2(n4880), .ZN(
        n5983) );
  ND4D1BWP12T U2147 ( .A1(n6088), .A2(n6029), .A3(n4881), .A4(n5983), .ZN(
        n4882) );
  NR4D0BWP12T U2148 ( .A1(n5853), .A2(n5931), .A3(n6161), .A4(n4882), .ZN(
        n4886) );
  INVD1BWP12T U2149 ( .I(n5752), .ZN(n4898) );
  MAOI22D0BWP12T U2150 ( .A1(n4883), .A2(n4898), .B1(n4883), .B2(n4898), .ZN(
        n5768) );
  MOAI22D0BWP12T U2151 ( .A1(n4884), .A2(n4897), .B1(n4884), .B2(n4897), .ZN(
        n5792) );
  MAOI22D0BWP12T U2152 ( .A1(n4885), .A2(n4896), .B1(n4885), .B2(n4896), .ZN(
        n5956) );
  ND4D1BWP12T U2153 ( .A1(n4886), .A2(n5768), .A3(n5792), .A4(n5956), .ZN(
        n4887) );
  NR4D0BWP12T U2154 ( .A1(n5908), .A2(n5616), .A3(n5743), .A4(n4887), .ZN(
        n4953) );
  OAI21D1BWP12T U2155 ( .A1(n5461), .A2(n4889), .B(n4888), .ZN(n4916) );
  MAOI222D1BWP12T U2156 ( .A(n5476), .B(n4916), .C(a[13]), .ZN(n4915) );
  MAOI222D1BWP12T U2157 ( .A(a[15]), .B(n4913), .C(n4890), .ZN(n4931) );
  INVD1BWP12T U2158 ( .I(n4893), .ZN(n4910) );
  AOI21D1BWP12T U2159 ( .A1(n4907), .A2(n5435), .B(n6134), .ZN(n4947) );
  MAOI22D0BWP12T U2160 ( .A1(n4899), .A2(n4900), .B1(n4899), .B2(n4900), .ZN(
        n5741) );
  MAOI22D0BWP12T U2161 ( .A1(n5580), .A2(n5457), .B1(n5580), .B2(n5457), .ZN(
        n5614) );
  MAOI22D0BWP12T U2162 ( .A1(n4903), .A2(n4902), .B1(n4903), .B2(n4902), .ZN(
        n5906) );
  MAOI22D0BWP12T U2163 ( .A1(n5917), .A2(n4904), .B1(n5917), .B2(n4904), .ZN(
        n5928) );
  MAOI22D0BWP12T U2164 ( .A1(n4906), .A2(n4905), .B1(n4906), .B2(n4905), .ZN(
        n5851) );
  MAOI22D0BWP12T U2165 ( .A1(n4908), .A2(n4907), .B1(n4908), .B2(n4907), .ZN(
        n6159) );
  MAOI22D0BWP12T U2166 ( .A1(n4910), .A2(n4909), .B1(n4910), .B2(n4909), .ZN(
        n6002) );
  MAOI22D0BWP12T U2167 ( .A1(n4912), .A2(n4911), .B1(n4912), .B2(n4911), .ZN(
        n5685) );
  MOAI22D0BWP12T U2168 ( .A1(n4914), .A2(n4913), .B1(n4914), .B2(n4913), .ZN(
        n6059) );
  MAOI22D0BWP12T U2169 ( .A1(n5858), .A2(n4915), .B1(n5858), .B2(n4915), .ZN(
        n5879) );
  MOAI22D0BWP12T U2170 ( .A1(n4917), .A2(n4916), .B1(n4917), .B2(n4916), .ZN(
        n5658) );
  ND4D1BWP12T U2171 ( .A1(n4919), .A2(n4918), .A3(n6160), .A4(n5798), .ZN(
        n4920) );
  NR4D0BWP12T U2172 ( .A1(n4923), .A2(n4922), .A3(n4921), .A4(n4920), .ZN(
        n4925) );
  ND4D1BWP12T U2173 ( .A1(n4927), .A2(n4926), .A3(n4925), .A4(n4924), .ZN(
        n4928) );
  INR4D0BWP12T U2174 ( .A1(n5658), .B1(n4930), .B2(n4929), .B3(n4928), .ZN(
        n4934) );
  MAOI22D0BWP12T U2175 ( .A1(n4932), .A2(n4931), .B1(n4932), .B2(n4931), .ZN(
        n5713) );
  ND4D1BWP12T U2176 ( .A1(n5879), .A2(n4934), .A3(n5713), .A4(n4933), .ZN(
        n4935) );
  NR4D0BWP12T U2177 ( .A1(n6002), .A2(n5685), .A3(n6059), .A4(n4935), .ZN(
        n4942) );
  MAOI22D0BWP12T U2178 ( .A1(n4937), .A2(n4936), .B1(n4937), .B2(n4936), .ZN(
        n6086) );
  MAOI22D0BWP12T U2179 ( .A1(n4939), .A2(n4938), .B1(n4939), .B2(n4938), .ZN(
        n5975) );
  MAOI22D0BWP12T U2180 ( .A1(n4941), .A2(n4940), .B1(n4941), .B2(n4940), .ZN(
        n6028) );
  ND4D1BWP12T U2181 ( .A1(n4942), .A2(n6086), .A3(n5975), .A4(n6028), .ZN(
        n4943) );
  NR4D0BWP12T U2182 ( .A1(n5928), .A2(n5851), .A3(n6159), .A4(n4943), .ZN(
        n4948) );
  MAOI22D0BWP12T U2183 ( .A1(n5752), .A2(n4944), .B1(n5752), .B2(n4944), .ZN(
        n5747) );
  MAOI22D0BWP12T U2184 ( .A1(n5772), .A2(n4945), .B1(n5772), .B2(n4945), .ZN(
        n5790) );
  MAOI22D0BWP12T U2185 ( .A1(n4947), .A2(n4946), .B1(n4947), .B2(n4946), .ZN(
        n5955) );
  ND4D1BWP12T U2186 ( .A1(n4948), .A2(n5747), .A3(n5790), .A4(n5955), .ZN(
        n4949) );
  NR4D0BWP12T U2187 ( .A1(n5741), .A2(n5614), .A3(n5906), .A4(n4949), .ZN(
        n4952) );
  MOAI22D0BWP12T U2188 ( .A1(n4951), .A2(n4950), .B1(n4951), .B2(n4950), .ZN(
        n6114) );
  AOI22D1BWP12T U2189 ( .A1(n6127), .A2(n4953), .B1(n4952), .B2(n6114), .ZN(
        n5574) );
  INVD1BWP12T U2190 ( .I(n5018), .ZN(n5287) );
  NR2D1BWP12T U2191 ( .A1(b[3]), .A2(n5703), .ZN(n5056) );
  AOI22D1BWP12T U2192 ( .A1(n5095), .A2(n5250), .B1(n5051), .B2(n5177), .ZN(
        n4955) );
  AOI22D1BWP12T U2193 ( .A1(n5057), .A2(n5249), .B1(n5178), .B2(n5052), .ZN(
        n4954) );
  ND2D1BWP12T U2194 ( .A1(n4955), .A2(n4954), .ZN(n5034) );
  AOI22D1BWP12T U2195 ( .A1(b[0]), .A2(a[16]), .B1(a[17]), .B2(n5379), .ZN(
        n5248) );
  NR2D1BWP12T U2196 ( .A1(n5150), .A2(n5128), .ZN(n4959) );
  ND2D1BWP12T U2197 ( .A1(n4957), .A2(n4956), .ZN(n5261) );
  OAI22D1BWP12T U2198 ( .A1(n4974), .A2(n5045), .B1(n5131), .B2(n5261), .ZN(
        n4958) );
  AOI211D1BWP12T U2199 ( .A1(n5052), .A2(n5248), .B(n4959), .C(n4958), .ZN(
        n5033) );
  INVD1BWP12T U2200 ( .I(n5079), .ZN(n5054) );
  INVD1BWP12T U2201 ( .I(n4960), .ZN(n5289) );
  INVD1BWP12T U2202 ( .I(n5770), .ZN(n5081) );
  NR2D1BWP12T U2203 ( .A1(n5379), .A2(n5131), .ZN(n5097) );
  INVD1BWP12T U2204 ( .I(n5097), .ZN(n4984) );
  AOI22D1BWP12T U2205 ( .A1(n5095), .A2(n5289), .B1(n5287), .B2(n5051), .ZN(
        n4962) );
  ND2D1BWP12T U2206 ( .A1(n5283), .A2(n5052), .ZN(n4961) );
  OAI211D1BWP12T U2207 ( .A1(a[30]), .A2(n4984), .B(n4962), .C(n4961), .ZN(
        n4965) );
  AOI22D1BWP12T U2208 ( .A1(n5178), .A2(n5051), .B1(n5052), .B2(n5250), .ZN(
        n4964) );
  AOI22D1BWP12T U2209 ( .A1(n5181), .A2(n5057), .B1(n5095), .B2(n5249), .ZN(
        n4963) );
  ND2D1BWP12T U2210 ( .A1(n4964), .A2(n4963), .ZN(n5038) );
  AOI22D1BWP12T U2211 ( .A1(n5770), .A2(n4965), .B1(n5056), .B2(n5038), .ZN(
        n4969) );
  AOI22D1BWP12T U2212 ( .A1(n5057), .A2(n5285), .B1(n5051), .B2(n5248), .ZN(
        n4967) );
  ND2D1BWP12T U2213 ( .A1(n5256), .A2(n5052), .ZN(n4966) );
  OAI211D1BWP12T U2214 ( .A1(n5261), .A2(n5128), .B(n4967), .C(n4966), .ZN(
        n5037) );
  NR2D1BWP12T U2215 ( .A1(n5632), .A2(b[4]), .ZN(n5268) );
  INVD1BWP12T U2216 ( .I(n5268), .ZN(n5165) );
  NR2D1BWP12T U2217 ( .A1(a[31]), .A2(n5165), .ZN(n5569) );
  AOI211D1BWP12T U2218 ( .A1(n5079), .A2(n5037), .B(n5569), .C(n5528), .ZN(
        n4968) );
  OAI211D1BWP12T U2219 ( .A1(n5024), .A2(n4995), .B(n4969), .C(n4968), .ZN(
        n5601) );
  AOI22D1BWP12T U2220 ( .A1(b[0]), .A2(a[21]), .B1(a[22]), .B2(n5379), .ZN(
        n5228) );
  INVD1BWP12T U2221 ( .I(n5208), .ZN(n5046) );
  NR2D1BWP12T U2222 ( .A1(n5046), .A2(n5047), .ZN(n4973) );
  NR2D1BWP12T U2223 ( .A1(n4971), .A2(n4970), .ZN(n4987) );
  MOAI22D0BWP12T U2224 ( .A1(n4987), .A2(n5131), .B1(n5188), .B2(n5095), .ZN(
        n4972) );
  AOI211D1BWP12T U2225 ( .A1(n5051), .A2(n5159), .B(n4973), .C(n4972), .ZN(
        n4996) );
  AOI22D1BWP12T U2226 ( .A1(b[0]), .A2(a[27]), .B1(a[28]), .B2(n5379), .ZN(
        n5231) );
  AOI22D1BWP12T U2227 ( .A1(b[0]), .A2(a[23]), .B1(a[24]), .B2(n5379), .ZN(
        n5230) );
  NR2D1BWP12T U2228 ( .A1(n4974), .A2(n5047), .ZN(n4976) );
  MOAI22D0BWP12T U2229 ( .A1(n5150), .A2(n5131), .B1(n5051), .B2(n5249), .ZN(
        n4975) );
  AOI211D1BWP12T U2230 ( .A1(n5248), .A2(n5095), .B(n4976), .C(n4975), .ZN(
        n5029) );
  AOI22D1BWP12T U2231 ( .A1(n5095), .A2(n5287), .B1(n5052), .B2(n5285), .ZN(
        n4978) );
  ND2D1BWP12T U2232 ( .A1(n5057), .A2(n5283), .ZN(n4977) );
  OAI211D1BWP12T U2233 ( .A1(n5261), .A2(n5045), .B(n4978), .C(n4977), .ZN(
        n4979) );
  AOI22D1BWP12T U2234 ( .A1(b[4]), .A2(n4980), .B1(n5770), .B2(n4979), .ZN(
        n4981) );
  OAI211D1BWP12T U2235 ( .A1(n5029), .A2(n5054), .B(n5570), .C(n4981), .ZN(
        n5756) );
  ND4D1BWP12T U2236 ( .A1(n5898), .A2(n5601), .A3(n5732), .A4(n5756), .ZN(
        n5077) );
  MAOI22D0BWP12T U2237 ( .A1(n4982), .A2(n5036), .B1(n5070), .B2(n5034), .ZN(
        n5648) );
  MOAI22D0BWP12T U2238 ( .A1(a[30]), .A2(n4983), .B1(n5230), .B2(n5051), .ZN(
        n4986) );
  MOAI22D0BWP12T U2239 ( .A1(a[29]), .A2(n4984), .B1(n5229), .B2(n5052), .ZN(
        n4985) );
  AOI211D1BWP12T U2240 ( .A1(n5095), .A2(n5231), .B(n4986), .C(n4985), .ZN(
        n4994) );
  INVD1BWP12T U2241 ( .I(n4987), .ZN(n5207) );
  AOI22D1BWP12T U2242 ( .A1(n5057), .A2(n5228), .B1(n5095), .B2(n5207), .ZN(
        n4989) );
  AOI22D1BWP12T U2243 ( .A1(n5051), .A2(n5208), .B1(n5052), .B2(n5188), .ZN(
        n4988) );
  ND2D1BWP12T U2244 ( .A1(n4989), .A2(n4988), .ZN(n5006) );
  AOI21D1BWP12T U2245 ( .A1(n5079), .A2(n5006), .B(n5528), .ZN(n4993) );
  AOI22D1BWP12T U2246 ( .A1(n5057), .A2(n5159), .B1(n5095), .B2(n5158), .ZN(
        n4991) );
  AOI22D1BWP12T U2247 ( .A1(n5122), .A2(n5051), .B1(n5052), .B2(n5123), .ZN(
        n4990) );
  ND2D1BWP12T U2248 ( .A1(n4991), .A2(n4990), .ZN(n5069) );
  AOI22D1BWP12T U2249 ( .A1(n5145), .A2(n5067), .B1(n5056), .B2(n5069), .ZN(
        n4992) );
  OAI211D1BWP12T U2250 ( .A1(n4994), .A2(n5081), .B(n4993), .C(n4992), .ZN(
        n6103) );
  ND2D1BWP12T U2251 ( .A1(n4995), .A2(n5570), .ZN(n5065) );
  INVD1BWP12T U2252 ( .I(n5065), .ZN(n5041) );
  MAOI22D0BWP12T U2253 ( .A1(b[3]), .A2(n4997), .B1(n5081), .B2(n4996), .ZN(
        n4998) );
  OAI211D1BWP12T U2254 ( .A1(n5703), .A2(n5014), .B(n5041), .C(n4998), .ZN(
        n6070) );
  ND4D1BWP12T U2255 ( .A1(n5648), .A2(n4999), .A3(n6103), .A4(n6070), .ZN(
        n5076) );
  AOI22D1BWP12T U2256 ( .A1(n5095), .A2(n5230), .B1(n5052), .B2(n5228), .ZN(
        n5001) );
  AOI22D1BWP12T U2257 ( .A1(n5057), .A2(n5229), .B1(n5051), .B2(n5207), .ZN(
        n5000) );
  ND2D1BWP12T U2258 ( .A1(n5001), .A2(n5000), .ZN(n5004) );
  OAI22D1BWP12T U2259 ( .A1(n5159), .A2(n5047), .B1(n5045), .B2(n5158), .ZN(
        n5003) );
  OAI22D1BWP12T U2260 ( .A1(n5208), .A2(n5128), .B1(n5131), .B2(n5188), .ZN(
        n5002) );
  NR2D1BWP12T U2261 ( .A1(n5003), .A2(n5002), .ZN(n5025) );
  AOI22D1BWP12T U2262 ( .A1(n5770), .A2(n5004), .B1(n5079), .B2(n5025), .ZN(
        n5005) );
  OAI211D1BWP12T U2263 ( .A1(n5703), .A2(n5011), .B(n5570), .C(n5005), .ZN(
        n5780) );
  AOI22D1BWP12T U2264 ( .A1(b[3]), .A2(n5069), .B1(n5770), .B2(n5006), .ZN(
        n5007) );
  OAI211D1BWP12T U2265 ( .A1(n5008), .A2(n5703), .B(n5041), .C(n5007), .ZN(
        n6139) );
  ND4D1BWP12T U2266 ( .A1(n6052), .A2(n5780), .A3(n6139), .A4(n5009), .ZN(
        n5075) );
  INVD1BWP12T U2267 ( .I(n5632), .ZN(n5275) );
  ND2D1BWP12T U2268 ( .A1(a[0]), .A2(n5275), .ZN(n5704) );
  IND4D1BWP12T U2269 ( .A1(n5032), .B1(n5067), .B2(n5010), .B3(n5704), .ZN(
        n5013) );
  OR4XD1BWP12T U2270 ( .A1(n5036), .A2(n5021), .A3(n5011), .A4(n5024), .Z(
        n5012) );
  NR4D0BWP12T U2271 ( .A1(n5015), .A2(n5014), .A3(n5013), .A4(n5012), .ZN(
        n5073) );
  INVD1BWP12T U2272 ( .I(n5670), .ZN(n5537) );
  AOI22D1BWP12T U2273 ( .A1(n5057), .A2(n5248), .B1(n5052), .B2(n5249), .ZN(
        n5017) );
  AOI22D1BWP12T U2274 ( .A1(n5181), .A2(n5095), .B1(n5051), .B2(n5250), .ZN(
        n5016) );
  ND2D1BWP12T U2275 ( .A1(n5017), .A2(n5016), .ZN(n5063) );
  NR2D1BWP12T U2276 ( .A1(n5047), .A2(n5261), .ZN(n5020) );
  OAI22D1BWP12T U2277 ( .A1(n5150), .A2(n5045), .B1(n5131), .B2(n5018), .ZN(
        n5019) );
  AOI211D1BWP12T U2278 ( .A1(n5285), .A2(n5095), .B(n5020), .C(n5019), .ZN(
        n5022) );
  OAI22D1BWP12T U2279 ( .A1(n5022), .A2(n5081), .B1(n5703), .B2(n5021), .ZN(
        n5023) );
  AOI211D1BWP12T U2280 ( .A1(n5079), .A2(n5063), .B(n5528), .C(n5023), .ZN(
        n5843) );
  INVD1BWP12T U2281 ( .I(n5024), .ZN(n5039) );
  OAI22D1BWP12T U2282 ( .A1(n5039), .A2(n5068), .B1(n5038), .B2(n5070), .ZN(
        n6051) );
  AOI22D1BWP12T U2283 ( .A1(b[3]), .A2(n5026), .B1(n5770), .B2(n5025), .ZN(
        n5027) );
  OAI211D1BWP12T U2284 ( .A1(n5703), .A2(n5028), .B(n5041), .C(n5027), .ZN(
        n6019) );
  MAOI22D0BWP12T U2285 ( .A1(b[3]), .A2(n5030), .B1(n5081), .B2(n5029), .ZN(
        n5031) );
  OAI211D1BWP12T U2286 ( .A1(n5703), .A2(n5032), .B(n5041), .C(n5031), .ZN(
        n5985) );
  MAOI22D0BWP12T U2287 ( .A1(b[3]), .A2(n5034), .B1(n5081), .B2(n5033), .ZN(
        n5035) );
  OAI211D1BWP12T U2288 ( .A1(n5703), .A2(n5036), .B(n5041), .C(n5035), .ZN(
        n5970) );
  INVD1BWP12T U2289 ( .I(n5037), .ZN(n5042) );
  AOI22D1BWP12T U2290 ( .A1(b[4]), .A2(n5039), .B1(b[3]), .B2(n5038), .ZN(
        n5040) );
  OAI211D1BWP12T U2291 ( .A1(n5042), .A2(n5081), .B(n5041), .C(n5040), .ZN(
        n5938) );
  ND4D1BWP12T U2292 ( .A1(n6019), .A2(n5985), .A3(n5970), .A4(n5938), .ZN(
        n5043) );
  NR4D0BWP12T U2293 ( .A1(n5843), .A2(n5044), .A3(n6051), .A4(n5043), .ZN(
        n5072) );
  NR2D1BWP12T U2294 ( .A1(n5045), .A2(n5191), .ZN(n5049) );
  OAI22D1BWP12T U2295 ( .A1(n5193), .A2(n5047), .B1(n5131), .B2(n5046), .ZN(
        n5048) );
  AOI211D1BWP12T U2296 ( .A1(n5095), .A2(n5159), .B(n5049), .C(n5048), .ZN(
        n5053) );
  MOAI22D0BWP12T U2297 ( .A1(n5053), .A2(n5081), .B1(n5055), .B2(b[3]), .ZN(
        n5050) );
  AOI211D1BWP12T U2298 ( .A1(b[4]), .A2(n5704), .B(n5528), .C(n5050), .ZN(
        n5699) );
  AOI22D1BWP12T U2299 ( .A1(n5052), .A2(n5207), .B1(n5051), .B2(n5188), .ZN(
        n5060) );
  MAOI22D0BWP12T U2300 ( .A1(n5056), .A2(n5055), .B1(n5054), .B2(n5053), .ZN(
        n5059) );
  AOI22D1BWP12T U2301 ( .A1(n5057), .A2(n5230), .B1(n5095), .B2(n5228), .ZN(
        n5058) );
  AOI32D1BWP12T U2302 ( .A1(n5060), .A2(n5059), .A3(n5058), .B1(n5081), .B2(
        n5059), .ZN(n5061) );
  AOI211D1BWP12T U2303 ( .A1(n5145), .A2(n5062), .B(n5528), .C(n5061), .ZN(
        n5922) );
  MOAI22D0BWP12T U2304 ( .A1(n5816), .A2(n5703), .B1(n5063), .B2(n5770), .ZN(
        n5064) );
  AOI211D1BWP12T U2305 ( .A1(n5079), .A2(n5066), .B(n5065), .C(n5064), .ZN(
        n5668) );
  OAI22D1BWP12T U2306 ( .A1(n5070), .A2(n5069), .B1(n5068), .B2(n5067), .ZN(
        n5861) );
  NR4D0BWP12T U2307 ( .A1(n5699), .A2(n5922), .A3(n5668), .A4(n5861), .ZN(
        n5071) );
  OAI211D1BWP12T U2308 ( .A1(n5073), .A2(n5537), .B(n5072), .C(n5071), .ZN(
        n5074) );
  NR4D0BWP12T U2309 ( .A1(n5077), .A2(n5076), .A3(n5075), .A4(n5074), .ZN(
        n5568) );
  MOAI22D0BWP12T U2310 ( .A1(n5081), .A2(n5080), .B1(n5079), .B2(n5078), .ZN(
        n6037) );
  IND4D1BWP12T U2311 ( .A1(n6037), .B1(n6071), .B2(n5083), .B3(n5082), .ZN(
        n5506) );
  INVD1BWP12T U2312 ( .I(n5084), .ZN(n5167) );
  ND2D1BWP12T U2313 ( .A1(n5086), .A2(n5085), .ZN(n5087) );
  OAI22D1BWP12T U2314 ( .A1(n5249), .A2(n5282), .B1(b[2]), .B2(n5087), .ZN(
        n5089) );
  OAI22D1BWP12T U2315 ( .A1(n5250), .A2(n5286), .B1(n5181), .B2(n5288), .ZN(
        n5088) );
  NR2D1BWP12T U2316 ( .A1(n5089), .A2(n5088), .ZN(n5223) );
  OAI22D1BWP12T U2317 ( .A1(n5090), .A2(n5280), .B1(n5223), .B2(n5263), .ZN(
        n6041) );
  AOI22D1BWP12T U2318 ( .A1(n5239), .A2(n5242), .B1(n5241), .B2(n5525), .ZN(
        n5530) );
  OAI21D1BWP12T U2319 ( .A1(n5136), .A2(n5138), .B(n5530), .ZN(n5665) );
  INVD1BWP12T U2320 ( .I(n5665), .ZN(n5515) );
  OAI21D1BWP12T U2321 ( .A1(n5171), .A2(n5269), .B(n5515), .ZN(n5824) );
  ND4D1BWP12T U2322 ( .A1(n5147), .A2(n5092), .A3(n6009), .A4(n5091), .ZN(
        n5093) );
  NR4D0BWP12T U2323 ( .A1(n5167), .A2(n6041), .A3(n5824), .A4(n5093), .ZN(
        n5115) );
  AOI222D1BWP12T U2324 ( .A1(a[2]), .A2(n5097), .B1(b[2]), .B2(n5096), .C1(
        n5095), .C2(n5094), .ZN(n5103) );
  AOI22D1BWP12T U2325 ( .A1(n5440), .A2(n5098), .B1(a[1]), .B2(n5275), .ZN(
        n5102) );
  AOI22D1BWP12T U2326 ( .A1(n5100), .A2(n5240), .B1(n5238), .B2(n5099), .ZN(
        n5101) );
  OAI211D1BWP12T U2327 ( .A1(b[3]), .A2(n5103), .B(n5102), .C(n5101), .ZN(
        n5814) );
  AOI22D1BWP12T U2328 ( .A1(n5238), .A2(n5278), .B1(n5240), .B2(n5104), .ZN(
        n5108) );
  AOI22D1BWP12T U2329 ( .A1(n5525), .A2(n5106), .B1(n5242), .B2(n5105), .ZN(
        n5107) );
  ND2D1BWP12T U2330 ( .A1(n5108), .A2(n5107), .ZN(n5707) );
  NR4D0BWP12T U2331 ( .A1(n5665), .A2(n5707), .A3(n5971), .A4(n5109), .ZN(
        n5111) );
  INVD1BWP12T U2332 ( .I(n5110), .ZN(n5986) );
  ND4D1BWP12T U2333 ( .A1(n5112), .A2(n5111), .A3(n5757), .A4(n5986), .ZN(
        n5496) );
  NR4D0BWP12T U2334 ( .A1(n5814), .A2(n5513), .A3(n5496), .A4(n5113), .ZN(
        n5114) );
  AOI32D1BWP12T U2335 ( .A1(n5116), .A2(n5115), .A3(n5114), .B1(b[4]), .B2(
        n5115), .ZN(n5303) );
  ND2D1BWP12T U2336 ( .A1(n5525), .A2(n5117), .ZN(n6109) );
  OAI22D1BWP12T U2337 ( .A1(n5119), .A2(n5136), .B1(n5118), .B2(n5245), .ZN(
        n5120) );
  AOI211D1BWP12T U2338 ( .A1(n5242), .A2(n5121), .B(b[4]), .C(n5120), .ZN(
        n5526) );
  AOI21D1BWP12T U2339 ( .A1(b[4]), .A2(n6109), .B(n5526), .ZN(n5871) );
  OAI22D1BWP12T U2340 ( .A1(n5122), .A2(n5284), .B1(n5282), .B2(n5158), .ZN(
        n5125) );
  OAI22D1BWP12T U2341 ( .A1(n5123), .A2(n5286), .B1(n5159), .B2(n5288), .ZN(
        n5124) );
  NR2D1BWP12T U2342 ( .A1(n5125), .A2(n5124), .ZN(n5216) );
  NR2D1BWP12T U2343 ( .A1(n5216), .A2(n5263), .ZN(n5126) );
  AOI211D1BWP12T U2344 ( .A1(n5258), .A2(n6111), .B(n5871), .C(n5126), .ZN(
        n5867) );
  NR2D1BWP12T U2345 ( .A1(a[0]), .A2(b[0]), .ZN(n5133) );
  NR2D1BWP12T U2346 ( .A1(a[1]), .A2(n5379), .ZN(n5132) );
  MAOI22D0BWP12T U2347 ( .A1(b[2]), .A2(n5129), .B1(n5128), .B2(n5127), .ZN(
        n5130) );
  OAI31D1BWP12T U2348 ( .A1(n5133), .A2(n5132), .A3(n5131), .B(n5130), .ZN(
        n5137) );
  AOI222D1BWP12T U2349 ( .A1(n5137), .A2(n5136), .B1(n5135), .B2(n5240), .C1(
        n5134), .C2(n5238), .ZN(n5510) );
  ND2D1BWP12T U2350 ( .A1(b[4]), .A2(n5707), .ZN(n5509) );
  ND4D1BWP12T U2351 ( .A1(n5510), .A2(n5146), .A3(n5138), .A4(n5509), .ZN(
        n5139) );
  NR4D0BWP12T U2352 ( .A1(n5769), .A2(n5172), .A3(n5140), .A4(n5139), .ZN(
        n5170) );
  NR2D1BWP12T U2353 ( .A1(n5188), .A2(n5286), .ZN(n5142) );
  OAI22D1BWP12T U2354 ( .A1(n5207), .A2(n5282), .B1(n5228), .B2(n5288), .ZN(
        n5141) );
  AOI211D1BWP12T U2355 ( .A1(n5144), .A2(n5143), .B(n5142), .C(n5141), .ZN(
        n5218) );
  NR2D1BWP12T U2356 ( .A1(n5145), .A2(n5201), .ZN(n5260) );
  ND2D1BWP12T U2357 ( .A1(n5260), .A2(n5165), .ZN(n5295) );
  OAI222D1BWP12T U2358 ( .A1(n5280), .A2(n5216), .B1(n5263), .B2(n5218), .C1(
        n5295), .C2(n5146), .ZN(n6144) );
  INVD1BWP12T U2359 ( .I(n5147), .ZN(n5155) );
  AOI22D1BWP12T U2360 ( .A1(n5248), .A2(n5254), .B1(n5249), .B2(n5255), .ZN(
        n5149) );
  ND2D1BWP12T U2361 ( .A1(n5181), .A2(n5192), .ZN(n5148) );
  OAI211D1BWP12T U2362 ( .A1(n5288), .A2(n5150), .B(n5149), .C(n5148), .ZN(
        n5175) );
  AOI22D1BWP12T U2363 ( .A1(n5287), .A2(n5254), .B1(n5285), .B2(n5192), .ZN(
        n5152) );
  ND2D1BWP12T U2364 ( .A1(n5283), .A2(n5262), .ZN(n5151) );
  OAI211D1BWP12T U2365 ( .A1(n5284), .A2(n5261), .B(n5152), .C(n5151), .ZN(
        n5153) );
  AOI22D1BWP12T U2366 ( .A1(n5258), .A2(n5175), .B1(n5290), .B2(n5153), .ZN(
        n5154) );
  OAI211D1BWP12T U2367 ( .A1(n5168), .A2(n5155), .B(n5154), .C(n5165), .ZN(
        n5755) );
  IND4D1BWP12T U2368 ( .A1(n5281), .B1(n5925), .B2(n6145), .B3(n5755), .ZN(
        n5156) );
  NR4D0BWP12T U2369 ( .A1(n5157), .A2(n6144), .A3(n5608), .A4(n5156), .ZN(
        n5169) );
  AOI22D1BWP12T U2370 ( .A1(n5208), .A2(n5254), .B1(n5255), .B2(n5158), .ZN(
        n5161) );
  AOI22D1BWP12T U2371 ( .A1(n5262), .A2(n5188), .B1(n5192), .B2(n5159), .ZN(
        n5160) );
  ND2D1BWP12T U2372 ( .A1(n5161), .A2(n5160), .ZN(n5203) );
  AOI22D1BWP12T U2373 ( .A1(n5254), .A2(n5230), .B1(n5255), .B2(n5207), .ZN(
        n5163) );
  AOI22D1BWP12T U2374 ( .A1(n5192), .A2(n5228), .B1(n5262), .B2(n5229), .ZN(
        n5162) );
  ND2D1BWP12T U2375 ( .A1(n5163), .A2(n5162), .ZN(n5164) );
  AOI22D1BWP12T U2376 ( .A1(n5258), .A2(n5203), .B1(n5290), .B2(n5164), .ZN(
        n5166) );
  OAI211D1BWP12T U2377 ( .A1(n5168), .A2(n5167), .B(n5166), .C(n5165), .ZN(
        n5771) );
  ND4D1BWP12T U2378 ( .A1(n5867), .A2(n5170), .A3(n5169), .A4(n5771), .ZN(
        n5302) );
  ND2D1BWP12T U2379 ( .A1(n5703), .A2(n5171), .ZN(n5199) );
  ND2D1BWP12T U2380 ( .A1(n5199), .A2(n5172), .ZN(n5176) );
  INVD1BWP12T U2381 ( .I(n5173), .ZN(n5174) );
  AOI222D1BWP12T U2382 ( .A1(n5176), .A2(n5204), .B1(n5175), .B2(n5290), .C1(
        n5174), .C2(n5201), .ZN(n5999) );
  ND2D1BWP12T U2383 ( .A1(n5199), .A2(n5281), .ZN(n5184) );
  OAI22D1BWP12T U2384 ( .A1(n5177), .A2(n5284), .B1(n5250), .B2(n5282), .ZN(
        n5180) );
  OAI22D1BWP12T U2385 ( .A1(n5249), .A2(n5288), .B1(n5178), .B2(n5286), .ZN(
        n5179) );
  NR2D1BWP12T U2386 ( .A1(n5180), .A2(n5179), .ZN(n5296) );
  AOI22D1BWP12T U2387 ( .A1(n5256), .A2(n5254), .B1(n5181), .B2(n5255), .ZN(
        n5183) );
  ND2D1BWP12T U2388 ( .A1(n5248), .A2(n5192), .ZN(n5182) );
  OAI211D1BWP12T U2389 ( .A1(n5288), .A2(n5261), .B(n5183), .C(n5182), .ZN(
        n5279) );
  AOI222D1BWP12T U2390 ( .A1(n5184), .A2(n5204), .B1(n5201), .B2(n5296), .C1(
        n5279), .C2(n5290), .ZN(n5978) );
  ND2D1BWP12T U2391 ( .A1(n5199), .A2(n5608), .ZN(n5187) );
  AOI22D1BWP12T U2392 ( .A1(n5256), .A2(n5192), .B1(n5248), .B2(n5255), .ZN(
        n5186) );
  ND2D1BWP12T U2393 ( .A1(n5285), .A2(n5262), .ZN(n5185) );
  OAI211D1BWP12T U2394 ( .A1(n5282), .A2(n5261), .B(n5186), .C(n5185), .ZN(
        n5225) );
  AOI222D1BWP12T U2395 ( .A1(n5187), .A2(n5204), .B1(n5201), .B2(n5223), .C1(
        n5225), .C2(n5290), .ZN(n5949) );
  INVD1BWP12T U2396 ( .I(n5199), .ZN(n5270) );
  AOI22D1BWP12T U2397 ( .A1(n5254), .A2(n5228), .B1(n5255), .B2(n5188), .ZN(
        n5190) );
  AOI22D1BWP12T U2398 ( .A1(n5262), .A2(n5230), .B1(n5192), .B2(n5207), .ZN(
        n5189) );
  AOI21D1BWP12T U2399 ( .A1(n5190), .A2(n5189), .B(n5263), .ZN(n5197) );
  AOI22D1BWP12T U2400 ( .A1(b[2]), .A2(n5211), .B1(n5255), .B2(n5191), .ZN(
        n5195) );
  ND2D1BWP12T U2401 ( .A1(n5193), .A2(n5192), .ZN(n5194) );
  OAI211D1BWP12T U2402 ( .A1(n5208), .A2(n5288), .B(n5195), .C(n5194), .ZN(
        n5697) );
  MOAI22D0BWP12T U2403 ( .A1(n5280), .A2(n5697), .B1(n5260), .B2(n5706), .ZN(
        n5196) );
  AOI211D1BWP12T U2404 ( .A1(n5270), .A2(n5198), .B(n5197), .C(n5196), .ZN(
        n5930) );
  NR4D0BWP12T U2405 ( .A1(n5999), .A2(n5978), .A3(n5949), .A4(n5930), .ZN(
        n5300) );
  ND2D1BWP12T U2406 ( .A1(n5200), .A2(n5199), .ZN(n5205) );
  AOI222D1BWP12T U2407 ( .A1(n5205), .A2(n5204), .B1(n5203), .B2(n5290), .C1(
        n5202), .C2(n5201), .ZN(n6022) );
  INVD1BWP12T U2408 ( .I(n5206), .ZN(n5226) );
  OAI22D1BWP12T U2409 ( .A1(n5208), .A2(n5286), .B1(n5288), .B2(n5207), .ZN(
        n5209) );
  AOI221D1BWP12T U2410 ( .A1(n5212), .A2(b[2]), .B1(n5211), .B2(n5210), .C(
        n5209), .ZN(n5236) );
  OAI222D1BWP12T U2411 ( .A1(n5280), .A2(n5226), .B1(n5263), .B2(n5236), .C1(
        n5295), .C2(n5213), .ZN(n6080) );
  NR2D1BWP12T U2412 ( .A1(n5229), .A2(n5286), .ZN(n5215) );
  OAI22D1BWP12T U2413 ( .A1(n5231), .A2(n5282), .B1(n5230), .B2(n5284), .ZN(
        n5214) );
  AOI211D1BWP12T U2414 ( .A1(n5262), .A2(a[29]), .B(n5215), .C(n5214), .ZN(
        n5217) );
  OAI222D1BWP12T U2415 ( .A1(n5280), .A2(n5218), .B1(n5263), .B2(n5217), .C1(
        n5295), .C2(n5216), .ZN(n6110) );
  NR4D0BWP12T U2416 ( .A1(n6022), .A2(n6080), .A3(n6110), .A4(n5219), .ZN(
        n5299) );
  NR2D1BWP12T U2417 ( .A1(n5283), .A2(n5286), .ZN(n5222) );
  OAI22D1BWP12T U2418 ( .A1(n5289), .A2(n5282), .B1(b[2]), .B2(n5220), .ZN(
        n5221) );
  AOI211D1BWP12T U2419 ( .A1(n5262), .A2(a[30]), .B(n5222), .C(n5221), .ZN(
        n5224) );
  OAI222D1BWP12T U2420 ( .A1(n5225), .A2(n5280), .B1(n5263), .B2(n5224), .C1(
        n5295), .C2(n5223), .ZN(n5607) );
  NR2D1BWP12T U2421 ( .A1(b[4]), .A2(n5705), .ZN(n6112) );
  MAOI22D0BWP12T U2422 ( .A1(n6112), .A2(n5227), .B1(n5295), .B2(n5226), .ZN(
        n5235) );
  OAI22D1BWP12T U2423 ( .A1(n5229), .A2(n5282), .B1(n5228), .B2(n5284), .ZN(
        n5233) );
  OAI22D1BWP12T U2424 ( .A1(n5231), .A2(n5288), .B1(n5230), .B2(n5286), .ZN(
        n5232) );
  OAI21D1BWP12T U2425 ( .A1(n5233), .A2(n5232), .B(n5290), .ZN(n5234) );
  OAI211D1BWP12T U2426 ( .A1(n5236), .A2(n5280), .B(n5235), .C(n5234), .ZN(
        n5729) );
  NR2D1BWP12T U2427 ( .A1(n5245), .A2(n5274), .ZN(n5886) );
  AOI21D1BWP12T U2428 ( .A1(n5238), .A2(n5237), .B(b[4]), .ZN(n5244) );
  AOI22D1BWP12T U2429 ( .A1(n5242), .A2(n5241), .B1(n5240), .B2(n5239), .ZN(
        n5243) );
  OAI211D1BWP12T U2430 ( .A1(n5246), .A2(n5245), .B(n5244), .C(n5243), .ZN(
        n5520) );
  OAI21D1BWP12T U2431 ( .A1(n5886), .A2(n5703), .B(n5520), .ZN(n5647) );
  ND2D1BWP12T U2432 ( .A1(n5258), .A2(n5281), .ZN(n5247) );
  OAI211D1BWP12T U2433 ( .A1(n5296), .A2(n5263), .B(n5647), .C(n5247), .ZN(
        n5653) );
  NR2D1BWP12T U2434 ( .A1(n5248), .A2(n5288), .ZN(n5252) );
  OAI22D1BWP12T U2435 ( .A1(n5250), .A2(n5284), .B1(n5249), .B2(n5286), .ZN(
        n5251) );
  AOI211D1BWP12T U2436 ( .A1(n5253), .A2(b[2]), .B(n5252), .C(n5251), .ZN(
        n5257) );
  OAI222D1BWP12T U2437 ( .A1(n5259), .A2(n5280), .B1(n5263), .B2(n5257), .C1(
        n5295), .C2(n5269), .ZN(n5667) );
  NR4D0BWP12T U2438 ( .A1(n5607), .A2(n5729), .A3(n5653), .A4(n5667), .ZN(
        n5298) );
  AOI22D1BWP12T U2439 ( .A1(n5256), .A2(n5255), .B1(n5285), .B2(n5254), .ZN(
        n5266) );
  AOI22D1BWP12T U2440 ( .A1(n5260), .A2(n5259), .B1(n5258), .B2(n5257), .ZN(
        n5265) );
  MAOI22D0BWP12T U2441 ( .A1(n5287), .A2(n5262), .B1(n5261), .B2(n5286), .ZN(
        n5264) );
  AOI32D1BWP12T U2442 ( .A1(n5266), .A2(n5265), .A3(n5264), .B1(n5263), .B2(
        n5265), .ZN(n5267) );
  AOI211D1BWP12T U2443 ( .A1(n5270), .A2(n5269), .B(n5268), .C(n5267), .ZN(
        n5844) );
  ND2D1BWP12T U2444 ( .A1(n5272), .A2(n5271), .ZN(n5501) );
  INR3D0BWP12T U2445 ( .A1(n5274), .B1(n5273), .B2(n5937), .ZN(n5276) );
  ND2D1BWP12T U2446 ( .A1(a[31]), .A2(n5275), .ZN(n5602) );
  IND4D1BWP12T U2447 ( .A1(n5278), .B1(n5277), .B2(n5276), .B3(n5602), .ZN(
        n5497) );
  MAOI22D0BWP12T U2448 ( .A1(n6112), .A2(n5281), .B1(n5280), .B2(n5279), .ZN(
        n5294) );
  OAI22D1BWP12T U2449 ( .A1(n5285), .A2(n5284), .B1(n5283), .B2(n5282), .ZN(
        n5292) );
  OAI22D1BWP12T U2450 ( .A1(n5289), .A2(n5288), .B1(n5287), .B2(n5286), .ZN(
        n5291) );
  OAI21D1BWP12T U2451 ( .A1(n5292), .A2(n5291), .B(n5290), .ZN(n5293) );
  OAI211D1BWP12T U2452 ( .A1(n5296), .A2(n5295), .B(n5294), .C(n5293), .ZN(
        n5895) );
  NR4D0BWP12T U2453 ( .A1(n5844), .A2(n5501), .A3(n5497), .A4(n5895), .ZN(
        n5297) );
  ND4D1BWP12T U2454 ( .A1(n5300), .A2(n5299), .A3(n5298), .A4(n5297), .ZN(
        n5301) );
  NR4D0BWP12T U2455 ( .A1(n5506), .A2(n5303), .A3(n5302), .A4(n5301), .ZN(
        n5567) );
  FA1D0BWP12T U2456 ( .A(n5306), .B(n5305), .CI(n5304), .CO(n5352), .S(n6049)
         );
  FA1D0BWP12T U2457 ( .A(n5309), .B(n5308), .CI(n5307), .CO(n5324), .S(n6011)
         );
  ND4D1BWP12T U2458 ( .A1(n5311), .A2(n5310), .A3(n6049), .A4(n6011), .ZN(
        n5378) );
  FA1D0BWP12T U2459 ( .A(n5314), .B(n5313), .CI(n5312), .CO(n5330), .S(n6131)
         );
  FA1D0BWP12T U2460 ( .A(n5317), .B(n5316), .CI(n5315), .CO(n5342), .S(n5724)
         );
  FA1D0BWP12T U2461 ( .A(n5320), .B(n5319), .CI(n5318), .CO(n4704), .S(n6098)
         );
  FA1D0BWP12T U2462 ( .A(n5323), .B(n5322), .CI(n5321), .CO(n5327), .S(n6069)
         );
  ND2D1BWP12T U2463 ( .A1(n6098), .A2(n6069), .ZN(n5337) );
  FA1D0BWP12T U2464 ( .A(n5326), .B(n5325), .CI(n5324), .CO(n5321), .S(n5991)
         );
  FA1D0BWP12T U2465 ( .A(n5329), .B(n5328), .CI(n5327), .CO(n5312), .S(n5966)
         );
  FA1D0BWP12T U2466 ( .A(n5332), .B(n5331), .CI(n5330), .CO(n5333), .S(n5946)
         );
  FA1D0BWP12T U2467 ( .A(n5335), .B(n5334), .CI(n5333), .CO(n5362), .S(n5919)
         );
  ND4D1BWP12T U2468 ( .A1(n5991), .A2(n5966), .A3(n5946), .A4(n5919), .ZN(
        n5336) );
  NR4D0BWP12T U2469 ( .A1(n5339), .A2(n5338), .A3(n5337), .A4(n5336), .ZN(
        n5340) );
  IND4D1BWP12T U2470 ( .A1(n5341), .B1(n6131), .B2(n5724), .B3(n5340), .ZN(
        n5377) );
  FA1D0BWP12T U2471 ( .A(n5344), .B(n5343), .CI(n5342), .CO(n5318), .S(n5888)
         );
  FA1D0BWP12T U2472 ( .A(n5347), .B(n5346), .CI(n5345), .CO(n5315), .S(n5748)
         );
  ND4D1BWP12T U2473 ( .A1(n5597), .A2(n5888), .A3(n5348), .A4(n5748), .ZN(
        n5376) );
  FA1D0BWP12T U2474 ( .A(n5351), .B(n5350), .CI(n5349), .CO(n5304), .S(n5864)
         );
  FA1D0BWP12T U2475 ( .A(n5354), .B(n5353), .CI(n5352), .CO(n5355), .S(n5691)
         );
  FA1D0BWP12T U2476 ( .A(n5357), .B(n5356), .CI(n5355), .CO(n5307), .S(n5677)
         );
  ND4D1BWP12T U2477 ( .A1(n5864), .A2(n5358), .A3(n5691), .A4(n5677), .ZN(
        n5370) );
  FA1D0BWP12T U2478 ( .A(n5361), .B(n5360), .CI(n5359), .CO(n5349), .S(n5644)
         );
  FA1D0BWP12T U2479 ( .A(n5364), .B(n5363), .CI(n5362), .CO(n5365), .S(n5836)
         );
  FA1D0BWP12T U2480 ( .A(n5367), .B(n5366), .CI(n5365), .CO(n5345), .S(n5775)
         );
  ND4D1BWP12T U2481 ( .A1(n5644), .A2(n5836), .A3(n5775), .A4(n5368), .ZN(
        n5369) );
  NR2D1BWP12T U2482 ( .A1(n5370), .A2(n5369), .ZN(n5371) );
  ND4D1BWP12T U2483 ( .A1(n5374), .A2(n5373), .A3(n5372), .A4(n5371), .ZN(
        n5375) );
  NR4D0BWP12T U2484 ( .A1(n5378), .A2(n5377), .A3(n5376), .A4(n5375), .ZN(
        n5411) );
  OAI21D1BWP12T U2485 ( .A1(n5804), .A2(n5380), .B(n5379), .ZN(n5382) );
  OAI22D1BWP12T U2486 ( .A1(n5492), .A2(n5805), .B1(n5633), .B2(n5798), .ZN(
        n5381) );
  ND2D1BWP12T U2487 ( .A1(n5382), .A2(n5381), .ZN(n5802) );
  NR2D1BWP12T U2488 ( .A1(n5989), .A2(n5988), .ZN(n5987) );
  NR4D0BWP12T U2489 ( .A1(n5987), .A2(n5385), .A3(n5384), .A4(n5383), .ZN(
        n5388) );
  ND4D1BWP12T U2490 ( .A1(n5389), .A2(n5388), .A3(n5387), .A4(n5386), .ZN(
        n5408) );
  NR2D1BWP12T U2491 ( .A1(n5390), .A2(n5874), .ZN(n5857) );
  ND2D1BWP12T U2492 ( .A1(b[22]), .A2(a[22]), .ZN(n6129) );
  ND2D1BWP12T U2493 ( .A1(b[12]), .A2(a[12]), .ZN(n5391) );
  IND4D1BWP12T U2494 ( .A1(n5857), .B1(n6129), .B2(n5645), .B3(n5391), .ZN(
        n5407) );
  NR2D1BWP12T U2495 ( .A1(n6010), .A2(n6024), .ZN(n6013) );
  ND2D1BWP12T U2496 ( .A1(b[16]), .A2(a[16]), .ZN(n5693) );
  IND4D1BWP12T U2497 ( .A1(n6013), .B1(n5673), .B2(n5693), .B3(n5392), .ZN(
        n5406) );
  NR4D0BWP12T U2498 ( .A1(n5396), .A2(n5395), .A3(n5394), .A4(n5393), .ZN(
        n5404) );
  ND2D1BWP12T U2499 ( .A1(b[26]), .A2(a[26]), .ZN(n5400) );
  ND2D1BWP12T U2500 ( .A1(b[25]), .A2(a[25]), .ZN(n5399) );
  ND2D1BWP12T U2501 ( .A1(b[24]), .A2(a[24]), .ZN(n5398) );
  ND2D1BWP12T U2502 ( .A1(b[23]), .A2(a[23]), .ZN(n5397) );
  ND4D1BWP12T U2503 ( .A1(n5400), .A2(n5399), .A3(n5398), .A4(n5397), .ZN(
        n5401) );
  AOI211D1BWP12T U2504 ( .A1(b[31]), .A2(a[31]), .B(n6128), .C(n5401), .ZN(
        n5403) );
  ND2D1BWP12T U2505 ( .A1(b[27]), .A2(a[27]), .ZN(n5402) );
  ND2D1BWP12T U2506 ( .A1(b[30]), .A2(a[30]), .ZN(n6095) );
  ND4D1BWP12T U2507 ( .A1(n5404), .A2(n5403), .A3(n5402), .A4(n6095), .ZN(
        n5405) );
  NR4D0BWP12T U2508 ( .A1(n5408), .A2(n5407), .A3(n5406), .A4(n5405), .ZN(
        n5409) );
  AOI31D1BWP12T U2509 ( .A1(n5411), .A2(n5802), .A3(n5410), .B(n5409), .ZN(
        n5491) );
  IND4D1BWP12T U2510 ( .A1(n5415), .B1(n5414), .B2(n5413), .B3(n5412), .ZN(
        n5428) );
  NR4D0BWP12T U2511 ( .A1(n5419), .A2(n5418), .A3(n5417), .A4(n5416), .ZN(
        n5427) );
  ND4D1BWP12T U2512 ( .A1(a[17]), .A2(a[16]), .A3(a[15]), .A4(a[31]), .ZN(
        n5420) );
  NR4D0BWP12T U2513 ( .A1(n5737), .A2(n5421), .A3(n5809), .A4(n5420), .ZN(
        n5426) );
  ND4D1BWP12T U2514 ( .A1(a[21]), .A2(a[18]), .A3(a[12]), .A4(a[11]), .ZN(
        n5422) );
  NR4D0BWP12T U2515 ( .A1(n6156), .A2(n5424), .A3(n5423), .A4(n5422), .ZN(
        n5425) );
  IND4D1BWP12T U2516 ( .A1(n5428), .B1(n5427), .B2(n5426), .B3(n5425), .ZN(
        n5490) );
  AN4XD1BWP12T U2517 ( .A1(n5431), .A2(n5430), .A3(n5916), .A4(n5429), .Z(
        n5488) );
  NR4D0BWP12T U2518 ( .A1(n5433), .A2(n5890), .A3(n5432), .A4(n6017), .ZN(
        n5487) );
  ND2D1BWP12T U2519 ( .A1(a[13]), .A2(n5476), .ZN(n5643) );
  IIND4D1BWP12T U2520 ( .A1(n5696), .A2(n5994), .B1(n5434), .B2(n5643), .ZN(
        n5451) );
  IND4D1BWP12T U2521 ( .A1(n5437), .B1(n5436), .B2(n5435), .B3(n5961), .ZN(
        n5450) );
  OR4XD1BWP12T U2522 ( .A1(n5440), .A2(n5439), .A3(n5438), .A4(n5804), .Z(
        n5449) );
  NR4D0BWP12T U2523 ( .A1(n5943), .A2(n5443), .A3(n5442), .A4(n5441), .ZN(
        n5445) );
  IND4D1BWP12T U2524 ( .A1(n5447), .B1(n5446), .B2(n5445), .B3(n5444), .ZN(
        n5448) );
  NR4D0BWP12T U2525 ( .A1(n5451), .A2(n5450), .A3(n5449), .A4(n5448), .ZN(
        n5486) );
  NR2D1BWP12T U2526 ( .A1(b[31]), .A2(n5593), .ZN(n5598) );
  ND4D1BWP12T U2527 ( .A1(n5455), .A2(n5454), .A3(n5453), .A4(n5452), .ZN(
        n5456) );
  NR4D0BWP12T U2528 ( .A1(n5459), .A2(n5458), .A3(n5457), .A4(n5456), .ZN(
        n5466) );
  IND4D1BWP12T U2529 ( .A1(n5461), .B1(n6135), .B2(n5460), .B3(n5840), .ZN(
        n5462) );
  AOI211D1BWP12T U2530 ( .A1(b[27]), .A2(n5758), .B(n5463), .C(n5462), .ZN(
        n5465) );
  ND4D1BWP12T U2531 ( .A1(n5467), .A2(n5466), .A3(n5465), .A4(n5464), .ZN(
        n5484) );
  IINR4D0BWP12T U2532 ( .A1(n5965), .A2(n5469), .B1(n6012), .B2(n5468), .ZN(
        n5482) );
  NR2D1BWP12T U2533 ( .A1(a[4]), .A2(n5703), .ZN(n5470) );
  NR4D0BWP12T U2534 ( .A1(n5472), .A2(n5471), .A3(n6134), .A4(n5470), .ZN(
        n5481) );
  NR4D0BWP12T U2535 ( .A1(n5475), .A2(n5474), .A3(n5473), .A4(n6068), .ZN(
        n5480) );
  NR2D1BWP12T U2536 ( .A1(a[13]), .A2(n5476), .ZN(n5477) );
  NR4D0BWP12T U2537 ( .A1(n5692), .A2(n5478), .A3(n6044), .A4(n5477), .ZN(
        n5479) );
  ND4D1BWP12T U2538 ( .A1(n5482), .A2(n5481), .A3(n5480), .A4(n5479), .ZN(
        n5483) );
  OAI22D1BWP12T U2539 ( .A1(n5598), .A2(n6093), .B1(n5484), .B2(n5483), .ZN(
        n5485) );
  ND4D1BWP12T U2540 ( .A1(n5488), .A2(n5487), .A3(n5486), .A4(n5485), .ZN(
        n5489) );
  OAI211D1BWP12T U2541 ( .A1(n5492), .A2(n5491), .B(n5490), .C(n5489), .ZN(
        n5566) );
  MAOI22D0BWP12T U2542 ( .A1(a[30]), .A2(n5493), .B1(a[30]), .B2(n5493), .ZN(
        n6119) );
  ND4D1BWP12T U2543 ( .A1(n5733), .A2(n6151), .A3(n5611), .A4(n5892), .ZN(
        n5563) );
  NR2D1BWP12T U2544 ( .A1(n5703), .A2(n5602), .ZN(n6038) );
  INR4D0BWP12T U2545 ( .A1(n5647), .B1(n5494), .B2(n6038), .B3(n5937), .ZN(
        n5505) );
  ND2D1BWP12T U2546 ( .A1(n5925), .A2(n5495), .ZN(n5535) );
  NR3D0BWP12T U2547 ( .A1(n5535), .A2(n5497), .A3(n5496), .ZN(n5499) );
  ND4D1BWP12T U2548 ( .A1(n5500), .A2(n5499), .A3(n5498), .A4(n6009), .ZN(
        n5502) );
  AOI211D1BWP12T U2549 ( .A1(n5703), .A2(n5502), .B(n5871), .C(n5501), .ZN(
        n5504) );
  INVD1BWP12T U2550 ( .I(n5845), .ZN(n5503) );
  IND4D1BWP12T U2551 ( .A1(n5506), .B1(n5505), .B2(n5504), .B3(n5503), .ZN(
        n5508) );
  AOI211D1BWP12T U2552 ( .A1(n5570), .A2(n5508), .B(n5507), .C(n5830), .ZN(
        n5561) );
  OA21D1BWP12T U2553 ( .A1(b[4]), .A2(n5510), .B(n5509), .Z(n5641) );
  ND2D1BWP12T U2554 ( .A1(n5641), .A2(n5511), .ZN(n5514) );
  AOI22D1BWP12T U2555 ( .A1(n5570), .A2(n5514), .B1(n5513), .B2(n5512), .ZN(
        n5560) );
  OAI21D1BWP12T U2556 ( .A1(n5814), .A2(b[4]), .B(n5570), .ZN(n5547) );
  AO21D1BWP12T U2557 ( .A1(b[4]), .A2(n5515), .B(n5547), .Z(n5831) );
  NR4D0BWP12T U2558 ( .A1(n5518), .A2(n5517), .A3(n6037), .A4(n5516), .ZN(
        n5529) );
  NR2D1BWP12T U2559 ( .A1(b[3]), .A2(n5519), .ZN(n5885) );
  OA21D1BWP12T U2560 ( .A1(n5521), .A2(n5885), .B(n5520), .Z(n5522) );
  MUX2ND0BWP12T U2561 ( .I0(n5522), .I1(a[31]), .S(n5528), .ZN(n5654) );
  AOI21D1BWP12T U2562 ( .A1(n5525), .A2(n5524), .B(n5523), .ZN(n5543) );
  NR2D1BWP12T U2563 ( .A1(n5543), .A2(n5528), .ZN(n6105) );
  INVD1BWP12T U2564 ( .I(n5526), .ZN(n5527) );
  OAI21D1BWP12T U2565 ( .A1(n5670), .A2(n6105), .B(n5527), .ZN(n5865) );
  OAI211D1BWP12T U2566 ( .A1(n5529), .A2(n5528), .B(n5654), .C(n5865), .ZN(
        n5556) );
  NR2D1BWP12T U2567 ( .A1(a[31]), .A2(n5670), .ZN(n5664) );
  IOA21D1BWP12T U2568 ( .A1(n5531), .A2(b[3]), .B(n5530), .ZN(n5666) );
  ND3D1BWP12T U2569 ( .A1(n5670), .A2(n5723), .A3(n5532), .ZN(n5728) );
  NR4D0BWP12T U2570 ( .A1(n5533), .A2(n5707), .A3(n5972), .A4(n5728), .ZN(
        n5534) );
  IND3D1BWP12T U2571 ( .A1(n5535), .B1(n5534), .B2(n5996), .ZN(n5546) );
  NR2D1BWP12T U2572 ( .A1(n5537), .A2(n5536), .ZN(n6065) );
  INVD1BWP12T U2573 ( .I(n5538), .ZN(n6142) );
  NR2D1BWP12T U2574 ( .A1(n5539), .A2(n6142), .ZN(n6149) );
  ND2D1BWP12T U2575 ( .A1(n5541), .A2(n5540), .ZN(n5783) );
  INR4D0BWP12T U2576 ( .A1(n5543), .B1(n5542), .B2(n5885), .B3(n5783), .ZN(
        n5544) );
  ND4D1BWP12T U2577 ( .A1(n6065), .A2(n6149), .A3(n5544), .A4(n5848), .ZN(
        n5545) );
  INR4D0BWP12T U2578 ( .A1(n6008), .B1(n5666), .B2(n5546), .B3(n5545), .ZN(
        n5554) );
  RCIAO21D0BWP12T U2579 ( .A1(n5703), .A2(n5666), .B(n5547), .ZN(n5827) );
  NR4D0BWP12T U2580 ( .A1(a[31]), .A2(n5827), .A3(n5548), .A4(n5866), .ZN(
        n5553) );
  AOI211D1BWP12T U2581 ( .A1(n5570), .A2(n5551), .B(n5550), .C(n5549), .ZN(
        n5552) );
  OAI211D1BWP12T U2582 ( .A1(n5664), .A2(n5554), .B(n5553), .C(n5552), .ZN(
        n5555) );
  NR4D0BWP12T U2583 ( .A1(n5558), .A2(n5557), .A3(n5556), .A4(n5555), .ZN(
        n5559) );
  AOI32D1BWP12T U2584 ( .A1(n5561), .A2(n5560), .A3(n5831), .B1(n5559), .B2(
        n5560), .ZN(n5562) );
  OAI31D1BWP12T U2585 ( .A1(n6119), .A2(n5564), .A3(n5563), .B(n5562), .ZN(
        n5565) );
  NR4D0BWP12T U2586 ( .A1(n5568), .A2(n5567), .A3(n5566), .A4(n5565), .ZN(
        n5572) );
  ND4D1BWP12T U2587 ( .A1(n5581), .A2(n5570), .A3(n6150), .A4(n5569), .ZN(
        n5571) );
  OAI211D1BWP12T U2588 ( .A1(n5574), .A2(n5573), .B(n5572), .C(n5571), .ZN(
        n5575) );
  AOI31D1BWP12T U2589 ( .A1(n6121), .A2(n5576), .A3(n5911), .B(n5575), .ZN(
        n5577) );
  OAI31D1BWP12T U2590 ( .A1(n6123), .A2(n5907), .A3(n5578), .B(n5577), .ZN(z)
         );
  NR2D1BWP12T U2591 ( .A1(a[31]), .A2(n5595), .ZN(n5591) );
  AOI22D1BWP12T U2592 ( .A1(n5580), .A2(n6160), .B1(n5579), .B2(n6122), .ZN(
        n5590) );
  NR3D1BWP12T U2593 ( .A1(a[31]), .A2(n5581), .A3(n6034), .ZN(n5613) );
  AOI22D1BWP12T U2594 ( .A1(n6162), .A2(n5583), .B1(n5595), .B2(n5582), .ZN(
        n5585) );
  OAI211D1BWP12T U2595 ( .A1(n6162), .A2(n6164), .B(a[31]), .C(b[31]), .ZN(
        n5584) );
  OAI211D1BWP12T U2596 ( .A1(n6120), .A2(n5586), .B(n5585), .C(n5584), .ZN(
        n5587) );
  OAI211D1BWP12T U2597 ( .A1(n5591), .A2(n5590), .B(n5589), .C(n5588), .ZN(
        c_out) );
  AOI211D1BWP12T U2598 ( .A1(n5595), .A2(n5594), .B(n5593), .C(n5592), .ZN(
        n5606) );
  OAI22D1BWP12T U2599 ( .A1(n5597), .A2(n6130), .B1(n5596), .B2(n6096), .ZN(
        n5605) );
  AOI21D1BWP12T U2600 ( .A1(b[31]), .A2(n5622), .B(n5598), .ZN(n5599) );
  OAI22D1BWP12T U2601 ( .A1(a[31]), .A2(n6156), .B1(n5599), .B2(n5671), .ZN(
        n5604) );
  NR2D1BWP12T U2602 ( .A1(b[4]), .A2(n5600), .ZN(n6143) );
  INVD1BWP12T U2603 ( .I(n6143), .ZN(n6108) );
  OAI22D1BWP12T U2604 ( .A1(n5602), .A2(n6108), .B1(n5601), .B2(n6138), .ZN(
        n5603) );
  NR4D0BWP12T U2605 ( .A1(n5606), .A2(n5605), .A3(n5604), .A4(n5603), .ZN(
        n5610) );
  AOI32D1BWP12T U2606 ( .A1(n6112), .A2(n6145), .A3(n5608), .B1(n5607), .B2(
        n6145), .ZN(n5609) );
  OAI211D1BWP12T U2607 ( .A1(n6034), .A2(n5611), .B(n5610), .C(n5609), .ZN(
        n5612) );
  AOI211D1BWP12T U2608 ( .A1(n6160), .A2(n5614), .B(n5613), .C(n5612), .ZN(
        n5618) );
  AOI22D1BWP12T U2609 ( .A1(n5616), .A2(n6162), .B1(n6164), .B2(n5615), .ZN(
        n5617) );
  OAI211D0BWP12T U2610 ( .A1(n5619), .A2(n6167), .B(n5618), .C(n5617), .ZN(
        result[31]) );
  BUFFXD0BWP12T U2611 ( .I(result[31]), .Z(n) );
  NR2D1BWP12T U2612 ( .A1(n5621), .A2(n5620), .ZN(n6040) );
  NR3D1BWP12T U2613 ( .A1(n5624), .A2(n5623), .A3(n5622), .ZN(n5629) );
  INVD1BWP12T U2614 ( .I(n5627), .ZN(n5626) );
  AOI32D1BWP12T U2615 ( .A1(n6135), .A2(b[0]), .A3(n5633), .B1(n6150), .B2(
        b[0]), .ZN(n5625) );
  OAI221D1BWP12T U2616 ( .A1(n5627), .A2(n6120), .B1(n5626), .B2(n6167), .C(
        n5625), .ZN(n5628) );
  AOI211D1BWP12T U2617 ( .A1(n6074), .A2(n5633), .B(n5629), .C(n5628), .ZN(
        n5640) );
  NR2D1BWP12T U2618 ( .A1(n6151), .A2(n6150), .ZN(n5630) );
  OAI32D1BWP12T U2619 ( .A1(n5633), .A2(n5632), .A3(n5631), .B1(n5630), .B2(
        n5633), .ZN(n5637) );
  AOI32D1BWP12T U2620 ( .A1(n6130), .A2(n5635), .A3(n6128), .B1(n5634), .B2(
        n5635), .ZN(n5636) );
  AOI211D1BWP12T U2621 ( .A1(n5638), .A2(n6133), .B(n5637), .C(n5636), .ZN(
        n5639) );
  OAI211D0BWP12T U2622 ( .A1(n5641), .A2(n6040), .B(n5640), .C(n5639), .ZN(
        result[0]) );
  AOI211D1BWP12T U2623 ( .A1(a[13]), .A2(n6092), .B(n5642), .C(n5939), .ZN(
        n5652) );
  OAI22D1BWP12T U2624 ( .A1(n5644), .A2(n6130), .B1(n6048), .B2(n5643), .ZN(
        n5651) );
  OAI22D1BWP12T U2625 ( .A1(a[13]), .A2(n6156), .B1(n6128), .B2(n5645), .ZN(
        n5650) );
  OAI22D1BWP12T U2626 ( .A1(n5648), .A2(n6138), .B1(n5647), .B2(n5646), .ZN(
        n5649) );
  NR4D0BWP12T U2627 ( .A1(n5652), .A2(n5651), .A3(n5650), .A4(n5649), .ZN(
        n5657) );
  MOAI22D0BWP12T U2628 ( .A1(n5654), .A2(n5866), .B1(n6145), .B2(n5653), .ZN(
        n5655) );
  AOI21D1BWP12T U2629 ( .A1(n5873), .A2(n5872), .B(n6034), .ZN(n5876) );
  OAI32D1BWP12T U2630 ( .A1(n5655), .A2(n5873), .A3(n5872), .B1(n5876), .B2(
        n5655), .ZN(n5656) );
  OAI211D1BWP12T U2631 ( .A1(n5658), .A2(n6113), .B(n5657), .C(n5656), .ZN(
        n5662) );
  OAI22D1BWP12T U2632 ( .A1(n5660), .A2(n6120), .B1(n5659), .B2(n6167), .ZN(
        n5661) );
  AO211D0BWP12T U2633 ( .A1(n6162), .A2(n5663), .B(n5662), .C(n5661), .Z(
        result[13]) );
  NR2D1BWP12T U2634 ( .A1(a[17]), .A2(n5709), .ZN(n6025) );
  AOI211D1BWP12T U2635 ( .A1(a[17]), .A2(n5709), .B(n6025), .C(n6034), .ZN(
        n5684) );
  NR2D1BWP12T U2636 ( .A1(n5664), .A2(n5866), .ZN(n6104) );
  AOI22D1BWP12T U2637 ( .A1(n6104), .A2(n5666), .B1(n6143), .B2(n5665), .ZN(
        n5682) );
  AOI22D1BWP12T U2638 ( .A1(n5668), .A2(n6052), .B1(n6145), .B2(n5667), .ZN(
        n5681) );
  NR2D1BWP12T U2639 ( .A1(n5670), .A2(n5669), .ZN(n6102) );
  NR2D1BWP12T U2640 ( .A1(b[17]), .A2(a[17]), .ZN(n5676) );
  AOI21D1BWP12T U2641 ( .A1(b[17]), .A2(op[1]), .B(n5671), .ZN(n5672) );
  AOI221D1BWP12T U2642 ( .A1(n6045), .A2(n5674), .B1(n6135), .B2(n5673), .C(
        n5672), .ZN(n5675) );
  OAI22D1BWP12T U2643 ( .A1(n5677), .A2(n6130), .B1(n5676), .B2(n5675), .ZN(
        n5678) );
  AOI211D1BWP12T U2644 ( .A1(n6074), .A2(n5679), .B(n6102), .C(n5678), .ZN(
        n5680) );
  ND3D1BWP12T U2645 ( .A1(n5682), .A2(n5681), .A3(n5680), .ZN(n5683) );
  AOI211D1BWP12T U2646 ( .A1(n6160), .A2(n5685), .B(n5684), .C(n5683), .ZN(
        n5689) );
  AOI22D1BWP12T U2647 ( .A1(n6164), .A2(n5687), .B1(n6162), .B2(n5686), .ZN(
        n5688) );
  OAI211D0BWP12T U2648 ( .A1(n5690), .A2(n6167), .B(n5689), .C(n5688), .ZN(
        result[17]) );
  NR2D1BWP12T U2649 ( .A1(b[16]), .A2(a[16]), .ZN(n5702) );
  OAI22D1BWP12T U2650 ( .A1(n5691), .A2(n6130), .B1(a[16]), .B2(n6156), .ZN(
        n5695) );
  MOAI22D0BWP12T U2651 ( .A1(n5693), .A2(n6128), .B1(n5692), .B2(n6135), .ZN(
        n5694) );
  AOI211D1BWP12T U2652 ( .A1(n5696), .A2(n6133), .B(n5695), .C(n5694), .ZN(
        n5701) );
  AOI22D1BWP12T U2653 ( .A1(n5699), .A2(n6052), .B1(n5698), .B2(n5697), .ZN(
        n5700) );
  OAI211D1BWP12T U2654 ( .A1(n5702), .A2(n6092), .B(n5701), .C(n5700), .ZN(
        n5718) );
  NR2D1BWP12T U2655 ( .A1(n5703), .A2(n6115), .ZN(n5825) );
  OAI21D1BWP12T U2656 ( .A1(n5706), .A2(n5705), .B(n5704), .ZN(n5708) );
  INVD1BWP12T U2657 ( .I(n6104), .ZN(n6148) );
  ND2D1BWP12T U2658 ( .A1(n6108), .A2(n6148), .ZN(n5936) );
  AOI22D1BWP12T U2659 ( .A1(n5825), .A2(n5708), .B1(n5707), .B2(n5936), .ZN(
        n5712) );
  OAI211D1BWP12T U2660 ( .A1(n6035), .A2(n5710), .B(n6151), .C(n5709), .ZN(
        n5711) );
  OAI211D1BWP12T U2661 ( .A1(n6113), .A2(n5713), .B(n5712), .C(n5711), .ZN(
        n5717) );
  OAI22D1BWP12T U2662 ( .A1(n5715), .A2(n6126), .B1(n6120), .B2(n5714), .ZN(
        n5716) );
  NR4D0BWP12T U2663 ( .A1(n6102), .A2(n5718), .A3(n5717), .A4(n5716), .ZN(
        n5719) );
  OAI21D0BWP12T U2664 ( .A1(n5720), .A2(n6167), .B(n5719), .ZN(result[16]) );
  OAI22D1BWP12T U2665 ( .A1(n5722), .A2(n6092), .B1(n5721), .B2(n6093), .ZN(
        n5726) );
  OAI22D1BWP12T U2666 ( .A1(n5724), .A2(n6130), .B1(n5723), .B2(n6108), .ZN(
        n5725) );
  AOI211D1BWP12T U2667 ( .A1(n6135), .A2(n5727), .B(n5726), .C(n5725), .ZN(
        n5731) );
  AOI22D1BWP12T U2668 ( .A1(n6145), .A2(n5729), .B1(n6104), .B2(n5728), .ZN(
        n5730) );
  OAI211D1BWP12T U2669 ( .A1(n5732), .A2(n6138), .B(n5731), .C(n5730), .ZN(
        n5740) );
  NR2D1BWP12T U2670 ( .A1(a[25]), .A2(a[24]), .ZN(n5735) );
  ND2D1BWP12T U2671 ( .A1(n5950), .A2(n6151), .ZN(n5914) );
  INR2D1BWP12T U2672 ( .A1(n5735), .B1(n5914), .ZN(n5899) );
  AOI22D1BWP12T U2673 ( .A1(b[28]), .A2(n6045), .B1(n5733), .B2(n5899), .ZN(
        n5738) );
  AOI21D1BWP12T U2674 ( .A1(n6151), .A2(n5734), .B(n6074), .ZN(n5913) );
  OAI21D1BWP12T U2675 ( .A1(n5735), .A2(n6034), .B(n5913), .ZN(n5785) );
  AOI21D1BWP12T U2676 ( .A1(n6151), .A2(n5736), .B(n5785), .ZN(n5902) );
  AOI32D1BWP12T U2677 ( .A1(n5738), .A2(a[28]), .A3(n6092), .B1(n5902), .B2(
        n5737), .ZN(n5739) );
  AOI211D1BWP12T U2678 ( .A1(n5741), .A2(n6160), .B(n5740), .C(n5739), .ZN(
        n5745) );
  MAOI22D0BWP12T U2679 ( .A1(n5743), .A2(n6162), .B1(n5742), .B2(n6167), .ZN(
        n5744) );
  OAI211D0BWP12T U2680 ( .A1(n5746), .A2(n6120), .B(n5745), .C(n5744), .ZN(
        result[28]) );
  NR2D1BWP12T U2681 ( .A1(n5747), .A2(n6113), .ZN(n5763) );
  OAI22D1BWP12T U2682 ( .A1(n5748), .A2(n6130), .B1(n5751), .B2(n6092), .ZN(
        n5749) );
  AOI211D1BWP12T U2683 ( .A1(n6104), .A2(n5750), .B(n6102), .C(n5749), .ZN(
        n5754) );
  AOI32D1BWP12T U2684 ( .A1(n5889), .A2(n5752), .A3(n5751), .B1(n6135), .B2(
        n5752), .ZN(n5753) );
  OAI211D1BWP12T U2685 ( .A1(n6115), .A2(n5755), .B(n5754), .C(n5753), .ZN(
        n5762) );
  OAI22D1BWP12T U2686 ( .A1(n5757), .A2(n6108), .B1(n5756), .B2(n6138), .ZN(
        n5761) );
  AOI22D1BWP12T U2687 ( .A1(b[27]), .A2(n6045), .B1(n5899), .B2(n5787), .ZN(
        n5759) );
  AOI32D1BWP12T U2688 ( .A1(n5759), .A2(a[27]), .A3(n6092), .B1(n5902), .B2(
        n5758), .ZN(n5760) );
  NR4D0BWP12T U2689 ( .A1(n5763), .A2(n5762), .A3(n5761), .A4(n5760), .ZN(
        n5767) );
  AOI22D1BWP12T U2690 ( .A1(n5765), .A2(n6122), .B1(n5764), .B2(n6164), .ZN(
        n5766) );
  OAI211D0BWP12T U2691 ( .A1(n5768), .A2(n6126), .B(n5767), .C(n5766), .ZN(
        result[27]) );
  ND2D1BWP12T U2692 ( .A1(n5770), .A2(n5769), .ZN(n5774) );
  AOI21D1BWP12T U2693 ( .A1(n5771), .A2(n5774), .B(n6115), .ZN(n5782) );
  AOI22D1BWP12T U2694 ( .A1(n5773), .A2(n5889), .B1(n6135), .B2(n5772), .ZN(
        n5779) );
  INVD1BWP12T U2695 ( .I(n5774), .ZN(n5777) );
  OAI22D1BWP12T U2696 ( .A1(n5775), .A2(n6130), .B1(n5784), .B2(n6092), .ZN(
        n5776) );
  AOI211D1BWP12T U2697 ( .A1(n5870), .A2(n5777), .B(n6102), .C(n5776), .ZN(
        n5778) );
  OAI211D1BWP12T U2698 ( .A1(n5780), .A2(n6138), .B(n5779), .C(n5778), .ZN(
        n5781) );
  AOI211D1BWP12T U2699 ( .A1(n6104), .A2(n5783), .B(n5782), .C(n5781), .ZN(
        n5789) );
  OAI21D1BWP12T U2700 ( .A1(n5784), .A2(n6128), .B(n6092), .ZN(n5786) );
  OAI32D1BWP12T U2701 ( .A1(n5787), .A2(n5899), .A3(n5786), .B1(a[26]), .B2(
        n5785), .ZN(n5788) );
  OAI211D1BWP12T U2702 ( .A1(n5790), .A2(n6113), .B(n5789), .C(n5788), .ZN(
        n5794) );
  OAI22D1BWP12T U2703 ( .A1(n5792), .A2(n6126), .B1(n5791), .B2(n6167), .ZN(
        n5793) );
  AO211D0BWP12T U2704 ( .A1(n6164), .A2(n5795), .B(n5794), .C(n5793), .Z(
        result[26]) );
  AOI22D1BWP12T U2705 ( .A1(n5799), .A2(n5798), .B1(n5797), .B2(n5796), .ZN(
        n5800) );
  OAI22D1BWP12T U2706 ( .A1(n6126), .A2(n5801), .B1(n6113), .B2(n5800), .ZN(
        n5823) );
  OAI22D1BWP12T U2707 ( .A1(n6120), .A2(n5803), .B1(n5802), .B2(n6130), .ZN(
        n5822) );
  AOI31D1BWP12T U2708 ( .A1(b[1]), .A2(n6135), .A3(n5805), .B(n5804), .ZN(
        n5820) );
  OAI22D1BWP12T U2709 ( .A1(n5807), .A2(n6092), .B1(n5806), .B2(n6128), .ZN(
        n5812) );
  ND2D1BWP12T U2710 ( .A1(n5809), .A2(n5808), .ZN(n5810) );
  OAI22D1BWP12T U2711 ( .A1(a[1]), .A2(n6156), .B1(n5810), .B2(n6034), .ZN(
        n5811) );
  AOI211D1BWP12T U2712 ( .A1(n6122), .A2(n5813), .B(n5812), .C(n5811), .ZN(
        n5819) );
  AOI22D1BWP12T U2713 ( .A1(n5817), .A2(n5816), .B1(n5815), .B2(n5814), .ZN(
        n5818) );
  OAI211D1BWP12T U2714 ( .A1(n6048), .A2(n5820), .B(n5819), .C(n5818), .ZN(
        n5821) );
  NR4D0BWP12T U2715 ( .A1(n5859), .A2(n5823), .A3(n5822), .A4(n5821), .ZN(
        n5829) );
  AOI22D1BWP12T U2716 ( .A1(n5827), .A2(n5826), .B1(n5825), .B2(n5824), .ZN(
        n5828) );
  OAI211D0BWP12T U2717 ( .A1(n5831), .A2(n5830), .B(n5829), .C(n5828), .ZN(
        result[1]) );
  NR2D1BWP12T U2718 ( .A1(a[24]), .A2(n5914), .ZN(n5832) );
  AOI211D1BWP12T U2719 ( .A1(b[25]), .A2(n6045), .B(n5832), .C(n5833), .ZN(
        n5834) );
  AOI22D1BWP12T U2720 ( .A1(n5834), .A2(n6092), .B1(n5913), .B2(n5833), .ZN(
        n5850) );
  ND2D1BWP12T U2721 ( .A1(a[24]), .A2(n6151), .ZN(n5835) );
  OAI22D1BWP12T U2722 ( .A1(n5836), .A2(n6130), .B1(a[25]), .B2(n5835), .ZN(
        n5842) );
  NR2D1BWP12T U2723 ( .A1(n6102), .A2(n5837), .ZN(n5945) );
  AOI22D1BWP12T U2724 ( .A1(b[25]), .A2(n6150), .B1(n5838), .B2(n6133), .ZN(
        n5839) );
  OAI211D1BWP12T U2725 ( .A1(n5840), .A2(n6096), .B(n5945), .C(n5839), .ZN(
        n5841) );
  AOI211D1BWP12T U2726 ( .A1(n5843), .A2(n6052), .B(n5842), .C(n5841), .ZN(
        n5847) );
  AOI22D1BWP12T U2727 ( .A1(n5845), .A2(n6143), .B1(n5844), .B2(n6145), .ZN(
        n5846) );
  OAI211D1BWP12T U2728 ( .A1(n5848), .A2(n6148), .B(n5847), .C(n5846), .ZN(
        n5849) );
  AOI211D1BWP12T U2729 ( .A1(n6160), .A2(n5851), .B(n5850), .C(n5849), .ZN(
        n5855) );
  AOI22D1BWP12T U2730 ( .A1(n5853), .A2(n6162), .B1(n6164), .B2(n5852), .ZN(
        n5854) );
  OAI211D0BWP12T U2731 ( .A1(n5856), .A2(n6167), .B(n5855), .C(n5854), .ZN(
        result[25]) );
  AOI22D1BWP12T U2732 ( .A1(b[14]), .A2(n6150), .B1(n5857), .B2(n6045), .ZN(
        n5863) );
  AOI211D1BWP12T U2733 ( .A1(n6052), .A2(n5861), .B(n5860), .C(n5859), .ZN(
        n5862) );
  OAI211D1BWP12T U2734 ( .A1(n5864), .A2(n6130), .B(n5863), .C(n5862), .ZN(
        n5869) );
  OAI22D1BWP12T U2735 ( .A1(n5867), .A2(n6115), .B1(n5866), .B2(n5865), .ZN(
        n5868) );
  AOI211D1BWP12T U2736 ( .A1(n5871), .A2(n5870), .B(n5869), .C(n5868), .ZN(
        n5878) );
  AO31D1BWP12T U2737 ( .A1(n5873), .A2(n6151), .A3(n5872), .B(n6150), .Z(n5875) );
  OAI32D1BWP12T U2738 ( .A1(a[14]), .A2(n6074), .A3(n5876), .B1(n5875), .B2(
        n5874), .ZN(n5877) );
  OA211D1BWP12T U2739 ( .A1(n5879), .A2(n6113), .B(n5878), .C(n5877), .Z(n5883) );
  AOI22D1BWP12T U2740 ( .A1(n5881), .A2(n6122), .B1(n6164), .B2(n5880), .ZN(
        n5882) );
  OAI211D0BWP12T U2741 ( .A1(n5884), .A2(n6126), .B(n5883), .C(n5882), .ZN(
        result[14]) );
  AOI22D1BWP12T U2742 ( .A1(n5886), .A2(n6143), .B1(n5885), .B2(n6104), .ZN(
        n5897) );
  OAI22D1BWP12T U2743 ( .A1(n5888), .A2(n6130), .B1(n5887), .B2(n6096), .ZN(
        n5894) );
  AOI22D1BWP12T U2744 ( .A1(b[29]), .A2(n6150), .B1(n5890), .B2(n5889), .ZN(
        n5891) );
  OAI211D1BWP12T U2745 ( .A1(n6034), .A2(n5892), .B(n5945), .C(n5891), .ZN(
        n5893) );
  AOI211D1BWP12T U2746 ( .A1(n6145), .A2(n5895), .B(n5894), .C(n5893), .ZN(
        n5896) );
  OAI211D1BWP12T U2747 ( .A1(n5898), .A2(n6138), .B(n5897), .C(n5896), .ZN(
        n5905) );
  AOI22D1BWP12T U2748 ( .A1(b[29]), .A2(n6045), .B1(n5900), .B2(n5899), .ZN(
        n5903) );
  AOI32D1BWP12T U2749 ( .A1(n5903), .A2(a[29]), .A3(n6092), .B1(n5902), .B2(
        n5901), .ZN(n5904) );
  AOI211D1BWP12T U2750 ( .A1(n6160), .A2(n5906), .B(n5905), .C(n5904), .ZN(
        n5910) );
  AOI22D1BWP12T U2751 ( .A1(n5908), .A2(n6162), .B1(n6122), .B2(n5907), .ZN(
        n5909) );
  OAI211D0BWP12T U2752 ( .A1(n5911), .A2(n6120), .B(n5910), .C(n5909), .ZN(
        result[29]) );
  AOI211D1BWP12T U2753 ( .A1(b[24]), .A2(n6045), .B(n6150), .C(n5912), .ZN(
        n5915) );
  AOI22D1BWP12T U2754 ( .A1(n5915), .A2(n5914), .B1(n5913), .B2(n5912), .ZN(
        n5927) );
  INVD1BWP12T U2755 ( .I(n5936), .ZN(n5924) );
  OAI22D1BWP12T U2756 ( .A1(n5917), .A2(n6096), .B1(n5916), .B2(n6093), .ZN(
        n5921) );
  OAI22D1BWP12T U2757 ( .A1(n5919), .A2(n6130), .B1(n5918), .B2(n6092), .ZN(
        n5920) );
  AOI211D1BWP12T U2758 ( .A1(n5922), .A2(n6052), .B(n5921), .C(n5920), .ZN(
        n5923) );
  OAI211D1BWP12T U2759 ( .A1(n5925), .A2(n5924), .B(n5945), .C(n5923), .ZN(
        n5926) );
  AO211D1BWP12T U2760 ( .A1(n6160), .A2(n5928), .B(n5927), .C(n5926), .Z(n5929) );
  AOI21D1BWP12T U2761 ( .A1(n5930), .A2(n6145), .B(n5929), .ZN(n5934) );
  AOI22D1BWP12T U2762 ( .A1(n6122), .A2(n5932), .B1(n6162), .B2(n5931), .ZN(
        n5933) );
  OAI211D0BWP12T U2763 ( .A1(n5935), .A2(n6120), .B(n5934), .C(n5933), .ZN(
        result[24]) );
  MOAI22D0BWP12T U2764 ( .A1(n6138), .A2(n5938), .B1(n5937), .B2(n5936), .ZN(
        n5948) );
  OAI211D1BWP12T U2765 ( .A1(n5939), .A2(n5940), .B(n6156), .C(n5951), .ZN(
        n5942) );
  OAI211D1BWP12T U2766 ( .A1(n5940), .A2(n6128), .B(a[23]), .C(n6092), .ZN(
        n5941) );
  AOI22D1BWP12T U2767 ( .A1(n5943), .A2(n6133), .B1(n5942), .B2(n5941), .ZN(
        n5944) );
  OAI211D1BWP12T U2768 ( .A1(n5946), .A2(n6130), .B(n5945), .C(n5944), .ZN(
        n5947) );
  AOI211D1BWP12T U2769 ( .A1(n5949), .A2(n6145), .B(n5948), .C(n5947), .ZN(
        n5954) );
  NR2D1BWP12T U2770 ( .A1(n5950), .A2(n6034), .ZN(n5952) );
  AOI32D1BWP12T U2771 ( .A1(n6152), .A2(n5952), .A3(n6155), .B1(n5951), .B2(
        n5952), .ZN(n5953) );
  OAI211D1BWP12T U2772 ( .A1(n6113), .A2(n5955), .B(n5954), .C(n5953), .ZN(
        n5959) );
  OAI22D1BWP12T U2773 ( .A1(n5957), .A2(n6120), .B1(n5956), .B2(n6126), .ZN(
        n5958) );
  AO211D0BWP12T U2774 ( .A1(n5960), .A2(n6122), .B(n5959), .C(n5958), .Z(
        result[23]) );
  IND2D1BWP12T U2775 ( .A1(n6152), .B1(n6151), .ZN(n6154) );
  AOI21D1BWP12T U2776 ( .A1(a[21]), .A2(n6081), .B(n6154), .ZN(n5977) );
  OAI22D1BWP12T U2777 ( .A1(n6045), .A2(n5962), .B1(n5961), .B2(n6133), .ZN(
        n5963) );
  AOI22D1BWP12T U2778 ( .A1(n5964), .A2(n6156), .B1(n6092), .B2(n5963), .ZN(
        n5968) );
  OAI22D1BWP12T U2779 ( .A1(n5966), .A2(n6130), .B1(n5965), .B2(n6096), .ZN(
        n5967) );
  AOI211D1BWP12T U2780 ( .A1(n6150), .A2(b[21]), .B(n5968), .C(n5967), .ZN(
        n5969) );
  INVD1BWP12T U2781 ( .I(n6102), .ZN(n6137) );
  OA211D1BWP12T U2782 ( .A1(n6138), .A2(n5970), .B(n5969), .C(n6137), .Z(n5974) );
  AOI22D1BWP12T U2783 ( .A1(n6104), .A2(n5972), .B1(n6143), .B2(n5971), .ZN(
        n5973) );
  OAI211D1BWP12T U2784 ( .A1(n5975), .A2(n6113), .B(n5974), .C(n5973), .ZN(
        n5976) );
  AOI211D1BWP12T U2785 ( .A1(n6145), .A2(n5978), .B(n5977), .C(n5976), .ZN(
        n5982) );
  MAOI22D0BWP12T U2786 ( .A1(n6122), .A2(n5980), .B1(n6120), .B2(n5979), .ZN(
        n5981) );
  OAI211D0BWP12T U2787 ( .A1(n5983), .A2(n6126), .B(n5982), .C(n5981), .ZN(
        result[21]) );
  INVD1BWP12T U2788 ( .I(n5984), .ZN(n6023) );
  NR2D1BWP12T U2789 ( .A1(a[19]), .A2(n6023), .ZN(n6083) );
  AOI211D1BWP12T U2790 ( .A1(a[19]), .A2(n6023), .B(n6083), .C(n6034), .ZN(
        n6001) );
  OAI22D1BWP12T U2791 ( .A1(n5986), .A2(n6108), .B1(n5985), .B2(n6138), .ZN(
        n5998) );
  AOI22D1BWP12T U2792 ( .A1(n6045), .A2(n5987), .B1(n6135), .B2(n5988), .ZN(
        n5990) );
  AOI22D1BWP12T U2793 ( .A1(n5990), .A2(n6092), .B1(n5989), .B2(n5988), .ZN(
        n5993) );
  OAI22D1BWP12T U2794 ( .A1(n5991), .A2(n6130), .B1(a[19]), .B2(n6156), .ZN(
        n5992) );
  AOI211D1BWP12T U2795 ( .A1(n5994), .A2(n6133), .B(n5993), .C(n5992), .ZN(
        n5995) );
  OAI211D1BWP12T U2796 ( .A1(n6148), .A2(n5996), .B(n5995), .C(n6137), .ZN(
        n5997) );
  AO211D1BWP12T U2797 ( .A1(n5999), .A2(n6145), .B(n5998), .C(n5997), .Z(n6000) );
  AOI211D1BWP12T U2798 ( .A1(n6160), .A2(n6002), .B(n6001), .C(n6000), .ZN(
        n6006) );
  AOI22D1BWP12T U2799 ( .A1(n6122), .A2(n6004), .B1(n6162), .B2(n6003), .ZN(
        n6005) );
  OAI211D0BWP12T U2800 ( .A1(n6007), .A2(n6120), .B(n6006), .C(n6005), .ZN(
        result[19]) );
  OAI22D1BWP12T U2801 ( .A1(n6009), .A2(n6108), .B1(n6008), .B2(n6148), .ZN(
        n6021) );
  OAI22D1BWP12T U2802 ( .A1(n6011), .A2(n6130), .B1(n6010), .B2(n6092), .ZN(
        n6016) );
  AOI22D1BWP12T U2803 ( .A1(n6013), .A2(n6045), .B1(n6012), .B2(n6135), .ZN(
        n6014) );
  OAI221D1BWP12T U2804 ( .A1(a[18]), .A2(n6156), .B1(n6024), .B2(n6092), .C(
        n6014), .ZN(n6015) );
  AOI211D1BWP12T U2805 ( .A1(n6017), .A2(n6133), .B(n6016), .C(n6015), .ZN(
        n6018) );
  OAI211D1BWP12T U2806 ( .A1(n6138), .A2(n6019), .B(n6018), .C(n6137), .ZN(
        n6020) );
  AOI211D1BWP12T U2807 ( .A1(n6022), .A2(n6145), .B(n6021), .C(n6020), .ZN(
        n6027) );
  OAI211D1BWP12T U2808 ( .A1(n6025), .A2(n6024), .B(n6151), .C(n6023), .ZN(
        n6026) );
  OAI211D1BWP12T U2809 ( .A1(n6113), .A2(n6028), .B(n6027), .C(n6026), .ZN(
        n6032) );
  OAI22D1BWP12T U2810 ( .A1(n6030), .A2(n6120), .B1(n6029), .B2(n6126), .ZN(
        n6031) );
  AO211D0BWP12T U2811 ( .A1(n6122), .A2(n6033), .B(n6032), .C(n6031), .Z(
        result[18]) );
  AOI211D1BWP12T U2812 ( .A1(a[15]), .A2(n6036), .B(n6035), .C(n6034), .ZN(
        n6058) );
  NR2D1BWP12T U2813 ( .A1(n6038), .A2(n6037), .ZN(n6039) );
  MAOI22D0BWP12T U2814 ( .A1(n6145), .A2(n6041), .B1(n6040), .B2(n6039), .ZN(
        n6056) );
  AOI22D1BWP12T U2815 ( .A1(n6150), .A2(n6043), .B1(n6074), .B2(n6042), .ZN(
        n6055) );
  AOI22D1BWP12T U2816 ( .A1(n6046), .A2(n6045), .B1(n6044), .B2(n6135), .ZN(
        n6054) );
  OAI22D1BWP12T U2817 ( .A1(n6049), .A2(n6130), .B1(n6048), .B2(n6047), .ZN(
        n6050) );
  AOI211D1BWP12T U2818 ( .A1(n6052), .A2(n6051), .B(n6102), .C(n6050), .ZN(
        n6053) );
  ND4D1BWP12T U2819 ( .A1(n6056), .A2(n6055), .A3(n6054), .A4(n6053), .ZN(
        n6057) );
  AOI211D1BWP12T U2820 ( .A1(n6160), .A2(n6059), .B(n6058), .C(n6057), .ZN(
        n6063) );
  AOI22D1BWP12T U2821 ( .A1(n6164), .A2(n6061), .B1(n6162), .B2(n6060), .ZN(
        n6062) );
  OAI211D0BWP12T U2822 ( .A1(n6064), .A2(n6167), .B(n6063), .C(n6062), .ZN(
        result[15]) );
  NR2D1BWP12T U2823 ( .A1(n6065), .A2(n6148), .ZN(n6079) );
  MAOI22D0BWP12T U2824 ( .A1(n6067), .A2(n6133), .B1(n6128), .B2(n6066), .ZN(
        n6077) );
  MOAI22D0BWP12T U2825 ( .A1(n6069), .A2(n6130), .B1(n6068), .B2(n6135), .ZN(
        n6073) );
  OAI22D1BWP12T U2826 ( .A1(n6071), .A2(n6108), .B1(n6138), .B2(n6070), .ZN(
        n6072) );
  AOI211D1BWP12T U2827 ( .A1(n6074), .A2(n6082), .B(n6073), .C(n6072), .ZN(
        n6076) );
  AOI32D1BWP12T U2828 ( .A1(n6077), .A2(n6076), .A3(n6092), .B1(n6075), .B2(
        n6076), .ZN(n6078) );
  AOI211D1BWP12T U2829 ( .A1(n6145), .A2(n6080), .B(n6079), .C(n6078), .ZN(
        n6085) );
  OAI211D1BWP12T U2830 ( .A1(n6083), .A2(n6082), .B(n6151), .C(n6081), .ZN(
        n6084) );
  OAI211D1BWP12T U2831 ( .A1(n6113), .A2(n6086), .B(n6085), .C(n6084), .ZN(
        n6090) );
  OAI22D1BWP12T U2832 ( .A1(n6088), .A2(n6126), .B1(n6167), .B2(n6087), .ZN(
        n6089) );
  AO211D0BWP12T U2833 ( .A1(n6091), .A2(n6164), .B(n6090), .C(n6089), .Z(
        result[20]) );
  NR2D1BWP12T U2834 ( .A1(b[30]), .A2(a[30]), .ZN(n6094) );
  OAI32D1BWP12T U2835 ( .A1(n6094), .A2(b[30]), .A3(n6093), .B1(n6092), .B2(
        n6094), .ZN(n6101) );
  OAI22D1BWP12T U2836 ( .A1(a[30]), .A2(n6156), .B1(n6128), .B2(n6095), .ZN(
        n6100) );
  OAI22D1BWP12T U2837 ( .A1(n6098), .A2(n6130), .B1(n6097), .B2(n6096), .ZN(
        n6099) );
  NR4D0BWP12T U2838 ( .A1(n6102), .A2(n6101), .A3(n6100), .A4(n6099), .ZN(
        n6107) );
  MAOI22D0BWP12T U2839 ( .A1(n6105), .A2(n6104), .B1(n6103), .B2(n6138), .ZN(
        n6106) );
  OAI211D1BWP12T U2840 ( .A1(n6109), .A2(n6108), .B(n6107), .C(n6106), .ZN(
        n6118) );
  AOI21D1BWP12T U2841 ( .A1(n6112), .A2(n6111), .B(n6110), .ZN(n6116) );
  OAI22D1BWP12T U2842 ( .A1(n6116), .A2(n6115), .B1(n6114), .B2(n6113), .ZN(
        n6117) );
  AOI211D1BWP12T U2843 ( .A1(n6119), .A2(n6151), .B(n6118), .C(n6117), .ZN(
        n6125) );
  MAOI22D0BWP12T U2844 ( .A1(n6123), .A2(n6122), .B1(n6121), .B2(n6120), .ZN(
        n6124) );
  OAI211D0BWP12T U2845 ( .A1(n6127), .A2(n6126), .B(n6125), .C(n6124), .ZN(
        result[30]) );
  OAI22D1BWP12T U2846 ( .A1(n6131), .A2(n6130), .B1(n6129), .B2(n6128), .ZN(
        n6141) );
  AOI22D1BWP12T U2847 ( .A1(n6135), .A2(n6134), .B1(n6133), .B2(n6132), .ZN(
        n6136) );
  OAI211D1BWP12T U2848 ( .A1(n6139), .A2(n6138), .B(n6137), .C(n6136), .ZN(
        n6140) );
  AOI211D1BWP12T U2849 ( .A1(b[22]), .A2(n6150), .B(n6141), .C(n6140), .ZN(
        n6147) );
  AOI22D1BWP12T U2850 ( .A1(n6145), .A2(n6144), .B1(n6143), .B2(n6142), .ZN(
        n6146) );
  OAI211D1BWP12T U2851 ( .A1(n6149), .A2(n6148), .B(n6147), .C(n6146), .ZN(
        n6158) );
  AOI21D1BWP12T U2852 ( .A1(n6152), .A2(n6151), .B(n6150), .ZN(n6153) );
  AOI32D1BWP12T U2853 ( .A1(n6156), .A2(n6155), .A3(n6154), .B1(a[22]), .B2(
        n6153), .ZN(n6157) );
  AOI211D1BWP12T U2854 ( .A1(n6160), .A2(n6159), .B(n6158), .C(n6157), .ZN(
        n6166) );
  AOI22D1BWP12T U2855 ( .A1(n6164), .A2(n6163), .B1(n6162), .B2(n6161), .ZN(
        n6165) );
  OAI211D0BWP12T U2856 ( .A1(n6168), .A2(n6167), .B(n6166), .C(n6165), .ZN(
        result[22]) );
endmodule


module memory_interface ( address, data_in, load, clk, reset, is_signed, 
        word_type, from_mem_data, to_mem_read_enable, to_mem_write_enable, 
        to_mem_mem_enable, to_mem_address, to_mem_data, data_out, write_ready, 
        output_valid, busy, store_BAR );
  input [11:0] address;
  input [31:0] data_in;
  input [1:0] word_type;
  input [15:0] from_mem_data;
  output [11:0] to_mem_address;
  output [15:0] to_mem_data;
  output [31:0] data_out;
  input load, clk, reset, is_signed, store_BAR;
  output to_mem_read_enable, to_mem_write_enable, to_mem_mem_enable,
         write_ready, output_valid, busy;
  wire   delayed_is_signed, fsm_N35, fsm_N34, fsm_N33, fsm_N32, fsm_state_0_,
         fsm_state_1_, fsm_state_2_, fsm_state_3_, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127;
  wire   [11:0] delay_addr_for_adder;
  wire   [11:0] delay_addr_single;
  wire   [31:0] delay_data_in32;
  wire   [15:0] delay_first_two_bytes_out;
  tri   [31:0] data_in;
  tri   clk;
  tri   reset;
  tri   [31:0] data_out;

  DFQD1BWP12T delay_first_two_bytes_out_reg_15_ ( .D(from_mem_data[7]), .CP(
        clk), .Q(delay_first_two_bytes_out[15]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_14_ ( .D(from_mem_data[6]), .CP(
        clk), .Q(delay_first_two_bytes_out[14]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_13_ ( .D(from_mem_data[5]), .CP(
        clk), .Q(delay_first_two_bytes_out[13]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_12_ ( .D(from_mem_data[4]), .CP(
        clk), .Q(delay_first_two_bytes_out[12]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_11_ ( .D(from_mem_data[3]), .CP(
        clk), .Q(delay_first_two_bytes_out[11]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_10_ ( .D(from_mem_data[2]), .CP(
        clk), .Q(delay_first_two_bytes_out[10]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_9_ ( .D(from_mem_data[1]), .CP(clk), .Q(delay_first_two_bytes_out[9]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_8_ ( .D(from_mem_data[0]), .CP(clk), .Q(delay_first_two_bytes_out[8]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_7_ ( .D(from_mem_data[15]), .CP(
        clk), .Q(delay_first_two_bytes_out[7]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_6_ ( .D(from_mem_data[14]), .CP(
        clk), .Q(delay_first_two_bytes_out[6]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_5_ ( .D(from_mem_data[13]), .CP(
        clk), .Q(delay_first_two_bytes_out[5]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_4_ ( .D(from_mem_data[12]), .CP(
        clk), .Q(delay_first_two_bytes_out[4]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_3_ ( .D(from_mem_data[11]), .CP(
        clk), .Q(delay_first_two_bytes_out[3]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_2_ ( .D(from_mem_data[10]), .CP(
        clk), .Q(delay_first_two_bytes_out[2]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_1_ ( .D(from_mem_data[9]), .CP(clk), .Q(delay_first_two_bytes_out[1]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_0_ ( .D(from_mem_data[8]), .CP(clk), .Q(delay_first_two_bytes_out[0]) );
  DFQD1BWP12T delay_data_in32_reg_31_ ( .D(data_in[31]), .CP(clk), .Q(
        delay_data_in32[31]) );
  DFQD1BWP12T delay_data_in32_reg_30_ ( .D(data_in[30]), .CP(clk), .Q(
        delay_data_in32[30]) );
  DFQD1BWP12T delay_data_in32_reg_29_ ( .D(data_in[29]), .CP(clk), .Q(
        delay_data_in32[29]) );
  DFQD1BWP12T delay_data_in32_reg_28_ ( .D(data_in[28]), .CP(clk), .Q(
        delay_data_in32[28]) );
  DFQD1BWP12T delay_data_in32_reg_27_ ( .D(data_in[27]), .CP(clk), .Q(
        delay_data_in32[27]) );
  DFQD1BWP12T delay_data_in32_reg_26_ ( .D(data_in[26]), .CP(clk), .Q(
        delay_data_in32[26]) );
  DFQD1BWP12T delay_data_in32_reg_25_ ( .D(data_in[25]), .CP(clk), .Q(
        delay_data_in32[25]) );
  DFQD1BWP12T delay_data_in32_reg_24_ ( .D(data_in[24]), .CP(clk), .Q(
        delay_data_in32[24]) );
  DFQD1BWP12T delay_data_in32_reg_23_ ( .D(data_in[23]), .CP(clk), .Q(
        delay_data_in32[23]) );
  DFQD1BWP12T delay_data_in32_reg_22_ ( .D(data_in[22]), .CP(clk), .Q(
        delay_data_in32[22]) );
  DFQD1BWP12T delay_data_in32_reg_21_ ( .D(data_in[21]), .CP(clk), .Q(
        delay_data_in32[21]) );
  DFQD1BWP12T delay_data_in32_reg_20_ ( .D(data_in[20]), .CP(clk), .Q(
        delay_data_in32[20]) );
  DFQD1BWP12T delay_data_in32_reg_19_ ( .D(data_in[19]), .CP(clk), .Q(
        delay_data_in32[19]) );
  DFQD1BWP12T delay_data_in32_reg_18_ ( .D(data_in[18]), .CP(clk), .Q(
        delay_data_in32[18]) );
  DFQD1BWP12T delay_data_in32_reg_17_ ( .D(data_in[17]), .CP(clk), .Q(
        delay_data_in32[17]) );
  DFQD1BWP12T delay_data_in32_reg_16_ ( .D(data_in[16]), .CP(clk), .Q(
        delay_data_in32[16]) );
  DFQD1BWP12T delay_data_in32_reg_15_ ( .D(data_in[15]), .CP(clk), .Q(
        delay_data_in32[15]) );
  DFQD1BWP12T delay_data_in32_reg_14_ ( .D(data_in[14]), .CP(clk), .Q(
        delay_data_in32[14]) );
  DFQD1BWP12T delay_data_in32_reg_13_ ( .D(data_in[13]), .CP(clk), .Q(
        delay_data_in32[13]) );
  DFQD1BWP12T delay_data_in32_reg_12_ ( .D(data_in[12]), .CP(clk), .Q(
        delay_data_in32[12]) );
  DFQD1BWP12T delay_data_in32_reg_11_ ( .D(data_in[11]), .CP(clk), .Q(
        delay_data_in32[11]) );
  DFQD1BWP12T delay_data_in32_reg_10_ ( .D(data_in[10]), .CP(clk), .Q(
        delay_data_in32[10]) );
  DFQD1BWP12T delay_data_in32_reg_9_ ( .D(data_in[9]), .CP(clk), .Q(
        delay_data_in32[9]) );
  DFQD1BWP12T delay_data_in32_reg_8_ ( .D(data_in[8]), .CP(clk), .Q(
        delay_data_in32[8]) );
  DFQD1BWP12T delay_data_in32_reg_7_ ( .D(data_in[7]), .CP(clk), .Q(
        delay_data_in32[7]) );
  DFQD1BWP12T delay_data_in32_reg_6_ ( .D(data_in[6]), .CP(clk), .Q(
        delay_data_in32[6]) );
  DFQD1BWP12T delay_data_in32_reg_5_ ( .D(data_in[5]), .CP(clk), .Q(
        delay_data_in32[5]) );
  DFQD1BWP12T delay_data_in32_reg_4_ ( .D(data_in[4]), .CP(clk), .Q(
        delay_data_in32[4]) );
  DFQD1BWP12T delay_data_in32_reg_3_ ( .D(data_in[3]), .CP(clk), .Q(
        delay_data_in32[3]) );
  DFQD1BWP12T delay_data_in32_reg_2_ ( .D(data_in[2]), .CP(clk), .Q(
        delay_data_in32[2]) );
  DFQD1BWP12T delay_data_in32_reg_1_ ( .D(data_in[1]), .CP(clk), .Q(
        delay_data_in32[1]) );
  DFQD1BWP12T delay_data_in32_reg_0_ ( .D(data_in[0]), .CP(clk), .Q(
        delay_data_in32[0]) );
  DFQD1BWP12T delay_addr_for_adder_reg_11_ ( .D(address[11]), .CP(clk), .Q(
        delay_addr_for_adder[11]) );
  DFQD1BWP12T delay_addr_for_adder_reg_10_ ( .D(address[10]), .CP(clk), .Q(
        delay_addr_for_adder[10]) );
  DFQD1BWP12T delay_addr_for_adder_reg_9_ ( .D(address[9]), .CP(clk), .Q(
        delay_addr_for_adder[9]) );
  DFQD1BWP12T delay_addr_for_adder_reg_8_ ( .D(address[8]), .CP(clk), .Q(
        delay_addr_for_adder[8]) );
  DFQD1BWP12T delay_addr_for_adder_reg_7_ ( .D(address[7]), .CP(clk), .Q(
        delay_addr_for_adder[7]) );
  DFQD1BWP12T delay_addr_for_adder_reg_6_ ( .D(address[6]), .CP(clk), .Q(
        delay_addr_for_adder[6]) );
  DFQD1BWP12T delay_addr_for_adder_reg_5_ ( .D(address[5]), .CP(clk), .Q(
        delay_addr_for_adder[5]) );
  DFQD1BWP12T delay_addr_for_adder_reg_4_ ( .D(address[4]), .CP(clk), .Q(
        delay_addr_for_adder[4]) );
  DFQD1BWP12T delay_addr_for_adder_reg_3_ ( .D(address[3]), .CP(clk), .Q(
        delay_addr_for_adder[3]) );
  DFQD1BWP12T delay_addr_for_adder_reg_2_ ( .D(address[2]), .CP(clk), .Q(
        delay_addr_for_adder[2]) );
  DFQD1BWP12T delay_addr_for_adder_reg_1_ ( .D(address[1]), .CP(clk), .Q(
        delay_addr_for_adder[1]) );
  DFQD1BWP12T delay_addr_for_adder_reg_0_ ( .D(address[0]), .CP(clk), .Q(
        delay_addr_for_adder[0]) );
  DFQD1BWP12T delay_addr_single_reg_11_ ( .D(address[11]), .CP(clk), .Q(
        delay_addr_single[11]) );
  DFQD1BWP12T delay_addr_single_reg_10_ ( .D(address[10]), .CP(clk), .Q(
        delay_addr_single[10]) );
  DFQD1BWP12T delay_addr_single_reg_9_ ( .D(address[9]), .CP(clk), .Q(
        delay_addr_single[9]) );
  DFQD1BWP12T delay_addr_single_reg_8_ ( .D(address[8]), .CP(clk), .Q(
        delay_addr_single[8]) );
  DFQD1BWP12T delay_addr_single_reg_7_ ( .D(address[7]), .CP(clk), .Q(
        delay_addr_single[7]) );
  DFQD1BWP12T delay_addr_single_reg_6_ ( .D(address[6]), .CP(clk), .Q(
        delay_addr_single[6]) );
  DFQD1BWP12T delay_addr_single_reg_5_ ( .D(address[5]), .CP(clk), .Q(
        delay_addr_single[5]) );
  DFQD1BWP12T delay_addr_single_reg_4_ ( .D(address[4]), .CP(clk), .Q(
        delay_addr_single[4]) );
  DFQD1BWP12T delay_addr_single_reg_3_ ( .D(address[3]), .CP(clk), .Q(
        delay_addr_single[3]) );
  DFQD1BWP12T delay_addr_single_reg_2_ ( .D(address[2]), .CP(clk), .Q(
        delay_addr_single[2]) );
  DFQD1BWP12T delay_addr_single_reg_1_ ( .D(address[1]), .CP(clk), .Q(
        delay_addr_single[1]) );
  DFQD1BWP12T delay_addr_single_reg_0_ ( .D(address[0]), .CP(clk), .Q(
        delay_addr_single[0]) );
  DFQD1BWP12T delayed_is_signed_reg ( .D(is_signed), .CP(clk), .Q(
        delayed_is_signed) );
  DFQD1BWP12T fsm_state_reg_3_ ( .D(fsm_N35), .CP(clk), .Q(fsm_state_3_) );
  DFQD1BWP12T fsm_state_reg_2_ ( .D(fsm_N34), .CP(clk), .Q(fsm_state_2_) );
  DFQD1BWP12T fsm_state_reg_1_ ( .D(fsm_N33), .CP(clk), .Q(fsm_state_1_) );
  DFQD1BWP12T fsm_state_reg_0_ ( .D(fsm_N32), .CP(clk), .Q(fsm_state_0_) );
  AOI21D1BWP12T U3 ( .A1(n2), .A2(n22), .B(n14), .ZN(write_ready) );
  ND2D1BWP12T U4 ( .A1(n15), .A2(n9), .ZN(n22) );
  INVD1BWP12T U5 ( .I(fsm_state_0_), .ZN(n9) );
  INVD1BWP12T U6 ( .I(fsm_state_1_), .ZN(n1) );
  INVD1BWP12T U7 ( .I(n105), .ZN(n100) );
  INVD1BWP12T U8 ( .I(n10), .ZN(n113) );
  OAI211D1BWP12T U9 ( .A1(fsm_state_3_), .A2(n22), .B(n124), .C(n111), .ZN(
        output_valid) );
  ND2D1BWP12T U10 ( .A1(n113), .A2(load), .ZN(n13) );
  NR2D1BWP12T U11 ( .A1(fsm_state_2_), .A2(n1), .ZN(n15) );
  INVD1BWP12T U12 ( .I(fsm_state_3_), .ZN(n14) );
  NR3D1BWP12T U13 ( .A1(load), .A2(store_BAR), .A3(n10), .ZN(n16) );
  MAOI22D0BWP12T U14 ( .A1(word_type[0]), .A2(n12), .B1(word_type[0]), .B2(n12), .ZN(n17) );
  OR2XD1BWP12T U15 ( .A1(n112), .A2(n23), .Z(n108) );
  INVD1BWP12T U16 ( .I(from_mem_data[8]), .ZN(n117) );
  INVD1BWP12T U17 ( .I(from_mem_data[9]), .ZN(n118) );
  INVD1BWP12T U18 ( .I(from_mem_data[10]), .ZN(n119) );
  INVD1BWP12T U19 ( .I(from_mem_data[11]), .ZN(n120) );
  INVD1BWP12T U20 ( .I(from_mem_data[12]), .ZN(n121) );
  INVD1BWP12T U21 ( .I(from_mem_data[13]), .ZN(n122) );
  INVD1BWP12T U22 ( .I(from_mem_data[14]), .ZN(n123) );
  INVD1BWP12T U23 ( .I(n127), .ZN(n124) );
  INVD1BWP12T U24 ( .I(from_mem_data[15]), .ZN(n125) );
  AN4XD1BWP12T U25 ( .A1(fsm_state_2_), .A2(n1), .A3(n9), .A4(n14), .Z(n127)
         );
  IOA21D0BWP12T U26 ( .A1(word_type[0]), .A2(word_type[1]), .B(n16), .ZN(n103)
         );
  MAOI22D0BWP12T U27 ( .A1(n16), .A2(n12), .B1(word_type[0]), .B2(n13), .ZN(
        n11) );
  ND4D1BWP12T U28 ( .A1(fsm_state_2_), .A2(fsm_state_0_), .A3(fsm_state_3_), 
        .A4(n1), .ZN(n105) );
  OAI221D0BWP12T U29 ( .A1(fsm_state_1_), .A2(n9), .B1(n1), .B2(fsm_state_0_), 
        .C(fsm_state_2_), .ZN(n2) );
  AO211D0BWP12T U30 ( .A1(fsm_state_0_), .A2(n15), .B(n100), .C(write_ready), 
        .Z(n112) );
  NR3D1BWP12T U31 ( .A1(fsm_state_1_), .A2(fsm_state_2_), .A3(fsm_state_3_), 
        .ZN(n23) );
  AOI22D0BWP12T U32 ( .A1(n127), .A2(delay_first_two_bytes_out[15]), .B1(
        from_mem_data[7]), .B2(n108), .ZN(n4) );
  TPNR3D0BWP12T U33 ( .A1(n23), .A2(n127), .A3(n112), .ZN(n3) );
  OAI211D1BWP12T U34 ( .A1(delayed_is_signed), .A2(n22), .B(n3), .C(n125), 
        .ZN(n109) );
  ND2D0BWP12T U35 ( .A1(n4), .A2(n109), .ZN(data_out[15]) );
  AOI22D0BWP12T U36 ( .A1(n127), .A2(delay_first_two_bytes_out[14]), .B1(
        from_mem_data[6]), .B2(n108), .ZN(n5) );
  CKND2D1BWP12T U37 ( .A1(n5), .A2(n109), .ZN(data_out[14]) );
  AOI22D0BWP12T U38 ( .A1(n127), .A2(delay_first_two_bytes_out[13]), .B1(
        from_mem_data[5]), .B2(n108), .ZN(n6) );
  ND2D0BWP12T U39 ( .A1(n6), .A2(n109), .ZN(data_out[13]) );
  AOI22D0BWP12T U40 ( .A1(n127), .A2(delay_first_two_bytes_out[12]), .B1(
        from_mem_data[4]), .B2(n108), .ZN(n7) );
  CKND2D1BWP12T U41 ( .A1(n7), .A2(n109), .ZN(data_out[12]) );
  AOI22D0BWP12T U42 ( .A1(n127), .A2(delay_first_two_bytes_out[11]), .B1(
        from_mem_data[3]), .B2(n108), .ZN(n8) );
  ND2D0BWP12T U43 ( .A1(n8), .A2(n109), .ZN(data_out[11]) );
  CKND2D1BWP12T U44 ( .A1(fsm_state_0_), .A2(n23), .ZN(n111) );
  TPNR2D0BWP12T U45 ( .A1(output_valid), .A2(n112), .ZN(n53) );
  OAI21D1BWP12T U46 ( .A1(word_type[0]), .A2(word_type[1]), .B(n53), .ZN(n51)
         );
  ND3D0BWP12T U47 ( .A1(fsm_state_0_), .A2(fsm_state_3_), .A3(n15), .ZN(n104)
         );
  OAI211D0BWP12T U48 ( .A1(n51), .A2(store_BAR), .B(n105), .C(n104), .ZN(
        to_mem_write_enable) );
  CKND2D0BWP12T U49 ( .A1(n9), .A2(n23), .ZN(n10) );
  INVD1BWP12T U50 ( .I(word_type[1]), .ZN(n12) );
  AOI21D1BWP12T U51 ( .A1(n11), .A2(n104), .B(reset), .ZN(fsm_N33) );
  OAI32D1BWP12T U52 ( .A1(reset), .A2(n13), .A3(n17), .B1(n103), .B2(reset), 
        .ZN(fsm_N32) );
  ND3D0BWP12T U53 ( .A1(fsm_state_0_), .A2(n15), .A3(n14), .ZN(n19) );
  IND2XD0BWP12T U54 ( .A1(n17), .B1(n16), .ZN(n18) );
  TPAOI31D0BWP12T U55 ( .A1(n105), .A2(n19), .A3(n18), .B(reset), .ZN(fsm_N34)
         );
  OAI32D0BWP12T U56 ( .A1(fsm_state_3_), .A2(fsm_state_1_), .A3(fsm_state_0_), 
        .B1(fsm_state_2_), .B2(fsm_state_3_), .ZN(n52) );
  NR2D0BWP12T U57 ( .A1(write_ready), .A2(n52), .ZN(n42) );
  AN2D1BWP12T U58 ( .A1(n42), .A2(n105), .Z(n99) );
  AOI21D1BWP12T U59 ( .A1(n42), .A2(n104), .B(n53), .ZN(n94) );
  INR2D1BWP12T U60 ( .A1(n94), .B1(n99), .ZN(n98) );
  AOI22D1BWP12T U61 ( .A1(n99), .A2(from_mem_data[7]), .B1(n98), .B2(
        delay_data_in32[15]), .ZN(n21) );
  AOI22D1BWP12T U62 ( .A1(n100), .A2(delay_data_in32[31]), .B1(n113), .B2(
        data_in[15]), .ZN(n20) );
  ND2D1BWP12T U63 ( .A1(n21), .A2(n20), .ZN(to_mem_data[7]) );
  CKND0BWP12T U64 ( .I(n22), .ZN(n114) );
  OR4D1BWP12T U65 ( .A1(write_ready), .A2(n114), .A3(n23), .A4(n127), .Z(n77)
         );
  AOI22D0BWP12T U66 ( .A1(n99), .A2(delay_addr_single[8]), .B1(address[8]), 
        .B2(n77), .ZN(n25) );
  AN2D1BWP12T U67 ( .A1(delay_addr_for_adder[1]), .A2(delay_addr_for_adder[0]), 
        .Z(n74) );
  ND2D1BWP12T U68 ( .A1(n74), .A2(delay_addr_for_adder[2]), .ZN(n68) );
  INVD1BWP12T U69 ( .I(delay_addr_for_adder[3]), .ZN(n48) );
  NR2D1BWP12T U70 ( .A1(n68), .A2(n48), .ZN(n47) );
  ND2D1BWP12T U71 ( .A1(n47), .A2(delay_addr_for_adder[4]), .ZN(n33) );
  INVD1BWP12T U72 ( .I(delay_addr_for_adder[5]), .ZN(n30) );
  NR2D1BWP12T U73 ( .A1(n33), .A2(n30), .ZN(n54) );
  ND2D1BWP12T U74 ( .A1(n54), .A2(delay_addr_for_adder[6]), .ZN(n59) );
  INVD1BWP12T U75 ( .I(delay_addr_for_adder[7]), .ZN(n58) );
  NR2D1BWP12T U76 ( .A1(n59), .A2(n58), .ZN(n57) );
  NR2D1BWP12T U77 ( .A1(n77), .A2(n99), .ZN(n75) );
  ND2D1BWP12T U78 ( .A1(n57), .A2(delay_addr_for_adder[8]), .ZN(n27) );
  OAI211D1BWP12T U79 ( .A1(n57), .A2(delay_addr_for_adder[8]), .B(n75), .C(n27), .ZN(n24) );
  ND2D1BWP12T U80 ( .A1(n25), .A2(n24), .ZN(to_mem_address[8]) );
  AOI22D0BWP12T U81 ( .A1(n99), .A2(delay_addr_single[9]), .B1(address[9]), 
        .B2(n77), .ZN(n29) );
  INVD1BWP12T U82 ( .I(delay_addr_for_adder[9]), .ZN(n26) );
  NR2D1BWP12T U83 ( .A1(n27), .A2(n26), .ZN(n63) );
  INVD1BWP12T U84 ( .I(n75), .ZN(n72) );
  AO211D1BWP12T U85 ( .A1(n27), .A2(n26), .B(n63), .C(n72), .Z(n28) );
  ND2D1BWP12T U86 ( .A1(n29), .A2(n28), .ZN(to_mem_address[9]) );
  AOI22D1BWP12T U87 ( .A1(n99), .A2(delay_addr_single[5]), .B1(address[5]), 
        .B2(n77), .ZN(n32) );
  AO211D1BWP12T U88 ( .A1(n33), .A2(n30), .B(n54), .C(n72), .Z(n31) );
  ND2D1BWP12T U89 ( .A1(n32), .A2(n31), .ZN(to_mem_address[5]) );
  AOI22D1BWP12T U90 ( .A1(n99), .A2(delay_addr_single[4]), .B1(address[4]), 
        .B2(n77), .ZN(n35) );
  OAI211D1BWP12T U91 ( .A1(n47), .A2(delay_addr_for_adder[4]), .B(n75), .C(n33), .ZN(n34) );
  ND2D1BWP12T U92 ( .A1(n35), .A2(n34), .ZN(to_mem_address[4]) );
  ND2D1BWP12T U93 ( .A1(n63), .A2(delay_addr_for_adder[10]), .ZN(n62) );
  MAOI22D0BWP12T U94 ( .A1(delay_addr_for_adder[11]), .A2(n62), .B1(
        delay_addr_for_adder[11]), .B2(n62), .ZN(n37) );
  AOI22D0BWP12T U95 ( .A1(n99), .A2(delay_addr_single[11]), .B1(address[11]), 
        .B2(n77), .ZN(n36) );
  OAI21D1BWP12T U96 ( .A1(n72), .A2(n37), .B(n36), .ZN(to_mem_address[11]) );
  AOI22D1BWP12T U97 ( .A1(n99), .A2(from_mem_data[0]), .B1(n98), .B2(
        delay_data_in32[8]), .ZN(n39) );
  AOI22D1BWP12T U98 ( .A1(n100), .A2(delay_data_in32[24]), .B1(n113), .B2(
        data_in[8]), .ZN(n38) );
  ND2D1BWP12T U99 ( .A1(n39), .A2(n38), .ZN(to_mem_data[0]) );
  AOI22D1BWP12T U100 ( .A1(n99), .A2(from_mem_data[2]), .B1(n98), .B2(
        delay_data_in32[10]), .ZN(n41) );
  AOI22D1BWP12T U101 ( .A1(n100), .A2(delay_data_in32[26]), .B1(n113), .B2(
        data_in[10]), .ZN(n40) );
  ND2D1BWP12T U102 ( .A1(n41), .A2(n40), .ZN(to_mem_data[2]) );
  AOI22D1BWP12T U103 ( .A1(n113), .A2(data_in[7]), .B1(n94), .B2(
        delay_data_in32[7]), .ZN(n44) );
  AN2D1BWP12T U104 ( .A1(n42), .A2(n53), .Z(n95) );
  AOI22D1BWP12T U105 ( .A1(n100), .A2(delay_data_in32[23]), .B1(n95), .B2(
        data_in[23]), .ZN(n43) );
  ND2D1BWP12T U106 ( .A1(n44), .A2(n43), .ZN(to_mem_data[15]) );
  AOI22D1BWP12T U107 ( .A1(n113), .A2(data_in[6]), .B1(n94), .B2(
        delay_data_in32[6]), .ZN(n46) );
  AOI22D1BWP12T U108 ( .A1(n100), .A2(delay_data_in32[22]), .B1(n95), .B2(
        data_in[22]), .ZN(n45) );
  ND2D1BWP12T U109 ( .A1(n46), .A2(n45), .ZN(to_mem_data[14]) );
  AOI22D1BWP12T U110 ( .A1(n99), .A2(delay_addr_single[3]), .B1(address[3]), 
        .B2(n77), .ZN(n50) );
  AO211D1BWP12T U111 ( .A1(n68), .A2(n48), .B(n47), .C(n72), .Z(n49) );
  ND2D1BWP12T U112 ( .A1(n50), .A2(n49), .ZN(to_mem_address[3]) );
  OA22D1BWP12T U113 ( .A1(n53), .A2(n52), .B1(load), .B2(n51), .Z(
        to_mem_read_enable) );
  AOI22D1BWP12T U114 ( .A1(n99), .A2(delay_addr_single[6]), .B1(address[6]), 
        .B2(n77), .ZN(n56) );
  OAI211D1BWP12T U115 ( .A1(n54), .A2(delay_addr_for_adder[6]), .B(n75), .C(
        n59), .ZN(n55) );
  ND2D1BWP12T U116 ( .A1(n56), .A2(n55), .ZN(to_mem_address[6]) );
  AOI22D0BWP12T U117 ( .A1(n99), .A2(delay_addr_single[7]), .B1(address[7]), 
        .B2(n77), .ZN(n61) );
  AO211D1BWP12T U118 ( .A1(n59), .A2(n58), .B(n57), .C(n72), .Z(n60) );
  ND2D1BWP12T U119 ( .A1(n61), .A2(n60), .ZN(to_mem_address[7]) );
  AOI22D0BWP12T U120 ( .A1(n99), .A2(delay_addr_single[10]), .B1(address[10]), 
        .B2(n77), .ZN(n65) );
  OAI211D1BWP12T U121 ( .A1(n63), .A2(delay_addr_for_adder[10]), .B(n75), .C(
        n62), .ZN(n64) );
  ND2D1BWP12T U122 ( .A1(n65), .A2(n64), .ZN(to_mem_address[10]) );
  AOI22D1BWP12T U123 ( .A1(n99), .A2(from_mem_data[1]), .B1(n98), .B2(
        delay_data_in32[9]), .ZN(n67) );
  AOI22D1BWP12T U124 ( .A1(n100), .A2(delay_data_in32[25]), .B1(n113), .B2(
        data_in[9]), .ZN(n66) );
  ND2D1BWP12T U125 ( .A1(n67), .A2(n66), .ZN(to_mem_data[1]) );
  AOI22D1BWP12T U126 ( .A1(n99), .A2(delay_addr_single[2]), .B1(address[2]), 
        .B2(n77), .ZN(n70) );
  OAI211D1BWP12T U127 ( .A1(n74), .A2(delay_addr_for_adder[2]), .B(n75), .C(
        n68), .ZN(n69) );
  ND2D1BWP12T U128 ( .A1(n70), .A2(n69), .ZN(to_mem_address[2]) );
  NR2D1BWP12T U129 ( .A1(delay_addr_for_adder[0]), .A2(delay_addr_for_adder[1]), .ZN(n73) );
  AOI22D1BWP12T U130 ( .A1(n99), .A2(delay_addr_single[1]), .B1(address[1]), 
        .B2(n77), .ZN(n71) );
  OAI31D1BWP12T U131 ( .A1(n74), .A2(n73), .A3(n72), .B(n71), .ZN(
        to_mem_address[1]) );
  INVD1BWP12T U132 ( .I(delay_addr_for_adder[0]), .ZN(n76) );
  AO222D1BWP12T U133 ( .A1(n77), .A2(address[0]), .B1(n76), .B2(n75), .C1(
        delay_addr_single[0]), .C2(n99), .Z(to_mem_address[0]) );
  AOI22D1BWP12T U134 ( .A1(n99), .A2(from_mem_data[3]), .B1(n98), .B2(
        delay_data_in32[11]), .ZN(n79) );
  AOI22D1BWP12T U135 ( .A1(n100), .A2(delay_data_in32[27]), .B1(n113), .B2(
        data_in[11]), .ZN(n78) );
  ND2D1BWP12T U136 ( .A1(n79), .A2(n78), .ZN(to_mem_data[3]) );
  AOI22D1BWP12T U137 ( .A1(n99), .A2(from_mem_data[5]), .B1(n98), .B2(
        delay_data_in32[13]), .ZN(n81) );
  AOI22D1BWP12T U138 ( .A1(n100), .A2(delay_data_in32[29]), .B1(n113), .B2(
        data_in[13]), .ZN(n80) );
  ND2D1BWP12T U139 ( .A1(n81), .A2(n80), .ZN(to_mem_data[5]) );
  AOI22D1BWP12T U140 ( .A1(n99), .A2(from_mem_data[4]), .B1(n98), .B2(
        delay_data_in32[12]), .ZN(n83) );
  AOI22D1BWP12T U141 ( .A1(n100), .A2(delay_data_in32[28]), .B1(n113), .B2(
        data_in[12]), .ZN(n82) );
  ND2D1BWP12T U142 ( .A1(n83), .A2(n82), .ZN(to_mem_data[4]) );
  AOI22D1BWP12T U143 ( .A1(n113), .A2(data_in[5]), .B1(n94), .B2(
        delay_data_in32[5]), .ZN(n85) );
  AOI22D1BWP12T U144 ( .A1(n100), .A2(delay_data_in32[21]), .B1(n95), .B2(
        data_in[21]), .ZN(n84) );
  ND2D1BWP12T U145 ( .A1(n85), .A2(n84), .ZN(to_mem_data[13]) );
  AOI22D1BWP12T U146 ( .A1(n113), .A2(data_in[1]), .B1(n94), .B2(
        delay_data_in32[1]), .ZN(n87) );
  AOI22D1BWP12T U147 ( .A1(n100), .A2(delay_data_in32[17]), .B1(n95), .B2(
        data_in[17]), .ZN(n86) );
  ND2D1BWP12T U148 ( .A1(n87), .A2(n86), .ZN(to_mem_data[9]) );
  AOI22D1BWP12T U149 ( .A1(n113), .A2(data_in[3]), .B1(n94), .B2(
        delay_data_in32[3]), .ZN(n89) );
  AOI22D1BWP12T U150 ( .A1(n100), .A2(delay_data_in32[19]), .B1(n95), .B2(
        data_in[19]), .ZN(n88) );
  ND2D1BWP12T U151 ( .A1(n89), .A2(n88), .ZN(to_mem_data[11]) );
  AOI22D1BWP12T U152 ( .A1(n113), .A2(data_in[4]), .B1(n94), .B2(
        delay_data_in32[4]), .ZN(n91) );
  AOI22D1BWP12T U153 ( .A1(n100), .A2(delay_data_in32[20]), .B1(n95), .B2(
        data_in[20]), .ZN(n90) );
  ND2D1BWP12T U154 ( .A1(n91), .A2(n90), .ZN(to_mem_data[12]) );
  AOI22D1BWP12T U155 ( .A1(n113), .A2(data_in[2]), .B1(n94), .B2(
        delay_data_in32[2]), .ZN(n93) );
  AOI22D1BWP12T U156 ( .A1(n100), .A2(delay_data_in32[18]), .B1(n95), .B2(
        data_in[18]), .ZN(n92) );
  ND2D1BWP12T U157 ( .A1(n93), .A2(n92), .ZN(to_mem_data[10]) );
  AOI22D1BWP12T U158 ( .A1(n113), .A2(data_in[0]), .B1(n94), .B2(
        delay_data_in32[0]), .ZN(n97) );
  AOI22D1BWP12T U159 ( .A1(n100), .A2(delay_data_in32[16]), .B1(n95), .B2(
        data_in[16]), .ZN(n96) );
  ND2D1BWP12T U160 ( .A1(n97), .A2(n96), .ZN(to_mem_data[8]) );
  AOI22D1BWP12T U161 ( .A1(n99), .A2(from_mem_data[6]), .B1(n98), .B2(
        delay_data_in32[14]), .ZN(n102) );
  AOI22D1BWP12T U162 ( .A1(n100), .A2(delay_data_in32[30]), .B1(n113), .B2(
        data_in[14]), .ZN(n101) );
  ND2D1BWP12T U163 ( .A1(n102), .A2(n101), .ZN(to_mem_data[6]) );
  AOI31D0BWP12T U164 ( .A1(n105), .A2(n104), .A3(n103), .B(reset), .ZN(fsm_N35) );
  MAOI22D0BWP12T U165 ( .A1(n124), .A2(n117), .B1(n124), .B2(
        delay_first_two_bytes_out[0]), .ZN(data_out[0]) );
  MAOI22D0BWP12T U166 ( .A1(n124), .A2(n118), .B1(n124), .B2(
        delay_first_two_bytes_out[1]), .ZN(data_out[1]) );
  MAOI22D0BWP12T U167 ( .A1(n124), .A2(n119), .B1(n124), .B2(
        delay_first_two_bytes_out[2]), .ZN(data_out[2]) );
  MAOI22D0BWP12T U168 ( .A1(n124), .A2(n120), .B1(n124), .B2(
        delay_first_two_bytes_out[3]), .ZN(data_out[3]) );
  MAOI22D0BWP12T U169 ( .A1(n124), .A2(n121), .B1(n124), .B2(
        delay_first_two_bytes_out[4]), .ZN(data_out[4]) );
  MAOI22D0BWP12T U170 ( .A1(n124), .A2(n122), .B1(n124), .B2(
        delay_first_two_bytes_out[5]), .ZN(data_out[5]) );
  MAOI22D0BWP12T U171 ( .A1(n124), .A2(n123), .B1(n124), .B2(
        delay_first_two_bytes_out[6]), .ZN(data_out[6]) );
  MAOI22D0BWP12T U172 ( .A1(n124), .A2(n125), .B1(n124), .B2(
        delay_first_two_bytes_out[7]), .ZN(data_out[7]) );
  AOI22D0BWP12T U173 ( .A1(n127), .A2(delay_first_two_bytes_out[8]), .B1(
        from_mem_data[0]), .B2(n108), .ZN(n106) );
  CKND2D0BWP12T U174 ( .A1(n106), .A2(n109), .ZN(data_out[8]) );
  AOI22D0BWP12T U175 ( .A1(n127), .A2(delay_first_two_bytes_out[9]), .B1(
        from_mem_data[1]), .B2(n108), .ZN(n107) );
  CKND2D0BWP12T U176 ( .A1(n107), .A2(n109), .ZN(data_out[9]) );
  AOI22D0BWP12T U177 ( .A1(n127), .A2(delay_first_two_bytes_out[10]), .B1(
        from_mem_data[2]), .B2(n108), .ZN(n110) );
  CKND2D0BWP12T U178 ( .A1(n110), .A2(n109), .ZN(data_out[10]) );
  IND3D1BWP12T U179 ( .A1(n111), .B1(from_mem_data[7]), .B2(delayed_is_signed), 
        .ZN(n116) );
  AOI211D0BWP12T U180 ( .A1(n114), .A2(delayed_is_signed), .B(n113), .C(n112), 
        .ZN(n115) );
  MUX2D1BWP12T U181 ( .I0(n125), .I1(n116), .S(n115), .Z(n126) );
  OAI21D0BWP12T U182 ( .A1(n124), .A2(n117), .B(n126), .ZN(data_out[16]) );
  OAI21D0BWP12T U183 ( .A1(n124), .A2(n118), .B(n126), .ZN(data_out[17]) );
  OAI21D0BWP12T U184 ( .A1(n124), .A2(n119), .B(n126), .ZN(data_out[18]) );
  OAI21D0BWP12T U185 ( .A1(n124), .A2(n120), .B(n126), .ZN(data_out[19]) );
  OAI21D0BWP12T U186 ( .A1(n124), .A2(n121), .B(n126), .ZN(data_out[20]) );
  OAI21D0BWP12T U187 ( .A1(n124), .A2(n122), .B(n126), .ZN(data_out[21]) );
  OAI21D0BWP12T U188 ( .A1(n124), .A2(n123), .B(n126), .ZN(data_out[22]) );
  OAI21D0BWP12T U189 ( .A1(n125), .A2(n124), .B(n126), .ZN(data_out[23]) );
  IOA21D0BWP12T U190 ( .A1(from_mem_data[0]), .A2(n127), .B(n126), .ZN(
        data_out[24]) );
  IOA21D0BWP12T U191 ( .A1(from_mem_data[1]), .A2(n127), .B(n126), .ZN(
        data_out[25]) );
  IOA21D0BWP12T U192 ( .A1(from_mem_data[2]), .A2(n127), .B(n126), .ZN(
        data_out[26]) );
  IOA21D0BWP12T U193 ( .A1(from_mem_data[3]), .A2(n127), .B(n126), .ZN(
        data_out[27]) );
  IOA21D0BWP12T U194 ( .A1(from_mem_data[4]), .A2(n127), .B(n126), .ZN(
        data_out[28]) );
  IOA21D0BWP12T U195 ( .A1(from_mem_data[5]), .A2(n127), .B(n126), .ZN(
        data_out[29]) );
  IOA21D0BWP12T U196 ( .A1(from_mem_data[6]), .A2(n127), .B(n126), .ZN(
        data_out[30]) );
  IOA21D0BWP12T U197 ( .A1(from_mem_data[7]), .A2(n127), .B(n126), .ZN(
        data_out[31]) );
endmodule


module Instruction_Fetch ( clk, reset, stall_decoder_in, memory_output_valid, 
        current_pc_in, instruction_in, memory_load_request, 
        incremented_pc_write_enable, instruction_valid, memory_address, 
        incremented_pc_out, instruction_out, finish_out );
  input [31:0] current_pc_in;
  input [15:0] instruction_in;
  output [11:0] memory_address;
  output [31:0] incremented_pc_out;
  output [15:0] instruction_out;
  input clk, reset, stall_decoder_in, memory_output_valid;
  output memory_load_request, incremented_pc_write_enable, instruction_valid,
         finish_out;
  wire   currentState_0_, first_instruction_fetched, N79, N80, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, n37,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98;
  wire   [15:0] fetched_instruction_reg;
  tri   clk;
  tri   reset;
  tri   [31:0] current_pc_in;
  tri   [15:0] instruction_in;
  tri   incremented_pc_write_enable;
  tri   [31:0] incremented_pc_out;

  DFQD1BWP12T first_instruction_fetched_reg ( .D(n37), .CP(clk), .Q(
        first_instruction_fetched) );
  DFQD1BWP12T currentState_reg_1_ ( .D(N80), .CP(clk), .Q(memory_load_request)
         );
  DFQD1BWP12T currentState_reg_0_ ( .D(N79), .CP(clk), .Q(currentState_0_) );
  DFQD1BWP12T fetched_instruction_reg_reg_0_ ( .D(N83), .CP(clk), .Q(
        fetched_instruction_reg[0]) );
  DFQD1BWP12T fetched_instruction_reg_reg_1_ ( .D(N84), .CP(clk), .Q(
        fetched_instruction_reg[1]) );
  DFQD1BWP12T fetched_instruction_reg_reg_2_ ( .D(N85), .CP(clk), .Q(
        fetched_instruction_reg[2]) );
  DFQD1BWP12T fetched_instruction_reg_reg_3_ ( .D(N86), .CP(clk), .Q(
        fetched_instruction_reg[3]) );
  DFQD1BWP12T fetched_instruction_reg_reg_4_ ( .D(N87), .CP(clk), .Q(
        fetched_instruction_reg[4]) );
  DFQD1BWP12T fetched_instruction_reg_reg_5_ ( .D(N88), .CP(clk), .Q(
        fetched_instruction_reg[5]) );
  DFQD1BWP12T fetched_instruction_reg_reg_6_ ( .D(N89), .CP(clk), .Q(
        fetched_instruction_reg[6]) );
  DFQD1BWP12T fetched_instruction_reg_reg_7_ ( .D(N90), .CP(clk), .Q(
        fetched_instruction_reg[7]) );
  DFQD1BWP12T fetched_instruction_reg_reg_8_ ( .D(N91), .CP(clk), .Q(
        fetched_instruction_reg[8]) );
  DFQD1BWP12T fetched_instruction_reg_reg_9_ ( .D(N92), .CP(clk), .Q(
        fetched_instruction_reg[9]) );
  DFQD1BWP12T fetched_instruction_reg_reg_10_ ( .D(N93), .CP(clk), .Q(
        fetched_instruction_reg[10]) );
  DFQD1BWP12T fetched_instruction_reg_reg_11_ ( .D(N94), .CP(clk), .Q(
        fetched_instruction_reg[11]) );
  DFQD1BWP12T fetched_instruction_reg_reg_12_ ( .D(N95), .CP(clk), .Q(
        fetched_instruction_reg[12]) );
  DFQD1BWP12T fetched_instruction_reg_reg_13_ ( .D(N96), .CP(clk), .Q(
        fetched_instruction_reg[13]) );
  DFQD1BWP12T fetched_instruction_reg_reg_14_ ( .D(N97), .CP(clk), .Q(
        fetched_instruction_reg[14]) );
  DFQD1BWP12T fetched_instruction_reg_reg_15_ ( .D(N98), .CP(clk), .Q(
        fetched_instruction_reg[15]) );
  NR2D1BWP12T U3 ( .A1(n89), .A2(n45), .ZN(n43) );
  ND2D1BWP12T U4 ( .A1(n47), .A2(n19), .ZN(instruction_out[13]) );
  ND2D1BWP12T U5 ( .A1(current_pc_in[1]), .A2(current_pc_in[2]), .ZN(n49) );
  INVD1BWP12T U6 ( .I(currentState_0_), .ZN(n1) );
  OR2XD1BWP12T U7 ( .A1(current_pc_in[1]), .A2(current_pc_in[2]), .Z(n40) );
  NR2D1BWP12T U8 ( .A1(current_pc_in[3]), .A2(n40), .ZN(n38) );
  OAI21D1BWP12T U9 ( .A1(n38), .A2(n52), .B(n42), .ZN(n36) );
  ND2D1BWP12T U10 ( .A1(n38), .A2(n52), .ZN(n42) );
  NR2D1BWP12T U11 ( .A1(current_pc_in[5]), .A2(n42), .ZN(n41) );
  ND2D1BWP12T U12 ( .A1(n41), .A2(n55), .ZN(n35) );
  NR2D1BWP12T U13 ( .A1(current_pc_in[7]), .A2(n35), .ZN(n33) );
  ND2D1BWP12T U14 ( .A1(n33), .A2(n58), .ZN(n32) );
  MAOI22D0BWP12T U15 ( .A1(current_pc_in[9]), .A2(n32), .B1(current_pc_in[9]), 
        .B2(n32), .ZN(n31) );
  MOAI22D0BWP12T U16 ( .A1(current_pc_in[10]), .A2(n20), .B1(current_pc_in[10]), .B2(n20), .ZN(n28) );
  ND2D1BWP12T U17 ( .A1(n20), .A2(n61), .ZN(n26) );
  ND2D1BWP12T U18 ( .A1(n47), .A2(n17), .ZN(instruction_out[10]) );
  ND2D1BWP12T U19 ( .A1(n47), .A2(n25), .ZN(instruction_out[12]) );
  ND2D1BWP12T U20 ( .A1(n47), .A2(n24), .ZN(instruction_out[11]) );
  ND2D1BWP12T U21 ( .A1(n47), .A2(n18), .ZN(instruction_out[8]) );
  NR2D1BWP12T U22 ( .A1(n1), .A2(memory_load_request), .ZN(n45) );
  ND2D1BWP12T U23 ( .A1(n89), .A2(memory_output_valid), .ZN(n96) );
  INVD1BWP12T U24 ( .I(current_pc_in[4]), .ZN(n52) );
  INVD1BWP12T U25 ( .I(current_pc_in[6]), .ZN(n55) );
  INVD1BWP12T U26 ( .I(current_pc_in[10]), .ZN(n61) );
  INVD1BWP12T U27 ( .I(current_pc_in[12]), .ZN(n64) );
  INVD1BWP12T U28 ( .I(current_pc_in[16]), .ZN(n70) );
  INVD1BWP12T U29 ( .I(n94), .ZN(n89) );
  ND2D1BWP12T U30 ( .A1(memory_load_request), .A2(n1), .ZN(n94) );
  AOI21D1BWP12T U31 ( .A1(current_pc_in[3]), .A2(n40), .B(n38), .ZN(n39) );
  INVD1BWP12T U32 ( .I(n96), .ZN(incremented_pc_write_enable) );
  AOI21D1BWP12T U33 ( .A1(current_pc_in[7]), .A2(n35), .B(n33), .ZN(n34) );
  ND2D1BWP12T U34 ( .A1(n47), .A2(n23), .ZN(instruction_out[9]) );
  AOI21D1BWP12T U35 ( .A1(current_pc_in[5]), .A2(n42), .B(n41), .ZN(n44) );
  NR2D1BWP12T U36 ( .A1(current_pc_in[11]), .A2(n26), .ZN(n21) );
  MAOI22D0BWP12T U37 ( .A1(n21), .A2(n64), .B1(n21), .B2(n64), .ZN(n22) );
  MAOI22D0BWP12T U38 ( .A1(current_pc_in[11]), .A2(n26), .B1(current_pc_in[11]), .B2(n26), .ZN(n27) );
  IIND4D1BWP12T U39 ( .A1(current_pc_in[2]), .A2(current_pc_in[3]), .B1(
        current_pc_in[1]), .B2(n70), .ZN(n7) );
  NR4D0BWP12T U40 ( .A1(current_pc_in[22]), .A2(current_pc_in[21]), .A3(
        current_pc_in[20]), .A4(current_pc_in[19]), .ZN(n2) );
  NR4D0BWP12T U41 ( .A1(current_pc_in[26]), .A2(current_pc_in[25]), .A3(
        current_pc_in[24]), .A4(current_pc_in[23]), .ZN(n3) );
  NR4D0BWP12T U42 ( .A1(current_pc_in[30]), .A2(current_pc_in[29]), .A3(
        current_pc_in[28]), .A4(current_pc_in[27]), .ZN(n4) );
  NR4D0BWP12T U43 ( .A1(current_pc_in[31]), .A2(current_pc_in[15]), .A3(
        current_pc_in[14]), .A4(current_pc_in[13]), .ZN(n5) );
  NR2D1BWP12T U44 ( .A1(current_pc_in[11]), .A2(n12), .ZN(n15) );
  ND4D1BWP12T U45 ( .A1(n5), .A2(n4), .A3(n3), .A4(n2), .ZN(n6) );
  ND2D1BWP12T U46 ( .A1(n64), .A2(n11), .ZN(n12) );
  OR3XD1BWP12T U47 ( .A1(n6), .A2(current_pc_in[5]), .A3(current_pc_in[7]), 
        .Z(n10) );
  IINR4D0BWP12T U48 ( .A1(n31), .A2(n28), .B1(n10), .B2(n9), .ZN(n11) );
  INVD1BWP12T U49 ( .I(current_pc_in[8]), .ZN(n58) );
  CKND0BWP12T U50 ( .I(n45), .ZN(n13) );
  IAO21D1BWP12T U51 ( .A1(n94), .A2(memory_output_valid), .B(n43), .ZN(n47) );
  NR2D1BWP12T U52 ( .A1(current_pc_in[9]), .A2(n32), .ZN(n20) );
  NR4D0BWP12T U53 ( .A1(current_pc_in[18]), .A2(current_pc_in[17]), .A3(n36), 
        .A4(n7), .ZN(n8) );
  ND3D0BWP12T U54 ( .A1(n55), .A2(n58), .A3(n8), .ZN(n9) );
  ND3D0BWP12T U55 ( .A1(n89), .A2(first_instruction_fetched), .A3(n15), .ZN(
        n97) );
  OA211D0BWP12T U56 ( .A1(stall_decoder_in), .A2(n13), .B(n47), .C(n97), .Z(
        n14) );
  NR2D1BWP12T U57 ( .A1(reset), .A2(n14), .ZN(N80) );
  AOI21D0BWP12T U58 ( .A1(memory_output_valid), .A2(n15), .B(
        first_instruction_fetched), .ZN(n16) );
  NR2D1BWP12T U59 ( .A1(reset), .A2(n16), .ZN(n37) );
  AOI22D0BWP12T U60 ( .A1(n89), .A2(instruction_in[10]), .B1(n45), .B2(
        fetched_instruction_reg[10]), .ZN(n17) );
  AOI22D0BWP12T U61 ( .A1(n89), .A2(instruction_in[8]), .B1(n45), .B2(
        fetched_instruction_reg[8]), .ZN(n18) );
  AOI22D0BWP12T U62 ( .A1(n89), .A2(instruction_in[13]), .B1(n45), .B2(
        fetched_instruction_reg[13]), .ZN(n19) );
  NR2D0BWP12T U63 ( .A1(n43), .A2(n22), .ZN(memory_address[11]) );
  AOI22D0BWP12T U64 ( .A1(n89), .A2(instruction_in[9]), .B1(n45), .B2(
        fetched_instruction_reg[9]), .ZN(n23) );
  AOI22D0BWP12T U65 ( .A1(n89), .A2(instruction_in[11]), .B1(n45), .B2(
        fetched_instruction_reg[11]), .ZN(n24) );
  AOI22D1BWP12T U66 ( .A1(n89), .A2(instruction_in[12]), .B1(n45), .B2(
        fetched_instruction_reg[12]), .ZN(n25) );
  NR2XD0BWP12T U67 ( .A1(reset), .A2(n96), .ZN(n30) );
  NR2D1BWP12T U68 ( .A1(reset), .A2(incremented_pc_write_enable), .ZN(n29) );
  AO22XD1BWP12T U69 ( .A1(n30), .A2(instruction_in[14]), .B1(n29), .B2(
        fetched_instruction_reg[14]), .Z(N97) );
  NR2D0BWP12T U70 ( .A1(n27), .A2(n43), .ZN(memory_address[10]) );
  AO22D1BWP12T U71 ( .A1(incremented_pc_write_enable), .A2(instruction_in[14]), 
        .B1(n45), .B2(fetched_instruction_reg[14]), .Z(instruction_out[14]) );
  AO22XD1BWP12T U72 ( .A1(n30), .A2(instruction_in[0]), .B1(n29), .B2(
        fetched_instruction_reg[0]), .Z(N83) );
  AO22XD1BWP12T U73 ( .A1(n30), .A2(instruction_in[1]), .B1(n29), .B2(
        fetched_instruction_reg[1]), .Z(N84) );
  AO22XD1BWP12T U74 ( .A1(n30), .A2(instruction_in[2]), .B1(n29), .B2(
        fetched_instruction_reg[2]), .Z(N85) );
  AO22XD1BWP12T U75 ( .A1(n30), .A2(instruction_in[6]), .B1(n29), .B2(
        fetched_instruction_reg[6]), .Z(N89) );
  NR2D0BWP12T U76 ( .A1(n28), .A2(n43), .ZN(memory_address[9]) );
  AO22XD1BWP12T U77 ( .A1(n30), .A2(instruction_in[4]), .B1(n29), .B2(
        fetched_instruction_reg[4]), .Z(N87) );
  AO22XD1BWP12T U78 ( .A1(n30), .A2(instruction_in[7]), .B1(n29), .B2(
        fetched_instruction_reg[7]), .Z(N90) );
  AO22XD1BWP12T U79 ( .A1(n30), .A2(instruction_in[3]), .B1(n29), .B2(
        fetched_instruction_reg[3]), .Z(N86) );
  AO22XD1BWP12T U80 ( .A1(n30), .A2(instruction_in[5]), .B1(n29), .B2(
        fetched_instruction_reg[5]), .Z(N88) );
  AO22XD1BWP12T U81 ( .A1(incremented_pc_write_enable), .A2(instruction_in[1]), 
        .B1(n45), .B2(fetched_instruction_reg[1]), .Z(instruction_out[1]) );
  AO22D1BWP12T U82 ( .A1(incremented_pc_write_enable), .A2(instruction_in[7]), 
        .B1(n45), .B2(fetched_instruction_reg[7]), .Z(instruction_out[7]) );
  AO22XD1BWP12T U83 ( .A1(incremented_pc_write_enable), .A2(instruction_in[3]), 
        .B1(n45), .B2(fetched_instruction_reg[3]), .Z(instruction_out[3]) );
  NR2D0BWP12T U84 ( .A1(n31), .A2(n43), .ZN(memory_address[8]) );
  AO22XD1BWP12T U85 ( .A1(incremented_pc_write_enable), .A2(instruction_in[4]), 
        .B1(n45), .B2(fetched_instruction_reg[4]), .Z(instruction_out[4]) );
  AO22XD1BWP12T U86 ( .A1(incremented_pc_write_enable), .A2(instruction_in[5]), 
        .B1(n45), .B2(fetched_instruction_reg[5]), .Z(instruction_out[5]) );
  AO22XD1BWP12T U87 ( .A1(incremented_pc_write_enable), .A2(instruction_in[6]), 
        .B1(n45), .B2(fetched_instruction_reg[6]), .Z(instruction_out[6]) );
  CKBD1BWP12T U88 ( .I(incremented_pc_write_enable), .Z(instruction_valid) );
  AO22XD1BWP12T U89 ( .A1(incremented_pc_write_enable), .A2(instruction_in[2]), 
        .B1(n45), .B2(fetched_instruction_reg[2]), .Z(instruction_out[2]) );
  AO22XD1BWP12T U90 ( .A1(incremented_pc_write_enable), .A2(instruction_in[0]), 
        .B1(n45), .B2(fetched_instruction_reg[0]), .Z(instruction_out[0]) );
  OAI32D0BWP12T U91 ( .A1(n43), .A2(n33), .A3(n58), .B1(n32), .B2(n43), .ZN(
        memory_address[7]) );
  NR2D0BWP12T U92 ( .A1(n34), .A2(n43), .ZN(memory_address[6]) );
  OAI32D0BWP12T U93 ( .A1(n43), .A2(n41), .A3(n55), .B1(n35), .B2(n43), .ZN(
        memory_address[5]) );
  INR2D0BWP12T U94 ( .A1(n36), .B1(n43), .ZN(memory_address[3]) );
  NR2D0BWP12T U95 ( .A1(current_pc_in[1]), .A2(n43), .ZN(memory_address[0]) );
  NR2D0BWP12T U96 ( .A1(n39), .A2(n43), .ZN(memory_address[2]) );
  CKND2D1BWP12T U97 ( .A1(n49), .A2(n40), .ZN(n48) );
  INR2D0BWP12T U98 ( .A1(n48), .B1(n43), .ZN(memory_address[1]) );
  NR2D0BWP12T U99 ( .A1(n44), .A2(n43), .ZN(memory_address[4]) );
  AOI22D0BWP12T U100 ( .A1(n89), .A2(instruction_in[15]), .B1(n45), .B2(
        fetched_instruction_reg[15]), .ZN(n46) );
  ND2D1BWP12T U101 ( .A1(n47), .A2(n46), .ZN(instruction_out[15]) );
  INR2D0BWP12T U102 ( .A1(current_pc_in[0]), .B1(n94), .ZN(
        incremented_pc_out[0]) );
  NR2D0BWP12T U103 ( .A1(current_pc_in[1]), .A2(n94), .ZN(
        incremented_pc_out[1]) );
  NR2D0BWP12T U104 ( .A1(n94), .A2(n48), .ZN(incremented_pc_out[2]) );
  INVD1BWP12T U105 ( .I(n49), .ZN(n50) );
  ND2D1BWP12T U106 ( .A1(current_pc_in[3]), .A2(n50), .ZN(n51) );
  OA211D0BWP12T U107 ( .A1(current_pc_in[3]), .A2(n50), .B(n89), .C(n51), .Z(
        incremented_pc_out[3]) );
  NR2D1BWP12T U108 ( .A1(n52), .A2(n51), .ZN(n53) );
  AOI211D0BWP12T U109 ( .A1(n52), .A2(n51), .B(n53), .C(n94), .ZN(
        incremented_pc_out[4]) );
  ND2D1BWP12T U110 ( .A1(current_pc_in[5]), .A2(n53), .ZN(n54) );
  OA211D0BWP12T U111 ( .A1(current_pc_in[5]), .A2(n53), .B(n89), .C(n54), .Z(
        incremented_pc_out[5]) );
  NR2D1BWP12T U112 ( .A1(n55), .A2(n54), .ZN(n56) );
  AOI211D0BWP12T U113 ( .A1(n55), .A2(n54), .B(n56), .C(n94), .ZN(
        incremented_pc_out[6]) );
  ND2D1BWP12T U114 ( .A1(current_pc_in[7]), .A2(n56), .ZN(n57) );
  OA211D0BWP12T U115 ( .A1(current_pc_in[7]), .A2(n56), .B(n89), .C(n57), .Z(
        incremented_pc_out[7]) );
  NR2D1BWP12T U116 ( .A1(n58), .A2(n57), .ZN(n59) );
  AOI211D0BWP12T U117 ( .A1(n58), .A2(n57), .B(n59), .C(n94), .ZN(
        incremented_pc_out[8]) );
  ND2D1BWP12T U118 ( .A1(current_pc_in[9]), .A2(n59), .ZN(n60) );
  OA211D0BWP12T U119 ( .A1(current_pc_in[9]), .A2(n59), .B(n89), .C(n60), .Z(
        incremented_pc_out[9]) );
  NR2D1BWP12T U120 ( .A1(n61), .A2(n60), .ZN(n62) );
  AOI211D0BWP12T U121 ( .A1(n61), .A2(n60), .B(n62), .C(n94), .ZN(
        incremented_pc_out[10]) );
  ND2D1BWP12T U122 ( .A1(current_pc_in[11]), .A2(n62), .ZN(n63) );
  OA211D0BWP12T U123 ( .A1(current_pc_in[11]), .A2(n62), .B(n89), .C(n63), .Z(
        incremented_pc_out[11]) );
  NR2D1BWP12T U124 ( .A1(n64), .A2(n63), .ZN(n65) );
  AOI211D0BWP12T U125 ( .A1(n64), .A2(n63), .B(n65), .C(n94), .ZN(
        incremented_pc_out[12]) );
  ND2D1BWP12T U126 ( .A1(current_pc_in[13]), .A2(n65), .ZN(n66) );
  OA211D0BWP12T U127 ( .A1(current_pc_in[13]), .A2(n65), .B(n89), .C(n66), .Z(
        incremented_pc_out[13]) );
  INVD1BWP12T U128 ( .I(current_pc_in[14]), .ZN(n67) );
  NR2D1BWP12T U129 ( .A1(n67), .A2(n66), .ZN(n68) );
  AOI211D0BWP12T U130 ( .A1(n67), .A2(n66), .B(n68), .C(n94), .ZN(
        incremented_pc_out[14]) );
  ND2D1BWP12T U131 ( .A1(current_pc_in[15]), .A2(n68), .ZN(n69) );
  OA211D0BWP12T U132 ( .A1(current_pc_in[15]), .A2(n68), .B(n89), .C(n69), .Z(
        incremented_pc_out[15]) );
  NR2D1BWP12T U133 ( .A1(n70), .A2(n69), .ZN(n71) );
  AOI211D0BWP12T U134 ( .A1(n70), .A2(n69), .B(n71), .C(n94), .ZN(
        incremented_pc_out[16]) );
  ND2D1BWP12T U135 ( .A1(current_pc_in[17]), .A2(n71), .ZN(n72) );
  OA211D0BWP12T U136 ( .A1(current_pc_in[17]), .A2(n71), .B(n89), .C(n72), .Z(
        incremented_pc_out[17]) );
  INVD1BWP12T U137 ( .I(current_pc_in[18]), .ZN(n73) );
  NR2D1BWP12T U138 ( .A1(n73), .A2(n72), .ZN(n74) );
  AOI211D0BWP12T U139 ( .A1(n73), .A2(n72), .B(n74), .C(n94), .ZN(
        incremented_pc_out[18]) );
  ND2D1BWP12T U140 ( .A1(current_pc_in[19]), .A2(n74), .ZN(n75) );
  OA211D0BWP12T U141 ( .A1(current_pc_in[19]), .A2(n74), .B(n89), .C(n75), .Z(
        incremented_pc_out[19]) );
  INVD1BWP12T U142 ( .I(current_pc_in[20]), .ZN(n76) );
  NR2D1BWP12T U143 ( .A1(n76), .A2(n75), .ZN(n77) );
  AOI211D0BWP12T U144 ( .A1(n76), .A2(n75), .B(n77), .C(n94), .ZN(
        incremented_pc_out[20]) );
  ND2D1BWP12T U145 ( .A1(current_pc_in[21]), .A2(n77), .ZN(n78) );
  OA211D0BWP12T U146 ( .A1(current_pc_in[21]), .A2(n77), .B(n89), .C(n78), .Z(
        incremented_pc_out[21]) );
  INVD1BWP12T U147 ( .I(current_pc_in[22]), .ZN(n79) );
  NR2D1BWP12T U148 ( .A1(n79), .A2(n78), .ZN(n80) );
  AOI211D0BWP12T U149 ( .A1(n79), .A2(n78), .B(n80), .C(n94), .ZN(
        incremented_pc_out[22]) );
  ND2D1BWP12T U150 ( .A1(current_pc_in[23]), .A2(n80), .ZN(n81) );
  OA211D0BWP12T U151 ( .A1(current_pc_in[23]), .A2(n80), .B(n89), .C(n81), .Z(
        incremented_pc_out[23]) );
  INVD1BWP12T U152 ( .I(current_pc_in[24]), .ZN(n82) );
  NR2D1BWP12T U153 ( .A1(n82), .A2(n81), .ZN(n83) );
  AOI211D0BWP12T U154 ( .A1(n82), .A2(n81), .B(n83), .C(n94), .ZN(
        incremented_pc_out[24]) );
  ND2D1BWP12T U155 ( .A1(current_pc_in[25]), .A2(n83), .ZN(n84) );
  OA211D0BWP12T U156 ( .A1(current_pc_in[25]), .A2(n83), .B(n89), .C(n84), .Z(
        incremented_pc_out[25]) );
  INVD1BWP12T U157 ( .I(current_pc_in[26]), .ZN(n85) );
  NR2D1BWP12T U158 ( .A1(n85), .A2(n84), .ZN(n86) );
  AOI211D0BWP12T U159 ( .A1(n85), .A2(n84), .B(n86), .C(n94), .ZN(
        incremented_pc_out[26]) );
  ND2D1BWP12T U160 ( .A1(current_pc_in[27]), .A2(n86), .ZN(n87) );
  OA211D0BWP12T U161 ( .A1(current_pc_in[27]), .A2(n86), .B(n89), .C(n87), .Z(
        incremented_pc_out[27]) );
  INVD1BWP12T U162 ( .I(current_pc_in[28]), .ZN(n88) );
  NR2D1BWP12T U163 ( .A1(n88), .A2(n87), .ZN(n90) );
  AOI211D0BWP12T U164 ( .A1(n88), .A2(n87), .B(n90), .C(n94), .ZN(
        incremented_pc_out[28]) );
  ND2D1BWP12T U165 ( .A1(current_pc_in[29]), .A2(n90), .ZN(n91) );
  OA211D0BWP12T U166 ( .A1(current_pc_in[29]), .A2(n90), .B(n89), .C(n91), .Z(
        incremented_pc_out[29]) );
  INVD1BWP12T U167 ( .I(current_pc_in[30]), .ZN(n92) );
  NR2D1BWP12T U168 ( .A1(n92), .A2(n91), .ZN(n95) );
  AOI211D0BWP12T U169 ( .A1(n92), .A2(n91), .B(n95), .C(n94), .ZN(
        incremented_pc_out[30]) );
  NR2D1BWP12T U170 ( .A1(current_pc_in[31]), .A2(n95), .ZN(n93) );
  AOI211D0BWP12T U171 ( .A1(current_pc_in[31]), .A2(n95), .B(n94), .C(n93), 
        .ZN(incremented_pc_out[31]) );
  AO221D0BWP12T U172 ( .A1(incremented_pc_write_enable), .A2(instruction_in[8]), .B1(n96), .B2(fetched_instruction_reg[8]), .C(reset), .Z(N91) );
  AO221D0BWP12T U173 ( .A1(incremented_pc_write_enable), .A2(instruction_in[9]), .B1(n96), .B2(fetched_instruction_reg[9]), .C(reset), .Z(N92) );
  AO221D0BWP12T U174 ( .A1(incremented_pc_write_enable), .A2(
        instruction_in[10]), .B1(n96), .B2(fetched_instruction_reg[10]), .C(
        reset), .Z(N93) );
  AO221D0BWP12T U175 ( .A1(incremented_pc_write_enable), .A2(
        instruction_in[11]), .B1(n96), .B2(fetched_instruction_reg[11]), .C(
        reset), .Z(N94) );
  AO221D0BWP12T U176 ( .A1(incremented_pc_write_enable), .A2(
        instruction_in[12]), .B1(n96), .B2(fetched_instruction_reg[12]), .C(
        reset), .Z(N95) );
  AO221D0BWP12T U177 ( .A1(incremented_pc_write_enable), .A2(
        instruction_in[13]), .B1(n96), .B2(fetched_instruction_reg[13]), .C(
        reset), .Z(N96) );
  AO221D0BWP12T U178 ( .A1(incremented_pc_write_enable), .A2(
        instruction_in[15]), .B1(n96), .B2(fetched_instruction_reg[15]), .C(
        reset), .Z(N98) );
  OAI21D0BWP12T U179 ( .A1(memory_load_request), .A2(stall_decoder_in), .B(
        currentState_0_), .ZN(n98) );
  AOI31D0BWP12T U180 ( .A1(n98), .A2(n97), .A3(n96), .B(reset), .ZN(N79) );
endmodule


module top7 ( clk, reset, MEM_MEMCTRL_from_mem_data, 
        MEMCTRL_MEM_to_mem_read_enable, MEMCTRL_MEM_to_mem_write_enable, 
        MEMCTRL_MEM_to_mem_mem_enable, MEMCTRL_MEM_to_mem_address, 
        MEMCTRL_MEM_to_mem_data );
  input [15:0] MEM_MEMCTRL_from_mem_data;
  output [11:0] MEMCTRL_MEM_to_mem_address;
  output [15:0] MEMCTRL_MEM_to_mem_data;
  input clk, reset;
  output MEMCTRL_MEM_to_mem_read_enable, MEMCTRL_MEM_to_mem_write_enable,
         MEMCTRL_MEM_to_mem_mem_enable;
  wire   DEC_CPSR_update_flag_n, ALU_OUT_n, DEC_CPSR_update_flag_c, ALU_OUT_c,
         DEC_CPSR_update_flag_z, ALU_OUT_z, DEC_CPSR_update_flag_v, ALU_OUT_v,
         IF_DEC_instruction_valid, MEMCTRL_write_finished,
         MEMCTRL_read_finished, DEC_MISC_OUT_memory_address_source_is_reg,
         DEC_MEMCTRL_memorycontroller_sign_extend,
         DEC_MEMCTRL_memory_load_request, DEC_MEMCTRL_memory_store_request,
         DEC_IF_stall_to_instructionfetch, ALU_IN_c, IF_memory_load_req,
         MEMCTRL_load_in, n2, n3, n4, n5, n6, n7, n8, n10, n11,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21;
  wire   [15:0] IF_DEC_instruction;
  wire   [4:0] DEC_ALU_alu_opcode;
  wire   [1:0] DEC_MEMCTRL_load_store_width;
  wire   [11:0] MEMCTRL_IN_address;
  wire   [11:0] IF_instruction_memory_address;
  tri   clk;
  tri   reset;
  tri   new_n;
  tri   RF_OUT_n;
  tri   new_c;
  tri   RF_OUT_c;
  tri   new_z;
  tri   RF_OUT_z;
  tri   new_v;
  tri   RF_OUT_v;
  tri   [4:0] DEC_RF_operand_a;
  tri   [4:0] DEC_RF_operand_b;
  tri   [31:0] DEC_RF_offset_a;
  tri   [31:0] DEC_RF_offset_b;
  tri   [4:0] DEC_RF_alu_write_to_reg;
  tri   DEC_RF_alu_write_to_reg_enable;
  tri   [4:0] DEC_RF_memory_write_to_reg;
  tri   DEC_RF_memory_write_to_reg_enable;
  tri   [4:0] DEC_RF_memory_store_data_reg;
  tri   [4:0] DEC_RF_memory_store_address_reg;
  tri   [31:0] ALU_MISC_OUT_result;
  tri   [31:0] MEMCTRL_RF_IF_data_in;
  tri   [31:0] IF_RF_incremented_pc_out;
  tri   [31:0] RF_next_sp;
  tri   IF_RF_incremented_pc_write_enable;
  tri   [31:0] RF_ALU_operand_a;
  tri   [31:0] RF_ALU_operand_b;
  tri   [31:0] RF_MEMCTRL_data_reg;
  tri   [12:2] RF_MEMCTRL_address_reg;
  tri   [31:0] RF_pc_out;

  irdecode irdecode_inst1 ( .clk(clk), .reset(reset), .instruction(
        IF_DEC_instruction), .instruction_valid(IF_DEC_instruction_valid), 
        .flag_n(RF_OUT_n), .flag_z(RF_OUT_z), .flag_c(RF_OUT_c), .flag_v(
        RF_OUT_v), .memory_write_finished(MEMCTRL_write_finished), 
        .memory_read_finished(MEMCTRL_read_finished), .operand_a(
        DEC_RF_operand_a), .operand_b(DEC_RF_operand_b), .offset_a(
        DEC_RF_offset_a), .offset_b(DEC_RF_offset_b), .alu_opcode(
        DEC_ALU_alu_opcode), .update_flag_n(DEC_CPSR_update_flag_n), 
        .update_flag_z(DEC_CPSR_update_flag_z), .update_flag_c(
        DEC_CPSR_update_flag_c), .update_flag_v(DEC_CPSR_update_flag_v), 
        .alu_write_to_reg(DEC_RF_alu_write_to_reg), .alu_write_to_reg_enable(
        DEC_RF_alu_write_to_reg_enable), .memory_write_to_reg(
        DEC_RF_memory_write_to_reg), .memory_write_to_reg_enable(
        DEC_RF_memory_write_to_reg_enable), .memory_store_data_reg(
        DEC_RF_memory_store_data_reg), .memory_store_address_reg(
        DEC_RF_memory_store_address_reg), .memory_address_source_is_reg(
        DEC_MISC_OUT_memory_address_source_is_reg), .load_store_width(
        DEC_MEMCTRL_load_store_width), .memorycontroller_sign_extend(
        DEC_MEMCTRL_memorycontroller_sign_extend), .memory_load_request(
        DEC_MEMCTRL_memory_load_request), .stall_to_instructionfetch(
        DEC_IF_stall_to_instructionfetch), .memory_store_request_BAR(
        DEC_MEMCTRL_memory_store_request) );
  register_file register_file_inst1 ( .readA_sel(DEC_RF_operand_a), 
        .readB_sel(DEC_RF_operand_b), .readC_sel(DEC_RF_memory_store_data_reg), 
        .readD_sel(DEC_RF_memory_store_address_reg), .write1_sel(
        DEC_RF_alu_write_to_reg), .write2_sel(DEC_RF_memory_write_to_reg), 
        .write1_en(DEC_RF_alu_write_to_reg_enable), .write2_en(
        DEC_RF_memory_write_to_reg_enable), .write1_in(ALU_MISC_OUT_result), 
        .write2_in(MEMCTRL_RF_IF_data_in), .immediate1_in(DEC_RF_offset_a), 
        .immediate2_in(DEC_RF_offset_b), .next_pc_in(IF_RF_incremented_pc_out), 
        .next_cpsr_in({new_n, new_c, new_z, new_v}), .next_sp_in(RF_next_sp), 
        .next_pc_en(IF_RF_incremented_pc_write_enable), .clk(clk), .reset(
        reset), .regA_out(RF_ALU_operand_a), .regB_out(RF_ALU_operand_b), 
        .regC_out(RF_MEMCTRL_data_reg), .regD_out({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        RF_MEMCTRL_address_reg, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21}), .pc_out(RF_pc_out), .cpsr_out({RF_OUT_n, 
        RF_OUT_c, RF_OUT_z, RF_OUT_v}), .sp_out(RF_next_sp) );
  ALU_VARIABLE ALU_VARIABLE_inst1 ( .a(RF_ALU_operand_a), .b(RF_ALU_operand_b), 
        .op(DEC_ALU_alu_opcode[3:0]), .c_in(ALU_IN_c), .result(
        ALU_MISC_OUT_result), .c_out(ALU_OUT_c), .z(ALU_OUT_z), .n(ALU_OUT_n), 
        .v(ALU_OUT_v) );
  memory_interface memory_interface_inst1 ( .address(MEMCTRL_IN_address), 
        .data_in(RF_MEMCTRL_data_reg), .load(MEMCTRL_load_in), .clk(clk), 
        .reset(reset), .is_signed(DEC_MEMCTRL_memorycontroller_sign_extend), 
        .word_type(DEC_MEMCTRL_load_store_width), .from_mem_data(
        MEM_MEMCTRL_from_mem_data), .to_mem_read_enable(
        MEMCTRL_MEM_to_mem_read_enable), .to_mem_write_enable(
        MEMCTRL_MEM_to_mem_write_enable), .to_mem_address(
        MEMCTRL_MEM_to_mem_address), .to_mem_data(MEMCTRL_MEM_to_mem_data), 
        .data_out(MEMCTRL_RF_IF_data_in), .write_ready(MEMCTRL_write_finished), 
        .output_valid(MEMCTRL_read_finished), .store_BAR(
        DEC_MEMCTRL_memory_store_request) );
  Instruction_Fetch Instruction_Fetch_inst1 ( .clk(clk), .reset(reset), 
        .stall_decoder_in(DEC_IF_stall_to_instructionfetch), 
        .memory_output_valid(MEMCTRL_read_finished), .current_pc_in(RF_pc_out), 
        .instruction_in(MEMCTRL_RF_IF_data_in[15:0]), .memory_load_request(
        IF_memory_load_req), .incremented_pc_write_enable(
        IF_RF_incremented_pc_write_enable), .instruction_valid(
        IF_DEC_instruction_valid), .memory_address(
        IF_instruction_memory_address), .incremented_pc_out(
        IF_RF_incremented_pc_out), .instruction_out(IF_DEC_instruction) );
  AO222D0BWP12T U12 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[11]), .B1(RF_MEMCTRL_address_reg[12]), 
        .B2(n3), .C1(ALU_MISC_OUT_result[12]), .C2(n4), .Z(
        MEMCTRL_IN_address[11]) );
  AO222D0BWP12T U13 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[10]), .B1(n4), .B2(
        ALU_MISC_OUT_result[11]), .C1(RF_MEMCTRL_address_reg[11]), .C2(n3), 
        .Z(MEMCTRL_IN_address[10]) );
  AO222D0BWP12T U14 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[9]), .B1(n4), .B2(
        ALU_MISC_OUT_result[10]), .C1(RF_MEMCTRL_address_reg[10]), .C2(n3), 
        .Z(MEMCTRL_IN_address[9]) );
  AO222D0BWP12T U15 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[8]), .B1(n4), .B2(ALU_MISC_OUT_result[9]), .C1(RF_MEMCTRL_address_reg[9]), .C2(n3), .Z(MEMCTRL_IN_address[8]) );
  AO222D0BWP12T U16 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[7]), .B1(n4), .B2(ALU_MISC_OUT_result[8]), .C1(RF_MEMCTRL_address_reg[8]), .C2(n3), .Z(MEMCTRL_IN_address[7]) );
  AO222D0BWP12T U17 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[6]), .B1(n4), .B2(ALU_MISC_OUT_result[7]), .C1(RF_MEMCTRL_address_reg[7]), .C2(n3), .Z(MEMCTRL_IN_address[6]) );
  AO222D0BWP12T U18 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[5]), .B1(n4), .B2(ALU_MISC_OUT_result[6]), .C1(RF_MEMCTRL_address_reg[6]), .C2(n3), .Z(MEMCTRL_IN_address[5]) );
  AO222D0BWP12T U19 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[4]), .B1(n4), .B2(ALU_MISC_OUT_result[5]), .C1(RF_MEMCTRL_address_reg[5]), .C2(n3), .Z(MEMCTRL_IN_address[4]) );
  AO222D0BWP12T U20 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[3]), .B1(n4), .B2(ALU_MISC_OUT_result[4]), .C1(RF_MEMCTRL_address_reg[4]), .C2(n3), .Z(MEMCTRL_IN_address[3]) );
  AO222D0BWP12T U21 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[2]), .B1(n4), .B2(ALU_MISC_OUT_result[3]), .C1(RF_MEMCTRL_address_reg[3]), .C2(n3), .Z(MEMCTRL_IN_address[2]) );
  AO222D0BWP12T U22 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[1]), .B1(n4), .B2(ALU_MISC_OUT_result[2]), .C1(RF_MEMCTRL_address_reg[2]), .C2(n3), .Z(MEMCTRL_IN_address[1]) );
  AO22D0BWP12T U25 ( .A1(ALU_OUT_v), .A2(DEC_CPSR_update_flag_v), .B1(n5), 
        .B2(RF_OUT_v), .Z(new_v) );
  AO22D0BWP12T U26 ( .A1(ALU_OUT_z), .A2(DEC_CPSR_update_flag_z), .B1(n7), 
        .B2(RF_OUT_z), .Z(new_z) );
  AO22D0BWP12T U27 ( .A1(ALU_OUT_c), .A2(DEC_CPSR_update_flag_c), .B1(n6), 
        .B2(RF_OUT_c), .Z(new_c) );
  AO22D0BWP12T U28 ( .A1(ALU_OUT_n), .A2(DEC_CPSR_update_flag_n), .B1(n8), 
        .B2(RF_OUT_n), .Z(new_n) );
  TIELBWP12T U29 ( .ZN(n10) );
  INVD1BWP12T U30 ( .I(n10), .ZN(MEMCTRL_MEM_to_mem_mem_enable) );
  NR2D1BWP12T U31 ( .A1(IF_memory_load_req), .A2(
        DEC_MISC_OUT_memory_address_source_is_reg), .ZN(n4) );
  INVD1BWP12T U32 ( .I(RF_OUT_c), .ZN(n2) );
  OAI22D1BWP12T U33 ( .A1(DEC_ALU_alu_opcode[4]), .A2(n2), .B1(
        DEC_ALU_alu_opcode[3]), .B2(n11), .ZN(ALU_IN_c) );
  AN2XD0BWP12T U34 ( .A1(IF_memory_load_req), .A2(
        IF_instruction_memory_address[0]), .Z(MEMCTRL_IN_address[0]) );
  IND4D1BWP12T U35 ( .A1(DEC_ALU_alu_opcode[0]), .B1(DEC_ALU_alu_opcode[4]), 
        .B2(DEC_ALU_alu_opcode[2]), .B3(DEC_ALU_alu_opcode[1]), .ZN(n11) );
  INR2XD0BWP12T U36 ( .A1(DEC_MISC_OUT_memory_address_source_is_reg), .B1(
        IF_memory_load_req), .ZN(n3) );
  OR2XD0BWP12T U37 ( .A1(IF_memory_load_req), .A2(
        DEC_MEMCTRL_memory_load_request), .Z(MEMCTRL_load_in) );
  INVD1BWP12T U38 ( .I(DEC_CPSR_update_flag_v), .ZN(n5) );
  INVD1BWP12T U39 ( .I(DEC_CPSR_update_flag_c), .ZN(n6) );
  INVD1BWP12T U40 ( .I(DEC_CPSR_update_flag_z), .ZN(n7) );
  INVD1BWP12T U41 ( .I(DEC_CPSR_update_flag_n), .ZN(n8) );
endmodule

