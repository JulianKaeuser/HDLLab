module memory (
  address,
  input_bus,
  output_bus,
  valid,
  rw,
  );


  endmodule
