// AUTHORS: Group 06 /Julian Käuser
// Friday 08/04/2017

module mem_cache (

  );

endmodule
