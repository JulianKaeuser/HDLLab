
module ALU_VARIABLE ( a, b, op, c_in, result, c_out, z, n, v );
  input [31:0] a;
  input [31:0] b;
  input [3:0] op;
  output [31:0] result;
  input c_in;
  output c_out, z, n, v;
  wire   n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
         n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234,
         n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
         n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
         n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
         n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
         n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
         n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282,
         n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
         n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
         n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306,
         n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314,
         n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
         n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
         n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338,
         n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346,
         n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354,
         n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
         n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
         n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378,
         n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386,
         n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
         n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
         n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410,
         n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418,
         n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426,
         n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434,
         n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
         n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450,
         n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
         n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466,
         n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474,
         n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482,
         n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490,
         n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498,
         n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506,
         n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
         n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522,
         n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530,
         n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538,
         n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546,
         n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554,
         n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562,
         n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570,
         n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578,
         n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
         n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594,
         n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602,
         n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610,
         n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618,
         n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626,
         n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634,
         n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642,
         n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650,
         n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658,
         n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666,
         n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674,
         n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682,
         n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690,
         n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698,
         n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706,
         n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714,
         n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
         n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730,
         n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738,
         n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746,
         n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754,
         n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762,
         n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770,
         n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778,
         n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786,
         n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794,
         n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802,
         n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810,
         n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818,
         n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826,
         n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834,
         n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842,
         n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850,
         n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858,
         n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866,
         n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874,
         n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882,
         n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890,
         n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898,
         n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906,
         n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914,
         n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922,
         n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930,
         n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938,
         n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946,
         n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954,
         n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962,
         n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970,
         n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978,
         n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986,
         n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994,
         n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002,
         n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010,
         n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018,
         n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026,
         n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034,
         n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042,
         n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050,
         n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058,
         n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066,
         n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074,
         n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082,
         n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090,
         n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098,
         n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106,
         n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114,
         n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122,
         n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130,
         n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138,
         n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146,
         n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154,
         n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162,
         n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170,
         n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178,
         n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186,
         n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194,
         n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202,
         n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210,
         n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218,
         n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226,
         n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234,
         n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242,
         n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250,
         n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258,
         n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266,
         n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274,
         n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282,
         n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290,
         n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298,
         n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306,
         n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314,
         n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322,
         n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330,
         n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338,
         n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346,
         n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354,
         n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362,
         n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370,
         n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378,
         n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386,
         n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394,
         n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402,
         n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410,
         n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418,
         n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426,
         n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434,
         n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442,
         n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450,
         n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458,
         n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466,
         n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474,
         n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482,
         n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490,
         n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498,
         n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506,
         n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514,
         n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522,
         n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530,
         n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538,
         n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546,
         n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554,
         n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562,
         n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570,
         n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578,
         n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586,
         n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594,
         n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602,
         n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610,
         n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618,
         n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626,
         n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634,
         n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642,
         n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650,
         n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658,
         n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666,
         n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674,
         n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682,
         n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690,
         n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698,
         n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706,
         n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714,
         n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722,
         n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730,
         n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738,
         n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746,
         n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754,
         n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762,
         n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770,
         n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778,
         n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786,
         n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794,
         n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802,
         n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810,
         n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818,
         n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826,
         n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834,
         n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842,
         n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850,
         n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858,
         n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866,
         n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874,
         n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882,
         n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890,
         n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898,
         n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906,
         n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914,
         n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922,
         n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930,
         n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938,
         n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946,
         n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954,
         n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962,
         n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970,
         n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978,
         n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986,
         n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994,
         n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002,
         n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010,
         n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018,
         n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026,
         n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034,
         n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042,
         n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050,
         n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058,
         n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066,
         n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074,
         n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082,
         n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090,
         n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098,
         n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106,
         n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114,
         n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122,
         n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130,
         n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138,
         n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146,
         n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154,
         n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162,
         n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170,
         n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178,
         n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186,
         n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194,
         n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202,
         n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210,
         n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218,
         n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226,
         n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234,
         n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242,
         n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250,
         n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258,
         n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266,
         n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274,
         n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282,
         n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290,
         n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298,
         n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306,
         n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314,
         n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322,
         n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330,
         n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338,
         n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346,
         n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354,
         n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362,
         n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370,
         n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378,
         n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386,
         n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394,
         n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402,
         n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410,
         n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418,
         n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426,
         n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434,
         n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442,
         n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450,
         n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458,
         n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466,
         n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474,
         n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482,
         n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490,
         n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498,
         n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506,
         n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514,
         n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522,
         n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530,
         n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538,
         n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546,
         n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554,
         n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562,
         n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570,
         n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578,
         n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586,
         n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594,
         n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602,
         n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610,
         n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618,
         n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626,
         n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634,
         n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642,
         n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650,
         n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658,
         n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666,
         n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674,
         n23675, n23676, n23677, n23678;

  AOI22D0BWP12T U10753 ( .A1(n21748), .A2(b[16]), .B1(n21076), .B2(n21585), 
        .ZN(n20323) );
  CKND2D0BWP12T U10754 ( .A1(b[15]), .A2(n21077), .ZN(n20324) );
  OAI211D0BWP12T U10755 ( .A1(n22547), .A2(n21745), .B(n20323), .C(n20324), 
        .ZN(n20325) );
  MOAI22D0BWP12T U10756 ( .A1(a[14]), .A2(n20325), .B1(a[14]), .B2(n20325), 
        .ZN(n20326) );
  MAOI22D0BWP12T U10757 ( .A1(n20999), .A2(n20326), .B1(n20999), .B2(n20326), 
        .ZN(n20327) );
  MAOI22D0BWP12T U10758 ( .A1(n21128), .A2(n20327), .B1(n21128), .B2(n20327), 
        .ZN(n21129) );
  CKND0BWP12T U10759 ( .I(n21128), .ZN(n20328) );
  MAOI222D0BWP12T U10760 ( .A(n20999), .B(n20326), .C(n20328), .ZN(n21121) );
  OAI22D0BWP12T U10761 ( .A1(n21757), .A2(n22612), .B1(n21887), .B2(n21207), 
        .ZN(n20329) );
  OAI22D0BWP12T U10762 ( .A1(n21760), .A2(n21934), .B1(n21758), .B2(n21595), 
        .ZN(n20330) );
  NR2D0BWP12T U10763 ( .A1(n20329), .A2(n20330), .ZN(n20331) );
  MOAI22D0BWP12T U10764 ( .A1(a[11]), .A2(n20331), .B1(a[11]), .B2(n20331), 
        .ZN(n20332) );
  MAOI22D0BWP12T U10765 ( .A1(n21152), .A2(n20332), .B1(n21152), .B2(n20332), 
        .ZN(n20333) );
  MAOI22D0BWP12T U10766 ( .A1(n21288), .A2(n20333), .B1(n21288), .B2(n20333), 
        .ZN(n21289) );
  CKND0BWP12T U10767 ( .I(n21288), .ZN(n20334) );
  MAOI222D0BWP12T U10768 ( .A(n21152), .B(n20334), .C(n20332), .ZN(n21286) );
  NR2D0BWP12T U10769 ( .A1(n21725), .A2(n21759), .ZN(n20335) );
  OAI22D0BWP12T U10770 ( .A1(n21727), .A2(n21932), .B1(n21724), .B2(n21886), 
        .ZN(n20336) );
  AOI211D0BWP12T U10771 ( .A1(b[21]), .A2(n21730), .B(n20335), .C(n20336), 
        .ZN(n20337) );
  MOAI22D0BWP12T U10772 ( .A1(n21966), .A2(n20337), .B1(n21966), .B2(n20337), 
        .ZN(n20338) );
  MAOI22D0BWP12T U10773 ( .A1(n21263), .A2(n20338), .B1(n21263), .B2(n20338), 
        .ZN(n20339) );
  MAOI22D0BWP12T U10774 ( .A1(n21377), .A2(n20339), .B1(n21377), .B2(n20339), 
        .ZN(n21378) );
  CKND0BWP12T U10775 ( .I(n21377), .ZN(n20340) );
  MAOI222D0BWP12T U10776 ( .A(n21263), .B(n20340), .C(n20338), .ZN(n21372) );
  NR4D0BWP12T U10777 ( .A1(n23494), .A2(n23496), .A3(n23495), .A4(n23497), 
        .ZN(n20341) );
  NR3D0BWP12T U10778 ( .A1(n23491), .A2(n23492), .A3(n23493), .ZN(n20342) );
  OA211D0BWP12T U10779 ( .A1(a[28]), .A2(n23490), .B(n20341), .C(n20342), .Z(
        n20343) );
  OAI211D0BWP12T U10780 ( .A1(a[20]), .A2(n23498), .B(n23501), .C(n20343), 
        .ZN(n20344) );
  NR4D0BWP12T U10781 ( .A1(n23499), .A2(n23500), .A3(n23503), .A4(n20344), 
        .ZN(n20345) );
  IND4D0BWP12T U10782 ( .A1(n23502), .B1(n23504), .B2(n23505), .B3(n20345), 
        .ZN(n20346) );
  ND4D0BWP12T U10783 ( .A1(n23487), .A2(n23486), .A3(n23488), .A4(n23489), 
        .ZN(n20347) );
  NR4D0BWP12T U10784 ( .A1(n23506), .A2(n23507), .A3(n20346), .A4(n20347), 
        .ZN(n20348) );
  INR4D0BWP12T U10785 ( .A1(n23482), .B1(n23481), .B2(n23479), .B3(n23480), 
        .ZN(n20349) );
  OAI211D0BWP12T U10786 ( .A1(n23484), .A2(a[15]), .B(n23483), .C(n20349), 
        .ZN(n20350) );
  AOI211D0BWP12T U10787 ( .A1(b[8]), .A2(n21966), .B(n23485), .C(n20350), .ZN(
        n20351) );
  AOI22D0BWP12T U10788 ( .A1(n23509), .A2(n23508), .B1(n20348), .B2(n20351), 
        .ZN(n23537) );
  OAI222D0BWP12T U10789 ( .A1(n23017), .A2(n21665), .B1(n22806), .B2(n21717), 
        .C1(n21667), .C2(n21666), .ZN(n20352) );
  NR2D0BWP12T U10790 ( .A1(n22941), .A2(n22939), .ZN(n20353) );
  MAOI22D0BWP12T U10791 ( .A1(n20352), .A2(n21882), .B1(n20352), .B2(n20353), 
        .ZN(n20354) );
  NR2D0BWP12T U10792 ( .A1(n22896), .A2(n22897), .ZN(n20355) );
  AOI31D0BWP12T U10793 ( .A1(n21663), .A2(a[2]), .A3(n21664), .B(n20355), .ZN(
        n20356) );
  AO31D0BWP12T U10794 ( .A1(n21670), .A2(n22955), .A3(n21669), .B(n21668), .Z(
        n20357) );
  MAOI222D0BWP12T U10795 ( .A(n20354), .B(n20356), .C(n20357), .ZN(n22839) );
  MOAI22D0BWP12T U10796 ( .A1(n20354), .A2(n20357), .B1(n20354), .B2(n20357), 
        .ZN(n20358) );
  MAOI22D0BWP12T U10797 ( .A1(n20356), .A2(n20358), .B1(n20356), .B2(n20358), 
        .ZN(n23305) );
  NR2D0BWP12T U10798 ( .A1(n21758), .A2(n21700), .ZN(n20359) );
  OAI22D0BWP12T U10799 ( .A1(n21757), .A2(n22418), .B1(n21760), .B2(n21944), 
        .ZN(n20360) );
  AOI211D0BWP12T U10800 ( .A1(n21763), .A2(b[17]), .B(n20359), .C(n20360), 
        .ZN(n20361) );
  MOAI22D0BWP12T U10801 ( .A1(a[11]), .A2(n20361), .B1(a[11]), .B2(n20361), 
        .ZN(n20362) );
  MAOI22D0BWP12T U10802 ( .A1(n21129), .A2(n20362), .B1(n21129), .B2(n20362), 
        .ZN(n20363) );
  MAOI22D0BWP12T U10803 ( .A1(n21264), .A2(n20363), .B1(n21264), .B2(n20363), 
        .ZN(n21265) );
  CKND0BWP12T U10804 ( .I(n21264), .ZN(n20364) );
  MAOI222D0BWP12T U10805 ( .A(n21129), .B(n20364), .C(n20362), .ZN(n21262) );
  NR2D0BWP12T U10806 ( .A1(n21725), .A2(n21765), .ZN(n20365) );
  OAI22D0BWP12T U10807 ( .A1(n22547), .A2(n21727), .B1(n21934), .B2(n21724), 
        .ZN(n20366) );
  AOI211D0BWP12T U10808 ( .A1(b[12]), .A2(n21730), .B(n20365), .C(n20366), 
        .ZN(n20367) );
  MOAI22D0BWP12T U10809 ( .A1(n21966), .A2(n20367), .B1(n21966), .B2(n20367), 
        .ZN(n20368) );
  MAOI22D0BWP12T U10810 ( .A1(n21504), .A2(n20368), .B1(n21504), .B2(n20368), 
        .ZN(n20369) );
  MAOI22D0BWP12T U10811 ( .A1(n21367), .A2(n20369), .B1(n21367), .B2(n20369), 
        .ZN(n21505) );
  CKND0BWP12T U10812 ( .I(n21504), .ZN(n20370) );
  MAOI222D0BWP12T U10813 ( .A(n21367), .B(n20368), .C(n20370), .ZN(n21403) );
  NR2D0BWP12T U10814 ( .A1(n21732), .A2(n21565), .ZN(n20371) );
  OAI22D0BWP12T U10815 ( .A1(n21731), .A2(n21886), .B1(n21734), .B2(n23498), 
        .ZN(n20372) );
  AOI211D0BWP12T U10816 ( .A1(b[21]), .A2(n21737), .B(n20371), .C(n20372), 
        .ZN(n20373) );
  MOAI22D0BWP12T U10817 ( .A1(a[5]), .A2(n20373), .B1(a[5]), .B2(n20373), .ZN(
        n20374) );
  MAOI22D0BWP12T U10818 ( .A1(n21390), .A2(n20374), .B1(n21390), .B2(n20374), 
        .ZN(n20375) );
  MAOI22D0BWP12T U10819 ( .A1(n21546), .A2(n20375), .B1(n21546), .B2(n20375), 
        .ZN(n21547) );
  CKND0BWP12T U10820 ( .I(n21546), .ZN(n20376) );
  MAOI222D0BWP12T U10821 ( .A(n21390), .B(n20376), .C(n20374), .ZN(n21544) );
  NR2D0BWP12T U10822 ( .A1(n22699), .A2(n21717), .ZN(n20377) );
  MAOI22D0BWP12T U10823 ( .A1(n22977), .A2(b[8]), .B1(n21716), .B2(n22675), 
        .ZN(n20378) );
  OAI21D0BWP12T U10824 ( .A1(n21711), .A2(n21678), .B(n20378), .ZN(n20379) );
  OAI22D0BWP12T U10825 ( .A1(n21716), .A2(n21678), .B1(n21711), .B2(n22675), 
        .ZN(n20380) );
  OAI21D0BWP12T U10826 ( .A1(n20377), .A2(n20379), .B(a[2]), .ZN(n20381) );
  OAI31D0BWP12T U10827 ( .A1(n20377), .A2(a[2]), .A3(n20380), .B(n20381), .ZN(
        n20382) );
  CKND0BWP12T U10828 ( .I(n22672), .ZN(n20383) );
  MAOI222D0BWP12T U10829 ( .A(n20382), .B(n21617), .C(n20383), .ZN(n22631) );
  MAOI22D0BWP12T U10830 ( .A1(n22672), .A2(n21617), .B1(n22672), .B2(n21617), 
        .ZN(n20384) );
  MAOI22D0BWP12T U10831 ( .A1(n20382), .A2(n20384), .B1(n20382), .B2(n20384), 
        .ZN(n23332) );
  AOI21D0BWP12T U10832 ( .A1(n20862), .A2(n20863), .B(n20861), .ZN(n20385) );
  NR2D0BWP12T U10833 ( .A1(n21237), .A2(n21667), .ZN(n20386) );
  OAI22D0BWP12T U10834 ( .A1(n23017), .A2(n21238), .B1(n22806), .B2(n21777), 
        .ZN(n20387) );
  AOI211D0BWP12T U10835 ( .A1(n21772), .A2(b[2]), .B(n20386), .C(n20387), .ZN(
        n20388) );
  MAOI22D0BWP12T U10836 ( .A1(a[23]), .A2(n20388), .B1(a[23]), .B2(n20388), 
        .ZN(n20389) );
  MAOI22D0BWP12T U10837 ( .A1(n20385), .A2(n20389), .B1(n20385), .B2(n20389), 
        .ZN(n20390) );
  IND2D0BWP12T U10838 ( .A1(n20890), .B1(n20891), .ZN(n20391) );
  OAI31D0BWP12T U10839 ( .A1(n22267), .A2(n20860), .A3(n20859), .B(n20391), 
        .ZN(n20392) );
  MAOI22D0BWP12T U10840 ( .A1(n20390), .A2(n20392), .B1(n20390), .B2(n20392), 
        .ZN(n20945) );
  MAOI222D0BWP12T U10841 ( .A(n20385), .B(n20392), .C(n20393), .ZN(n20878) );
  CKND0BWP12T U10842 ( .I(n20389), .ZN(n20393) );
  OAI22D0BWP12T U10843 ( .A1(n22699), .A2(n21757), .B1(n21758), .B2(n21678), 
        .ZN(n20394) );
  OAI22D0BWP12T U10844 ( .A1(n22675), .A2(n21760), .B1(n21207), .B2(n22741), 
        .ZN(n20395) );
  NR2D0BWP12T U10845 ( .A1(n20394), .A2(n20395), .ZN(n20396) );
  MOAI22D0BWP12T U10846 ( .A1(a[11]), .A2(n20396), .B1(a[11]), .B2(n20396), 
        .ZN(n20397) );
  MAOI22D0BWP12T U10847 ( .A1(n21161), .A2(n21364), .B1(n21161), .B2(n21364), 
        .ZN(n20398) );
  MAOI22D0BWP12T U10848 ( .A1(n20397), .A2(n20398), .B1(n20397), .B2(n20398), 
        .ZN(n21365) );
  CKND0BWP12T U10849 ( .I(n21364), .ZN(n20399) );
  MAOI222D0BWP12T U10850 ( .A(n21161), .B(n20397), .C(n20399), .ZN(n21366) );
  NR2D0BWP12T U10851 ( .A1(n21725), .A2(n21751), .ZN(n20400) );
  OAI22D0BWP12T U10852 ( .A1(n21750), .A2(n21727), .B1(n21724), .B2(n21753), 
        .ZN(n20401) );
  AOI211D0BWP12T U10853 ( .A1(b[15]), .A2(n21730), .B(n20400), .C(n20401), 
        .ZN(n20402) );
  MOAI22D0BWP12T U10854 ( .A1(n21966), .A2(n20402), .B1(n21966), .B2(n20402), 
        .ZN(n20403) );
  MAOI22D0BWP12T U10855 ( .A1(n21287), .A2(n20403), .B1(n21287), .B2(n20403), 
        .ZN(n20404) );
  MAOI22D0BWP12T U10856 ( .A1(n21396), .A2(n20404), .B1(n21396), .B2(n20404), 
        .ZN(n21397) );
  CKND0BWP12T U10857 ( .I(n21396), .ZN(n20405) );
  MAOI222D0BWP12T U10858 ( .A(n21287), .B(n20405), .C(n20403), .ZN(n21391) );
  NR2D0BWP12T U10859 ( .A1(n21732), .A2(n21759), .ZN(n20406) );
  OAI22D0BWP12T U10860 ( .A1(n21731), .A2(n21932), .B1(n21734), .B2(n22293), 
        .ZN(n20407) );
  AOI211D0BWP12T U10861 ( .A1(b[22]), .A2(n21737), .B(n20406), .C(n20407), 
        .ZN(n20408) );
  MOAI22D0BWP12T U10862 ( .A1(a[5]), .A2(n20408), .B1(a[5]), .B2(n20408), .ZN(
        n20409) );
  MAOI22D0BWP12T U10863 ( .A1(n21388), .A2(n20409), .B1(n21388), .B2(n20409), 
        .ZN(n20410) );
  MAOI22D0BWP12T U10864 ( .A1(n21544), .A2(n20410), .B1(n21544), .B2(n20410), 
        .ZN(n21545) );
  CKND0BWP12T U10865 ( .I(n21544), .ZN(n20411) );
  MAOI222D0BWP12T U10866 ( .A(n21388), .B(n20411), .C(n20409), .ZN(n21536) );
  NR2D0BWP12T U10867 ( .A1(n21717), .A2(n21887), .ZN(n20412) );
  AOI22D0BWP12T U10868 ( .A1(b[10]), .A2(n22977), .B1(n21719), .B2(n21684), 
        .ZN(n20413) );
  OAI21D0BWP12T U10869 ( .A1(n21716), .A2(n22612), .B(n20413), .ZN(n20414) );
  OAI22D0BWP12T U10870 ( .A1(n21683), .A2(n21716), .B1(n21711), .B2(n22612), 
        .ZN(n20415) );
  OAI21D0BWP12T U10871 ( .A1(n20412), .A2(n20414), .B(a[2]), .ZN(n20416) );
  OAI31D0BWP12T U10872 ( .A1(n20412), .A2(a[2]), .A3(n20415), .B(n20416), .ZN(
        n20417) );
  CKND0BWP12T U10873 ( .I(n22614), .ZN(n20418) );
  MAOI222D0BWP12T U10874 ( .A(n21682), .B(n20417), .C(n20418), .ZN(n22591) );
  MAOI22D0BWP12T U10875 ( .A1(n21682), .A2(n22614), .B1(n21682), .B2(n22614), 
        .ZN(n20419) );
  MAOI22D0BWP12T U10876 ( .A1(n20417), .A2(n20419), .B1(n20417), .B2(n20419), 
        .ZN(n23323) );
  NR2D0BWP12T U10877 ( .A1(n21636), .A2(n21237), .ZN(n20420) );
  OAI22D0BWP12T U10878 ( .A1(n21935), .A2(n21238), .B1(n23370), .B2(n21777), 
        .ZN(n20421) );
  AOI211D0BWP12T U10879 ( .A1(n21772), .A2(b[5]), .B(n20420), .C(n20421), .ZN(
        n20422) );
  MOAI22D0BWP12T U10880 ( .A1(a[23]), .A2(n20422), .B1(a[23]), .B2(n20422), 
        .ZN(n20423) );
  MAOI22D0BWP12T U10881 ( .A1(n20838), .A2(n20423), .B1(n20838), .B2(n20423), 
        .ZN(n20424) );
  MAOI22D0BWP12T U10882 ( .A1(n20870), .A2(n20424), .B1(n20870), .B2(n20424), 
        .ZN(n20918) );
  CKND0BWP12T U10883 ( .I(n20870), .ZN(n20425) );
  MAOI222D0BWP12T U10884 ( .A(n20838), .B(n20425), .C(n20423), .ZN(n21101) );
  AOI22D0BWP12T U10885 ( .A1(b[11]), .A2(n21748), .B1(b[10]), .B2(n21077), 
        .ZN(n20426) );
  CKND2D0BWP12T U10886 ( .A1(n21076), .A2(n21773), .ZN(n20427) );
  OAI211D0BWP12T U10887 ( .A1(n22699), .A2(n21745), .B(n20426), .C(n20427), 
        .ZN(n20428) );
  MOAI22D0BWP12T U10888 ( .A1(a[14]), .A2(n20428), .B1(a[14]), .B2(n20428), 
        .ZN(n20429) );
  MAOI22D0BWP12T U10889 ( .A1(n21026), .A2(n20429), .B1(n21026), .B2(n20429), 
        .ZN(n20430) );
  MAOI22D0BWP12T U10890 ( .A1(n21147), .A2(n20430), .B1(n21147), .B2(n20430), 
        .ZN(n21148) );
  CKND0BWP12T U10891 ( .I(n21147), .ZN(n20431) );
  MAOI222D0BWP12T U10892 ( .A(n21026), .B(n20429), .C(n20431), .ZN(n21145) );
  NR2D0BWP12T U10893 ( .A1(n21758), .A2(n21744), .ZN(n20432) );
  OAI22D0BWP12T U10894 ( .A1(n21757), .A2(n21944), .B1(n21760), .B2(n23498), 
        .ZN(n20433) );
  AOI211D0BWP12T U10895 ( .A1(n21763), .A2(b[18]), .B(n20432), .C(n20433), 
        .ZN(n20434) );
  MOAI22D0BWP12T U10896 ( .A1(a[11]), .A2(n20434), .B1(a[11]), .B2(n20434), 
        .ZN(n20435) );
  MAOI22D0BWP12T U10897 ( .A1(n21124), .A2(n20435), .B1(n21124), .B2(n20435), 
        .ZN(n20436) );
  MAOI22D0BWP12T U10898 ( .A1(n21262), .A2(n20436), .B1(n21262), .B2(n20436), 
        .ZN(n21263) );
  CKND0BWP12T U10899 ( .I(n21262), .ZN(n20437) );
  MAOI222D0BWP12T U10900 ( .A(n21124), .B(n20437), .C(n20435), .ZN(n21257) );
  NR2D0BWP12T U10901 ( .A1(n21725), .A2(n21573), .ZN(n20438) );
  OAI22D0BWP12T U10902 ( .A1(n21727), .A2(n22418), .B1(n21750), .B2(n21724), 
        .ZN(n20439) );
  AOI211D0BWP12T U10903 ( .A1(b[16]), .A2(n21730), .B(n20438), .C(n20439), 
        .ZN(n20440) );
  MOAI22D0BWP12T U10904 ( .A1(n21966), .A2(n20440), .B1(n21966), .B2(n20440), 
        .ZN(n20441) );
  MAOI22D0BWP12T U10905 ( .A1(n21285), .A2(n20441), .B1(n21285), .B2(n20441), 
        .ZN(n20442) );
  MAOI22D0BWP12T U10906 ( .A1(n21391), .A2(n20442), .B1(n21391), .B2(n20442), 
        .ZN(n21392) );
  CKND0BWP12T U10907 ( .I(n21391), .ZN(n20443) );
  MAOI222D0BWP12T U10908 ( .A(n21285), .B(n20443), .C(n20441), .ZN(n21389) );
  NR2D0BWP12T U10909 ( .A1(n21732), .A2(n21555), .ZN(n20444) );
  OAI22D0BWP12T U10910 ( .A1(n21731), .A2(n21556), .B1(n21734), .B2(n21886), 
        .ZN(n20445) );
  AOI211D0BWP12T U10911 ( .A1(b[23]), .A2(n21737), .B(n20444), .C(n20445), 
        .ZN(n20446) );
  MOAI22D0BWP12T U10912 ( .A1(a[5]), .A2(n20446), .B1(a[5]), .B2(n20446), .ZN(
        n20447) );
  MAOI22D0BWP12T U10913 ( .A1(n21384), .A2(n20447), .B1(n21384), .B2(n20447), 
        .ZN(n20448) );
  MAOI22D0BWP12T U10914 ( .A1(n21536), .A2(n20448), .B1(n21536), .B2(n20448), 
        .ZN(n21537) );
  CKND0BWP12T U10915 ( .I(n21536), .ZN(n20449) );
  MAOI222D0BWP12T U10916 ( .A(n21384), .B(n20449), .C(n20447), .ZN(n21533) );
  NR2D0BWP12T U10917 ( .A1(n22547), .A2(n21717), .ZN(n20450) );
  AOI22D0BWP12T U10918 ( .A1(a[2]), .A2(n20450), .B1(b[13]), .B2(n21738), .ZN(
        n20451) );
  AOI22D0BWP12T U10919 ( .A1(n21720), .A2(b[14]), .B1(n22978), .B2(n21689), 
        .ZN(n20452) );
  OAI211D0BWP12T U10920 ( .A1(n21711), .A2(n23484), .B(n21882), .C(n20452), 
        .ZN(n20453) );
  OAI211D0BWP12T U10921 ( .A1(n23484), .A2(n23559), .B(n20451), .C(n20453), 
        .ZN(n20454) );
  AO21D0BWP12T U10922 ( .A1(n21689), .A2(n21690), .B(n20454), .Z(n20455) );
  CKND0BWP12T U10923 ( .I(n22511), .ZN(n20456) );
  MAOI222D0BWP12T U10924 ( .A(n21688), .B(n20455), .C(n20456), .ZN(n22471) );
  MAOI22D0BWP12T U10925 ( .A1(n21688), .A2(n20455), .B1(n21688), .B2(n20455), 
        .ZN(n20457) );
  MAOI22D0BWP12T U10926 ( .A1(n22511), .A2(n20457), .B1(n22511), .B2(n20457), 
        .ZN(n23304) );
  AOI22D0BWP12T U10927 ( .A1(b[6]), .A2(n21772), .B1(n21781), .B2(n21774), 
        .ZN(n20458) );
  AOI22D0BWP12T U10928 ( .A1(b[7]), .A2(n22291), .B1(b[8]), .B2(n21771), .ZN(
        n20459) );
  CKND2D0BWP12T U10929 ( .A1(n20458), .A2(n20459), .ZN(n20460) );
  MOAI22D0BWP12T U10930 ( .A1(n22267), .A2(n20460), .B1(n22267), .B2(n20460), 
        .ZN(n20461) );
  MAOI22D0BWP12T U10931 ( .A1(n20461), .A2(n20837), .B1(n20461), .B2(n20837), 
        .ZN(n20462) );
  MAOI22D0BWP12T U10932 ( .A1(n21101), .A2(n20462), .B1(n21101), .B2(n20462), 
        .ZN(n21103) );
  CKND0BWP12T U10933 ( .I(n21101), .ZN(n20463) );
  MAOI222D0BWP12T U10934 ( .A(n20461), .B(n20837), .C(n20463), .ZN(n21239) );
  AOI22D0BWP12T U10935 ( .A1(n21748), .A2(b[12]), .B1(n21076), .B2(n21684), 
        .ZN(n20464) );
  CKND2D0BWP12T U10936 ( .A1(b[11]), .A2(n21077), .ZN(n20465) );
  OAI211D0BWP12T U10937 ( .A1(n22675), .A2(n21745), .B(n20464), .C(n20465), 
        .ZN(n20466) );
  MOAI22D0BWP12T U10938 ( .A1(a[14]), .A2(n20466), .B1(a[14]), .B2(n20466), 
        .ZN(n20467) );
  MAOI22D0BWP12T U10939 ( .A1(n21022), .A2(n20467), .B1(n21022), .B2(n20467), 
        .ZN(n20468) );
  MAOI22D0BWP12T U10940 ( .A1(n21145), .A2(n20468), .B1(n21145), .B2(n20468), 
        .ZN(n21146) );
  CKND0BWP12T U10941 ( .I(n21145), .ZN(n20469) );
  MAOI222D0BWP12T U10942 ( .A(n21022), .B(n20467), .C(n20469), .ZN(n21140) );
  NR2D0BWP12T U10943 ( .A1(n21758), .A2(n21710), .ZN(n20470) );
  OAI22D0BWP12T U10944 ( .A1(n21757), .A2(n23498), .B1(n21760), .B2(n22293), 
        .ZN(n20471) );
  AOI211D0BWP12T U10945 ( .A1(n21763), .A2(b[19]), .B(n20470), .C(n20471), 
        .ZN(n20472) );
  MOAI22D0BWP12T U10946 ( .A1(a[11]), .A2(n20472), .B1(a[11]), .B2(n20472), 
        .ZN(n20473) );
  MAOI22D0BWP12T U10947 ( .A1(n21112), .A2(n20473), .B1(n21112), .B2(n20473), 
        .ZN(n20474) );
  MAOI22D0BWP12T U10948 ( .A1(n21257), .A2(n20474), .B1(n21257), .B2(n20474), 
        .ZN(n21258) );
  CKND0BWP12T U10949 ( .I(n21257), .ZN(n20475) );
  MAOI222D0BWP12T U10950 ( .A(n21112), .B(n20475), .C(n20473), .ZN(n21814) );
  NR2D0BWP12T U10951 ( .A1(n21725), .A2(n21700), .ZN(n20476) );
  OAI22D0BWP12T U10952 ( .A1(n21727), .A2(n21944), .B1(n21724), .B2(n22418), 
        .ZN(n20477) );
  AOI211D0BWP12T U10953 ( .A1(b[17]), .A2(n21730), .B(n20476), .C(n20477), 
        .ZN(n20478) );
  MOAI22D0BWP12T U10954 ( .A1(n21966), .A2(n20478), .B1(n21966), .B2(n20478), 
        .ZN(n20479) );
  CKND0BWP12T U10955 ( .I(n21389), .ZN(n20480) );
  MAOI222D0BWP12T U10956 ( .A(n21283), .B(n20479), .C(n20480), .ZN(n21385) );
  MAOI22D0BWP12T U10957 ( .A1(n21283), .A2(n20479), .B1(n21283), .B2(n20479), 
        .ZN(n20481) );
  MAOI22D0BWP12T U10958 ( .A1(n21389), .A2(n20481), .B1(n21389), .B2(n20481), 
        .ZN(n21390) );
  NR2D0BWP12T U10959 ( .A1(n21732), .A2(n21549), .ZN(n20482) );
  OAI22D0BWP12T U10960 ( .A1(n21731), .A2(n22150), .B1(n21734), .B2(n21932), 
        .ZN(n20483) );
  AOI211D0BWP12T U10961 ( .A1(b[24]), .A2(n21737), .B(n20482), .C(n20483), 
        .ZN(n20484) );
  MOAI22D0BWP12T U10962 ( .A1(a[5]), .A2(n20484), .B1(a[5]), .B2(n20484), .ZN(
        n20485) );
  MAOI22D0BWP12T U10963 ( .A1(n21380), .A2(n20485), .B1(n21380), .B2(n20485), 
        .ZN(n20486) );
  MAOI22D0BWP12T U10964 ( .A1(n21533), .A2(n20486), .B1(n21533), .B2(n20486), 
        .ZN(n21534) );
  CKND0BWP12T U10965 ( .I(n21533), .ZN(n20487) );
  MAOI222D0BWP12T U10966 ( .A(n21380), .B(n20487), .C(n20485), .ZN(n21523) );
  NR2D0BWP12T U10967 ( .A1(n21717), .A2(n21753), .ZN(n20488) );
  OAI22D0BWP12T U10968 ( .A1(n21750), .A2(n21716), .B1(n23484), .B2(n21868), 
        .ZN(n20489) );
  NR3D0BWP12T U10969 ( .A1(n21882), .A2(n20488), .A3(n20489), .ZN(n20490) );
  OAI22D0BWP12T U10970 ( .A1(n21750), .A2(n21711), .B1(n21716), .B2(n21751), 
        .ZN(n20491) );
  IAO21D0BWP12T U10971 ( .A1(n20488), .A2(n20491), .B(a[2]), .ZN(n20492) );
  OAI22D0BWP12T U10972 ( .A1(n22992), .A2(n21751), .B1(n20490), .B2(n20492), 
        .ZN(n20493) );
  CKND0BWP12T U10973 ( .I(n22445), .ZN(n20494) );
  MAOI222D0BWP12T U10974 ( .A(n21694), .B(n20493), .C(n20494), .ZN(n22410) );
  MAOI22D0BWP12T U10975 ( .A1(n21694), .A2(n20493), .B1(n21694), .B2(n20493), 
        .ZN(n20495) );
  MAOI22D0BWP12T U10976 ( .A1(n22445), .A2(n20495), .B1(n22445), .B2(n20495), 
        .ZN(n23331) );
  AOI22D0BWP12T U10977 ( .A1(b[7]), .A2(n21772), .B1(n21623), .B2(n21774), 
        .ZN(n20496) );
  AOI22D0BWP12T U10978 ( .A1(b[8]), .A2(n22291), .B1(b[9]), .B2(n21771), .ZN(
        n20497) );
  CKND2D0BWP12T U10979 ( .A1(n20496), .A2(n20497), .ZN(n20498) );
  MOAI22D0BWP12T U10980 ( .A1(n22267), .A2(n20498), .B1(n22267), .B2(n20498), 
        .ZN(n20499) );
  MAOI22D0BWP12T U10981 ( .A1(n21100), .A2(n20499), .B1(n21100), .B2(n20499), 
        .ZN(n20500) );
  MAOI22D0BWP12T U10982 ( .A1(n21239), .A2(n20500), .B1(n21239), .B2(n20500), 
        .ZN(n21217) );
  CKND0BWP12T U10983 ( .I(n21239), .ZN(n20501) );
  MAOI222D0BWP12T U10984 ( .A(n21100), .B(n20499), .C(n20501), .ZN(n21829) );
  OAI22D0BWP12T U10985 ( .A1(n22612), .A2(n21742), .B1(n21745), .B2(n21887), 
        .ZN(n20502) );
  OAI22D0BWP12T U10986 ( .A1(n21934), .A2(n21072), .B1(n21743), .B2(n21595), 
        .ZN(n20503) );
  NR2D0BWP12T U10987 ( .A1(n20502), .A2(n20503), .ZN(n20504) );
  MOAI22D0BWP12T U10988 ( .A1(n21933), .A2(n20504), .B1(n21933), .B2(n20504), 
        .ZN(n20505) );
  MAOI22D0BWP12T U10989 ( .A1(n21018), .A2(n20505), .B1(n21018), .B2(n20505), 
        .ZN(n20506) );
  MAOI22D0BWP12T U10990 ( .A1(n21140), .A2(n20506), .B1(n21140), .B2(n20506), 
        .ZN(n21141) );
  CKND0BWP12T U10991 ( .I(n21140), .ZN(n20507) );
  MAOI222D0BWP12T U10992 ( .A(n21018), .B(n20507), .C(n20505), .ZN(n21138) );
  NR2D0BWP12T U10993 ( .A1(n21758), .A2(n21565), .ZN(n20508) );
  OAI22D0BWP12T U10994 ( .A1(n21757), .A2(n22293), .B1(n21760), .B2(n21886), 
        .ZN(n20509) );
  AOI211D0BWP12T U10995 ( .A1(b[20]), .A2(n21763), .B(n20508), .C(n20509), 
        .ZN(n20510) );
  MOAI22D0BWP12T U10996 ( .A1(a[11]), .A2(n20510), .B1(a[11]), .B2(n20510), 
        .ZN(n20511) );
  MAOI22D0BWP12T U10997 ( .A1(n21814), .A2(n20511), .B1(n21814), .B2(n20511), 
        .ZN(n20512) );
  MAOI22D0BWP12T U10998 ( .A1(n21252), .A2(n20512), .B1(n21252), .B2(n20512), 
        .ZN(n21253) );
  CKND0BWP12T U10999 ( .I(n21814), .ZN(n20513) );
  MAOI222D0BWP12T U11000 ( .A(n21252), .B(n20513), .C(n20511), .ZN(n21819) );
  AOI22D0BWP12T U11001 ( .A1(b[15]), .A2(n21346), .B1(n21347), .B2(n21585), 
        .ZN(n20514) );
  CKND2D0BWP12T U11002 ( .A1(n21730), .A2(b[14]), .ZN(n20515) );
  OAI211D0BWP12T U11003 ( .A1(n21753), .A2(n21727), .B(n20514), .C(n20515), 
        .ZN(n20516) );
  MOAI22D0BWP12T U11004 ( .A1(a[8]), .A2(n20516), .B1(a[8]), .B2(n20516), .ZN(
        n20517) );
  CKND0BWP12T U11005 ( .I(n21401), .ZN(n20518) );
  MAOI222D0BWP12T U11006 ( .A(n21289), .B(n20517), .C(n20518), .ZN(n21396) );
  MAOI22D0BWP12T U11007 ( .A1(n20517), .A2(n21289), .B1(n20517), .B2(n21289), 
        .ZN(n20519) );
  MAOI22D0BWP12T U11008 ( .A1(n21401), .A2(n20519), .B1(n21401), .B2(n20519), 
        .ZN(n21402) );
  CKND0BWP12T U11009 ( .I(n23349), .ZN(n20520) );
  AOI21D0BWP12T U11010 ( .A1(n22937), .A2(n22936), .B(n20520), .ZN(n22916) );
  NR2D0BWP12T U11011 ( .A1(n22220), .A2(n22100), .ZN(n20521) );
  OAI22D0BWP12T U11012 ( .A1(n22223), .A2(n22721), .B1(n22224), .B2(n22865), 
        .ZN(n20522) );
  AOI211D0BWP12T U11013 ( .A1(n22198), .A2(n22227), .B(n20521), .C(n20522), 
        .ZN(n22402) );
  IOA21D0BWP12T U11014 ( .A1(n22465), .A2(n22433), .B(n23086), .ZN(n22394) );
  NR2D0BWP12T U11015 ( .A1(n21732), .A2(n21726), .ZN(n20523) );
  OAI22D0BWP12T U11016 ( .A1(n21731), .A2(n22088), .B1(n21734), .B2(n21556), 
        .ZN(n20524) );
  AOI211D0BWP12T U11017 ( .A1(b[25]), .A2(n21737), .B(n20523), .C(n20524), 
        .ZN(n20525) );
  MOAI22D0BWP12T U11018 ( .A1(a[5]), .A2(n20525), .B1(a[5]), .B2(n20525), .ZN(
        n20526) );
  MAOI22D0BWP12T U11019 ( .A1(n21378), .A2(n20526), .B1(n21378), .B2(n20526), 
        .ZN(n20527) );
  MAOI22D0BWP12T U11020 ( .A1(n21523), .A2(n20527), .B1(n21523), .B2(n20527), 
        .ZN(n21524) );
  CKND0BWP12T U11021 ( .I(n21523), .ZN(n20528) );
  MAOI222D0BWP12T U11022 ( .A(n21378), .B(n20528), .C(n20526), .ZN(n21515) );
  NR2D0BWP12T U11023 ( .A1(n21717), .A2(n21944), .ZN(n20529) );
  MAOI22D0BWP12T U11024 ( .A1(b[18]), .A2(n22977), .B1(n21716), .B2(n23498), 
        .ZN(n20530) );
  OAI21D0BWP12T U11025 ( .A1(n21711), .A2(n21744), .B(n20530), .ZN(n20531) );
  OAI22D0BWP12T U11026 ( .A1(n21716), .A2(n21744), .B1(n21711), .B2(n23498), 
        .ZN(n20532) );
  OAI21D0BWP12T U11027 ( .A1(n20529), .A2(n20531), .B(a[2]), .ZN(n20533) );
  OAI31D0BWP12T U11028 ( .A1(n20529), .A2(a[2]), .A3(n20532), .B(n20533), .ZN(
        n20534) );
  CKND0BWP12T U11029 ( .I(n22340), .ZN(n20535) );
  MAOI222D0BWP12T U11030 ( .A(n20534), .B(n21571), .C(n20535), .ZN(n22315) );
  MAOI22D0BWP12T U11031 ( .A1(n22340), .A2(n21571), .B1(n22340), .B2(n21571), 
        .ZN(n20536) );
  MAOI22D0BWP12T U11032 ( .A1(n20534), .A2(n20536), .B1(n20534), .B2(n20536), 
        .ZN(n23314) );
  OAI22D0BWP12T U11033 ( .A1(n21934), .A2(n21742), .B1(n22612), .B2(n21745), 
        .ZN(n20537) );
  OAI22D0BWP12T U11034 ( .A1(n22547), .A2(n21072), .B1(n21743), .B2(n21765), 
        .ZN(n20538) );
  NR2D0BWP12T U11035 ( .A1(n20537), .A2(n20538), .ZN(n20539) );
  MOAI22D0BWP12T U11036 ( .A1(n21933), .A2(n20539), .B1(n21933), .B2(n20539), 
        .ZN(n20540) );
  MAOI22D0BWP12T U11037 ( .A1(n21014), .A2(n20540), .B1(n21014), .B2(n20540), 
        .ZN(n20541) );
  MAOI22D0BWP12T U11038 ( .A1(n21138), .A2(n20541), .B1(n21138), .B2(n20541), 
        .ZN(n21139) );
  CKND0BWP12T U11039 ( .I(n21138), .ZN(n20542) );
  MAOI222D0BWP12T U11040 ( .A(n21014), .B(n20542), .C(n20540), .ZN(n21130) );
  AOI22D0BWP12T U11041 ( .A1(b[7]), .A2(n21779), .B1(n21780), .B2(n21638), 
        .ZN(n20543) );
  CKND2D0BWP12T U11042 ( .A1(b[6]), .A2(n21778), .ZN(n20544) );
  OAI211D0BWP12T U11043 ( .A1(n21885), .A2(n21784), .B(n20543), .C(n20544), 
        .ZN(n20545) );
  MOAI22D0BWP12T U11044 ( .A1(a[26]), .A2(n20545), .B1(a[26]), .B2(n20545), 
        .ZN(n20546) );
  MAOI22D0BWP12T U11045 ( .A1(n21232), .A2(n20546), .B1(n21232), .B2(n20546), 
        .ZN(n20547) );
  MAOI22D0BWP12T U11046 ( .A1(n21820), .A2(n20547), .B1(n21820), .B2(n20547), 
        .ZN(n21236) );
  CKND0BWP12T U11047 ( .I(n21820), .ZN(n20548) );
  MAOI222D0BWP12T U11048 ( .A(n21232), .B(n20546), .C(n20548), .ZN(n21825) );
  CKND0BWP12T U11049 ( .I(n21359), .ZN(n20549) );
  NR2D0BWP12T U11050 ( .A1(n21757), .A2(n22741), .ZN(n20550) );
  OAI22D0BWP12T U11051 ( .A1(n22699), .A2(n21760), .B1(n21935), .B2(n21207), 
        .ZN(n20551) );
  AOI211D0BWP12T U11052 ( .A1(n21208), .A2(n21623), .B(n20550), .C(n20551), 
        .ZN(n20552) );
  MOAI22D0BWP12T U11053 ( .A1(a[11]), .A2(n20552), .B1(a[11]), .B2(n20552), 
        .ZN(n20553) );
  MAOI222D0BWP12T U11054 ( .A(n21206), .B(n20549), .C(n20553), .ZN(n21364) );
  MAOI22D0BWP12T U11055 ( .A1(n21359), .A2(n20553), .B1(n21359), .B2(n20553), 
        .ZN(n20554) );
  MAOI22D0BWP12T U11056 ( .A1(n21206), .A2(n20554), .B1(n21206), .B2(n20554), 
        .ZN(n21360) );
  INR2D0BWP12T U11057 ( .A1(n20806), .B1(n20805), .ZN(n21771) );
  AOI22D0BWP12T U11058 ( .A1(b[14]), .A2(n21346), .B1(n21347), .B2(n21689), 
        .ZN(n20555) );
  CKND2D0BWP12T U11059 ( .A1(n21730), .A2(b[13]), .ZN(n20556) );
  OAI211D0BWP12T U11060 ( .A1(n21727), .A2(n23484), .B(n20555), .C(n20556), 
        .ZN(n20557) );
  MOAI22D0BWP12T U11061 ( .A1(a[8]), .A2(n20557), .B1(a[8]), .B2(n20557), .ZN(
        n20558) );
  MAOI22D0BWP12T U11062 ( .A1(n20558), .A2(n21293), .B1(n20558), .B2(n21293), 
        .ZN(n20559) );
  MAOI22D0BWP12T U11063 ( .A1(n21403), .A2(n20559), .B1(n21403), .B2(n20559), 
        .ZN(n21404) );
  CKND0BWP12T U11064 ( .I(n21403), .ZN(n20560) );
  MAOI222D0BWP12T U11065 ( .A(n20558), .B(n21293), .C(n20560), .ZN(n21401) );
  IAO21D0BWP12T U11066 ( .A1(n22917), .A2(n22903), .B(n23496), .ZN(n22881) );
  IAO21D0BWP12T U11067 ( .A1(n22503), .A2(n23167), .B(n23521), .ZN(n22498) );
  CKND2D0BWP12T U11068 ( .A1(n20991), .A2(n20992), .ZN(n20561) );
  MOAI22D0BWP12T U11069 ( .A1(n21750), .A2(n20561), .B1(n21750), .B2(n20561), 
        .ZN(n21751) );
  IOA21D0BWP12T U11070 ( .A1(n22425), .A2(n22394), .B(n21943), .ZN(n22357) );
  IAO21D0BWP12T U11071 ( .A1(n22114), .A2(n22075), .B(n23185), .ZN(n22063) );
  NR2D0BWP12T U11072 ( .A1(n21732), .A2(n21539), .ZN(n20562) );
  OAI22D0BWP12T U11073 ( .A1(n21731), .A2(n22032), .B1(n21734), .B2(n22150), 
        .ZN(n20563) );
  AOI211D0BWP12T U11074 ( .A1(b[26]), .A2(n21737), .B(n20562), .C(n20563), 
        .ZN(n20564) );
  MOAI22D0BWP12T U11075 ( .A1(a[5]), .A2(n20564), .B1(a[5]), .B2(n20564), .ZN(
        n20565) );
  MAOI22D0BWP12T U11076 ( .A1(n21373), .A2(n20565), .B1(n21373), .B2(n20565), 
        .ZN(n20566) );
  MAOI22D0BWP12T U11077 ( .A1(n21515), .A2(n20566), .B1(n21515), .B2(n20566), 
        .ZN(n21516) );
  CKND0BWP12T U11078 ( .I(n21515), .ZN(n20567) );
  MAOI222D0BWP12T U11079 ( .A(n21373), .B(n20567), .C(n20565), .ZN(n21833) );
  IAO21D0BWP12T U11080 ( .A1(n21984), .A2(n21983), .B(n21947), .ZN(n23045) );
  AOI22D0BWP12T U11081 ( .A1(n22447), .A2(n22236), .B1(n22174), .B2(n22235), 
        .ZN(n20568) );
  OAI21D0BWP12T U11082 ( .A1(n22220), .A2(n22239), .B(n20568), .ZN(n20569) );
  AOI21D0BWP12T U11083 ( .A1(n22687), .A2(n22227), .B(n20569), .ZN(n23456) );
  NR2D0BWP12T U11084 ( .A1(n21717), .A2(n22293), .ZN(n20570) );
  OAI22D0BWP12T U11085 ( .A1(n21716), .A2(n21886), .B1(n23498), .B2(n21868), 
        .ZN(n20571) );
  NR3D0BWP12T U11086 ( .A1(n21882), .A2(n20570), .A3(n20571), .ZN(n20572) );
  OAI22D0BWP12T U11087 ( .A1(n21716), .A2(n21565), .B1(n21711), .B2(n21886), 
        .ZN(n20573) );
  IAO21D0BWP12T U11088 ( .A1(n20570), .A2(n20573), .B(a[2]), .ZN(n20574) );
  OAI22D0BWP12T U11089 ( .A1(n22992), .A2(n21565), .B1(n20572), .B2(n20574), 
        .ZN(n20575) );
  CKND0BWP12T U11090 ( .I(n22279), .ZN(n20576) );
  MAOI222D0BWP12T U11091 ( .A(n21564), .B(n20575), .C(n20576), .ZN(n22230) );
  MAOI22D0BWP12T U11092 ( .A1(n21564), .A2(n20575), .B1(n21564), .B2(n20575), 
        .ZN(n20577) );
  MAOI22D0BWP12T U11093 ( .A1(n22279), .A2(n20577), .B1(n22279), .B2(n20577), 
        .ZN(n23311) );
  AOI21D0BWP12T U11094 ( .A1(n20899), .A2(n20900), .B(n20898), .ZN(n20578) );
  INR2D0BWP12T U11095 ( .A1(n20963), .B1(n20962), .ZN(n20579) );
  AOI31D0BWP12T U11096 ( .A1(a[20]), .A2(n20909), .A3(n20967), .B(n20579), 
        .ZN(n20580) );
  NR2D0BWP12T U11097 ( .A1(n21766), .A2(n21667), .ZN(n20581) );
  OAI22D0BWP12T U11098 ( .A1(n23017), .A2(n21764), .B1(n22806), .B2(n21767), 
        .ZN(n20582) );
  AOI211D0BWP12T U11099 ( .A1(b[2]), .A2(n21770), .B(n20581), .C(n20582), .ZN(
        n20583) );
  MOAI22D0BWP12T U11100 ( .A1(a[20]), .A2(n20583), .B1(a[20]), .B2(n20583), 
        .ZN(n20584) );
  MAOI22D0BWP12T U11101 ( .A1(n20580), .A2(n20584), .B1(n20580), .B2(n20584), 
        .ZN(n20585) );
  MAOI22D0BWP12T U11102 ( .A1(n20578), .A2(n20585), .B1(n20578), .B2(n20585), 
        .ZN(n21029) );
  CKND0BWP12T U11103 ( .I(n20580), .ZN(n20586) );
  MAOI222D0BWP12T U11104 ( .A(n20578), .B(n20586), .C(n20584), .ZN(n20953) );
  NR2D0BWP12T U11105 ( .A1(n21743), .A2(n21700), .ZN(n20587) );
  OAI22D0BWP12T U11106 ( .A1(n21745), .A2(n21750), .B1(n22418), .B2(n21742), 
        .ZN(n20588) );
  AOI211D0BWP12T U11107 ( .A1(n21748), .A2(b[19]), .B(n20587), .C(n20588), 
        .ZN(n20589) );
  MOAI22D0BWP12T U11108 ( .A1(n21933), .A2(n20589), .B1(n21933), .B2(n20589), 
        .ZN(n20590) );
  MAOI22D0BWP12T U11109 ( .A1(n21248), .A2(n20590), .B1(n21248), .B2(n20590), 
        .ZN(n20591) );
  MAOI22D0BWP12T U11110 ( .A1(n21809), .A2(n20591), .B1(n21809), .B2(n20591), 
        .ZN(n21252) );
  CKND0BWP12T U11111 ( .I(n21809), .ZN(n20592) );
  MAOI222D0BWP12T U11112 ( .A(n21248), .B(n20592), .C(n20590), .ZN(n21810) );
  OAI22D0BWP12T U11113 ( .A1(n21757), .A2(n21934), .B1(n22612), .B2(n21207), 
        .ZN(n20593) );
  OAI22D0BWP12T U11114 ( .A1(n22547), .A2(n21760), .B1(n21758), .B2(n21765), 
        .ZN(n20594) );
  NR2D0BWP12T U11115 ( .A1(n20593), .A2(n20594), .ZN(n20595) );
  MOAI22D0BWP12T U11116 ( .A1(a[11]), .A2(n20595), .B1(a[11]), .B2(n20595), 
        .ZN(n20596) );
  MAOI22D0BWP12T U11117 ( .A1(n21148), .A2(n20596), .B1(n21148), .B2(n20596), 
        .ZN(n20597) );
  MAOI22D0BWP12T U11118 ( .A1(n21286), .A2(n20597), .B1(n21286), .B2(n20597), 
        .ZN(n21287) );
  CKND0BWP12T U11119 ( .I(n21286), .ZN(n20598) );
  MAOI222D0BWP12T U11120 ( .A(n21148), .B(n20598), .C(n20596), .ZN(n21284) );
  OAI22D0BWP12T U11121 ( .A1(a[16]), .A2(n22605), .B1(a[13]), .B2(b[0]), .ZN(
        n20599) );
  OAI22D0BWP12T U11122 ( .A1(n22864), .A2(n20599), .B1(n22574), .B2(n22867), 
        .ZN(n22690) );
  NR2D0BWP12T U11123 ( .A1(n21725), .A2(n21565), .ZN(n20600) );
  OAI22D0BWP12T U11124 ( .A1(n21727), .A2(n21886), .B1(n21724), .B2(n22293), 
        .ZN(n20601) );
  AOI211D0BWP12T U11125 ( .A1(b[20]), .A2(n21730), .B(n20600), .C(n20601), 
        .ZN(n20602) );
  MOAI22D0BWP12T U11126 ( .A1(n21966), .A2(n20602), .B1(n21966), .B2(n20602), 
        .ZN(n20603) );
  CKND0BWP12T U11127 ( .I(n21379), .ZN(n20604) );
  MAOI222D0BWP12T U11128 ( .A(n21265), .B(n20603), .C(n20604), .ZN(n21377) );
  MAOI22D0BWP12T U11129 ( .A1(n21265), .A2(n20603), .B1(n21265), .B2(n20603), 
        .ZN(n20605) );
  MAOI22D0BWP12T U11130 ( .A1(n21379), .A2(n20605), .B1(n21379), .B2(n20605), 
        .ZN(n21380) );
  NR3D0BWP12T U11131 ( .A1(n23222), .A2(n23223), .A3(n23221), .ZN(n20606) );
  ND4D0BWP12T U11132 ( .A1(n23225), .A2(n23226), .A3(n23224), .A4(n20606), 
        .ZN(n23411) );
  IOA21D0BWP12T U11133 ( .A1(n22990), .A2(n22970), .B(n23347), .ZN(n22929) );
  OA21D0BWP12T U11134 ( .A1(n22901), .A2(n22916), .B(n23350), .Z(n22871) );
  IOA21D0BWP12T U11135 ( .A1(n22560), .A2(n22561), .B(n22549), .ZN(n22525) );
  IOA21D0BWP12T U11136 ( .A1(n22558), .A2(n23518), .B(n22526), .ZN(n22470) );
  OAI21D0BWP12T U11137 ( .A1(n22497), .A2(n22469), .B(n23084), .ZN(n22433) );
  IAO21D0BWP12T U11138 ( .A1(n21984), .A2(n21985), .B(n21947), .ZN(n23042) );
  NR2D0BWP12T U11139 ( .A1(n21732), .A2(n21535), .ZN(n20607) );
  OAI22D0BWP12T U11140 ( .A1(n21731), .A2(n23490), .B1(n21734), .B2(n22088), 
        .ZN(n20608) );
  AOI211D0BWP12T U11141 ( .A1(b[27]), .A2(n21737), .B(n20607), .C(n20608), 
        .ZN(n20609) );
  MOAI22D0BWP12T U11142 ( .A1(a[5]), .A2(n20609), .B1(a[5]), .B2(n20609), .ZN(
        n20610) );
  MAOI22D0BWP12T U11143 ( .A1(n21368), .A2(n20610), .B1(n21368), .B2(n20610), 
        .ZN(n20611) );
  MAOI22D0BWP12T U11144 ( .A1(n21833), .A2(n20611), .B1(n21833), .B2(n20611), 
        .ZN(n21506) );
  CKND0BWP12T U11145 ( .I(n21833), .ZN(n20612) );
  MAOI222D0BWP12T U11146 ( .A(n21368), .B(n20612), .C(n20610), .ZN(n21834) );
  CKND0BWP12T U11147 ( .I(n22478), .ZN(n20613) );
  AOI21D0BWP12T U11148 ( .A1(n22806), .A2(n20613), .B(n22197), .ZN(n20614) );
  AOI21D0BWP12T U11149 ( .A1(n22479), .A2(n23008), .B(n20614), .ZN(n23280) );
  CKND0BWP12T U11150 ( .I(n21781), .ZN(n20615) );
  OAI22D0BWP12T U11151 ( .A1(n23370), .A2(n21645), .B1(n22992), .B2(n20615), 
        .ZN(n20616) );
  NR2D0BWP12T U11152 ( .A1(n21717), .A2(n21935), .ZN(n20617) );
  OAI22D0BWP12T U11153 ( .A1(n21711), .A2(n22741), .B1(n21716), .B2(n20615), 
        .ZN(n20618) );
  CKND0BWP12T U11154 ( .I(n20617), .ZN(n20619) );
  OAI32D0BWP12T U11155 ( .A1(n20617), .A2(a[2]), .A3(n20618), .B1(n21882), 
        .B2(n20619), .ZN(n20620) );
  AO211D0BWP12T U11156 ( .A1(b[8]), .A2(n21651), .B(n20616), .C(n20620), .Z(
        n20621) );
  CKND0BWP12T U11157 ( .I(n22730), .ZN(n20622) );
  MAOI222D0BWP12T U11158 ( .A(n21631), .B(n20621), .C(n20622), .ZN(n22695) );
  MAOI22D0BWP12T U11159 ( .A1(n21631), .A2(n20621), .B1(n21631), .B2(n20621), 
        .ZN(n20623) );
  MAOI22D0BWP12T U11160 ( .A1(n22730), .A2(n20623), .B1(n22730), .B2(n20623), 
        .ZN(n23328) );
  IOA21D0BWP12T U11161 ( .A1(n22353), .A2(n22354), .B(n22341), .ZN(n22329) );
  NR2D0BWP12T U11162 ( .A1(n21717), .A2(n21932), .ZN(n20624) );
  MAOI22D0BWP12T U11163 ( .A1(b[22]), .A2(n22977), .B1(n21716), .B2(n21556), 
        .ZN(n20625) );
  OAI21D0BWP12T U11164 ( .A1(n21711), .A2(n21555), .B(n20625), .ZN(n20626) );
  OAI22D0BWP12T U11165 ( .A1(n21716), .A2(n21555), .B1(n21711), .B2(n21556), 
        .ZN(n20627) );
  OAI21D0BWP12T U11166 ( .A1(n20624), .A2(n20626), .B(a[2]), .ZN(n20628) );
  OAI31D0BWP12T U11167 ( .A1(n20624), .A2(a[2]), .A3(n20627), .B(n20628), .ZN(
        n20629) );
  CKND0BWP12T U11168 ( .I(n22184), .ZN(n20630) );
  MAOI222D0BWP12T U11169 ( .A(n21554), .B(n20629), .C(n20630), .ZN(n22147) );
  MAOI22D0BWP12T U11170 ( .A1(n20629), .A2(n21554), .B1(n20629), .B2(n21554), 
        .ZN(n20631) );
  MAOI22D0BWP12T U11171 ( .A1(n22184), .A2(n20631), .B1(n22184), .B2(n20631), 
        .ZN(n23312) );
  MOAI22D0BWP12T U11172 ( .A1(n20985), .A2(n20984), .B1(n20985), .B2(n20984), 
        .ZN(n21050) );
  AOI22D0BWP12T U11173 ( .A1(b[15]), .A2(n21748), .B1(n21076), .B2(n21689), 
        .ZN(n20632) );
  CKND2D0BWP12T U11174 ( .A1(b[14]), .A2(n21077), .ZN(n20633) );
  OAI211D0BWP12T U11175 ( .A1(n21934), .A2(n21745), .B(n20632), .C(n20633), 
        .ZN(n20634) );
  MOAI22D0BWP12T U11176 ( .A1(a[14]), .A2(n20634), .B1(a[14]), .B2(n20634), 
        .ZN(n20635) );
  CKND0BWP12T U11177 ( .I(n21130), .ZN(n20636) );
  MAOI222D0BWP12T U11178 ( .A(n20635), .B(n21010), .C(n20636), .ZN(n21128) );
  MAOI22D0BWP12T U11179 ( .A1(n21010), .A2(n20635), .B1(n21010), .B2(n20635), 
        .ZN(n20637) );
  MAOI22D0BWP12T U11180 ( .A1(n21130), .A2(n20637), .B1(n21130), .B2(n20637), 
        .ZN(n21131) );
  NR2D0BWP12T U11181 ( .A1(n22699), .A2(n21777), .ZN(n20638) );
  OAI22D0BWP12T U11182 ( .A1(n22675), .A2(n21238), .B1(n21678), .B2(n21237), 
        .ZN(n20639) );
  AOI211D0BWP12T U11183 ( .A1(n21772), .A2(b[8]), .B(n20638), .C(n20639), .ZN(
        n20640) );
  MOAI22D0BWP12T U11184 ( .A1(a[23]), .A2(n20640), .B1(a[23]), .B2(n20640), 
        .ZN(n20641) );
  MAOI22D0BWP12T U11185 ( .A1(n21236), .A2(n20641), .B1(n21236), .B2(n20641), 
        .ZN(n20642) );
  MAOI22D0BWP12T U11186 ( .A1(n21829), .A2(n20642), .B1(n21829), .B2(n20642), 
        .ZN(n21826) );
  CKND0BWP12T U11187 ( .I(n21829), .ZN(n20643) );
  MAOI222D0BWP12T U11188 ( .A(n21236), .B(n20643), .C(n20641), .ZN(n21830) );
  NR2D0BWP12T U11189 ( .A1(n21760), .A2(n21887), .ZN(n20644) );
  OAI22D0BWP12T U11190 ( .A1(n22675), .A2(n21757), .B1(n22699), .B2(n21207), 
        .ZN(n20645) );
  AOI211D0BWP12T U11191 ( .A1(n21208), .A2(n21773), .B(n20644), .C(n20645), 
        .ZN(n20646) );
  MOAI22D0BWP12T U11192 ( .A1(a[11]), .A2(n20646), .B1(a[11]), .B2(n20646), 
        .ZN(n20647) );
  CKND0BWP12T U11193 ( .I(n21366), .ZN(n20648) );
  MAOI222D0BWP12T U11194 ( .A(n21212), .B(n20647), .C(n20648), .ZN(n21290) );
  MAOI22D0BWP12T U11195 ( .A1(n21366), .A2(n20647), .B1(n21366), .B2(n20647), 
        .ZN(n20649) );
  MAOI22D0BWP12T U11196 ( .A1(n21212), .A2(n20649), .B1(n21212), .B2(n20649), 
        .ZN(n21367) );
  NR2D0BWP12T U11197 ( .A1(n21725), .A2(n21555), .ZN(n20650) );
  OAI22D0BWP12T U11198 ( .A1(n21727), .A2(n21556), .B1(n21724), .B2(n21932), 
        .ZN(n20651) );
  AOI211D0BWP12T U11199 ( .A1(b[22]), .A2(n21730), .B(n20650), .C(n20651), 
        .ZN(n20652) );
  MOAI22D0BWP12T U11200 ( .A1(n21966), .A2(n20652), .B1(n21966), .B2(n20652), 
        .ZN(n20653) );
  MAOI22D0BWP12T U11201 ( .A1(n21258), .A2(n20653), .B1(n21258), .B2(n20653), 
        .ZN(n20654) );
  MAOI22D0BWP12T U11202 ( .A1(n21372), .A2(n20654), .B1(n21372), .B2(n20654), 
        .ZN(n21373) );
  CKND0BWP12T U11203 ( .I(n21372), .ZN(n20655) );
  MAOI222D0BWP12T U11204 ( .A(n21258), .B(n20655), .C(n20653), .ZN(n21832) );
  IOA21D0BWP12T U11205 ( .A1(n22937), .A2(n22929), .B(n23349), .ZN(n22895) );
  AO21D0BWP12T U11206 ( .A1(n22886), .A2(n22881), .B(n23477), .Z(n22837) );
  OAI22D0BWP12T U11207 ( .A1(b[0]), .A2(a[23]), .B1(n22605), .B2(a[26]), .ZN(
        n20656) );
  OAI22D0BWP12T U11208 ( .A1(n22864), .A2(n20656), .B1(n22867), .B2(n22218), 
        .ZN(n22362) );
  MOAI22D0BWP12T U11209 ( .A1(a[15]), .A2(b[15]), .B1(n22525), .B2(n23167), 
        .ZN(n22500) );
  NR2D0BWP12T U11210 ( .A1(n21732), .A2(n21573), .ZN(n20657) );
  OAI22D0BWP12T U11211 ( .A1(n21731), .A2(n22418), .B1(n21734), .B2(n21753), 
        .ZN(n20658) );
  AOI211D0BWP12T U11212 ( .A1(b[17]), .A2(n21737), .B(n20657), .C(n20658), 
        .ZN(n20659) );
  MOAI22D0BWP12T U11213 ( .A1(a[5]), .A2(n20659), .B1(a[5]), .B2(n20659), .ZN(
        n20660) );
  CKND0BWP12T U11214 ( .I(n21566), .ZN(n20661) );
  MAOI222D0BWP12T U11215 ( .A(n21404), .B(n20660), .C(n20661), .ZN(n21561) );
  MAOI22D0BWP12T U11216 ( .A1(n21404), .A2(n20660), .B1(n21404), .B2(n20660), 
        .ZN(n20662) );
  MAOI22D0BWP12T U11217 ( .A1(n21566), .A2(n20662), .B1(n21566), .B2(n20662), 
        .ZN(n21567) );
  MOAI22D0BWP12T U11218 ( .A1(a[19]), .A2(b[19]), .B1(n22357), .B2(n23099), 
        .ZN(n22354) );
  IAO21D0BWP12T U11219 ( .A1(n22070), .A2(n22063), .B(n23170), .ZN(n21989) );
  IAO21D0BWP12T U11220 ( .A1(n21988), .A2(n23169), .B(n23517), .ZN(n21951) );
  IAO21D0BWP12T U11221 ( .A1(n23044), .A2(n23042), .B(n23541), .ZN(n23062) );
  IOA21D0BWP12T U11222 ( .A1(b[11]), .A2(n22642), .B(n22610), .ZN(n20663) );
  MAOI22D0BWP12T U11223 ( .A1(n22611), .A2(n20663), .B1(n22611), .B2(n20663), 
        .ZN(n23142) );
  CKND2D0BWP12T U11224 ( .A1(n21720), .A2(b[13]), .ZN(n20664) );
  OAI22D0BWP12T U11225 ( .A1(n22612), .A2(n21645), .B1(n21882), .B2(n20664), 
        .ZN(n20665) );
  OAI211D0BWP12T U11226 ( .A1(n22547), .A2(n21711), .B(n21882), .C(n20664), 
        .ZN(n20666) );
  NR2D0BWP12T U11227 ( .A1(n21765), .A2(n21716), .ZN(n20667) );
  OAI22D0BWP12T U11228 ( .A1(n20667), .A2(n20666), .B1(n21765), .B2(n22992), 
        .ZN(n20668) );
  AO211D0BWP12T U11229 ( .A1(b[14]), .A2(n21651), .B(n20665), .C(n20668), .Z(
        n20669) );
  CKND0BWP12T U11230 ( .I(n22548), .ZN(n20670) );
  MAOI222D0BWP12T U11231 ( .A(n21593), .B(n20669), .C(n20670), .ZN(n22511) );
  MAOI22D0BWP12T U11232 ( .A1(n21593), .A2(n20669), .B1(n21593), .B2(n20669), 
        .ZN(n20671) );
  MAOI22D0BWP12T U11233 ( .A1(n22548), .A2(n20671), .B1(n22548), .B2(n20671), 
        .ZN(n23302) );
  OA222D0BWP12T U11234 ( .A1(n22223), .A2(n22100), .B1(n22242), .B2(n23516), 
        .C1(n22168), .C2(n22177), .Z(n23424) );
  OAI21D0BWP12T U11235 ( .A1(n22352), .A2(n22334), .B(n22341), .ZN(n22304) );
  NR2D0BWP12T U11236 ( .A1(n21717), .A2(n22150), .ZN(n20672) );
  MAOI22D0BWP12T U11237 ( .A1(b[24]), .A2(n22977), .B1(n21716), .B2(n22088), 
        .ZN(n20673) );
  OAI21D0BWP12T U11238 ( .A1(n21711), .A2(n21726), .B(n20673), .ZN(n20674) );
  OAI22D0BWP12T U11239 ( .A1(n21716), .A2(n21726), .B1(n21711), .B2(n22088), 
        .ZN(n20675) );
  OAI21D0BWP12T U11240 ( .A1(n20672), .A2(n20674), .B(a[2]), .ZN(n20676) );
  OAI31D0BWP12T U11241 ( .A1(n20672), .A2(a[2]), .A3(n20675), .B(n20676), .ZN(
        n20677) );
  CKND0BWP12T U11242 ( .I(n22086), .ZN(n20678) );
  MAOI222D0BWP12T U11243 ( .A(n21545), .B(n20677), .C(n20678), .ZN(n22055) );
  MAOI22D0BWP12T U11244 ( .A1(n20677), .A2(n21545), .B1(n20677), .B2(n21545), 
        .ZN(n20679) );
  MAOI22D0BWP12T U11245 ( .A1(n22086), .A2(n20679), .B1(n22086), .B2(n20679), 
        .ZN(n23326) );
  AOI22D0BWP12T U11246 ( .A1(n22686), .A2(n23027), .B1(n22712), .B2(n22945), 
        .ZN(n20680) );
  CKND2D0BWP12T U11247 ( .A1(n22694), .A2(n22668), .ZN(n20681) );
  AOI22D0BWP12T U11248 ( .A1(n23658), .A2(n23332), .B1(n22674), .B2(n22673), 
        .ZN(n20682) );
  MOAI22D0BWP12T U11249 ( .A1(n23647), .A2(n23522), .B1(n22974), .B2(n23480), 
        .ZN(n20683) );
  AOI211D0BWP12T U11250 ( .A1(n22677), .A2(n22676), .B(n23037), .C(n20683), 
        .ZN(n20684) );
  OAI211D0BWP12T U11251 ( .A1(n22887), .A2(n23246), .B(n20682), .C(n20684), 
        .ZN(n20685) );
  CKND2D0BWP12T U11252 ( .A1(n22700), .A2(n22670), .ZN(n20686) );
  AOI32D0BWP12T U11253 ( .A1(n22812), .A2(n20686), .A3(n22675), .B1(n23030), 
        .B2(n20686), .ZN(n20687) );
  AOI22D0BWP12T U11254 ( .A1(a[10]), .A2(n20687), .B1(n23281), .B2(n22671), 
        .ZN(n20688) );
  MAOI22D0BWP12T U11255 ( .A1(n22848), .A2(n23238), .B1(n22737), .B2(n23426), 
        .ZN(n20689) );
  OAI211D0BWP12T U11256 ( .A1(n22948), .A2(n23129), .B(n20688), .C(n20689), 
        .ZN(n20690) );
  AOI211D0BWP12T U11257 ( .A1(n22945), .A2(n22678), .B(n20685), .C(n20690), 
        .ZN(n20691) );
  AOI22D0BWP12T U11258 ( .A1(n23027), .A2(n22681), .B1(n23601), .B2(n23631), 
        .ZN(n20692) );
  OAI211D0BWP12T U11259 ( .A1(n20680), .A2(n20681), .B(n20691), .C(n20692), 
        .ZN(result[10]) );
  CKND0BWP12T U11260 ( .I(n20845), .ZN(n20693) );
  NR3D0BWP12T U11261 ( .A1(n22087), .A2(n20836), .A3(n20835), .ZN(n20694) );
  AOI21D0BWP12T U11262 ( .A1(n20846), .A2(n20693), .B(n20694), .ZN(n20695) );
  AO21D0BWP12T U11263 ( .A1(n20824), .A2(n20825), .B(n20823), .Z(n20696) );
  OAI22D0BWP12T U11264 ( .A1(n21784), .A2(n22342), .B1(n22806), .B2(n20826), 
        .ZN(n20697) );
  OAI22D0BWP12T U11265 ( .A1(n23017), .A2(n20828), .B1(n21667), .B2(n20827), 
        .ZN(n20698) );
  NR2D0BWP12T U11266 ( .A1(n20697), .A2(n20698), .ZN(n20699) );
  MOAI22D0BWP12T U11267 ( .A1(n22087), .A2(n20699), .B1(n22087), .B2(n20699), 
        .ZN(n20700) );
  MAOI222D0BWP12T U11268 ( .A(n20695), .B(n20696), .C(n20700), .ZN(n21090) );
  MOAI22D0BWP12T U11269 ( .A1(n20695), .A2(n20696), .B1(n20695), .B2(n20696), 
        .ZN(n20701) );
  MAOI22D0BWP12T U11270 ( .A1(n20701), .A2(n20700), .B1(n20701), .B2(n20700), 
        .ZN(n20838) );
  OR3D0BWP12T U11271 ( .A1(n22009), .A2(n21933), .A3(n21184), .Z(n21197) );
  AOI22D0BWP12T U11272 ( .A1(b[8]), .A2(n21077), .B1(b[9]), .B2(n21748), .ZN(
        n20702) );
  CKND2D0BWP12T U11273 ( .A1(n21076), .A2(n21623), .ZN(n20703) );
  OAI211D0BWP12T U11274 ( .A1(n21935), .A2(n21745), .B(n20702), .C(n20703), 
        .ZN(n20704) );
  MOAI22D0BWP12T U11275 ( .A1(a[14]), .A2(n20704), .B1(a[14]), .B2(n20704), 
        .ZN(n20705) );
  CKND0BWP12T U11276 ( .I(n21156), .ZN(n20706) );
  MAOI222D0BWP12T U11277 ( .A(n21037), .B(n20705), .C(n20706), .ZN(n21149) );
  MAOI22D0BWP12T U11278 ( .A1(n20705), .A2(n21037), .B1(n20705), .B2(n21037), 
        .ZN(n20707) );
  MAOI22D0BWP12T U11279 ( .A1(n21156), .A2(n20707), .B1(n21156), .B2(n20707), 
        .ZN(n21157) );
  NR2D0BWP12T U11280 ( .A1(n21760), .A2(n23484), .ZN(n20708) );
  OAI22D0BWP12T U11281 ( .A1(n22547), .A2(n21757), .B1(n21934), .B2(n21207), 
        .ZN(n20709) );
  AOI211D0BWP12T U11282 ( .A1(n21208), .A2(n21689), .B(n20708), .C(n20709), 
        .ZN(n20710) );
  MOAI22D0BWP12T U11283 ( .A1(a[11]), .A2(n20710), .B1(a[11]), .B2(n20710), 
        .ZN(n20711) );
  CKND0BWP12T U11284 ( .I(n21284), .ZN(n20712) );
  MAOI222D0BWP12T U11285 ( .A(n21146), .B(n20711), .C(n20712), .ZN(n21280) );
  MAOI22D0BWP12T U11286 ( .A1(n21146), .A2(n20711), .B1(n21146), .B2(n20711), 
        .ZN(n20713) );
  MAOI22D0BWP12T U11287 ( .A1(n21284), .A2(n20713), .B1(n21284), .B2(n20713), 
        .ZN(n21285) );
  OAI22D0BWP12T U11288 ( .A1(b[0]), .A2(a[19]), .B1(n22009), .B2(a[20]), .ZN(
        n20714) );
  OAI22D0BWP12T U11289 ( .A1(n22485), .A2(n20714), .B1(b[1]), .B2(n22516), 
        .ZN(n22575) );
  NR2D0BWP12T U11290 ( .A1(n21725), .A2(n21549), .ZN(n20715) );
  OAI22D0BWP12T U11291 ( .A1(n21727), .A2(n22150), .B1(n21724), .B2(n21556), 
        .ZN(n20716) );
  AOI211D0BWP12T U11292 ( .A1(b[23]), .A2(n21730), .B(n20715), .C(n20716), 
        .ZN(n20717) );
  MOAI22D0BWP12T U11293 ( .A1(n21966), .A2(n20717), .B1(n21966), .B2(n20717), 
        .ZN(n20718) );
  MAOI22D0BWP12T U11294 ( .A1(n21253), .A2(n20718), .B1(n21253), .B2(n20718), 
        .ZN(n20719) );
  MAOI22D0BWP12T U11295 ( .A1(n21832), .A2(n20719), .B1(n21832), .B2(n20719), 
        .ZN(n21368) );
  CKND0BWP12T U11296 ( .I(n21832), .ZN(n20720) );
  MAOI222D0BWP12T U11297 ( .A(n21253), .B(n20720), .C(n20718), .ZN(n21835) );
  AOI22D0BWP12T U11298 ( .A1(a[17]), .A2(b[17]), .B1(a[18]), .B2(b[18]), .ZN(
        n20721) );
  ND3D0BWP12T U11299 ( .A1(n23341), .A2(n23340), .A3(n20721), .ZN(n23342) );
  IOA21D0BWP12T U11300 ( .A1(c_in), .A2(n23639), .B(n23382), .ZN(n22970) );
  IAO21D0BWP12T U11301 ( .A1(n22932), .A2(n22937), .B(n23495), .ZN(n22903) );
  IOA21D0BWP12T U11302 ( .A1(n23088), .A2(n22824), .B(n23482), .ZN(n22753) );
  IOA21D0BWP12T U11303 ( .A1(n23180), .A2(n22568), .B(n23179), .ZN(n22561) );
  IOA21D0BWP12T U11304 ( .A1(n22393), .A2(n23085), .B(n20771), .ZN(n22355) );
  NR2D0BWP12T U11305 ( .A1(n21732), .A2(n21710), .ZN(n20722) );
  OAI22D0BWP12T U11306 ( .A1(n21731), .A2(n22293), .B1(n21734), .B2(n21944), 
        .ZN(n20723) );
  AOI211D0BWP12T U11307 ( .A1(b[20]), .A2(n21737), .B(n20722), .C(n20723), 
        .ZN(n20724) );
  MOAI22D0BWP12T U11308 ( .A1(a[5]), .A2(n20724), .B1(a[5]), .B2(n20724), .ZN(
        n20725) );
  CKND0BWP12T U11309 ( .I(n21553), .ZN(n20726) );
  MAOI222D0BWP12T U11310 ( .A(n21392), .B(n20725), .C(n20726), .ZN(n21546) );
  MAOI22D0BWP12T U11311 ( .A1(n21392), .A2(n20725), .B1(n21392), .B2(n20725), 
        .ZN(n20727) );
  MAOI22D0BWP12T U11312 ( .A1(n21553), .A2(n20727), .B1(n21553), .B2(n20727), 
        .ZN(n21554) );
  IAO21D0BWP12T U11313 ( .A1(n23182), .A2(n22118), .B(n23174), .ZN(n22075) );
  IAO21D0BWP12T U11314 ( .A1(n21989), .A2(n22028), .B(n23540), .ZN(n21985) );
  IAO21D0BWP12T U11315 ( .A1(n23044), .A2(n23045), .B(n23541), .ZN(n23206) );
  IOA21D0BWP12T U11316 ( .A1(n22917), .A2(n22895), .B(n23350), .ZN(n22885) );
  IOA21D0BWP12T U11317 ( .A1(n22499), .A2(n22500), .B(n23084), .ZN(n22463) );
  NR2D0BWP12T U11318 ( .A1(n22220), .A2(n22198), .ZN(n20728) );
  MOAI22D0BWP12T U11319 ( .A1(n22168), .A2(n22081), .B1(n22174), .B2(n22721), 
        .ZN(n20729) );
  AOI211D0BWP12T U11320 ( .A1(n22200), .A2(n22447), .B(n20728), .C(n20729), 
        .ZN(n23437) );
  IOA21D0BWP12T U11321 ( .A1(n22009), .A2(a[18]), .B(n22535), .ZN(n22196) );
  NR2D0BWP12T U11322 ( .A1(n21717), .A2(n22032), .ZN(n20730) );
  MAOI22D0BWP12T U11323 ( .A1(b[26]), .A2(n22977), .B1(n21716), .B2(n23490), 
        .ZN(n20731) );
  OAI21D0BWP12T U11324 ( .A1(n21666), .A2(n21535), .B(n20731), .ZN(n20732) );
  OAI22D0BWP12T U11325 ( .A1(n21716), .A2(n21535), .B1(n21711), .B2(n23490), 
        .ZN(n20733) );
  OAI21D0BWP12T U11326 ( .A1(n20730), .A2(n20732), .B(a[2]), .ZN(n20734) );
  OAI31D0BWP12T U11327 ( .A1(n20730), .A2(a[2]), .A3(n20733), .B(n20734), .ZN(
        n20735) );
  CKND0BWP12T U11328 ( .I(n22014), .ZN(n20736) );
  MAOI222D0BWP12T U11329 ( .A(n21534), .B(n20735), .C(n20736), .ZN(n21953) );
  MAOI22D0BWP12T U11330 ( .A1(n20735), .A2(n21534), .B1(n20735), .B2(n21534), 
        .ZN(n20737) );
  MAOI22D0BWP12T U11331 ( .A1(n22014), .A2(n20737), .B1(n22014), .B2(n20737), 
        .ZN(n23324) );
  CKND2D0BWP12T U11332 ( .A1(n22403), .A2(n23299), .ZN(n20738) );
  OAI31D0BWP12T U11333 ( .A1(n22404), .A2(n22417), .A3(n22339), .B(n20738), 
        .ZN(n20739) );
  OAI31D0BWP12T U11334 ( .A1(a[20]), .A2(n22858), .A3(n22344), .B(n22426), 
        .ZN(n20740) );
  CKND0BWP12T U11335 ( .I(n22870), .ZN(n20741) );
  OAI22D0BWP12T U11336 ( .A1(n22343), .A2(n20741), .B1(n22888), .B2(n22345), 
        .ZN(n20742) );
  AOI211D0BWP12T U11337 ( .A1(n22461), .A2(n23438), .B(n20740), .C(n20742), 
        .ZN(n20743) );
  AOI22D0BWP12T U11338 ( .A1(n23498), .A2(n23509), .B1(n23652), .B2(n23355), 
        .ZN(n20744) );
  OAI211D0BWP12T U11339 ( .A1(n23499), .A2(n23355), .B(n23645), .C(n20744), 
        .ZN(n20745) );
  AOI22D0BWP12T U11340 ( .A1(n23658), .A2(n23314), .B1(n22341), .B2(n20745), 
        .ZN(n20746) );
  OAI211D0BWP12T U11341 ( .A1(n22449), .A2(n23424), .B(n20743), .C(n20746), 
        .ZN(n20747) );
  OAI22D0BWP12T U11342 ( .A1(n22948), .A2(n23147), .B1(n23211), .B2(n22350), 
        .ZN(n20748) );
  OAI22D0BWP12T U11343 ( .A1(n23669), .A2(n23201), .B1(n23653), .B2(n23636), 
        .ZN(n20749) );
  NR4D0BWP12T U11344 ( .A1(n20739), .A2(n20747), .A3(n20748), .A4(n20749), 
        .ZN(n20750) );
  OAI21D0BWP12T U11345 ( .A1(n23670), .A2(n23114), .B(n20750), .ZN(result[20])
         );
  INVD1BWP12T U11346 ( .I(b[31]), .ZN(n23043) );
  ND2D1BWP12T U11347 ( .A1(a[31]), .A2(n23043), .ZN(n23508) );
  INVD1BWP12T U11348 ( .I(n23508), .ZN(n21875) );
  INVD1BWP12T U11349 ( .I(op[2]), .ZN(n22812) );
  ND2D1BWP12T U11350 ( .A1(n22812), .A2(op[3]), .ZN(n23021) );
  INVD1BWP12T U11351 ( .I(op[1]), .ZN(n23020) );
  NR2D1BWP12T U11352 ( .A1(n23020), .A2(op[0]), .ZN(n21920) );
  IND2D1BWP12T U11353 ( .A1(n23021), .B1(n21920), .ZN(n22948) );
  INVD1BWP12T U11354 ( .I(b[30]), .ZN(n21921) );
  INVD1BWP12T U11355 ( .I(b[29]), .ZN(n23375) );
  NR2D1BWP12T U11356 ( .A1(a[29]), .A2(n23375), .ZN(n23492) );
  INVD1BWP12T U11357 ( .I(a[28]), .ZN(n21962) );
  NR2D1BWP12T U11358 ( .A1(b[28]), .A2(n21962), .ZN(n23517) );
  AOI21D1BWP12T U11359 ( .A1(b[28]), .A2(n21962), .B(n23517), .ZN(n22028) );
  INVD1BWP12T U11360 ( .I(n22028), .ZN(n23169) );
  INVD1BWP12T U11361 ( .I(b[27]), .ZN(n22032) );
  ND2D1BWP12T U11362 ( .A1(n22032), .A2(a[27]), .ZN(n23514) );
  INVD1BWP12T U11363 ( .I(a[26]), .ZN(n22087) );
  INVD1BWP12T U11364 ( .I(b[25]), .ZN(n22150) );
  INVD1BWP12T U11365 ( .I(b[23]), .ZN(n21932) );
  INVD1BWP12T U11366 ( .I(a[20]), .ZN(n22404) );
  INVD1BWP12T U11367 ( .I(b[19]), .ZN(n21944) );
  INVD1BWP12T U11368 ( .I(b[18]), .ZN(n22418) );
  NR2D1BWP12T U11369 ( .A1(a[18]), .A2(n22418), .ZN(n23506) );
  INVD1BWP12T U11370 ( .I(a[17]), .ZN(n22441) );
  NR2D1BWP12T U11371 ( .A1(b[17]), .A2(n22441), .ZN(n23520) );
  INVD1BWP12T U11372 ( .I(a[15]), .ZN(n22514) );
  NR2D1BWP12T U11373 ( .A1(b[15]), .A2(n22514), .ZN(n23521) );
  AOI21D1BWP12T U11374 ( .A1(b[15]), .A2(n22514), .B(n23521), .ZN(n22528) );
  INVD1BWP12T U11375 ( .I(n22528), .ZN(n23167) );
  INVD1BWP12T U11376 ( .I(a[14]), .ZN(n21933) );
  INVD1BWP12T U11377 ( .I(b[14]), .ZN(n22547) );
  INVD1BWP12T U11378 ( .I(b[13]), .ZN(n21934) );
  NR2D1BWP12T U11379 ( .A1(a[13]), .A2(n21934), .ZN(n23481) );
  INVD1BWP12T U11380 ( .I(a[12]), .ZN(n22689) );
  INVD1BWP12T U11381 ( .I(a[11]), .ZN(n22642) );
  AOI22D1BWP12T U11382 ( .A1(b[12]), .A2(n22689), .B1(b[11]), .B2(n22642), 
        .ZN(n23501) );
  INVD1BWP12T U11383 ( .I(b[10]), .ZN(n22675) );
  INVD1BWP12T U11384 ( .I(b[9]), .ZN(n22699) );
  INVD1BWP12T U11385 ( .I(a[8]), .ZN(n21966) );
  INVD1BWP12T U11386 ( .I(b[7]), .ZN(n21935) );
  NR2D1BWP12T U11387 ( .A1(a[7]), .A2(n21935), .ZN(n23479) );
  INVD1BWP12T U11388 ( .I(a[6]), .ZN(n23369) );
  ND2D1BWP12T U11389 ( .A1(b[6]), .A2(n23369), .ZN(n23482) );
  NR2D1BWP12T U11390 ( .A1(b[6]), .A2(n23369), .ZN(n22813) );
  INVD1BWP12T U11391 ( .I(n22813), .ZN(n23474) );
  ND2D1BWP12T U11392 ( .A1(n23482), .A2(n23474), .ZN(n22823) );
  INVD1BWP12T U11393 ( .I(n22823), .ZN(n23088) );
  INVD1BWP12T U11394 ( .I(b[5]), .ZN(n21885) );
  NR2D1BWP12T U11395 ( .A1(a[5]), .A2(n21885), .ZN(n23494) );
  INVD1BWP12T U11396 ( .I(n23494), .ZN(n20751) );
  INVD1BWP12T U11397 ( .I(a[4]), .ZN(n22873) );
  NR2D1BWP12T U11398 ( .A1(b[4]), .A2(n22873), .ZN(n23477) );
  NR2D1BWP12T U11399 ( .A1(a[4]), .A2(n23017), .ZN(n23497) );
  NR2D1BWP12T U11400 ( .A1(n23477), .A2(n23497), .ZN(n22886) );
  INVD1BWP12T U11401 ( .I(b[3]), .ZN(n22806) );
  NR2D1BWP12T U11402 ( .A1(a[3]), .A2(n22806), .ZN(n23496) );
  INVD1BWP12T U11403 ( .I(b[2]), .ZN(n22342) );
  NR2D1BWP12T U11404 ( .A1(n22342), .A2(a[2]), .ZN(n23495) );
  ND2D1BWP12T U11405 ( .A1(a[2]), .A2(n22342), .ZN(n23473) );
  IND2D1BWP12T U11406 ( .A1(n23495), .B1(n23473), .ZN(n22937) );
  INVD1BWP12T U11407 ( .I(a[1]), .ZN(n23011) );
  NR2D1BWP12T U11408 ( .A1(b[1]), .A2(n23011), .ZN(n22999) );
  INVD1BWP12T U11409 ( .I(n22999), .ZN(n23472) );
  NR2D1BWP12T U11410 ( .A1(n22009), .A2(a[0]), .ZN(n22973) );
  NR2D1BWP12T U11411 ( .A1(a[1]), .A2(n22485), .ZN(n22975) );
  NR2D1BWP12T U11412 ( .A1(n22973), .A2(n22975), .ZN(n22972) );
  INVD1BWP12T U11413 ( .I(n22972), .ZN(n23500) );
  ND2D1BWP12T U11414 ( .A1(n23472), .A2(n23500), .ZN(n22932) );
  ND2D1BWP12T U11415 ( .A1(a[3]), .A2(n22806), .ZN(n23515) );
  INR2D1BWP12T U11416 ( .A1(n23515), .B1(n23496), .ZN(n22901) );
  INVD1BWP12T U11417 ( .I(n22901), .ZN(n22917) );
  ND2D1BWP12T U11418 ( .A1(a[5]), .A2(n21885), .ZN(n22854) );
  INVD1BWP12T U11419 ( .I(n22854), .ZN(n23475) );
  AOI21D1BWP12T U11420 ( .A1(n20751), .A2(n22837), .B(n23475), .ZN(n22824) );
  ND2D1BWP12T U11421 ( .A1(a[7]), .A2(n21935), .ZN(n23471) );
  OAI21D1BWP12T U11422 ( .A1(n23479), .A2(n22753), .B(n23471), .ZN(n22738) );
  INVD1BWP12T U11423 ( .I(n22738), .ZN(n22746) );
  MAOI222D1BWP12T U11424 ( .A(n21966), .B(b[8]), .C(n22746), .ZN(n22711) );
  MAOI222D1BWP12T U11425 ( .A(n22699), .B(a[9]), .C(n22711), .ZN(n22669) );
  INVD1BWP12T U11426 ( .I(n22669), .ZN(n22667) );
  MAOI222D1BWP12T U11427 ( .A(a[10]), .B(n22675), .C(n22667), .ZN(n22630) );
  NR2D1BWP12T U11428 ( .A1(b[11]), .A2(n22642), .ZN(n20762) );
  INVD1BWP12T U11429 ( .I(n20762), .ZN(n23523) );
  ND2D1BWP12T U11430 ( .A1(n22630), .A2(n23523), .ZN(n22610) );
  NR2D1BWP12T U11431 ( .A1(b[12]), .A2(n22689), .ZN(n23525) );
  AOI21D1BWP12T U11432 ( .A1(n23501), .A2(n22610), .B(n23525), .ZN(n22583) );
  ND2D1BWP12T U11433 ( .A1(a[13]), .A2(n21934), .ZN(n23524) );
  OAI21D1BWP12T U11434 ( .A1(n23481), .A2(n22583), .B(n23524), .ZN(n22545) );
  MAOI222D1BWP12T U11435 ( .A(a[14]), .B(n22547), .C(n22545), .ZN(n22503) );
  INVD1BWP12T U11436 ( .I(a[16]), .ZN(n22515) );
  MAOI222D1BWP12T U11437 ( .A(b[16]), .B(n22498), .C(n22515), .ZN(n22464) );
  INVD1BWP12T U11438 ( .I(b[17]), .ZN(n21750) );
  OAI22D1BWP12T U11439 ( .A1(n23520), .A2(n22464), .B1(a[17]), .B2(n21750), 
        .ZN(n22424) );
  ND2D1BWP12T U11440 ( .A1(a[18]), .A2(n22418), .ZN(n22408) );
  OAI21D1BWP12T U11441 ( .A1(n23506), .A2(n22424), .B(n22408), .ZN(n22384) );
  MAOI222D1BWP12T U11442 ( .A(a[19]), .B(n21944), .C(n22384), .ZN(n22349) );
  INVD1BWP12T U11443 ( .I(b[20]), .ZN(n23498) );
  ND2D1BWP12T U11444 ( .A1(a[20]), .A2(n23498), .ZN(n23530) );
  AOI22D1BWP12T U11445 ( .A1(b[20]), .A2(n22404), .B1(n22349), .B2(n23530), 
        .ZN(n22302) );
  INVD1BWP12T U11446 ( .I(b[21]), .ZN(n22293) );
  ND2D1BWP12T U11447 ( .A1(a[21]), .A2(n22293), .ZN(n23510) );
  IND2D1BWP12T U11448 ( .A1(n22302), .B1(n23510), .ZN(n22292) );
  INVD1BWP12T U11449 ( .I(a[22]), .ZN(n20804) );
  INVD1BWP12T U11450 ( .I(a[21]), .ZN(n22406) );
  AOI22D1BWP12T U11451 ( .A1(n20804), .A2(b[22]), .B1(n22406), .B2(b[21]), 
        .ZN(n23489) );
  INVD1BWP12T U11452 ( .I(b[22]), .ZN(n21886) );
  ND2D1BWP12T U11453 ( .A1(a[22]), .A2(n21886), .ZN(n23511) );
  IOA21D1BWP12T U11454 ( .A1(n22292), .A2(n23489), .B(n23511), .ZN(n22258) );
  MAOI222D1BWP12T U11455 ( .A(a[23]), .B(n21932), .C(n22258), .ZN(n22213) );
  INVD1BWP12T U11456 ( .I(b[24]), .ZN(n21556) );
  NR2D1BWP12T U11457 ( .A1(a[24]), .A2(n21556), .ZN(n23502) );
  NR2D1BWP12T U11458 ( .A1(n22213), .A2(n23502), .ZN(n22119) );
  INVD1BWP12T U11459 ( .I(a[25]), .ZN(n22151) );
  NR2D1BWP12T U11460 ( .A1(n22151), .A2(b[25]), .ZN(n20777) );
  ND2D1BWP12T U11461 ( .A1(a[24]), .A2(n21556), .ZN(n22187) );
  IND2D1BWP12T U11462 ( .A1(n20777), .B1(n22187), .ZN(n23527) );
  OAI22D1BWP12T U11463 ( .A1(a[25]), .A2(n22150), .B1(n22119), .B2(n23527), 
        .ZN(n22074) );
  MAOI222D1BWP12T U11464 ( .A(b[26]), .B(n22087), .C(n22074), .ZN(n22065) );
  INVD1BWP12T U11465 ( .I(n22065), .ZN(n22064) );
  NR2D1BWP12T U11466 ( .A1(n22032), .A2(a[27]), .ZN(n23491) );
  AO21D1BWP12T U11467 ( .A1(n23514), .A2(n22064), .B(n23491), .Z(n21988) );
  NR2D1BWP12T U11468 ( .A1(n23492), .A2(n21951), .ZN(n21876) );
  ND2D1BWP12T U11469 ( .A1(a[30]), .A2(n21921), .ZN(n20781) );
  INVD1BWP12T U11470 ( .I(a[29]), .ZN(n23376) );
  NR2D1BWP12T U11471 ( .A1(b[29]), .A2(n23376), .ZN(n21909) );
  INVD1BWP12T U11472 ( .I(n21909), .ZN(n21958) );
  ND2D1BWP12T U11473 ( .A1(n20781), .A2(n21958), .ZN(n23533) );
  OAI22D1BWP12T U11474 ( .A1(a[30]), .A2(n21921), .B1(n21876), .B2(n23533), 
        .ZN(n23121) );
  OAI22D1BWP12T U11475 ( .A1(a[31]), .A2(n23043), .B1(n21875), .B2(n23121), 
        .ZN(n20785) );
  NR2D1BWP12T U11476 ( .A1(op[3]), .A2(n22812), .ZN(n21931) );
  ND2D1BWP12T U11477 ( .A1(n21920), .A2(n21931), .ZN(n23653) );
  AOI22D1BWP12T U11478 ( .A1(b[29]), .A2(n23376), .B1(a[29]), .B2(n23375), 
        .ZN(n21984) );
  INVD1BWP12T U11479 ( .I(b[26]), .ZN(n22088) );
  ND2D1BWP12T U11480 ( .A1(a[26]), .A2(n22088), .ZN(n23512) );
  INVD1BWP12T U11481 ( .I(n23512), .ZN(n20779) );
  ND2D1BWP12T U11482 ( .A1(b[26]), .A2(a[26]), .ZN(n23356) );
  NR2D1BWP12T U11483 ( .A1(b[26]), .A2(a[26]), .ZN(n23185) );
  INR2D1BWP12T U11484 ( .A1(n23356), .B1(n23185), .ZN(n23173) );
  INVD1BWP12T U11485 ( .I(a[23]), .ZN(n22267) );
  NR2D1BWP12T U11486 ( .A1(n22267), .A2(b[23]), .ZN(n23513) );
  NR2D1BWP12T U11487 ( .A1(b[22]), .A2(a[22]), .ZN(n23066) );
  NR2D1BWP12T U11488 ( .A1(n21886), .A2(n20804), .ZN(n23353) );
  NR2D1BWP12T U11489 ( .A1(n23066), .A2(n23353), .ZN(n23077) );
  ND2D1BWP12T U11490 ( .A1(n23498), .A2(n22404), .ZN(n22341) );
  INVD1BWP12T U11491 ( .I(n22341), .ZN(n23070) );
  NR2D1BWP12T U11492 ( .A1(n23498), .A2(n22404), .ZN(n23355) );
  NR2D1BWP12T U11493 ( .A1(n23070), .A2(n23355), .ZN(n22353) );
  INVD1BWP12T U11494 ( .I(n22353), .ZN(n22352) );
  ND2D1BWP12T U11495 ( .A1(a[19]), .A2(n21944), .ZN(n22376) );
  NR2D1BWP12T U11496 ( .A1(b[16]), .A2(n22515), .ZN(n23519) );
  NR2D1BWP12T U11497 ( .A1(b[14]), .A2(n21933), .ZN(n23518) );
  ND2D1BWP12T U11498 ( .A1(a[10]), .A2(n22675), .ZN(n23522) );
  NR2D1BWP12T U11499 ( .A1(a[9]), .A2(n22699), .ZN(n23485) );
  NR2D1BWP12T U11500 ( .A1(b[8]), .A2(n21966), .ZN(n23476) );
  NR2D1BWP12T U11501 ( .A1(n22999), .A2(n22975), .ZN(n22971) );
  ND2D1BWP12T U11502 ( .A1(a[0]), .A2(n22605), .ZN(n23516) );
  INVD1BWP12T U11503 ( .I(n23516), .ZN(n23029) );
  NR2D1BWP12T U11504 ( .A1(n22973), .A2(n23029), .ZN(n23025) );
  AOI21D1BWP12T U11505 ( .A1(n23025), .A2(c_in), .B(n23029), .ZN(n22969) );
  ND2D1BWP12T U11506 ( .A1(b[1]), .A2(a[1]), .ZN(n23347) );
  OA21D1BWP12T U11507 ( .A1(n22971), .A2(n22969), .B(n23347), .Z(n22938) );
  NR2D1BWP12T U11508 ( .A1(n20753), .A2(n23473), .ZN(n22898) );
  INVD1BWP12T U11509 ( .I(n22898), .ZN(n20752) );
  AN2D1BWP12T U11510 ( .A1(n20753), .A2(n23473), .Z(n22899) );
  AOI22D1BWP12T U11511 ( .A1(n23496), .A2(n20752), .B1(n22899), .B2(n23515), 
        .ZN(n20754) );
  OAI31D1BWP12T U11512 ( .A1(n20753), .A2(n23515), .A3(n23473), .B(n20754), 
        .ZN(n22880) );
  NR2D1BWP12T U11513 ( .A1(n22886), .A2(n22880), .ZN(n22879) );
  INR2D1BWP12T U11514 ( .A1(n20754), .B1(n22879), .ZN(n20755) );
  ND2D1BWP12T U11515 ( .A1(n23477), .A2(n20755), .ZN(n22830) );
  NR2D1BWP12T U11516 ( .A1(n22854), .A2(n22830), .ZN(n20757) );
  ND2D1BWP12T U11517 ( .A1(n22813), .A2(n20757), .ZN(n22786) );
  NR2D1BWP12T U11518 ( .A1(n23477), .A2(n20755), .ZN(n22829) );
  OAI211D1BWP12T U11519 ( .A1(n23494), .A2(n22829), .B(n22830), .C(n22854), 
        .ZN(n20756) );
  OAI21D1BWP12T U11520 ( .A1(n22854), .A2(n22830), .B(n20756), .ZN(n22798) );
  NR2D1BWP12T U11521 ( .A1(n22823), .A2(n22798), .ZN(n22797) );
  NR3D1BWP12T U11522 ( .A1(n22813), .A2(n20757), .A3(n22797), .ZN(n22785) );
  AOI22D1BWP12T U11523 ( .A1(n23479), .A2(n22786), .B1(n22785), .B2(n23471), 
        .ZN(n20758) );
  NR2D1BWP12T U11524 ( .A1(a[8]), .A2(b[8]), .ZN(n22740) );
  ND2D1BWP12T U11525 ( .A1(a[8]), .A2(b[8]), .ZN(n23344) );
  INVD1BWP12T U11526 ( .I(n23344), .ZN(n21937) );
  NR2D1BWP12T U11527 ( .A1(n22740), .A2(n21937), .ZN(n23067) );
  INVD1BWP12T U11528 ( .I(n23067), .ZN(n23122) );
  OAI21D1BWP12T U11529 ( .A1(n23471), .A2(n22786), .B(n20758), .ZN(n22720) );
  NR2D1BWP12T U11530 ( .A1(n23122), .A2(n22720), .ZN(n22719) );
  INR2D1BWP12T U11531 ( .A1(n20758), .B1(n22719), .ZN(n20759) );
  ND2D1BWP12T U11532 ( .A1(n23476), .A2(n20759), .ZN(n22684) );
  NR2D1BWP12T U11533 ( .A1(n23476), .A2(n20759), .ZN(n22683) );
  ND2D1BWP12T U11534 ( .A1(a[9]), .A2(n22699), .ZN(n23478) );
  AOI22D1BWP12T U11535 ( .A1(n23485), .A2(n22684), .B1(n22683), .B2(n23478), 
        .ZN(n20760) );
  NR2D1BWP12T U11536 ( .A1(b[10]), .A2(a[10]), .ZN(n22629) );
  AOI21D1BWP12T U11537 ( .A1(a[10]), .A2(b[10]), .B(n22629), .ZN(n23063) );
  OA21D1BWP12T U11538 ( .A1(n23478), .A2(n22684), .B(n20760), .Z(n22680) );
  ND2D1BWP12T U11539 ( .A1(n23063), .A2(n22680), .ZN(n22679) );
  ND2D1BWP12T U11540 ( .A1(n20760), .A2(n22679), .ZN(n20761) );
  NR2D1BWP12T U11541 ( .A1(n23522), .A2(n20761), .ZN(n20763) );
  NR2D1BWP12T U11542 ( .A1(b[11]), .A2(a[11]), .ZN(n22645) );
  INVD1BWP12T U11543 ( .I(b[11]), .ZN(n21887) );
  NR2D1BWP12T U11544 ( .A1(n21887), .A2(n22642), .ZN(n23343) );
  NR2D1BWP12T U11545 ( .A1(n22645), .A2(n23343), .ZN(n22655) );
  MOAI22D0BWP12T U11546 ( .A1(n23522), .A2(n20761), .B1(n23522), .B2(n20761), 
        .ZN(n22654) );
  NR2D1BWP12T U11547 ( .A1(n22655), .A2(n22654), .ZN(n22653) );
  NR3D1BWP12T U11548 ( .A1(n20762), .A2(n20763), .A3(n22653), .ZN(n20764) );
  INVD1BWP12T U11549 ( .I(b[12]), .ZN(n22612) );
  NR2D1BWP12T U11550 ( .A1(n22612), .A2(n22689), .ZN(n23351) );
  NR2D1BWP12T U11551 ( .A1(b[12]), .A2(a[12]), .ZN(n23181) );
  NR2D1BWP12T U11552 ( .A1(n23351), .A2(n23181), .ZN(n22626) );
  INVD1BWP12T U11553 ( .I(n22626), .ZN(n22611) );
  AO21D1BWP12T U11554 ( .A1(n20763), .A2(n20762), .B(n20764), .Z(n22602) );
  NR2D1BWP12T U11555 ( .A1(n22611), .A2(n22602), .ZN(n22601) );
  NR2D1BWP12T U11556 ( .A1(n20764), .A2(n22601), .ZN(n20765) );
  ND2D1BWP12T U11557 ( .A1(n23525), .A2(n20765), .ZN(n22572) );
  NR2D1BWP12T U11558 ( .A1(n23524), .A2(n22572), .ZN(n22558) );
  NR2D1BWP12T U11559 ( .A1(n23525), .A2(n20765), .ZN(n22571) );
  AOI22D1BWP12T U11560 ( .A1(n23481), .A2(n22572), .B1(n22571), .B2(n23524), 
        .ZN(n22557) );
  ND2D1BWP12T U11561 ( .A1(b[14]), .A2(n21933), .ZN(n23483) );
  AOI21D1BWP12T U11562 ( .A1(n22557), .A2(n23483), .B(n22558), .ZN(n20766) );
  MUX2ND0BWP12T U11563 ( .I0(n20766), .I1(n22558), .S(n23518), .ZN(n22527) );
  ND2D1BWP12T U11564 ( .A1(n22528), .A2(n22527), .ZN(n22526) );
  ND4D1BWP12T U11565 ( .A1(n23520), .A2(n23521), .A3(n23519), .A4(n22470), 
        .ZN(n20771) );
  INVD1BWP12T U11566 ( .I(n22376), .ZN(n23529) );
  NR2D1BWP12T U11567 ( .A1(n21944), .A2(a[19]), .ZN(n23507) );
  NR2D1BWP12T U11568 ( .A1(n23529), .A2(n23507), .ZN(n22385) );
  INVD1BWP12T U11569 ( .I(b[16]), .ZN(n21753) );
  ND2D1BWP12T U11570 ( .A1(n21753), .A2(n22515), .ZN(n23084) );
  ND2D1BWP12T U11571 ( .A1(b[16]), .A2(a[16]), .ZN(n23340) );
  ND2D1BWP12T U11572 ( .A1(n23084), .A2(n23340), .ZN(n22497) );
  ND2D1BWP12T U11573 ( .A1(n22441), .A2(n21750), .ZN(n23086) );
  OAI21D1BWP12T U11574 ( .A1(n21750), .A2(n22441), .B(n23086), .ZN(n23083) );
  MAOI222D1BWP12T U11575 ( .A(n23519), .B(n22443), .C(n23083), .ZN(n20768) );
  INVD1BWP12T U11576 ( .I(n23520), .ZN(n22442) );
  INVD1BWP12T U11577 ( .I(n20771), .ZN(n20767) );
  AOI21D1BWP12T U11578 ( .A1(n20768), .A2(n22442), .B(n20767), .ZN(n22393) );
  INVD1BWP12T U11579 ( .I(a[18]), .ZN(n22421) );
  ND2D1BWP12T U11580 ( .A1(n22418), .A2(n22421), .ZN(n21943) );
  INVD1BWP12T U11581 ( .I(n21943), .ZN(n23100) );
  AOI21D1BWP12T U11582 ( .A1(a[18]), .A2(b[18]), .B(n23100), .ZN(n22425) );
  INVD1BWP12T U11583 ( .I(n22425), .ZN(n23085) );
  NR2D1BWP12T U11584 ( .A1(n22385), .A2(n22355), .ZN(n20770) );
  ND2D1BWP12T U11585 ( .A1(n22385), .A2(n22355), .ZN(n20769) );
  OAI211D1BWP12T U11586 ( .A1(n20770), .A2(n22408), .B(n22376), .C(n20769), 
        .ZN(n20772) );
  OAI31D1BWP12T U11587 ( .A1(n22408), .A2(n22376), .A3(n20771), .B(n20772), 
        .ZN(n22351) );
  OAI21D1BWP12T U11588 ( .A1(n22352), .A2(n22351), .B(n20772), .ZN(n22313) );
  NR2D1BWP12T U11589 ( .A1(b[21]), .A2(a[21]), .ZN(n23078) );
  NR2D1BWP12T U11590 ( .A1(n22293), .A2(n22406), .ZN(n23354) );
  NR2D1BWP12T U11591 ( .A1(n23078), .A2(n23354), .ZN(n23069) );
  NR2D1BWP12T U11592 ( .A1(n22233), .A2(n23511), .ZN(n22232) );
  ND2D1BWP12T U11593 ( .A1(n23513), .A2(n22232), .ZN(n20776) );
  NR2D1BWP12T U11594 ( .A1(n22187), .A2(n20776), .ZN(n22122) );
  ND2D1BWP12T U11595 ( .A1(n20777), .A2(n22122), .ZN(n22107) );
  ND2D1BWP12T U11596 ( .A1(n22267), .A2(b[23]), .ZN(n23505) );
  ND2D1BWP12T U11597 ( .A1(n22233), .A2(n23511), .ZN(n20773) );
  OAI22D1BWP12T U11598 ( .A1(n22232), .A2(n23505), .B1(n23513), .B2(n20773), 
        .ZN(n20774) );
  AOI21D1BWP12T U11599 ( .A1(n22232), .A2(n23513), .B(n20774), .ZN(n22167) );
  NR2D1BWP12T U11600 ( .A1(b[24]), .A2(a[24]), .ZN(n21946) );
  INVD1BWP12T U11601 ( .I(n21946), .ZN(n23183) );
  ND2D1BWP12T U11602 ( .A1(b[24]), .A2(a[24]), .ZN(n23358) );
  ND2D1BWP12T U11603 ( .A1(n23183), .A2(n23358), .ZN(n23092) );
  ND2D1BWP12T U11604 ( .A1(n22167), .A2(n23092), .ZN(n20775) );
  ND3D1BWP12T U11605 ( .A1(n22187), .A2(n20776), .A3(n20775), .ZN(n22121) );
  ND2D1BWP12T U11606 ( .A1(n22151), .A2(b[25]), .ZN(n23504) );
  OAI22D1BWP12T U11607 ( .A1(n20777), .A2(n22121), .B1(n22122), .B2(n23504), 
        .ZN(n22106) );
  AOI21D1BWP12T U11608 ( .A1(n23173), .A2(n22107), .B(n22106), .ZN(n20778) );
  ND2D1BWP12T U11609 ( .A1(n20779), .A2(n20778), .ZN(n22052) );
  NR2D1BWP12T U11610 ( .A1(n20779), .A2(n20778), .ZN(n22051) );
  AOI22D1BWP12T U11611 ( .A1(n22051), .A2(n23514), .B1(n23491), .B2(n22052), 
        .ZN(n20780) );
  OAI21D1BWP12T U11612 ( .A1(n23514), .A2(n22052), .B(n20780), .ZN(n22021) );
  OAI22D1BWP12T U11613 ( .A1(n23169), .A2(n22021), .B1(n23514), .B2(n22052), 
        .ZN(n21952) );
  ND2D1BWP12T U11614 ( .A1(n21909), .A2(n21908), .ZN(n21907) );
  NR2D1BWP12T U11615 ( .A1(n20781), .A2(n21907), .ZN(n20784) );
  NR2D1BWP12T U11616 ( .A1(a[30]), .A2(n21921), .ZN(n23493) );
  NR2D1BWP12T U11617 ( .A1(n21908), .A2(n23533), .ZN(n20782) );
  AOI211D1BWP12T U11618 ( .A1(n23493), .A2(n21907), .B(n20784), .C(n20782), 
        .ZN(n23593) );
  INVD1BWP12T U11619 ( .I(a[31]), .ZN(n23642) );
  ND2D1BWP12T U11620 ( .A1(b[31]), .A2(n23642), .ZN(n21872) );
  AOI22D1BWP12T U11621 ( .A1(n23593), .A2(n21872), .B1(n20784), .B2(n23508), 
        .ZN(n20783) );
  OAI21D1BWP12T U11622 ( .A1(n20784), .A2(n23508), .B(n20783), .ZN(n20786) );
  OAI22D1BWP12T U11623 ( .A1(n22948), .A2(n20785), .B1(n23653), .B2(n20786), 
        .ZN(n23058) );
  INVD1BWP12T U11624 ( .I(n23653), .ZN(n23601) );
  INVD1BWP12T U11625 ( .I(n22948), .ZN(n23674) );
  AOI21D1BWP12T U11626 ( .A1(n23601), .A2(n20786), .B(n23674), .ZN(n21873) );
  ND2D1BWP12T U11627 ( .A1(n23020), .A2(op[0]), .ZN(n21918) );
  ND2D1BWP12T U11628 ( .A1(op[2]), .A2(op[3]), .ZN(n21899) );
  NR2D1BWP12T U11629 ( .A1(n21918), .A2(n21899), .ZN(n23658) );
  INVD1BWP12T U11630 ( .I(a[3]), .ZN(n22911) );
  NR2D1BWP12T U11631 ( .A1(n22873), .A2(n22911), .ZN(n23552) );
  INVD1BWP12T U11632 ( .I(a[2]), .ZN(n21882) );
  AOI22D1BWP12T U11633 ( .A1(a[3]), .A2(a[2]), .B1(n21882), .B2(n22911), .ZN(
        n21670) );
  NR2D1BWP12T U11634 ( .A1(a[4]), .A2(a[3]), .ZN(n21901) );
  NR3D1BWP12T U11635 ( .A1(n23552), .A2(n21670), .A3(n21901), .ZN(n21737) );
  INVD1BWP12T U11636 ( .I(b[28]), .ZN(n23490) );
  OAI22D1BWP12T U11637 ( .A1(n21803), .A2(a[4]), .B1(n22873), .B2(a[5]), .ZN(
        n20787) );
  IND2D1BWP12T U11638 ( .A1(n20787), .B1(n21670), .ZN(n21731) );
  INVD1BWP12T U11639 ( .I(a[5]), .ZN(n21803) );
  AOI33D1BWP12T U11640 ( .A1(a[2]), .A2(n23552), .A3(n21803), .B1(a[5]), .B2(
        n21901), .B3(n21882), .ZN(n21734) );
  AN2D1BWP12T U11641 ( .A1(n21670), .A2(n20787), .Z(n21502) );
  INVD1BWP12T U11642 ( .I(n21502), .ZN(n21732) );
  NR2D1BWP12T U11643 ( .A1(n22342), .A2(n22485), .ZN(n22951) );
  INVD1BWP12T U11644 ( .I(n22951), .ZN(n22244) );
  INVD1BWP12T U11645 ( .I(b[4]), .ZN(n23017) );
  AOI21D1BWP12T U11646 ( .A1(n22806), .A2(n22244), .B(n23017), .ZN(n22673) );
  INVD1BWP12T U11647 ( .I(b[6]), .ZN(n23370) );
  NR2D1BWP12T U11648 ( .A1(n22605), .A2(n22485), .ZN(n22842) );
  INVD1BWP12T U11649 ( .I(n22842), .ZN(n22993) );
  ND2D1BWP12T U11650 ( .A1(n22342), .A2(n22993), .ZN(n20831) );
  AOI21D1BWP12T U11651 ( .A1(b[3]), .A2(n20831), .B(b[4]), .ZN(n20840) );
  OAI33D1BWP12T U11652 ( .A1(b[5]), .A2(n22673), .A3(n23370), .B1(n21885), 
        .B2(n20840), .B3(b[6]), .ZN(n20839) );
  OAI21D1BWP12T U11653 ( .A1(b[5]), .A2(n22673), .B(b[6]), .ZN(n20788) );
  IOA21D1BWP12T U11654 ( .A1(b[7]), .A2(n20839), .B(n20788), .ZN(n20807) );
  NR2D1BWP12T U11655 ( .A1(b[9]), .A2(n20789), .ZN(n20865) );
  NR2D1BWP12T U11656 ( .A1(n20865), .A2(n22675), .ZN(n20798) );
  IND2D1BWP12T U11657 ( .A1(n20798), .B1(n21887), .ZN(n20930) );
  ND2D1BWP12T U11658 ( .A1(n20930), .A2(b[12]), .ZN(n20921) );
  ND2D1BWP12T U11659 ( .A1(n21934), .A2(n20921), .ZN(n21004) );
  INVD1BWP12T U11660 ( .I(n21004), .ZN(n21003) );
  INVD1BWP12T U11661 ( .I(b[15]), .ZN(n23484) );
  OAI21D1BWP12T U11662 ( .A1(n21003), .A2(n22547), .B(n23484), .ZN(n21000) );
  ND2D1BWP12T U11663 ( .A1(b[16]), .A2(n21000), .ZN(n20992) );
  ND2D1BWP12T U11664 ( .A1(n21750), .A2(n20992), .ZN(n21107) );
  ND2D1BWP12T U11665 ( .A1(b[18]), .A2(n21107), .ZN(n21126) );
  ND2D1BWP12T U11666 ( .A1(n21944), .A2(n21126), .ZN(n21119) );
  ND2D1BWP12T U11667 ( .A1(b[20]), .A2(n21119), .ZN(n21116) );
  ND2D1BWP12T U11668 ( .A1(n22293), .A2(n21116), .ZN(n21214) );
  ND2D1BWP12T U11669 ( .A1(b[22]), .A2(n21214), .ZN(n21260) );
  ND2D1BWP12T U11670 ( .A1(n21932), .A2(n21260), .ZN(n21255) );
  ND2D1BWP12T U11671 ( .A1(b[24]), .A2(n21255), .ZN(n20794) );
  ND2D1BWP12T U11672 ( .A1(n22150), .A2(n20794), .ZN(n21375) );
  ND2D1BWP12T U11673 ( .A1(b[26]), .A2(n21375), .ZN(n21370) );
  ND2D1BWP12T U11674 ( .A1(n22032), .A2(n21370), .ZN(n21508) );
  ND2D1BWP12T U11675 ( .A1(b[9]), .A2(n20789), .ZN(n20864) );
  ND2D1BWP12T U11676 ( .A1(n22675), .A2(n20864), .ZN(n20799) );
  ND2D1BWP12T U11677 ( .A1(b[11]), .A2(n20799), .ZN(n20929) );
  ND2D1BWP12T U11678 ( .A1(n22612), .A2(n20929), .ZN(n20920) );
  ND2D1BWP12T U11679 ( .A1(b[13]), .A2(n20920), .ZN(n20912) );
  ND2D1BWP12T U11680 ( .A1(n22547), .A2(n20912), .ZN(n21005) );
  ND2D1BWP12T U11681 ( .A1(b[15]), .A2(n21005), .ZN(n21002) );
  ND2D1BWP12T U11682 ( .A1(n21753), .A2(n21002), .ZN(n20991) );
  ND2D1BWP12T U11683 ( .A1(b[17]), .A2(n20991), .ZN(n21106) );
  ND2D1BWP12T U11684 ( .A1(n22418), .A2(n21106), .ZN(n21125) );
  ND2D1BWP12T U11685 ( .A1(b[19]), .A2(n21125), .ZN(n21118) );
  ND2D1BWP12T U11686 ( .A1(n23498), .A2(n21118), .ZN(n21115) );
  ND2D1BWP12T U11687 ( .A1(b[21]), .A2(n21115), .ZN(n21213) );
  ND2D1BWP12T U11688 ( .A1(n21886), .A2(n21213), .ZN(n21259) );
  ND2D1BWP12T U11689 ( .A1(b[23]), .A2(n21259), .ZN(n21254) );
  ND2D1BWP12T U11690 ( .A1(n21556), .A2(n21254), .ZN(n20793) );
  ND2D1BWP12T U11691 ( .A1(b[25]), .A2(n20793), .ZN(n21374) );
  ND2D1BWP12T U11692 ( .A1(n22088), .A2(n21374), .ZN(n21369) );
  ND2D1BWP12T U11693 ( .A1(b[27]), .A2(n21369), .ZN(n21507) );
  ND2D1BWP12T U11694 ( .A1(n21508), .A2(n21507), .ZN(n20790) );
  MAOI22D0BWP12T U11695 ( .A1(b[28]), .A2(n20790), .B1(b[28]), .B2(n20790), 
        .ZN(n21535) );
  INVD1BWP12T U11696 ( .I(a[7]), .ZN(n22776) );
  NR2D1BWP12T U11697 ( .A1(a[6]), .A2(a[5]), .ZN(n22775) );
  NR2D1BWP12T U11698 ( .A1(n23369), .A2(n21803), .ZN(n20791) );
  AO33D1BWP12T U11699 ( .A1(n22776), .A2(n22775), .A3(a[8]), .B1(a[7]), .B2(
        n20791), .B3(n21966), .Z(n21730) );
  INR2D1BWP12T U11700 ( .A1(n22775), .B1(n22776), .ZN(n22768) );
  ND2D1BWP12T U11701 ( .A1(a[7]), .A2(a[6]), .ZN(n23557) );
  OAI21D1BWP12T U11702 ( .A1(n20791), .A2(n22768), .B(n23557), .ZN(n21724) );
  OAI22D1BWP12T U11703 ( .A1(n21966), .A2(a[7]), .B1(n22776), .B2(a[8]), .ZN(
        n20792) );
  NR2D1BWP12T U11704 ( .A1(n22775), .A2(n20791), .ZN(n21342) );
  IND2D1BWP12T U11705 ( .A1(n20792), .B1(n21342), .ZN(n21727) );
  ND2D1BWP12T U11706 ( .A1(n21342), .A2(n20792), .ZN(n21725) );
  ND2D1BWP12T U11707 ( .A1(n20794), .A2(n20793), .ZN(n20795) );
  MAOI22D0BWP12T U11708 ( .A1(b[25]), .A2(n20795), .B1(b[25]), .B2(n20795), 
        .ZN(n21549) );
  AOI22D1BWP12T U11709 ( .A1(a[18]), .A2(a[17]), .B1(n22441), .B2(n22421), 
        .ZN(n20903) );
  INVD1BWP12T U11710 ( .I(a[19]), .ZN(n22383) );
  AOI22D1BWP12T U11711 ( .A1(a[20]), .A2(n22383), .B1(a[19]), .B2(n22404), 
        .ZN(n20797) );
  ND2D1BWP12T U11712 ( .A1(n20903), .A2(n20797), .ZN(n21764) );
  ND2D1BWP12T U11713 ( .A1(n22383), .A2(n22421), .ZN(n22339) );
  ND2D1BWP12T U11714 ( .A1(a[19]), .A2(a[18]), .ZN(n23551) );
  INVD1BWP12T U11715 ( .I(n20903), .ZN(n20796) );
  ND3D1BWP12T U11716 ( .A1(n22339), .A2(n23551), .A3(n20796), .ZN(n21767) );
  INVD1BWP12T U11717 ( .I(n21767), .ZN(n20904) );
  AOI211D1BWP12T U11718 ( .A1(n22339), .A2(n23551), .B(n20903), .C(n20797), 
        .ZN(n21770) );
  AOI22D1BWP12T U11719 ( .A1(b[10]), .A2(n20904), .B1(b[9]), .B2(n21770), .ZN(
        n20802) );
  NR2D1BWP12T U11720 ( .A1(n20797), .A2(n20796), .ZN(n20905) );
  INR2D1BWP12T U11721 ( .A1(n20799), .B1(n20798), .ZN(n20800) );
  MAOI22D0BWP12T U11722 ( .A1(b[11]), .A2(n20800), .B1(b[11]), .B2(n20800), 
        .ZN(n21773) );
  ND2D1BWP12T U11723 ( .A1(n20905), .A2(n21773), .ZN(n20801) );
  OAI211D1BWP12T U11724 ( .A1(n21764), .A2(n21887), .B(n20802), .C(n20801), 
        .ZN(n20803) );
  MAOI22D0BWP12T U11725 ( .A1(n22404), .A2(n20803), .B1(n22404), .B2(n20803), 
        .ZN(n21104) );
  AOI22D1BWP12T U11726 ( .A1(a[23]), .A2(n20804), .B1(a[22]), .B2(n22267), 
        .ZN(n20806) );
  AOI22D1BWP12T U11727 ( .A1(a[21]), .A2(n22404), .B1(a[20]), .B2(n22406), 
        .ZN(n20805) );
  ND2D1BWP12T U11728 ( .A1(n20804), .A2(n22406), .ZN(n23046) );
  ND2D1BWP12T U11729 ( .A1(a[22]), .A2(a[21]), .ZN(n23555) );
  ND3D1BWP12T U11730 ( .A1(n23046), .A2(n23555), .A3(n20805), .ZN(n21777) );
  INVD1BWP12T U11731 ( .I(n21777), .ZN(n22291) );
  INVD1BWP12T U11732 ( .I(n20805), .ZN(n20853) );
  AOI211D1BWP12T U11733 ( .A1(n23046), .A2(n23555), .B(n20853), .C(n20806), 
        .ZN(n21772) );
  NR2D1BWP12T U11734 ( .A1(n20806), .A2(n20805), .ZN(n21774) );
  FA1D0BWP12T U11735 ( .A(b[7]), .B(b[8]), .CI(n20807), .CO(n20871), .S(n21781) );
  INVD1BWP12T U11736 ( .I(a[27]), .ZN(n22190) );
  AOI22D1BWP12T U11737 ( .A1(a[27]), .A2(a[26]), .B1(n22087), .B2(n22190), 
        .ZN(n20810) );
  ND2D1BWP12T U11738 ( .A1(b[0]), .A2(n20810), .ZN(n20845) );
  NR2D1BWP12T U11739 ( .A1(n23376), .A2(n20845), .ZN(n20825) );
  INVD1BWP12T U11740 ( .I(n20810), .ZN(n20808) );
  AOI22D1BWP12T U11741 ( .A1(a[29]), .A2(n21962), .B1(a[28]), .B2(n23376), 
        .ZN(n20809) );
  NR2D1BWP12T U11742 ( .A1(n20808), .A2(n20809), .ZN(n20811) );
  INVD1BWP12T U11743 ( .I(n20811), .ZN(n21798) );
  NR2D1BWP12T U11744 ( .A1(b[0]), .A2(b[1]), .ZN(n22757) );
  NR2D1BWP12T U11745 ( .A1(n22842), .A2(n22757), .ZN(n22864) );
  INVD1BWP12T U11746 ( .I(n22864), .ZN(n22867) );
  ND2D1BWP12T U11747 ( .A1(n21962), .A2(n22190), .ZN(n21895) );
  ND2D1BWP12T U11748 ( .A1(a[28]), .A2(a[27]), .ZN(n23554) );
  ND3D1BWP12T U11749 ( .A1(n21895), .A2(n23554), .A3(n20808), .ZN(n21799) );
  INVD1BWP12T U11750 ( .I(b[0]), .ZN(n22009) );
  INVD1BWP12T U11751 ( .I(b[1]), .ZN(n22485) );
  ND2D1BWP12T U11752 ( .A1(n20810), .A2(n20809), .ZN(n21796) );
  OAI222D1BWP12T U11753 ( .A1(n21798), .A2(n22867), .B1(n21799), .B2(n22009), 
        .C1(n22485), .C2(n21796), .ZN(n20824) );
  NR2D1BWP12T U11754 ( .A1(n20825), .A2(n20824), .ZN(n20823) );
  NR2D1BWP12T U11755 ( .A1(n20823), .A2(n23376), .ZN(n20815) );
  AOI211D1BWP12T U11756 ( .A1(n21895), .A2(n23554), .B(n20810), .C(n20809), 
        .ZN(n21802) );
  MAOI22D0BWP12T U11757 ( .A1(b[0]), .A2(n21802), .B1(n22485), .B2(n21799), 
        .ZN(n20813) );
  ND2D1BWP12T U11758 ( .A1(b[1]), .A2(n22342), .ZN(n22245) );
  NR2D1BWP12T U11759 ( .A1(n22485), .A2(b[0]), .ZN(n22843) );
  OAI22D1BWP12T U11760 ( .A1(b[0]), .A2(n22245), .B1(n22843), .B2(n22342), 
        .ZN(n21655) );
  ND2D1BWP12T U11761 ( .A1(n20811), .A2(n21655), .ZN(n20812) );
  OAI211D1BWP12T U11762 ( .A1(n21796), .A2(n22342), .B(n20813), .C(n20812), 
        .ZN(n20814) );
  NR2D1BWP12T U11763 ( .A1(n20815), .A2(n20814), .ZN(n21098) );
  AOI21D1BWP12T U11764 ( .A1(n20815), .A2(n20814), .B(n21098), .ZN(n21092) );
  ND2D1BWP12T U11765 ( .A1(n22087), .A2(n22151), .ZN(n21896) );
  ND2D1BWP12T U11766 ( .A1(a[26]), .A2(a[25]), .ZN(n23553) );
  INVD1BWP12T U11767 ( .I(a[24]), .ZN(n23560) );
  ND2D1BWP12T U11768 ( .A1(n23560), .A2(n22267), .ZN(n23047) );
  OAI21D1BWP12T U11769 ( .A1(n22267), .A2(n23560), .B(n23047), .ZN(n20858) );
  AOI21D1BWP12T U11770 ( .A1(n21896), .A2(n23553), .B(n20858), .ZN(n21779) );
  INVD1BWP12T U11771 ( .I(n21779), .ZN(n20828) );
  ND2D1BWP12T U11772 ( .A1(n21896), .A2(n23553), .ZN(n20816) );
  NR2D1BWP12T U11773 ( .A1(n20816), .A2(n20858), .ZN(n21780) );
  INVD1BWP12T U11774 ( .I(n21780), .ZN(n20827) );
  NR2D1BWP12T U11775 ( .A1(n22673), .A2(n20840), .ZN(n20817) );
  MAOI22D0BWP12T U11776 ( .A1(n20817), .A2(n21885), .B1(n20817), .B2(n21885), 
        .ZN(n21797) );
  OAI22D1BWP12T U11777 ( .A1(n21885), .A2(n20828), .B1(n20827), .B2(n21797), 
        .ZN(n20820) );
  OAI33D1BWP12T U11778 ( .A1(a[25]), .A2(n23560), .A3(n22267), .B1(n22151), 
        .B2(a[24]), .B3(a[23]), .ZN(n21778) );
  INVD1BWP12T U11779 ( .I(n21778), .ZN(n20826) );
  OAI33D1BWP12T U11780 ( .A1(a[24]), .A2(a[23]), .A3(n22087), .B1(n23560), 
        .B2(n22151), .B3(n22267), .ZN(n20818) );
  ND2D1BWP12T U11781 ( .A1(n20818), .A2(n23553), .ZN(n21784) );
  OAI22D1BWP12T U11782 ( .A1(n23017), .A2(n20826), .B1(n22806), .B2(n21784), 
        .ZN(n20819) );
  NR2D1BWP12T U11783 ( .A1(n20820), .A2(n20819), .ZN(n20821) );
  MAOI22D0BWP12T U11784 ( .A1(n20821), .A2(n22087), .B1(n20821), .B2(n22087), 
        .ZN(n21091) );
  AOI22D1BWP12T U11785 ( .A1(b[3]), .A2(n20831), .B1(n22244), .B2(n22806), 
        .ZN(n20822) );
  MAOI22D0BWP12T U11786 ( .A1(n20822), .A2(n23017), .B1(n20822), .B2(n23017), 
        .ZN(n21667) );
  OAI32D1BWP12T U11787 ( .A1(n22009), .A2(n22087), .A3(n20858), .B1(n20826), 
        .B2(n22009), .ZN(n20863) );
  OAI22D1BWP12T U11788 ( .A1(n22485), .A2(n20828), .B1(n22867), .B2(n20827), 
        .ZN(n20862) );
  NR2D1BWP12T U11789 ( .A1(n20863), .A2(n20862), .ZN(n20861) );
  NR2D1BWP12T U11790 ( .A1(n20861), .A2(n22087), .ZN(n20849) );
  AOI22D1BWP12T U11791 ( .A1(b[2]), .A2(n21779), .B1(n21780), .B2(n21655), 
        .ZN(n20830) );
  ND2D1BWP12T U11792 ( .A1(b[1]), .A2(n21778), .ZN(n20829) );
  OAI211D1BWP12T U11793 ( .A1(n21784), .A2(n22605), .B(n20830), .C(n20829), 
        .ZN(n20848) );
  NR2D1BWP12T U11794 ( .A1(n20849), .A2(n20848), .ZN(n20847) );
  NR2D1BWP12T U11795 ( .A1(n20847), .A2(n22087), .ZN(n20836) );
  ND2D1BWP12T U11796 ( .A1(n22244), .A2(n20831), .ZN(n20832) );
  MAOI22D0BWP12T U11797 ( .A1(b[3]), .A2(n20832), .B1(b[3]), .B2(n20832), .ZN(
        n21659) );
  INVD1BWP12T U11798 ( .I(n21659), .ZN(n21348) );
  AOI22D1BWP12T U11799 ( .A1(b[3]), .A2(n21779), .B1(n21348), .B2(n21780), 
        .ZN(n20834) );
  ND2D1BWP12T U11800 ( .A1(b[2]), .A2(n21778), .ZN(n20833) );
  OAI211D1BWP12T U11801 ( .A1(n21784), .A2(n22485), .B(n20834), .C(n20833), 
        .ZN(n20835) );
  MAOI22D0BWP12T U11802 ( .A1(n20836), .A2(n20835), .B1(n20836), .B2(n20835), 
        .ZN(n20846) );
  INVD1BWP12T U11803 ( .I(n21771), .ZN(n21238) );
  INVD1BWP12T U11804 ( .I(n21774), .ZN(n21237) );
  MAOI22D0BWP12T U11805 ( .A1(n20839), .A2(n21935), .B1(n20839), .B2(n21935), 
        .ZN(n21636) );
  NR2D1BWP12T U11806 ( .A1(n23370), .A2(n21238), .ZN(n20843) );
  AOI22D1BWP12T U11807 ( .A1(b[5]), .A2(n20840), .B1(n22673), .B2(n21885), 
        .ZN(n20841) );
  MAOI22D0BWP12T U11808 ( .A1(b[6]), .A2(n20841), .B1(b[6]), .B2(n20841), .ZN(
        n21671) );
  OAI22D1BWP12T U11809 ( .A1(n21885), .A2(n21777), .B1(n21237), .B2(n21671), 
        .ZN(n20842) );
  AOI211D1BWP12T U11810 ( .A1(n21772), .A2(b[4]), .B(n20843), .C(n20842), .ZN(
        n20844) );
  MAOI22D0BWP12T U11811 ( .A1(a[23]), .A2(n20844), .B1(a[23]), .B2(n20844), 
        .ZN(n20877) );
  MAOI22D0BWP12T U11812 ( .A1(n20846), .A2(n20845), .B1(n20846), .B2(n20845), 
        .ZN(n20876) );
  AO21D1BWP12T U11813 ( .A1(n20849), .A2(n20848), .B(n20847), .Z(n20880) );
  NR2D1BWP12T U11814 ( .A1(n21885), .A2(n21238), .ZN(n20851) );
  OAI22D1BWP12T U11815 ( .A1(n23017), .A2(n21777), .B1(n21237), .B2(n21797), 
        .ZN(n20850) );
  AOI211D1BWP12T U11816 ( .A1(n21772), .A2(b[3]), .B(n20851), .C(n20850), .ZN(
        n20852) );
  MAOI22D0BWP12T U11817 ( .A1(a[23]), .A2(n20852), .B1(a[23]), .B2(n20852), 
        .ZN(n20879) );
  ND2D1BWP12T U11818 ( .A1(b[0]), .A2(n20853), .ZN(n20962) );
  NR2D1BWP12T U11819 ( .A1(n22267), .A2(n20962), .ZN(n20900) );
  OAI222D1BWP12T U11820 ( .A1(n21237), .A2(n22867), .B1(n21777), .B2(n22009), 
        .C1(n22485), .C2(n21238), .ZN(n20899) );
  NR2D1BWP12T U11821 ( .A1(n20900), .A2(n20899), .ZN(n20898) );
  NR2D1BWP12T U11822 ( .A1(n20898), .A2(n22267), .ZN(n20894) );
  AOI22D1BWP12T U11823 ( .A1(b[0]), .A2(n21772), .B1(b[2]), .B2(n21771), .ZN(
        n20855) );
  AOI22D1BWP12T U11824 ( .A1(b[1]), .A2(n22291), .B1(n21774), .B2(n21655), 
        .ZN(n20854) );
  ND2D1BWP12T U11825 ( .A1(n20855), .A2(n20854), .ZN(n20893) );
  NR2D1BWP12T U11826 ( .A1(n20894), .A2(n20893), .ZN(n20892) );
  NR2D1BWP12T U11827 ( .A1(n20892), .A2(n22267), .ZN(n20860) );
  AOI22D1BWP12T U11828 ( .A1(b[3]), .A2(n21771), .B1(b[2]), .B2(n22291), .ZN(
        n20857) );
  ND2D1BWP12T U11829 ( .A1(b[1]), .A2(n21772), .ZN(n20856) );
  OAI211D1BWP12T U11830 ( .A1(n21237), .A2(n21659), .B(n20857), .C(n20856), 
        .ZN(n20859) );
  MOAI22D0BWP12T U11831 ( .A1(n20860), .A2(n20859), .B1(n20860), .B2(n20859), 
        .ZN(n20890) );
  NR2D1BWP12T U11832 ( .A1(n22605), .A2(n20858), .ZN(n20891) );
  INVD1BWP12T U11833 ( .I(n20905), .ZN(n21766) );
  IND2D1BWP12T U11834 ( .A1(n20865), .B1(n20864), .ZN(n20866) );
  MAOI22D0BWP12T U11835 ( .A1(b[10]), .A2(n20866), .B1(b[10]), .B2(n20866), 
        .ZN(n21678) );
  NR2D1BWP12T U11836 ( .A1(n21766), .A2(n21678), .ZN(n20868) );
  OAI22D1BWP12T U11837 ( .A1(n22675), .A2(n21764), .B1(n22699), .B2(n21767), 
        .ZN(n20867) );
  AOI211D1BWP12T U11838 ( .A1(n21770), .A2(b[8]), .B(n20868), .C(n20867), .ZN(
        n20869) );
  MAOI22D0BWP12T U11839 ( .A1(a[20]), .A2(n20869), .B1(a[20]), .B2(n20869), 
        .ZN(n20919) );
  AOI22D1BWP12T U11840 ( .A1(b[8]), .A2(n20904), .B1(b[7]), .B2(n21770), .ZN(
        n20873) );
  FA1D0BWP12T U11841 ( .A(b[8]), .B(b[9]), .CI(n20871), .CO(n20789), .S(n21623) );
  ND2D1BWP12T U11842 ( .A1(n20905), .A2(n21623), .ZN(n20872) );
  OAI211D1BWP12T U11843 ( .A1(n21764), .A2(n22699), .B(n20873), .C(n20872), 
        .ZN(n20874) );
  MAOI22D0BWP12T U11844 ( .A1(n22404), .A2(n20874), .B1(n22404), .B2(n20874), 
        .ZN(n20928) );
  FA1D0BWP12T U11845 ( .A(n20877), .B(n20876), .CI(n20875), .CO(n20870), .S(
        n20927) );
  FA1D0BWP12T U11846 ( .A(n20880), .B(n20879), .CI(n20878), .CO(n20875), .S(
        n20937) );
  INVD1BWP12T U11847 ( .I(b[8]), .ZN(n22741) );
  AOI22D1BWP12T U11848 ( .A1(b[7]), .A2(n20904), .B1(b[6]), .B2(n21770), .ZN(
        n20882) );
  ND2D1BWP12T U11849 ( .A1(n20905), .A2(n21781), .ZN(n20881) );
  OAI211D1BWP12T U11850 ( .A1(n21764), .A2(n22741), .B(n20882), .C(n20881), 
        .ZN(n20883) );
  MAOI22D0BWP12T U11851 ( .A1(n22404), .A2(n20883), .B1(n22404), .B2(n20883), 
        .ZN(n20936) );
  NR2D1BWP12T U11852 ( .A1(n21935), .A2(n21764), .ZN(n20885) );
  OAI22D1BWP12T U11853 ( .A1(n23370), .A2(n21767), .B1(n21766), .B2(n21636), 
        .ZN(n20884) );
  AOI211D1BWP12T U11854 ( .A1(n21770), .A2(b[5]), .B(n20885), .C(n20884), .ZN(
        n20886) );
  MAOI22D0BWP12T U11855 ( .A1(a[20]), .A2(n20886), .B1(a[20]), .B2(n20886), 
        .ZN(n20946) );
  NR2D1BWP12T U11856 ( .A1(n23370), .A2(n21764), .ZN(n20888) );
  OAI22D1BWP12T U11857 ( .A1(n21885), .A2(n21767), .B1(n21766), .B2(n21671), 
        .ZN(n20887) );
  AOI211D1BWP12T U11858 ( .A1(n21770), .A2(b[4]), .B(n20888), .C(n20887), .ZN(
        n20889) );
  MAOI22D0BWP12T U11859 ( .A1(a[20]), .A2(n20889), .B1(a[20]), .B2(n20889), 
        .ZN(n20952) );
  MAOI22D0BWP12T U11860 ( .A1(n20891), .A2(n20890), .B1(n20891), .B2(n20890), 
        .ZN(n20951) );
  AO21D1BWP12T U11861 ( .A1(n20894), .A2(n20893), .B(n20892), .Z(n20955) );
  NR2D1BWP12T U11862 ( .A1(n21885), .A2(n21764), .ZN(n20896) );
  OAI22D1BWP12T U11863 ( .A1(n23017), .A2(n21767), .B1(n21766), .B2(n21797), 
        .ZN(n20895) );
  AOI211D1BWP12T U11864 ( .A1(n21770), .A2(b[3]), .B(n20896), .C(n20895), .ZN(
        n20897) );
  MAOI22D0BWP12T U11865 ( .A1(a[20]), .A2(n20897), .B1(a[20]), .B2(n20897), 
        .ZN(n20954) );
  NR2D1BWP12T U11866 ( .A1(n22806), .A2(n21764), .ZN(n20902) );
  OAI22D1BWP12T U11867 ( .A1(n22342), .A2(n21767), .B1(n21659), .B2(n21766), 
        .ZN(n20901) );
  AOI211D1BWP12T U11868 ( .A1(n21770), .A2(b[1]), .B(n20902), .C(n20901), .ZN(
        n20909) );
  ND2D1BWP12T U11869 ( .A1(b[0]), .A2(n20903), .ZN(n21051) );
  NR2D1BWP12T U11870 ( .A1(n22404), .A2(n21051), .ZN(n20975) );
  OAI22D1BWP12T U11871 ( .A1(n22485), .A2(n21764), .B1(n22867), .B2(n21766), 
        .ZN(n20974) );
  AOI211D1BWP12T U11872 ( .A1(n20904), .A2(b[0]), .B(n20975), .C(n20974), .ZN(
        n20973) );
  NR2D1BWP12T U11873 ( .A1(n20973), .A2(n22404), .ZN(n20969) );
  AOI22D1BWP12T U11874 ( .A1(b[0]), .A2(n21770), .B1(b[1]), .B2(n20904), .ZN(
        n20907) );
  ND2D1BWP12T U11875 ( .A1(n20905), .A2(n21655), .ZN(n20906) );
  OAI211D1BWP12T U11876 ( .A1(n21764), .A2(n22342), .B(n20907), .C(n20906), 
        .ZN(n20968) );
  NR2D1BWP12T U11877 ( .A1(n20969), .A2(n20968), .ZN(n20967) );
  NR2D1BWP12T U11878 ( .A1(n20967), .A2(n22404), .ZN(n20908) );
  MOAI22D0BWP12T U11879 ( .A1(n20909), .A2(n20908), .B1(n20909), .B2(n20908), 
        .ZN(n20963) );
  ND2D1BWP12T U11880 ( .A1(n22515), .A2(n22514), .ZN(n21897) );
  ND2D1BWP12T U11881 ( .A1(a[16]), .A2(a[15]), .ZN(n23550) );
  AOI22D1BWP12T U11882 ( .A1(a[15]), .A2(a[14]), .B1(n21933), .B2(n22514), 
        .ZN(n20911) );
  ND2D1BWP12T U11883 ( .A1(a[17]), .A2(a[14]), .ZN(n23549) );
  OAI21D1BWP12T U11884 ( .A1(a[17]), .A2(a[14]), .B(n23549), .ZN(n21813) );
  AOI211D1BWP12T U11885 ( .A1(n21897), .A2(n23550), .B(n20911), .C(n21813), 
        .ZN(n21756) );
  INVD1BWP12T U11886 ( .I(n20911), .ZN(n21070) );
  OAI22D1BWP12T U11887 ( .A1(n22441), .A2(a[16]), .B1(n22515), .B2(a[17]), 
        .ZN(n20910) );
  NR2D1BWP12T U11888 ( .A1(n21070), .A2(n20910), .ZN(n20981) );
  INVD1BWP12T U11889 ( .I(n20981), .ZN(n21749) );
  NR2D1BWP12T U11890 ( .A1(n22547), .A2(n21749), .ZN(n20915) );
  ND3D1BWP12T U11891 ( .A1(n21897), .A2(n23550), .A3(n21070), .ZN(n22477) );
  ND2D1BWP12T U11892 ( .A1(n20911), .A2(n20910), .ZN(n21752) );
  INR2D1BWP12T U11893 ( .A1(n20912), .B1(n21003), .ZN(n20913) );
  MAOI22D0BWP12T U11894 ( .A1(n20913), .A2(n22547), .B1(n20913), .B2(n22547), 
        .ZN(n21765) );
  OAI22D1BWP12T U11895 ( .A1(n21934), .A2(n22477), .B1(n21752), .B2(n21765), 
        .ZN(n20914) );
  AOI211D1BWP12T U11896 ( .A1(n21756), .A2(b[12]), .B(n20915), .C(n20914), 
        .ZN(n20916) );
  MAOI22D0BWP12T U11897 ( .A1(a[17]), .A2(n20916), .B1(a[17]), .B2(n20916), 
        .ZN(n21082) );
  FA1D0BWP12T U11898 ( .A(n20919), .B(n20918), .CI(n20917), .CO(n21102), .S(
        n20998) );
  NR2D1BWP12T U11899 ( .A1(n21934), .A2(n21749), .ZN(n20924) );
  ND2D1BWP12T U11900 ( .A1(n20921), .A2(n20920), .ZN(n20922) );
  MAOI22D0BWP12T U11901 ( .A1(b[13]), .A2(n20922), .B1(b[13]), .B2(n20922), 
        .ZN(n21595) );
  OAI22D1BWP12T U11902 ( .A1(n22612), .A2(n22477), .B1(n21752), .B2(n21595), 
        .ZN(n20923) );
  AOI211D1BWP12T U11903 ( .A1(n21756), .A2(b[11]), .B(n20924), .C(n20923), 
        .ZN(n20925) );
  MAOI22D0BWP12T U11904 ( .A1(a[17]), .A2(n20925), .B1(a[17]), .B2(n20925), 
        .ZN(n20997) );
  FA1D0BWP12T U11905 ( .A(n20928), .B(n20927), .CI(n20926), .CO(n20917), .S(
        n21009) );
  NR2D1BWP12T U11906 ( .A1(n21887), .A2(n22477), .ZN(n20933) );
  ND2D1BWP12T U11907 ( .A1(n20930), .A2(n20929), .ZN(n20931) );
  MAOI22D0BWP12T U11908 ( .A1(b[12]), .A2(n20931), .B1(b[12]), .B2(n20931), 
        .ZN(n21683) );
  OAI22D1BWP12T U11909 ( .A1(n22612), .A2(n21749), .B1(n21752), .B2(n21683), 
        .ZN(n20932) );
  AOI211D1BWP12T U11910 ( .A1(n21756), .A2(b[10]), .B(n20933), .C(n20932), 
        .ZN(n20934) );
  MAOI22D0BWP12T U11911 ( .A1(a[17]), .A2(n20934), .B1(a[17]), .B2(n20934), 
        .ZN(n21008) );
  FA1D0BWP12T U11912 ( .A(n20937), .B(n20936), .CI(n20935), .CO(n20926), .S(
        n21013) );
  INVD1BWP12T U11913 ( .I(n22477), .ZN(n21241) );
  AOI22D1BWP12T U11914 ( .A1(b[10]), .A2(n21241), .B1(b[11]), .B2(n20981), 
        .ZN(n20939) );
  INVD1BWP12T U11915 ( .I(n21752), .ZN(n21240) );
  AOI22D1BWP12T U11916 ( .A1(b[9]), .A2(n21756), .B1(n21240), .B2(n21773), 
        .ZN(n20938) );
  ND2D1BWP12T U11917 ( .A1(n20939), .A2(n20938), .ZN(n20940) );
  MAOI22D0BWP12T U11918 ( .A1(n22441), .A2(n20940), .B1(n22441), .B2(n20940), 
        .ZN(n21012) );
  NR2D1BWP12T U11919 ( .A1(n21752), .A2(n21678), .ZN(n20942) );
  OAI22D1BWP12T U11920 ( .A1(n22675), .A2(n21749), .B1(n22699), .B2(n22477), 
        .ZN(n20941) );
  AOI211D1BWP12T U11921 ( .A1(n21756), .A2(b[8]), .B(n20942), .C(n20941), .ZN(
        n20943) );
  MAOI22D0BWP12T U11922 ( .A1(a[17]), .A2(n20943), .B1(a[17]), .B2(n20943), 
        .ZN(n21017) );
  FA1D0BWP12T U11923 ( .A(n20946), .B(n20945), .CI(n20944), .CO(n20935), .S(
        n21016) );
  AOI22D1BWP12T U11924 ( .A1(b[9]), .A2(n20981), .B1(b[8]), .B2(n21241), .ZN(
        n20948) );
  AOI22D1BWP12T U11925 ( .A1(b[7]), .A2(n21756), .B1(n21240), .B2(n21623), 
        .ZN(n20947) );
  ND2D1BWP12T U11926 ( .A1(n20948), .A2(n20947), .ZN(n20949) );
  MAOI22D0BWP12T U11927 ( .A1(n22441), .A2(n20949), .B1(n22441), .B2(n20949), 
        .ZN(n21021) );
  FA1D0BWP12T U11928 ( .A(n20952), .B(n20951), .CI(n20950), .CO(n20944), .S(
        n21020) );
  FA1D0BWP12T U11929 ( .A(n20955), .B(n20954), .CI(n20953), .CO(n20950), .S(
        n21025) );
  AOI22D1BWP12T U11930 ( .A1(b[8]), .A2(n20981), .B1(b[7]), .B2(n21241), .ZN(
        n20957) );
  AOI22D1BWP12T U11931 ( .A1(b[6]), .A2(n21756), .B1(n21240), .B2(n21781), 
        .ZN(n20956) );
  ND2D1BWP12T U11932 ( .A1(n20957), .A2(n20956), .ZN(n20958) );
  MAOI22D0BWP12T U11933 ( .A1(n22441), .A2(n20958), .B1(n22441), .B2(n20958), 
        .ZN(n21024) );
  NR2D1BWP12T U11934 ( .A1(n21935), .A2(n21749), .ZN(n20960) );
  OAI22D1BWP12T U11935 ( .A1(n23370), .A2(n22477), .B1(n21752), .B2(n21636), 
        .ZN(n20959) );
  AOI211D1BWP12T U11936 ( .A1(n21756), .A2(b[5]), .B(n20960), .C(n20959), .ZN(
        n20961) );
  MAOI22D0BWP12T U11937 ( .A1(a[17]), .A2(n20961), .B1(a[17]), .B2(n20961), 
        .ZN(n21028) );
  MAOI22D0BWP12T U11938 ( .A1(n20963), .A2(n20962), .B1(n20963), .B2(n20962), 
        .ZN(n21036) );
  NR2D1BWP12T U11939 ( .A1(n21885), .A2(n22477), .ZN(n20965) );
  OAI22D1BWP12T U11940 ( .A1(n23370), .A2(n21749), .B1(n21752), .B2(n21671), 
        .ZN(n20964) );
  AOI211D1BWP12T U11941 ( .A1(n21756), .A2(b[4]), .B(n20965), .C(n20964), .ZN(
        n20966) );
  MAOI22D0BWP12T U11942 ( .A1(a[17]), .A2(n20966), .B1(a[17]), .B2(n20966), 
        .ZN(n21035) );
  AO21D1BWP12T U11943 ( .A1(n20969), .A2(n20968), .B(n20967), .Z(n21040) );
  NR2D1BWP12T U11944 ( .A1(n21885), .A2(n21749), .ZN(n20971) );
  OAI22D1BWP12T U11945 ( .A1(n23017), .A2(n22477), .B1(n21752), .B2(n21797), 
        .ZN(n20970) );
  AOI211D1BWP12T U11946 ( .A1(n21756), .A2(b[3]), .B(n20971), .C(n20970), .ZN(
        n20972) );
  MAOI22D0BWP12T U11947 ( .A1(a[17]), .A2(n20972), .B1(a[17]), .B2(n20972), 
        .ZN(n21039) );
  AO21D1BWP12T U11948 ( .A1(n20975), .A2(n20974), .B(n20973), .Z(n21047) );
  NR2D1BWP12T U11949 ( .A1(n23017), .A2(n21749), .ZN(n20977) );
  OAI22D1BWP12T U11950 ( .A1(n22806), .A2(n22477), .B1(n21752), .B2(n21667), 
        .ZN(n20976) );
  AOI211D1BWP12T U11951 ( .A1(n21756), .A2(b[2]), .B(n20977), .C(n20976), .ZN(
        n20978) );
  MAOI22D0BWP12T U11952 ( .A1(a[17]), .A2(n20978), .B1(a[17]), .B2(n20978), 
        .ZN(n21046) );
  ND2D1BWP12T U11953 ( .A1(b[0]), .A2(a[17]), .ZN(n22535) );
  NR2D1BWP12T U11954 ( .A1(n22535), .A2(n21070), .ZN(n21063) );
  OAI222D1BWP12T U11955 ( .A1(n21752), .A2(n22867), .B1(n22477), .B2(n22009), 
        .C1(n22485), .C2(n21749), .ZN(n21062) );
  NR2D1BWP12T U11956 ( .A1(n21063), .A2(n21062), .ZN(n21061) );
  NR2D1BWP12T U11957 ( .A1(n21061), .A2(n22441), .ZN(n21057) );
  AOI22D1BWP12T U11958 ( .A1(b[1]), .A2(n21241), .B1(n21240), .B2(n21655), 
        .ZN(n20980) );
  ND2D1BWP12T U11959 ( .A1(b[0]), .A2(n21756), .ZN(n20979) );
  OAI211D1BWP12T U11960 ( .A1(n21749), .A2(n22342), .B(n20980), .C(n20979), 
        .ZN(n21056) );
  NR2D1BWP12T U11961 ( .A1(n21057), .A2(n21056), .ZN(n21055) );
  NR2D1BWP12T U11962 ( .A1(n21055), .A2(n22441), .ZN(n20985) );
  AOI22D1BWP12T U11963 ( .A1(b[3]), .A2(n20981), .B1(b[1]), .B2(n21756), .ZN(
        n20983) );
  ND2D1BWP12T U11964 ( .A1(b[2]), .A2(n21241), .ZN(n20982) );
  OAI211D1BWP12T U11965 ( .A1(n21752), .A2(n21659), .B(n20983), .C(n20982), 
        .ZN(n20984) );
  NR2D1BWP12T U11966 ( .A1(n20985), .A2(n20984), .ZN(n20986) );
  NR2D1BWP12T U11967 ( .A1(n21051), .A2(n21050), .ZN(n21049) );
  AOI21D1BWP12T U11968 ( .A1(n20986), .A2(a[17]), .B(n21049), .ZN(n21045) );
  INVD1BWP12T U11969 ( .I(n20987), .ZN(n21123) );
  NR2D1BWP12T U11970 ( .A1(n21933), .A2(a[13]), .ZN(n22544) );
  ND2D1BWP12T U11971 ( .A1(a[12]), .A2(a[11]), .ZN(n23566) );
  IND2D1BWP12T U11972 ( .A1(n22544), .B1(n23566), .ZN(n20989) );
  INVD1BWP12T U11973 ( .I(a[13]), .ZN(n22588) );
  ND2D1BWP12T U11974 ( .A1(n22689), .A2(n22642), .ZN(n21869) );
  OAI21D1BWP12T U11975 ( .A1(a[14]), .A2(n22588), .B(n21869), .ZN(n20988) );
  NR2D1BWP12T U11976 ( .A1(n20989), .A2(n20988), .ZN(n21748) );
  ND2D1BWP12T U11977 ( .A1(n21869), .A2(n23566), .ZN(n21184) );
  OAI221D1BWP12T U11978 ( .A1(a[12]), .A2(a[13]), .B1(n22689), .B2(n22588), 
        .C(n21184), .ZN(n21742) );
  NR2D1BWP12T U11979 ( .A1(n21753), .A2(n21742), .ZN(n20994) );
  ND2D1BWP12T U11980 ( .A1(n20989), .A2(n20988), .ZN(n21745) );
  NR2D1BWP12T U11981 ( .A1(a[14]), .A2(n22588), .ZN(n20990) );
  OAI211D1BWP12T U11982 ( .A1(n22544), .A2(n20990), .B(n21869), .C(n23566), 
        .ZN(n21743) );
  OAI22D1BWP12T U11983 ( .A1(n23484), .A2(n21745), .B1(n21743), .B2(n21751), 
        .ZN(n20993) );
  AOI211D1BWP12T U11984 ( .A1(n21748), .A2(b[17]), .B(n20994), .C(n20993), 
        .ZN(n20995) );
  MAOI22D0BWP12T U11985 ( .A1(n20995), .A2(n21933), .B1(n20995), .B2(n21933), 
        .ZN(n21122) );
  FA1D0BWP12T U11986 ( .A(n20998), .B(n20997), .CI(n20996), .CO(n21081), .S(
        n20999) );
  INVD1BWP12T U11987 ( .I(n21743), .ZN(n21076) );
  ND2D1BWP12T U11988 ( .A1(n21000), .A2(n21002), .ZN(n21001) );
  MAOI22D0BWP12T U11989 ( .A1(n21753), .A2(n21001), .B1(n21753), .B2(n21001), 
        .ZN(n21585) );
  INVD1BWP12T U11990 ( .I(n21742), .ZN(n21077) );
  OAI222D1BWP12T U11991 ( .A1(b[15]), .A2(n21005), .B1(b[15]), .B2(n21004), 
        .C1(n21003), .C2(n21002), .ZN(n21006) );
  MAOI22D0BWP12T U11992 ( .A1(n22547), .A2(n21006), .B1(n22547), .B2(n21006), 
        .ZN(n21689) );
  FA1D0BWP12T U11993 ( .A(n21009), .B(n21008), .CI(n21007), .CO(n20996), .S(
        n21010) );
  FA1D0BWP12T U11994 ( .A(n21013), .B(n21012), .CI(n21011), .CO(n21007), .S(
        n21014) );
  INVD1BWP12T U11995 ( .I(n21748), .ZN(n21072) );
  FA1D0BWP12T U11996 ( .A(n21017), .B(n21016), .CI(n21015), .CO(n21011), .S(
        n21018) );
  FA1D0BWP12T U11997 ( .A(n21021), .B(n21020), .CI(n21019), .CO(n21015), .S(
        n21022) );
  INVD1BWP12T U11998 ( .I(n21683), .ZN(n21684) );
  FA1D0BWP12T U11999 ( .A(n21025), .B(n21024), .CI(n21023), .CO(n21019), .S(
        n21026) );
  FA1D0BWP12T U12000 ( .A(n21029), .B(n21028), .CI(n21027), .CO(n21023), .S(
        n21030) );
  INVD1BWP12T U12001 ( .I(n21030), .ZN(n21151) );
  OAI22D1BWP12T U12002 ( .A1(n22675), .A2(n21072), .B1(n22699), .B2(n21742), 
        .ZN(n21032) );
  OAI22D1BWP12T U12003 ( .A1(n22741), .A2(n21745), .B1(n21743), .B2(n21678), 
        .ZN(n21031) );
  NR2D1BWP12T U12004 ( .A1(n21032), .A2(n21031), .ZN(n21033) );
  MAOI22D0BWP12T U12005 ( .A1(n21033), .A2(n21933), .B1(n21033), .B2(n21933), 
        .ZN(n21150) );
  FA1D0BWP12T U12006 ( .A(n21036), .B(n21035), .CI(n21034), .CO(n21027), .S(
        n21037) );
  FA1D0BWP12T U12007 ( .A(n21040), .B(n21039), .CI(n21038), .CO(n21034), .S(
        n21041) );
  INVD1BWP12T U12008 ( .I(n21041), .ZN(n21211) );
  AOI22D1BWP12T U12009 ( .A1(b[8]), .A2(n21748), .B1(b[7]), .B2(n21077), .ZN(
        n21043) );
  ND2D1BWP12T U12010 ( .A1(n21076), .A2(n21781), .ZN(n21042) );
  OAI211D1BWP12T U12011 ( .A1(n21745), .A2(n23370), .B(n21043), .C(n21042), 
        .ZN(n21044) );
  MAOI22D0BWP12T U12012 ( .A1(a[14]), .A2(n21044), .B1(a[14]), .B2(n21044), 
        .ZN(n21210) );
  FA1D0BWP12T U12013 ( .A(n21047), .B(n21046), .CI(n21045), .CO(n21038), .S(
        n21048) );
  INVD1BWP12T U12014 ( .I(n21048), .ZN(n21160) );
  AOI21D1BWP12T U12015 ( .A1(n21051), .A2(n21050), .B(n21049), .ZN(n21205) );
  INVD1BWP12T U12016 ( .I(n21671), .ZN(n21673) );
  AOI22D1BWP12T U12017 ( .A1(b[6]), .A2(n21748), .B1(n21076), .B2(n21673), 
        .ZN(n21053) );
  ND2D1BWP12T U12018 ( .A1(b[5]), .A2(n21077), .ZN(n21052) );
  OAI211D1BWP12T U12019 ( .A1(n21745), .A2(n23017), .B(n21053), .C(n21052), 
        .ZN(n21054) );
  MAOI22D0BWP12T U12020 ( .A1(a[14]), .A2(n21054), .B1(a[14]), .B2(n21054), 
        .ZN(n21204) );
  AOI21D1BWP12T U12021 ( .A1(n21057), .A2(n21056), .B(n21055), .ZN(n21201) );
  OAI22D1BWP12T U12022 ( .A1(n21885), .A2(n21072), .B1(n21743), .B2(n21797), 
        .ZN(n21059) );
  OAI22D1BWP12T U12023 ( .A1(n23017), .A2(n21742), .B1(n22806), .B2(n21745), 
        .ZN(n21058) );
  NR2D1BWP12T U12024 ( .A1(n21059), .A2(n21058), .ZN(n21060) );
  MAOI22D0BWP12T U12025 ( .A1(n21060), .A2(n21933), .B1(n21060), .B2(n21933), 
        .ZN(n21200) );
  AOI21D1BWP12T U12026 ( .A1(n21063), .A2(n21062), .B(n21061), .ZN(n21167) );
  NR2D1BWP12T U12027 ( .A1(n22342), .A2(n21742), .ZN(n21065) );
  OAI22D1BWP12T U12028 ( .A1(n22485), .A2(n21745), .B1(n21659), .B2(n21743), 
        .ZN(n21064) );
  AOI211D1BWP12T U12029 ( .A1(n21748), .A2(b[3]), .B(n21065), .C(n21064), .ZN(
        n21068) );
  NR2D1BWP12T U12030 ( .A1(n22009), .A2(n21745), .ZN(n21067) );
  OAI22D1BWP12T U12031 ( .A1(n22342), .A2(n21072), .B1(n22485), .B2(n21742), 
        .ZN(n21066) );
  AOI211D1BWP12T U12032 ( .A1(n21076), .A2(n21655), .B(n21067), .C(n21066), 
        .ZN(n21180) );
  AOI22D1BWP12T U12033 ( .A1(b[1]), .A2(n21748), .B1(n22864), .B2(n21076), 
        .ZN(n21198) );
  OAI211D1BWP12T U12034 ( .A1(n21742), .A2(n22605), .B(n21198), .C(n21197), 
        .ZN(n21196) );
  ND2D1BWP12T U12035 ( .A1(a[14]), .A2(n21196), .ZN(n21179) );
  ND2D1BWP12T U12036 ( .A1(n21180), .A2(n21179), .ZN(n21178) );
  ND2D1BWP12T U12037 ( .A1(a[14]), .A2(n21178), .ZN(n21069) );
  ND2D1BWP12T U12038 ( .A1(n21068), .A2(n21069), .ZN(n21071) );
  MAOI22D0BWP12T U12039 ( .A1(n21069), .A2(n21068), .B1(n21069), .B2(n21068), 
        .ZN(n21174) );
  NR2D1BWP12T U12040 ( .A1(n22009), .A2(n21070), .ZN(n21173) );
  ND2D1BWP12T U12041 ( .A1(n21174), .A2(n21173), .ZN(n21172) );
  OAI21D1BWP12T U12042 ( .A1(n21071), .A2(n21933), .B(n21172), .ZN(n21166) );
  OAI22D1BWP12T U12043 ( .A1(n23017), .A2(n21072), .B1(n21743), .B2(n21667), 
        .ZN(n21074) );
  OAI22D1BWP12T U12044 ( .A1(n22806), .A2(n21742), .B1(n22342), .B2(n21745), 
        .ZN(n21073) );
  NR2D1BWP12T U12045 ( .A1(n21074), .A2(n21073), .ZN(n21075) );
  MAOI22D0BWP12T U12046 ( .A1(n21075), .A2(n21933), .B1(n21075), .B2(n21933), 
        .ZN(n21165) );
  INVD1BWP12T U12047 ( .I(n21636), .ZN(n21638) );
  AOI22D1BWP12T U12048 ( .A1(b[7]), .A2(n21748), .B1(n21076), .B2(n21638), 
        .ZN(n21079) );
  ND2D1BWP12T U12049 ( .A1(b[6]), .A2(n21077), .ZN(n21078) );
  OAI211D1BWP12T U12050 ( .A1(n21745), .A2(n21885), .B(n21079), .C(n21078), 
        .ZN(n21080) );
  MAOI22D0BWP12T U12051 ( .A1(a[14]), .A2(n21080), .B1(a[14]), .B2(n21080), 
        .ZN(n21158) );
  FA1D0BWP12T U12052 ( .A(n21083), .B(n21082), .CI(n21081), .CO(n21247), .S(
        n20987) );
  AOI22D1BWP12T U12053 ( .A1(b[13]), .A2(n21756), .B1(n21240), .B2(n21689), 
        .ZN(n21085) );
  ND2D1BWP12T U12054 ( .A1(b[14]), .A2(n21241), .ZN(n21084) );
  OAI211D1BWP12T U12055 ( .A1(n21749), .A2(n23484), .B(n21085), .C(n21084), 
        .ZN(n21086) );
  MAOI22D0BWP12T U12056 ( .A1(n22441), .A2(n21086), .B1(n22441), .B2(n21086), 
        .ZN(n21246) );
  NR2D1BWP12T U12057 ( .A1(n22612), .A2(n21764), .ZN(n21088) );
  OAI22D1BWP12T U12058 ( .A1(n21887), .A2(n21767), .B1(n21766), .B2(n21683), 
        .ZN(n21087) );
  AOI211D1BWP12T U12059 ( .A1(n21770), .A2(b[10]), .B(n21088), .C(n21087), 
        .ZN(n21089) );
  MAOI22D0BWP12T U12060 ( .A1(a[20]), .A2(n21089), .B1(a[20]), .B2(n21089), 
        .ZN(n21218) );
  FA1D0BWP12T U12061 ( .A(n21092), .B(n21091), .CI(n21090), .CO(n21235), .S(
        n20837) );
  AOI22D1BWP12T U12062 ( .A1(b[6]), .A2(n21779), .B1(n21780), .B2(n21673), 
        .ZN(n21094) );
  ND2D1BWP12T U12063 ( .A1(b[5]), .A2(n21778), .ZN(n21093) );
  OAI211D1BWP12T U12064 ( .A1(n21784), .A2(n23017), .B(n21094), .C(n21093), 
        .ZN(n21095) );
  MAOI22D0BWP12T U12065 ( .A1(a[26]), .A2(n21095), .B1(a[26]), .B2(n21095), 
        .ZN(n21234) );
  NR2D1BWP12T U12066 ( .A1(a[30]), .A2(a[29]), .ZN(n23050) );
  INVD1BWP12T U12067 ( .I(a[30]), .ZN(n21903) );
  NR2D1BWP12T U12068 ( .A1(n21903), .A2(n23376), .ZN(n23556) );
  NR2D1BWP12T U12069 ( .A1(n23050), .A2(n23556), .ZN(n21789) );
  ND2D1BWP12T U12070 ( .A1(b[0]), .A2(n21789), .ZN(n21222) );
  OAI22D1BWP12T U12071 ( .A1(n22342), .A2(n21799), .B1(n21659), .B2(n21798), 
        .ZN(n21096) );
  AOI21D1BWP12T U12072 ( .A1(b[1]), .A2(n21802), .B(n21096), .ZN(n21097) );
  OAI21D1BWP12T U12073 ( .A1(n22806), .A2(n21796), .B(n21097), .ZN(n21225) );
  NR2D1BWP12T U12074 ( .A1(n21098), .A2(n23376), .ZN(n21226) );
  MOAI22D0BWP12T U12075 ( .A1(n21225), .A2(n21226), .B1(n21225), .B2(n21226), 
        .ZN(n21099) );
  NR2D1BWP12T U12076 ( .A1(n21222), .A2(n21099), .ZN(n21227) );
  AOI21D1BWP12T U12077 ( .A1(n21222), .A2(n21099), .B(n21227), .ZN(n21233) );
  FA1D0BWP12T U12078 ( .A(n21104), .B(n21103), .CI(n21102), .CO(n21216), .S(
        n21083) );
  INVD1BWP12T U12079 ( .I(n21105), .ZN(n21250) );
  NR2D1BWP12T U12080 ( .A1(n21753), .A2(n21745), .ZN(n21110) );
  ND2D1BWP12T U12081 ( .A1(n21107), .A2(n21106), .ZN(n21108) );
  MAOI22D0BWP12T U12082 ( .A1(b[18]), .A2(n21108), .B1(b[18]), .B2(n21108), 
        .ZN(n21573) );
  OAI22D1BWP12T U12083 ( .A1(n21750), .A2(n21742), .B1(n21743), .B2(n21573), 
        .ZN(n21109) );
  AOI211D1BWP12T U12084 ( .A1(n21748), .A2(b[18]), .B(n21110), .C(n21109), 
        .ZN(n21111) );
  MAOI22D0BWP12T U12085 ( .A1(n21111), .A2(n21933), .B1(n21111), .B2(n21933), 
        .ZN(n21249) );
  ND2D1BWP12T U12086 ( .A1(a[10]), .A2(a[9]), .ZN(n23565) );
  INVD1BWP12T U12087 ( .I(a[10]), .ZN(n22677) );
  INVD1BWP12T U12088 ( .I(a[9]), .ZN(n22700) );
  ND2D1BWP12T U12089 ( .A1(n22677), .A2(n22700), .ZN(n22634) );
  OAI33D1BWP12T U12090 ( .A1(a[11]), .A2(n23565), .A3(n21966), .B1(n22642), 
        .B2(n22634), .B3(a[8]), .ZN(n21763) );
  AOI22D1BWP12T U12091 ( .A1(a[9]), .A2(n21966), .B1(a[8]), .B2(n22700), .ZN(
        n21189) );
  ND3D1BWP12T U12092 ( .A1(n22634), .A2(n23565), .A3(n21189), .ZN(n21757) );
  OAI22D1BWP12T U12093 ( .A1(n22677), .A2(a[11]), .B1(n22642), .B2(a[10]), 
        .ZN(n21113) );
  INVD1BWP12T U12094 ( .I(n21189), .ZN(n21114) );
  IND2D1BWP12T U12095 ( .A1(n21113), .B1(n21114), .ZN(n21760) );
  ND2D1BWP12T U12096 ( .A1(n21114), .A2(n21113), .ZN(n21758) );
  ND2D1BWP12T U12097 ( .A1(n21116), .A2(n21115), .ZN(n21117) );
  MAOI22D0BWP12T U12098 ( .A1(b[21]), .A2(n21117), .B1(b[21]), .B2(n21117), 
        .ZN(n21710) );
  ND2D1BWP12T U12099 ( .A1(n21119), .A2(n21118), .ZN(n21120) );
  MAOI22D0BWP12T U12100 ( .A1(b[20]), .A2(n21120), .B1(b[20]), .B2(n21120), 
        .ZN(n21744) );
  FA1D0BWP12T U12101 ( .A(n21123), .B(n21122), .CI(n21121), .CO(n21251), .S(
        n21124) );
  ND2D1BWP12T U12102 ( .A1(n21126), .A2(n21125), .ZN(n21127) );
  MAOI22D0BWP12T U12103 ( .A1(b[19]), .A2(n21127), .B1(b[19]), .B2(n21127), 
        .ZN(n21700) );
  INVD1BWP12T U12104 ( .I(n21131), .ZN(n21271) );
  NR2D1BWP12T U12105 ( .A1(n21750), .A2(n21757), .ZN(n21133) );
  OAI22D1BWP12T U12106 ( .A1(n22418), .A2(n21760), .B1(n21758), .B2(n21573), 
        .ZN(n21132) );
  AOI211D1BWP12T U12107 ( .A1(b[16]), .A2(n21763), .B(n21133), .C(n21132), 
        .ZN(n21134) );
  MAOI22D0BWP12T U12108 ( .A1(a[11]), .A2(n21134), .B1(a[11]), .B2(n21134), 
        .ZN(n21270) );
  NR2D1BWP12T U12109 ( .A1(n21753), .A2(n21757), .ZN(n21136) );
  OAI22D1BWP12T U12110 ( .A1(n21750), .A2(n21760), .B1(n21751), .B2(n21758), 
        .ZN(n21135) );
  AOI211D1BWP12T U12111 ( .A1(b[15]), .A2(n21763), .B(n21136), .C(n21135), 
        .ZN(n21137) );
  MAOI22D0BWP12T U12112 ( .A1(a[11]), .A2(n21137), .B1(a[11]), .B2(n21137), 
        .ZN(n21278) );
  INVD1BWP12T U12113 ( .I(n21139), .ZN(n21277) );
  INVD1BWP12T U12114 ( .I(n21141), .ZN(n21282) );
  INVD1BWP12T U12115 ( .I(n21758), .ZN(n21208) );
  INVD1BWP12T U12116 ( .I(n21763), .ZN(n21207) );
  NR2D1BWP12T U12117 ( .A1(n21207), .A2(n22547), .ZN(n21143) );
  OAI22D1BWP12T U12118 ( .A1(n21753), .A2(n21760), .B1(n23484), .B2(n21757), 
        .ZN(n21142) );
  AOI211D1BWP12T U12119 ( .A1(n21585), .A2(n21208), .B(n21143), .C(n21142), 
        .ZN(n21144) );
  MAOI22D0BWP12T U12120 ( .A1(a[11]), .A2(n21144), .B1(a[11]), .B2(n21144), 
        .ZN(n21281) );
  FA1D0BWP12T U12121 ( .A(n21151), .B(n21150), .CI(n21149), .CO(n21147), .S(
        n21152) );
  OAI22D1BWP12T U12122 ( .A1(n22612), .A2(n21760), .B1(n21758), .B2(n21683), 
        .ZN(n21154) );
  OAI22D1BWP12T U12123 ( .A1(n21207), .A2(n22675), .B1(n21887), .B2(n21757), 
        .ZN(n21153) );
  NR2D1BWP12T U12124 ( .A1(n21154), .A2(n21153), .ZN(n21155) );
  MAOI22D0BWP12T U12125 ( .A1(a[11]), .A2(n21155), .B1(a[11]), .B2(n21155), 
        .ZN(n21292) );
  INVD1BWP12T U12126 ( .I(n21157), .ZN(n21291) );
  FA1D0BWP12T U12127 ( .A(n21160), .B(n21159), .CI(n21158), .CO(n21209), .S(
        n21161) );
  NR2D1BWP12T U12128 ( .A1(n22741), .A2(n21760), .ZN(n21163) );
  OAI22D1BWP12T U12129 ( .A1(n21207), .A2(n23370), .B1(n21935), .B2(n21757), 
        .ZN(n21162) );
  AOI211D1BWP12T U12130 ( .A1(n21781), .A2(n21208), .B(n21163), .C(n21162), 
        .ZN(n21164) );
  MAOI22D0BWP12T U12131 ( .A1(a[11]), .A2(n21164), .B1(a[11]), .B2(n21164), 
        .ZN(n21357) );
  FA1D0BWP12T U12132 ( .A(n21167), .B(n21166), .CI(n21165), .CO(n21199), .S(
        n21168) );
  INVD1BWP12T U12133 ( .I(n21168), .ZN(n21305) );
  OAI22D1BWP12T U12134 ( .A1(n21935), .A2(n21760), .B1(n21758), .B2(n21636), 
        .ZN(n21170) );
  OAI22D1BWP12T U12135 ( .A1(n21207), .A2(n21885), .B1(n23370), .B2(n21757), 
        .ZN(n21169) );
  NR2D1BWP12T U12136 ( .A1(n21170), .A2(n21169), .ZN(n21171) );
  MAOI22D0BWP12T U12137 ( .A1(a[11]), .A2(n21171), .B1(a[11]), .B2(n21171), 
        .ZN(n21304) );
  OAI21D1BWP12T U12138 ( .A1(n21174), .A2(n21173), .B(n21172), .ZN(n21309) );
  OAI22D1BWP12T U12139 ( .A1(n23370), .A2(n21760), .B1(n21758), .B2(n21671), 
        .ZN(n21176) );
  OAI22D1BWP12T U12140 ( .A1(n21207), .A2(n23017), .B1(n21885), .B2(n21757), 
        .ZN(n21175) );
  NR2D1BWP12T U12141 ( .A1(n21176), .A2(n21175), .ZN(n21177) );
  MAOI22D0BWP12T U12142 ( .A1(a[11]), .A2(n21177), .B1(a[11]), .B2(n21177), 
        .ZN(n21308) );
  OAI21D1BWP12T U12143 ( .A1(n21180), .A2(n21179), .B(n21178), .ZN(n21316) );
  OAI22D1BWP12T U12144 ( .A1(n21885), .A2(n21760), .B1(n21758), .B2(n21797), 
        .ZN(n21182) );
  OAI22D1BWP12T U12145 ( .A1(n21207), .A2(n22806), .B1(n23017), .B2(n21757), 
        .ZN(n21181) );
  NR2D1BWP12T U12146 ( .A1(n21182), .A2(n21181), .ZN(n21183) );
  MAOI22D0BWP12T U12147 ( .A1(a[11]), .A2(n21183), .B1(a[11]), .B2(n21183), 
        .ZN(n21315) );
  NR2D1BWP12T U12148 ( .A1(n22009), .A2(n21184), .ZN(n21328) );
  OAI22D1BWP12T U12149 ( .A1(n22806), .A2(n21760), .B1(n21659), .B2(n21758), 
        .ZN(n21186) );
  OAI22D1BWP12T U12150 ( .A1(n21207), .A2(n22485), .B1(n22342), .B2(n21757), 
        .ZN(n21185) );
  NR2D1BWP12T U12151 ( .A1(n21186), .A2(n21185), .ZN(n21191) );
  NR2D1BWP12T U12152 ( .A1(n22485), .A2(n21757), .ZN(n21188) );
  OAI22D1BWP12T U12153 ( .A1(n21207), .A2(n22009), .B1(n22342), .B2(n21760), 
        .ZN(n21187) );
  AOI211D1BWP12T U12154 ( .A1(n21208), .A2(n21655), .B(n21188), .C(n21187), 
        .ZN(n21335) );
  OA222D1BWP12T U12155 ( .A1(n22605), .A2(n21757), .B1(n22485), .B2(n21760), 
        .C1(n22867), .C2(n21758), .Z(n21341) );
  NR2D1BWP12T U12156 ( .A1(n22009), .A2(n21189), .ZN(n21469) );
  ND2D1BWP12T U12157 ( .A1(a[11]), .A2(n21469), .ZN(n21340) );
  ND2D1BWP12T U12158 ( .A1(n21341), .A2(n21340), .ZN(n21339) );
  ND2D1BWP12T U12159 ( .A1(a[11]), .A2(n21339), .ZN(n21334) );
  ND2D1BWP12T U12160 ( .A1(n21335), .A2(n21334), .ZN(n21333) );
  ND2D1BWP12T U12161 ( .A1(a[11]), .A2(n21333), .ZN(n21190) );
  MAOI22D0BWP12T U12162 ( .A1(n21191), .A2(n21190), .B1(n21191), .B2(n21190), 
        .ZN(n21329) );
  INR3D0BWP12T U12163 ( .A1(n21191), .B1(n22642), .B2(n21333), .ZN(n21192) );
  AOI21D1BWP12T U12164 ( .A1(n21328), .A2(n21329), .B(n21192), .ZN(n21326) );
  OAI22D1BWP12T U12165 ( .A1(n23017), .A2(n21760), .B1(n21758), .B2(n21667), 
        .ZN(n21194) );
  OAI22D1BWP12T U12166 ( .A1(n21207), .A2(n22342), .B1(n22806), .B2(n21757), 
        .ZN(n21193) );
  NR2D1BWP12T U12167 ( .A1(n21194), .A2(n21193), .ZN(n21195) );
  MAOI22D0BWP12T U12168 ( .A1(a[11]), .A2(n21195), .B1(a[11]), .B2(n21195), 
        .ZN(n21325) );
  OAI21D1BWP12T U12169 ( .A1(n21198), .A2(n21197), .B(n21196), .ZN(n21324) );
  FA1D0BWP12T U12170 ( .A(n21201), .B(n21200), .CI(n21199), .CO(n21203), .S(
        n21202) );
  INVD1BWP12T U12171 ( .I(n21202), .ZN(n21355) );
  FA1D0BWP12T U12172 ( .A(n21205), .B(n21204), .CI(n21203), .CO(n21159), .S(
        n21206) );
  FA1D0BWP12T U12173 ( .A(n21211), .B(n21210), .CI(n21209), .CO(n21156), .S(
        n21212) );
  ND2D1BWP12T U12174 ( .A1(n21214), .A2(n21213), .ZN(n21215) );
  MAOI22D0BWP12T U12175 ( .A1(b[22]), .A2(n21215), .B1(b[22]), .B2(n21215), 
        .ZN(n21565) );
  FA1D0BWP12T U12176 ( .A(n21218), .B(n21217), .CI(n21216), .CO(n21828), .S(
        n21245) );
  NR2D1BWP12T U12177 ( .A1(n21934), .A2(n21764), .ZN(n21220) );
  OAI22D1BWP12T U12178 ( .A1(n22612), .A2(n21767), .B1(n21766), .B2(n21595), 
        .ZN(n21219) );
  AOI211D1BWP12T U12179 ( .A1(n21770), .A2(b[11]), .B(n21220), .C(n21219), 
        .ZN(n21221) );
  MAOI22D0BWP12T U12180 ( .A1(a[20]), .A2(n21221), .B1(a[20]), .B2(n21221), 
        .ZN(n21827) );
  NR2D1BWP12T U12181 ( .A1(n23642), .A2(n21222), .ZN(n21224) );
  AOI22D1BWP12T U12182 ( .A1(a[31]), .A2(n23050), .B1(n23642), .B2(n23556), 
        .ZN(n21788) );
  MOAI22D0BWP12T U12183 ( .A1(n21788), .A2(n22009), .B1(b[1]), .B2(n21789), 
        .ZN(n21223) );
  NR2D1BWP12T U12184 ( .A1(n21224), .A2(n21223), .ZN(n21787) );
  AO21D1BWP12T U12185 ( .A1(n21224), .A2(n21223), .B(n21787), .Z(n21817) );
  NR2D1BWP12T U12186 ( .A1(n21226), .A2(n21225), .ZN(n21228) );
  AOI21D1BWP12T U12187 ( .A1(n21228), .A2(a[29]), .B(n21227), .ZN(n21816) );
  NR2D1BWP12T U12188 ( .A1(n23017), .A2(n21796), .ZN(n21230) );
  OAI22D1BWP12T U12189 ( .A1(n22806), .A2(n21799), .B1(n21798), .B2(n21667), 
        .ZN(n21229) );
  AOI211D1BWP12T U12190 ( .A1(n21802), .A2(b[2]), .B(n21230), .C(n21229), .ZN(
        n21231) );
  MAOI22D0BWP12T U12191 ( .A1(a[29]), .A2(n21231), .B1(a[29]), .B2(n21231), 
        .ZN(n21815) );
  FA1D0BWP12T U12192 ( .A(n21235), .B(n21234), .CI(n21233), .CO(n21820), .S(
        n21100) );
  AOI22D1BWP12T U12193 ( .A1(b[14]), .A2(n21756), .B1(n21240), .B2(n21585), 
        .ZN(n21243) );
  ND2D1BWP12T U12194 ( .A1(b[15]), .A2(n21241), .ZN(n21242) );
  OAI211D1BWP12T U12195 ( .A1(n21749), .A2(n21753), .B(n21243), .C(n21242), 
        .ZN(n21244) );
  MAOI22D0BWP12T U12196 ( .A1(n22441), .A2(n21244), .B1(n22441), .B2(n21244), 
        .ZN(n21822) );
  FA1D0BWP12T U12197 ( .A(n21247), .B(n21246), .CI(n21245), .CO(n21821), .S(
        n21105) );
  FA1D0BWP12T U12198 ( .A(n21251), .B(n21250), .CI(n21249), .CO(n21809), .S(
        n21112) );
  ND2D1BWP12T U12199 ( .A1(n21255), .A2(n21254), .ZN(n21256) );
  MAOI22D0BWP12T U12200 ( .A1(b[24]), .A2(n21256), .B1(b[24]), .B2(n21256), 
        .ZN(n21555) );
  ND2D1BWP12T U12201 ( .A1(n21260), .A2(n21259), .ZN(n21261) );
  MAOI22D0BWP12T U12202 ( .A1(b[23]), .A2(n21261), .B1(b[23]), .B2(n21261), 
        .ZN(n21759) );
  NR2D1BWP12T U12203 ( .A1(n23498), .A2(n21724), .ZN(n21267) );
  OAI22D1BWP12T U12204 ( .A1(n22293), .A2(n21727), .B1(n21725), .B2(n21710), 
        .ZN(n21266) );
  AOI211D1BWP12T U12205 ( .A1(b[19]), .A2(n21730), .B(n21267), .C(n21266), 
        .ZN(n21268) );
  MAOI22D0BWP12T U12206 ( .A1(n21268), .A2(n21966), .B1(n21268), .B2(n21966), 
        .ZN(n21383) );
  FA1D0BWP12T U12207 ( .A(n21271), .B(n21270), .CI(n21269), .CO(n21264), .S(
        n21272) );
  INVD1BWP12T U12208 ( .I(n21272), .ZN(n21382) );
  NR2D1BWP12T U12209 ( .A1(n21944), .A2(n21724), .ZN(n21274) );
  OAI22D1BWP12T U12210 ( .A1(n23498), .A2(n21727), .B1(n21725), .B2(n21744), 
        .ZN(n21273) );
  AOI211D1BWP12T U12211 ( .A1(b[18]), .A2(n21730), .B(n21274), .C(n21273), 
        .ZN(n21275) );
  MAOI22D0BWP12T U12212 ( .A1(n21275), .A2(n21966), .B1(n21275), .B2(n21966), 
        .ZN(n21387) );
  FA1D0BWP12T U12213 ( .A(n21278), .B(n21277), .CI(n21276), .CO(n21269), .S(
        n21279) );
  INVD1BWP12T U12214 ( .I(n21279), .ZN(n21386) );
  FA1D0BWP12T U12215 ( .A(n21282), .B(n21281), .CI(n21280), .CO(n21276), .S(
        n21283) );
  INVD1BWP12T U12216 ( .I(n21724), .ZN(n21346) );
  INVD1BWP12T U12217 ( .I(n21725), .ZN(n21347) );
  FA1D0BWP12T U12218 ( .A(n21292), .B(n21291), .CI(n21290), .CO(n21288), .S(
        n21293) );
  AOI22D1BWP12T U12219 ( .A1(b[10]), .A2(n21730), .B1(b[11]), .B2(n21346), 
        .ZN(n21295) );
  ND2D1BWP12T U12220 ( .A1(n21347), .A2(n21684), .ZN(n21294) );
  OAI211D1BWP12T U12221 ( .A1(n21727), .A2(n22612), .B(n21295), .C(n21294), 
        .ZN(n21296) );
  MAOI22D0BWP12T U12222 ( .A1(a[8]), .A2(n21296), .B1(a[8]), .B2(n21296), .ZN(
        n21497) );
  AOI22D1BWP12T U12223 ( .A1(b[10]), .A2(n21346), .B1(b[9]), .B2(n21730), .ZN(
        n21298) );
  ND2D1BWP12T U12224 ( .A1(n21347), .A2(n21773), .ZN(n21297) );
  OAI211D1BWP12T U12225 ( .A1(n21727), .A2(n21887), .B(n21298), .C(n21297), 
        .ZN(n21299) );
  MAOI22D0BWP12T U12226 ( .A1(a[8]), .A2(n21299), .B1(a[8]), .B2(n21299), .ZN(
        n21493) );
  NR2D1BWP12T U12227 ( .A1(n21725), .A2(n21678), .ZN(n21301) );
  OAI22D1BWP12T U12228 ( .A1(n22675), .A2(n21727), .B1(n22699), .B2(n21724), 
        .ZN(n21300) );
  AOI211D1BWP12T U12229 ( .A1(b[8]), .A2(n21730), .B(n21301), .C(n21300), .ZN(
        n21302) );
  MAOI22D0BWP12T U12230 ( .A1(n21302), .A2(n21966), .B1(n21302), .B2(n21966), 
        .ZN(n21423) );
  FA1D0BWP12T U12231 ( .A(n21305), .B(n21304), .CI(n21303), .CO(n21356), .S(
        n21306) );
  INVD1BWP12T U12232 ( .I(n21306), .ZN(n21422) );
  FA1D0BWP12T U12233 ( .A(n21309), .B(n21308), .CI(n21307), .CO(n21303), .S(
        n21310) );
  INVD1BWP12T U12234 ( .I(n21310), .ZN(n21427) );
  AOI22D1BWP12T U12235 ( .A1(b[8]), .A2(n21346), .B1(b[7]), .B2(n21730), .ZN(
        n21312) );
  ND2D1BWP12T U12236 ( .A1(n21347), .A2(n21623), .ZN(n21311) );
  OAI211D1BWP12T U12237 ( .A1(n21727), .A2(n22699), .B(n21312), .C(n21311), 
        .ZN(n21313) );
  MAOI22D0BWP12T U12238 ( .A1(a[8]), .A2(n21313), .B1(a[8]), .B2(n21313), .ZN(
        n21426) );
  FA1D0BWP12T U12239 ( .A(n21316), .B(n21315), .CI(n21314), .CO(n21307), .S(
        n21317) );
  INVD1BWP12T U12240 ( .I(n21317), .ZN(n21434) );
  AOI22D1BWP12T U12241 ( .A1(b[7]), .A2(n21346), .B1(b[6]), .B2(n21730), .ZN(
        n21319) );
  ND2D1BWP12T U12242 ( .A1(n21347), .A2(n21781), .ZN(n21318) );
  OAI211D1BWP12T U12243 ( .A1(n21727), .A2(n22741), .B(n21319), .C(n21318), 
        .ZN(n21320) );
  MAOI22D0BWP12T U12244 ( .A1(a[8]), .A2(n21320), .B1(a[8]), .B2(n21320), .ZN(
        n21433) );
  AOI22D1BWP12T U12245 ( .A1(b[5]), .A2(n21730), .B1(n21347), .B2(n21638), 
        .ZN(n21322) );
  ND2D1BWP12T U12246 ( .A1(b[6]), .A2(n21346), .ZN(n21321) );
  OAI211D1BWP12T U12247 ( .A1(n21727), .A2(n21935), .B(n21322), .C(n21321), 
        .ZN(n21323) );
  MAOI22D0BWP12T U12248 ( .A1(a[8]), .A2(n21323), .B1(a[8]), .B2(n21323), .ZN(
        n21441) );
  FA1D0BWP12T U12249 ( .A(n21326), .B(n21325), .CI(n21324), .CO(n21314), .S(
        n21327) );
  INVD1BWP12T U12250 ( .I(n21327), .ZN(n21440) );
  MAOI22D0BWP12T U12251 ( .A1(n21329), .A2(n21328), .B1(n21329), .B2(n21328), 
        .ZN(n21451) );
  AOI22D1BWP12T U12252 ( .A1(b[4]), .A2(n21730), .B1(n21347), .B2(n21673), 
        .ZN(n21331) );
  ND2D1BWP12T U12253 ( .A1(b[5]), .A2(n21346), .ZN(n21330) );
  OAI211D1BWP12T U12254 ( .A1(n21727), .A2(n23370), .B(n21331), .C(n21330), 
        .ZN(n21332) );
  MAOI22D0BWP12T U12255 ( .A1(a[8]), .A2(n21332), .B1(a[8]), .B2(n21332), .ZN(
        n21450) );
  OA21D1BWP12T U12256 ( .A1(n21335), .A2(n21334), .B(n21333), .Z(n21458) );
  NR2D1BWP12T U12257 ( .A1(n23017), .A2(n21724), .ZN(n21337) );
  OAI22D1BWP12T U12258 ( .A1(n21885), .A2(n21727), .B1(n21725), .B2(n21797), 
        .ZN(n21336) );
  AOI211D1BWP12T U12259 ( .A1(b[3]), .A2(n21730), .B(n21337), .C(n21336), .ZN(
        n21338) );
  MAOI22D0BWP12T U12260 ( .A1(n21338), .A2(n21966), .B1(n21338), .B2(n21966), 
        .ZN(n21457) );
  OA21D1BWP12T U12261 ( .A1(n21341), .A2(n21340), .B(n21339), .Z(n21465) );
  OAI22D1BWP12T U12262 ( .A1(n22485), .A2(n21727), .B1(n22867), .B2(n21725), 
        .ZN(n21490) );
  ND2D1BWP12T U12263 ( .A1(b[0]), .A2(n21342), .ZN(n21644) );
  OAI22D1BWP12T U12264 ( .A1(n22605), .A2(n21724), .B1(n21966), .B2(n21644), 
        .ZN(n21343) );
  NR2D1BWP12T U12265 ( .A1(n21490), .A2(n21343), .ZN(n21489) );
  NR2D1BWP12T U12266 ( .A1(n21489), .A2(n21966), .ZN(n21475) );
  AOI22D1BWP12T U12267 ( .A1(b[1]), .A2(n21346), .B1(n21347), .B2(n21655), 
        .ZN(n21345) );
  ND2D1BWP12T U12268 ( .A1(b[0]), .A2(n21730), .ZN(n21344) );
  OAI211D1BWP12T U12269 ( .A1(n21727), .A2(n22342), .B(n21345), .C(n21344), 
        .ZN(n21474) );
  NR3D1BWP12T U12270 ( .A1(n21475), .A2(n21966), .A3(n21474), .ZN(n21468) );
  AOI22D1BWP12T U12271 ( .A1(b[2]), .A2(n21346), .B1(b[1]), .B2(n21730), .ZN(
        n21350) );
  ND2D1BWP12T U12272 ( .A1(n21348), .A2(n21347), .ZN(n21349) );
  OAI211D1BWP12T U12273 ( .A1(n21727), .A2(n22806), .B(n21350), .C(n21349), 
        .ZN(n21351) );
  MAOI22D0BWP12T U12274 ( .A1(a[8]), .A2(n21351), .B1(a[8]), .B2(n21351), .ZN(
        n21467) );
  NR2D1BWP12T U12275 ( .A1(n22806), .A2(n21724), .ZN(n21353) );
  OAI22D1BWP12T U12276 ( .A1(n23017), .A2(n21727), .B1(n21725), .B2(n21667), 
        .ZN(n21352) );
  AOI211D1BWP12T U12277 ( .A1(b[2]), .A2(n21730), .B(n21353), .C(n21352), .ZN(
        n21354) );
  MAOI22D0BWP12T U12278 ( .A1(n21354), .A2(n21966), .B1(n21354), .B2(n21966), 
        .ZN(n21463) );
  FA1D0BWP12T U12279 ( .A(n21357), .B(n21356), .CI(n21355), .CO(n21359), .S(
        n21358) );
  INVD1BWP12T U12280 ( .I(n21358), .ZN(n21491) );
  INVD1BWP12T U12281 ( .I(n21360), .ZN(n21495) );
  NR2D1BWP12T U12282 ( .A1(n22612), .A2(n21724), .ZN(n21362) );
  OAI22D1BWP12T U12283 ( .A1(n21934), .A2(n21727), .B1(n21725), .B2(n21595), 
        .ZN(n21361) );
  AOI211D1BWP12T U12284 ( .A1(b[11]), .A2(n21730), .B(n21362), .C(n21361), 
        .ZN(n21363) );
  MAOI22D0BWP12T U12285 ( .A1(n21363), .A2(n21966), .B1(n21363), .B2(n21966), 
        .ZN(n21409) );
  INVD1BWP12T U12286 ( .I(n21365), .ZN(n21408) );
  ND2D1BWP12T U12287 ( .A1(n21370), .A2(n21369), .ZN(n21371) );
  MAOI22D0BWP12T U12288 ( .A1(b[27]), .A2(n21371), .B1(b[27]), .B2(n21371), 
        .ZN(n21539) );
  ND2D1BWP12T U12289 ( .A1(n21375), .A2(n21374), .ZN(n21376) );
  MAOI22D0BWP12T U12290 ( .A1(b[26]), .A2(n21376), .B1(b[26]), .B2(n21376), 
        .ZN(n21726) );
  FA1D0BWP12T U12291 ( .A(n21383), .B(n21382), .CI(n21381), .CO(n21379), .S(
        n21384) );
  FA1D0BWP12T U12292 ( .A(n21387), .B(n21386), .CI(n21385), .CO(n21381), .S(
        n21388) );
  NR2D1BWP12T U12293 ( .A1(n23498), .A2(n21731), .ZN(n21394) );
  OAI22D1BWP12T U12294 ( .A1(n21734), .A2(n22418), .B1(n21732), .B2(n21744), 
        .ZN(n21393) );
  AOI211D1BWP12T U12295 ( .A1(n21737), .A2(b[19]), .B(n21394), .C(n21393), 
        .ZN(n21395) );
  MAOI22D0BWP12T U12296 ( .A1(a[5]), .A2(n21395), .B1(a[5]), .B2(n21395), .ZN(
        n21559) );
  INVD1BWP12T U12297 ( .I(n21397), .ZN(n21558) );
  NR2D1BWP12T U12298 ( .A1(n21944), .A2(n21731), .ZN(n21399) );
  OAI22D1BWP12T U12299 ( .A1(n21734), .A2(n21750), .B1(n21732), .B2(n21700), 
        .ZN(n21398) );
  AOI211D1BWP12T U12300 ( .A1(n21737), .A2(b[18]), .B(n21399), .C(n21398), 
        .ZN(n21400) );
  MAOI22D0BWP12T U12301 ( .A1(a[5]), .A2(n21400), .B1(a[5]), .B2(n21400), .ZN(
        n21563) );
  INVD1BWP12T U12302 ( .I(n21402), .ZN(n21562) );
  NR2D1BWP12T U12303 ( .A1(n21750), .A2(n21731), .ZN(n21406) );
  OAI22D1BWP12T U12304 ( .A1(n21734), .A2(n23484), .B1(n21732), .B2(n21751), 
        .ZN(n21405) );
  AOI211D1BWP12T U12305 ( .A1(n21737), .A2(b[16]), .B(n21406), .C(n21405), 
        .ZN(n21407) );
  MAOI22D0BWP12T U12306 ( .A1(a[5]), .A2(n21407), .B1(a[5]), .B2(n21407), .ZN(
        n21570) );
  FA1D0BWP12T U12307 ( .A(n21410), .B(n21409), .CI(n21408), .CO(n21504), .S(
        n21411) );
  INVD1BWP12T U12308 ( .I(n21411), .ZN(n21707) );
  INVD1BWP12T U12309 ( .I(n21737), .ZN(n21499) );
  NR2D1BWP12T U12310 ( .A1(n22547), .A2(n21499), .ZN(n21413) );
  OAI22D1BWP12T U12311 ( .A1(n21734), .A2(n21934), .B1(n23484), .B2(n21731), 
        .ZN(n21412) );
  AOI211D1BWP12T U12312 ( .A1(n21689), .A2(n21502), .B(n21413), .C(n21412), 
        .ZN(n21414) );
  MAOI22D0BWP12T U12313 ( .A1(a[5]), .A2(n21414), .B1(a[5]), .B2(n21414), .ZN(
        n21697) );
  OAI22D1BWP12T U12314 ( .A1(n21734), .A2(n22612), .B1(n21732), .B2(n21765), 
        .ZN(n21416) );
  OAI22D1BWP12T U12315 ( .A1(n22547), .A2(n21731), .B1(n21934), .B2(n21499), 
        .ZN(n21415) );
  NR2D1BWP12T U12316 ( .A1(n21416), .A2(n21415), .ZN(n21417) );
  MAOI22D0BWP12T U12317 ( .A1(a[5]), .A2(n21417), .B1(a[5]), .B2(n21417), .ZN(
        n21693) );
  OAI22D1BWP12T U12318 ( .A1(n21734), .A2(n21887), .B1(n21732), .B2(n21595), 
        .ZN(n21419) );
  OAI22D1BWP12T U12319 ( .A1(n21934), .A2(n21731), .B1(n22612), .B2(n21499), 
        .ZN(n21418) );
  NR2D1BWP12T U12320 ( .A1(n21419), .A2(n21418), .ZN(n21420) );
  MAOI22D0BWP12T U12321 ( .A1(a[5]), .A2(n21420), .B1(a[5]), .B2(n21420), .ZN(
        n21581) );
  FA1D0BWP12T U12322 ( .A(n21423), .B(n21422), .CI(n21421), .CO(n21492), .S(
        n21424) );
  INVD1BWP12T U12323 ( .I(n21424), .ZN(n21580) );
  FA1D0BWP12T U12324 ( .A(n21427), .B(n21426), .CI(n21425), .CO(n21421), .S(
        n21428) );
  INVD1BWP12T U12325 ( .I(n21428), .ZN(n21687) );
  OAI22D1BWP12T U12326 ( .A1(n21734), .A2(n22675), .B1(n21732), .B2(n21683), 
        .ZN(n21430) );
  OAI22D1BWP12T U12327 ( .A1(n22612), .A2(n21731), .B1(n21887), .B2(n21499), 
        .ZN(n21429) );
  NR2D1BWP12T U12328 ( .A1(n21430), .A2(n21429), .ZN(n21431) );
  MAOI22D0BWP12T U12329 ( .A1(a[5]), .A2(n21431), .B1(a[5]), .B2(n21431), .ZN(
        n21686) );
  FA1D0BWP12T U12330 ( .A(n21434), .B(n21433), .CI(n21432), .CO(n21425), .S(
        n21435) );
  INVD1BWP12T U12331 ( .I(n21435), .ZN(n21592) );
  OAI22D1BWP12T U12332 ( .A1(n21734), .A2(n22699), .B1(n21887), .B2(n21731), 
        .ZN(n21437) );
  INVD1BWP12T U12333 ( .I(n21773), .ZN(n21608) );
  OAI22D1BWP12T U12334 ( .A1(n22675), .A2(n21499), .B1(n21732), .B2(n21608), 
        .ZN(n21436) );
  NR2D1BWP12T U12335 ( .A1(n21437), .A2(n21436), .ZN(n21438) );
  MAOI22D0BWP12T U12336 ( .A1(a[5]), .A2(n21438), .B1(a[5]), .B2(n21438), .ZN(
        n21591) );
  FA1D0BWP12T U12337 ( .A(n21441), .B(n21440), .CI(n21439), .CO(n21432), .S(
        n21442) );
  INVD1BWP12T U12338 ( .I(n21442), .ZN(n21602) );
  OAI22D1BWP12T U12339 ( .A1(n21734), .A2(n22741), .B1(n22699), .B2(n21499), 
        .ZN(n21444) );
  OAI22D1BWP12T U12340 ( .A1(n22675), .A2(n21731), .B1(n21732), .B2(n21678), 
        .ZN(n21443) );
  NR2D1BWP12T U12341 ( .A1(n21444), .A2(n21443), .ZN(n21445) );
  MAOI22D0BWP12T U12342 ( .A1(a[5]), .A2(n21445), .B1(a[5]), .B2(n21445), .ZN(
        n21601) );
  NR2D1BWP12T U12343 ( .A1(n21734), .A2(n21935), .ZN(n21447) );
  OAI22D1BWP12T U12344 ( .A1(n22699), .A2(n21731), .B1(n22741), .B2(n21499), 
        .ZN(n21446) );
  AOI211D1BWP12T U12345 ( .A1(n21623), .A2(n21502), .B(n21447), .C(n21446), 
        .ZN(n21448) );
  MAOI22D0BWP12T U12346 ( .A1(a[5]), .A2(n21448), .B1(a[5]), .B2(n21448), .ZN(
        n21681) );
  FA1D0BWP12T U12347 ( .A(n21451), .B(n21450), .CI(n21449), .CO(n21439), .S(
        n21452) );
  INVD1BWP12T U12348 ( .I(n21452), .ZN(n21680) );
  NR2D1BWP12T U12349 ( .A1(n21734), .A2(n23370), .ZN(n21454) );
  OAI22D1BWP12T U12350 ( .A1(n22741), .A2(n21731), .B1(n21935), .B2(n21499), 
        .ZN(n21453) );
  AOI211D1BWP12T U12351 ( .A1(n21781), .A2(n21502), .B(n21454), .C(n21453), 
        .ZN(n21455) );
  MAOI22D0BWP12T U12352 ( .A1(a[5]), .A2(n21455), .B1(a[5]), .B2(n21455), .ZN(
        n21606) );
  FA1D0BWP12T U12353 ( .A(n21458), .B(n21457), .CI(n21456), .CO(n21449), .S(
        n21459) );
  INVD1BWP12T U12354 ( .I(n21459), .ZN(n21605) );
  OAI22D1BWP12T U12355 ( .A1(n21734), .A2(n21885), .B1(n21732), .B2(n21636), 
        .ZN(n21461) );
  OAI22D1BWP12T U12356 ( .A1(n21935), .A2(n21731), .B1(n23370), .B2(n21499), 
        .ZN(n21460) );
  NR2D1BWP12T U12357 ( .A1(n21461), .A2(n21460), .ZN(n21462) );
  MAOI22D0BWP12T U12358 ( .A1(a[5]), .A2(n21462), .B1(a[5]), .B2(n21462), .ZN(
        n21616) );
  FA1D0BWP12T U12359 ( .A(n21465), .B(n21464), .CI(n21463), .CO(n21456), .S(
        n21466) );
  INVD1BWP12T U12360 ( .I(n21466), .ZN(n21615) );
  FA1D0BWP12T U12361 ( .A(n21469), .B(n21468), .CI(n21467), .CO(n21464), .S(
        n21470) );
  INVD1BWP12T U12362 ( .I(n21470), .ZN(n21620) );
  OAI22D1BWP12T U12363 ( .A1(n21734), .A2(n23017), .B1(n21732), .B2(n21671), 
        .ZN(n21472) );
  OAI22D1BWP12T U12364 ( .A1(n23370), .A2(n21731), .B1(n21885), .B2(n21499), 
        .ZN(n21471) );
  NR2D1BWP12T U12365 ( .A1(n21472), .A2(n21471), .ZN(n21473) );
  MAOI22D0BWP12T U12366 ( .A1(a[5]), .A2(n21473), .B1(a[5]), .B2(n21473), .ZN(
        n21619) );
  MOAI22D0BWP12T U12367 ( .A1(n21475), .A2(n21474), .B1(n21475), .B2(n21474), 
        .ZN(n21630) );
  OAI22D1BWP12T U12368 ( .A1(n21734), .A2(n22806), .B1(n21732), .B2(n21797), 
        .ZN(n21477) );
  OAI22D1BWP12T U12369 ( .A1(n21885), .A2(n21731), .B1(n23017), .B2(n21499), 
        .ZN(n21476) );
  NR2D1BWP12T U12370 ( .A1(n21477), .A2(n21476), .ZN(n21478) );
  MAOI22D0BWP12T U12371 ( .A1(a[5]), .A2(n21478), .B1(a[5]), .B2(n21478), .ZN(
        n21629) );
  OAI22D1BWP12T U12372 ( .A1(n21734), .A2(n22342), .B1(n21732), .B2(n21667), 
        .ZN(n21480) );
  OAI22D1BWP12T U12373 ( .A1(n23017), .A2(n21731), .B1(n22806), .B2(n21499), 
        .ZN(n21479) );
  NR2D1BWP12T U12374 ( .A1(n21480), .A2(n21479), .ZN(n21481) );
  MAOI22D0BWP12T U12375 ( .A1(a[5]), .A2(n21481), .B1(a[5]), .B2(n21481), .ZN(
        n21634) );
  OAI22D1BWP12T U12376 ( .A1(n21734), .A2(n22485), .B1(n21659), .B2(n21732), 
        .ZN(n21483) );
  OAI22D1BWP12T U12377 ( .A1(n22806), .A2(n21731), .B1(n22342), .B2(n21499), 
        .ZN(n21482) );
  NR2D1BWP12T U12378 ( .A1(n21483), .A2(n21482), .ZN(n21486) );
  NR2D1BWP12T U12379 ( .A1(n22485), .A2(n21499), .ZN(n21485) );
  OAI22D1BWP12T U12380 ( .A1(n21734), .A2(n22009), .B1(n22342), .B2(n21731), 
        .ZN(n21484) );
  AOI211D1BWP12T U12381 ( .A1(n21502), .A2(n21655), .B(n21485), .C(n21484), 
        .ZN(n21653) );
  NR2D1BWP12T U12382 ( .A1(n22605), .A2(n21803), .ZN(n22955) );
  OAI222D1BWP12T U12383 ( .A1(n21732), .A2(n22867), .B1(n21499), .B2(n22009), 
        .C1(n22485), .C2(n21731), .ZN(n21669) );
  AOI21D1BWP12T U12384 ( .A1(n22955), .A2(n21670), .B(n21669), .ZN(n21668) );
  AOI21D1BWP12T U12385 ( .A1(n21653), .A2(n21668), .B(n21803), .ZN(n21487) );
  MAOI22D0BWP12T U12386 ( .A1(n21486), .A2(n21487), .B1(n21486), .B2(n21487), 
        .ZN(n21643) );
  IND3D1BWP12T U12387 ( .A1(n21487), .B1(n21486), .B2(a[5]), .ZN(n21488) );
  OA21D1BWP12T U12388 ( .A1(n21643), .A2(n21644), .B(n21488), .Z(n21633) );
  AO31D1BWP12T U12389 ( .A1(a[8]), .A2(b[0]), .A3(n21490), .B(n21489), .Z(
        n21632) );
  FA1D0BWP12T U12390 ( .A(n21493), .B(n21492), .CI(n21491), .CO(n21496), .S(
        n21494) );
  INVD1BWP12T U12391 ( .I(n21494), .ZN(n21691) );
  FA1D0BWP12T U12392 ( .A(n21497), .B(n21496), .CI(n21495), .CO(n21410), .S(
        n21498) );
  INVD1BWP12T U12393 ( .I(n21498), .ZN(n21695) );
  NR2D1BWP12T U12394 ( .A1(n23484), .A2(n21499), .ZN(n21501) );
  OAI22D1BWP12T U12395 ( .A1(n21734), .A2(n22547), .B1(n21753), .B2(n21731), 
        .ZN(n21500) );
  AOI211D1BWP12T U12396 ( .A1(n21585), .A2(n21502), .B(n21501), .C(n21500), 
        .ZN(n21503) );
  MAOI22D0BWP12T U12397 ( .A1(a[5]), .A2(n21503), .B1(a[5]), .B2(n21503), .ZN(
        n21705) );
  INVD1BWP12T U12398 ( .I(n21505), .ZN(n21568) );
  INVD1BWP12T U12399 ( .I(n21506), .ZN(n21808) );
  NR2D1BWP12T U12400 ( .A1(a[0]), .A2(n23011), .ZN(n21720) );
  ND2D1BWP12T U12401 ( .A1(a[0]), .A2(n23011), .ZN(n21711) );
  INVD1BWP12T U12402 ( .I(n21711), .ZN(n21719) );
  NR2D1BWP12T U12403 ( .A1(a[2]), .A2(n21711), .ZN(n21584) );
  ND2D1BWP12T U12404 ( .A1(a[0]), .A2(a[1]), .ZN(n21716) );
  NR2D1BWP12T U12405 ( .A1(n21882), .A2(n21716), .ZN(n21651) );
  NR2D1BWP12T U12406 ( .A1(n21584), .A2(n21651), .ZN(n21665) );
  NR2D1BWP12T U12407 ( .A1(a[2]), .A2(n21716), .ZN(n21583) );
  NR2D1BWP12T U12408 ( .A1(n21882), .A2(n21711), .ZN(n21690) );
  NR2D1BWP12T U12409 ( .A1(n21583), .A2(n21690), .ZN(n21666) );
  INVD1BWP12T U12410 ( .I(n21666), .ZN(n21656) );
  ND2D1BWP12T U12411 ( .A1(n23490), .A2(n21507), .ZN(n21525) );
  ND2D1BWP12T U12412 ( .A1(b[29]), .A2(n21525), .ZN(n21517) );
  AN2D1BWP12T U12413 ( .A1(n21517), .A2(n21921), .Z(n21510) );
  ND2D1BWP12T U12414 ( .A1(n21656), .A2(n21510), .ZN(n21518) );
  ND2D1BWP12T U12415 ( .A1(b[28]), .A2(n21508), .ZN(n21526) );
  ND2D1BWP12T U12416 ( .A1(n23375), .A2(n21526), .ZN(n21519) );
  INR2D1BWP12T U12417 ( .A1(n21519), .B1(n21921), .ZN(n21509) );
  ND2D1BWP12T U12418 ( .A1(n21509), .A2(n21656), .ZN(n21740) );
  AOI31D1BWP12T U12419 ( .A1(n21665), .A2(n21518), .A3(n21740), .B(n23043), 
        .ZN(n21512) );
  NR4D0BWP12T U12420 ( .A1(b[31]), .A2(n21666), .A3(n21510), .A4(n21509), .ZN(
        n21511) );
  AOI211D1BWP12T U12421 ( .A1(n21720), .A2(b[30]), .B(n21512), .C(n21511), 
        .ZN(n21514) );
  INVD1BWP12T U12422 ( .I(a[0]), .ZN(n23034) );
  ND2D1BWP12T U12423 ( .A1(n23034), .A2(n23011), .ZN(n21868) );
  OAI211D1BWP12T U12424 ( .A1(n21868), .A2(n23375), .B(a[2]), .C(n21514), .ZN(
        n21513) );
  OAI21D1BWP12T U12425 ( .A1(n21514), .A2(a[2]), .B(n21513), .ZN(n21807) );
  INVD1BWP12T U12426 ( .I(n21516), .ZN(n21906) );
  AOI32D1BWP12T U12427 ( .A1(n21517), .A2(n21665), .A3(n21519), .B1(n21666), 
        .B2(n21665), .ZN(n21520) );
  INVD1BWP12T U12428 ( .I(n21518), .ZN(n21739) );
  AOI222D1BWP12T U12429 ( .A1(n21520), .A2(b[30]), .B1(b[29]), .B2(n21720), 
        .C1(n21519), .C2(n21739), .ZN(n21522) );
  OAI211D1BWP12T U12430 ( .A1(n21868), .A2(n23490), .B(a[2]), .C(n21522), .ZN(
        n21521) );
  OAI21D1BWP12T U12431 ( .A1(n21522), .A2(a[2]), .B(n21521), .ZN(n21905) );
  INVD1BWP12T U12432 ( .I(n21524), .ZN(n21955) );
  INVD1BWP12T U12433 ( .I(n21720), .ZN(n21717) );
  NR2D1BWP12T U12434 ( .A1(n23490), .A2(n21717), .ZN(n21530) );
  ND2D1BWP12T U12435 ( .A1(n21526), .A2(n21525), .ZN(n21527) );
  MAOI22D0BWP12T U12436 ( .A1(b[29]), .A2(n21527), .B1(b[29]), .B2(n21527), 
        .ZN(n21733) );
  OAI22D1BWP12T U12437 ( .A1(n23375), .A2(n21711), .B1(n21716), .B2(n21733), 
        .ZN(n21528) );
  NR2D1BWP12T U12438 ( .A1(n21530), .A2(n21528), .ZN(n21532) );
  INVD1BWP12T U12439 ( .I(n21716), .ZN(n22978) );
  OAI22D1BWP12T U12440 ( .A1(n22032), .A2(n21868), .B1(n21711), .B2(n21733), 
        .ZN(n21529) );
  AO211D1BWP12T U12441 ( .A1(b[29]), .A2(n22978), .B(n21882), .C(n21529), .Z(
        n21531) );
  OAI22D1BWP12T U12442 ( .A1(n21532), .A2(a[2]), .B1(n21531), .B2(n21530), 
        .ZN(n21954) );
  INVD1BWP12T U12443 ( .I(n21868), .ZN(n22977) );
  INVD1BWP12T U12444 ( .I(n21537), .ZN(n22057) );
  NR2D1BWP12T U12445 ( .A1(n22088), .A2(n21717), .ZN(n21541) );
  OAI22D1BWP12T U12446 ( .A1(n22032), .A2(n21711), .B1(n21716), .B2(n21539), 
        .ZN(n21538) );
  NR2D1BWP12T U12447 ( .A1(n21541), .A2(n21538), .ZN(n21543) );
  MAOI22D0BWP12T U12448 ( .A1(b[25]), .A2(n22977), .B1(n21711), .B2(n21539), 
        .ZN(n21540) );
  OAI211D1BWP12T U12449 ( .A1(n22032), .A2(n21716), .B(a[2]), .C(n21540), .ZN(
        n21542) );
  OAI22D1BWP12T U12450 ( .A1(n21543), .A2(a[2]), .B1(n21542), .B2(n21541), 
        .ZN(n22056) );
  INVD1BWP12T U12451 ( .I(n21547), .ZN(n22149) );
  OAI22D1BWP12T U12452 ( .A1(n21556), .A2(n21717), .B1(n21716), .B2(n21549), 
        .ZN(n21548) );
  AOI22D1BWP12T U12453 ( .A1(b[25]), .A2(n21584), .B1(n21882), .B2(n21548), 
        .ZN(n21552) );
  MAOI22D0BWP12T U12454 ( .A1(b[23]), .A2(n22977), .B1(n21711), .B2(n21549), 
        .ZN(n21550) );
  OAI211D1BWP12T U12455 ( .A1(n22150), .A2(n21716), .B(a[2]), .C(n21550), .ZN(
        n21551) );
  AOI32D1BWP12T U12456 ( .A1(n21720), .A2(n21552), .A3(b[24]), .B1(n21551), 
        .B2(n21552), .ZN(n22148) );
  FA1D0BWP12T U12457 ( .A(n21559), .B(n21558), .CI(n21557), .CO(n21553), .S(
        n21560) );
  INVD1BWP12T U12458 ( .I(n21560), .ZN(n22231) );
  FA1D0BWP12T U12459 ( .A(n21563), .B(n21562), .CI(n21561), .CO(n21557), .S(
        n21564) );
  INVD1BWP12T U12460 ( .I(n21690), .ZN(n22992) );
  INVD1BWP12T U12461 ( .I(n21567), .ZN(n22316) );
  FA1D0BWP12T U12462 ( .A(n21570), .B(n21569), .CI(n21568), .CO(n21566), .S(
        n21571) );
  OAI22D1BWP12T U12463 ( .A1(n21753), .A2(n21868), .B1(n21711), .B2(n21573), 
        .ZN(n21578) );
  ND2D1BWP12T U12464 ( .A1(b[17]), .A2(n21720), .ZN(n21572) );
  OAI211D1BWP12T U12465 ( .A1(n22418), .A2(n21716), .B(a[2]), .C(n21572), .ZN(
        n21577) );
  INVD1BWP12T U12466 ( .I(n21573), .ZN(n21575) );
  OAI22D1BWP12T U12467 ( .A1(n22418), .A2(n21711), .B1(n21750), .B2(n21717), 
        .ZN(n21574) );
  AOI22D1BWP12T U12468 ( .A1(n21575), .A2(n21583), .B1(n21882), .B2(n21574), 
        .ZN(n21576) );
  OAI21D1BWP12T U12469 ( .A1(n21578), .A2(n21577), .B(n21576), .ZN(n22411) );
  FA1D0BWP12T U12470 ( .A(n21581), .B(n21580), .CI(n21579), .CO(n21692), .S(
        n21582) );
  INVD1BWP12T U12471 ( .I(n21582), .ZN(n22473) );
  AOI22D1BWP12T U12472 ( .A1(b[16]), .A2(n21584), .B1(n21583), .B2(n21585), 
        .ZN(n21589) );
  AOI22D1BWP12T U12473 ( .A1(b[15]), .A2(n21720), .B1(n21719), .B2(n21585), 
        .ZN(n21586) );
  AOI32D1BWP12T U12474 ( .A1(b[15]), .A2(n21882), .A3(n21720), .B1(n21586), 
        .B2(a[2]), .ZN(n21588) );
  INVD1BWP12T U12475 ( .I(n21651), .ZN(n23559) );
  NR2D1BWP12T U12476 ( .A1(n21882), .A2(n21868), .ZN(n21738) );
  INVD1BWP12T U12477 ( .I(n21738), .ZN(n21645) );
  OAI22D1BWP12T U12478 ( .A1(n21753), .A2(n23559), .B1(n22547), .B2(n21645), 
        .ZN(n21587) );
  AOI21D1BWP12T U12479 ( .A1(n21589), .A2(n21588), .B(n21587), .ZN(n22472) );
  FA1D0BWP12T U12480 ( .A(n21592), .B(n21591), .CI(n21590), .CO(n21685), .S(
        n21593) );
  ND2D1BWP12T U12481 ( .A1(b[12]), .A2(n21720), .ZN(n21594) );
  OAI22D1BWP12T U12482 ( .A1(n21934), .A2(n23559), .B1(n21882), .B2(n21594), 
        .ZN(n21599) );
  NR2D1BWP12T U12483 ( .A1(n21595), .A2(n21716), .ZN(n21597) );
  OAI211D1BWP12T U12484 ( .A1(n21934), .A2(n21711), .B(n21882), .C(n21594), 
        .ZN(n21596) );
  OAI22D1BWP12T U12485 ( .A1(n21597), .A2(n21596), .B1(n22992), .B2(n21595), 
        .ZN(n21598) );
  AOI211D1BWP12T U12486 ( .A1(b[11]), .A2(n21738), .B(n21599), .C(n21598), 
        .ZN(n22593) );
  FA1D0BWP12T U12487 ( .A(n21602), .B(n21601), .CI(n21600), .CO(n21590), .S(
        n21603) );
  INVD1BWP12T U12488 ( .I(n21603), .ZN(n22592) );
  FA1D0BWP12T U12489 ( .A(n21606), .B(n21605), .CI(n21604), .CO(n21679), .S(
        n21607) );
  INVD1BWP12T U12490 ( .I(n21607), .ZN(n22633) );
  NR2D1BWP12T U12491 ( .A1(n22675), .A2(n21717), .ZN(n21611) );
  OAI22D1BWP12T U12492 ( .A1(n21887), .A2(n21711), .B1(n21716), .B2(n21608), 
        .ZN(n21609) );
  NR2D1BWP12T U12493 ( .A1(n21611), .A2(n21609), .ZN(n21613) );
  AOI22D1BWP12T U12494 ( .A1(b[9]), .A2(n22977), .B1(n21719), .B2(n21773), 
        .ZN(n21610) );
  OAI211D1BWP12T U12495 ( .A1(n21716), .A2(n21887), .B(a[2]), .C(n21610), .ZN(
        n21612) );
  OAI22D1BWP12T U12496 ( .A1(n21613), .A2(a[2]), .B1(n21612), .B2(n21611), 
        .ZN(n22632) );
  FA1D0BWP12T U12497 ( .A(n21616), .B(n21615), .CI(n21614), .CO(n21604), .S(
        n21617) );
  FA1D0BWP12T U12498 ( .A(n21620), .B(n21619), .CI(n21618), .CO(n21614), .S(
        n21621) );
  INVD1BWP12T U12499 ( .I(n21621), .ZN(n22697) );
  NR2D1BWP12T U12500 ( .A1(n22741), .A2(n21717), .ZN(n21627) );
  AOI22D1BWP12T U12501 ( .A1(b[7]), .A2(n22977), .B1(n21719), .B2(n21623), 
        .ZN(n21622) );
  OAI21D1BWP12T U12502 ( .A1(n22699), .A2(n21716), .B(n21622), .ZN(n21626) );
  MOAI22D0BWP12T U12503 ( .A1(n22699), .A2(n21711), .B1(n22978), .B2(n21623), 
        .ZN(n21624) );
  NR2D1BWP12T U12504 ( .A1(n21627), .A2(n21624), .ZN(n21625) );
  OAI32D1BWP12T U12505 ( .A1(n21882), .A2(n21627), .A3(n21626), .B1(n21625), 
        .B2(a[2]), .ZN(n22696) );
  FA1D0BWP12T U12506 ( .A(n21630), .B(n21629), .CI(n21628), .CO(n21618), .S(
        n21631) );
  FA1D0BWP12T U12507 ( .A(n21634), .B(n21633), .CI(n21632), .CO(n21628), .S(
        n21635) );
  INVD1BWP12T U12508 ( .I(n21635), .ZN(n22771) );
  NR2D1BWP12T U12509 ( .A1(n23370), .A2(n21717), .ZN(n21640) );
  OAI22D1BWP12T U12510 ( .A1(n21935), .A2(n21711), .B1(n21716), .B2(n21636), 
        .ZN(n21637) );
  NR2D1BWP12T U12511 ( .A1(n21640), .A2(n21637), .ZN(n21642) );
  AOI22D1BWP12T U12512 ( .A1(b[5]), .A2(n22977), .B1(n21719), .B2(n21638), 
        .ZN(n21639) );
  OAI211D1BWP12T U12513 ( .A1(n21935), .A2(n21716), .B(a[2]), .C(n21639), .ZN(
        n21641) );
  OAI22D1BWP12T U12514 ( .A1(n21642), .A2(a[2]), .B1(n21641), .B2(n21640), 
        .ZN(n22770) );
  MAOI22D0BWP12T U12515 ( .A1(n21644), .A2(n21643), .B1(n21644), .B2(n21643), 
        .ZN(n22801) );
  ND2D1BWP12T U12516 ( .A1(b[4]), .A2(n21720), .ZN(n21646) );
  OAI22D1BWP12T U12517 ( .A1(n22806), .A2(n21645), .B1(n21882), .B2(n21646), 
        .ZN(n21650) );
  NR2D1BWP12T U12518 ( .A1(n21797), .A2(n21716), .ZN(n21648) );
  OAI211D1BWP12T U12519 ( .A1(n21885), .A2(n21711), .B(n21882), .C(n21646), 
        .ZN(n21647) );
  OAI22D1BWP12T U12520 ( .A1(n21648), .A2(n21647), .B1(n22992), .B2(n21797), 
        .ZN(n21649) );
  AOI211D1BWP12T U12521 ( .A1(b[5]), .A2(n21651), .B(n21650), .C(n21649), .ZN(
        n22841) );
  NR2D1BWP12T U12522 ( .A1(n21668), .A2(n21803), .ZN(n21652) );
  MOAI22D0BWP12T U12523 ( .A1(n21653), .A2(n21652), .B1(n21653), .B2(n21652), 
        .ZN(n22840) );
  ND2D1BWP12T U12524 ( .A1(b[0]), .A2(n21670), .ZN(n22896) );
  ND2D1BWP12T U12525 ( .A1(a[0]), .A2(b[0]), .ZN(n23382) );
  NR2D1BWP12T U12526 ( .A1(n22971), .A2(n23382), .ZN(n21940) );
  OAI22D1BWP12T U12527 ( .A1(n21665), .A2(n22485), .B1(n21666), .B2(n22867), 
        .ZN(n21654) );
  AOI211D1BWP12T U12528 ( .A1(b[0]), .A2(n21720), .B(n21940), .C(n21654), .ZN(
        n22995) );
  NR2D1BWP12T U12529 ( .A1(n22995), .A2(n21882), .ZN(n22931) );
  MAOI22D0BWP12T U12530 ( .A1(n21656), .A2(n21655), .B1(n22342), .B2(n21665), 
        .ZN(n21658) );
  ND2D1BWP12T U12531 ( .A1(b[0]), .A2(n21738), .ZN(n21657) );
  OAI211D1BWP12T U12532 ( .A1(a[0]), .A2(n23347), .B(n21658), .C(n21657), .ZN(
        n22930) );
  NR2D1BWP12T U12533 ( .A1(n22931), .A2(n22930), .ZN(n21664) );
  NR2D1BWP12T U12534 ( .A1(n21664), .A2(n21882), .ZN(n21662) );
  NR2D1BWP12T U12535 ( .A1(n22342), .A2(n21717), .ZN(n21661) );
  OAI22D1BWP12T U12536 ( .A1(n21665), .A2(n22806), .B1(n21666), .B2(n21659), 
        .ZN(n21660) );
  AOI211D1BWP12T U12537 ( .A1(n21738), .A2(b[1]), .B(n21661), .C(n21660), .ZN(
        n21663) );
  MAOI22D0BWP12T U12538 ( .A1(n21662), .A2(n21663), .B1(n21662), .B2(n21663), 
        .ZN(n22897) );
  NR2D1BWP12T U12539 ( .A1(n22977), .A2(n21882), .ZN(n22941) );
  INVD1BWP12T U12540 ( .I(n23473), .ZN(n22939) );
  NR2D1BWP12T U12541 ( .A1(n21885), .A2(n21717), .ZN(n21675) );
  OAI22D1BWP12T U12542 ( .A1(n23370), .A2(n21711), .B1(n21716), .B2(n21671), 
        .ZN(n21672) );
  NR2D1BWP12T U12543 ( .A1(n21675), .A2(n21672), .ZN(n21677) );
  AOI22D1BWP12T U12544 ( .A1(b[4]), .A2(n22977), .B1(n21719), .B2(n21673), 
        .ZN(n21674) );
  OAI211D1BWP12T U12545 ( .A1(n23370), .A2(n21716), .B(a[2]), .C(n21674), .ZN(
        n21676) );
  OAI22D1BWP12T U12546 ( .A1(n21677), .A2(a[2]), .B1(n21676), .B2(n21675), 
        .ZN(n22799) );
  FA1D0BWP12T U12547 ( .A(n21681), .B(n21680), .CI(n21679), .CO(n21600), .S(
        n21682) );
  FA1D0BWP12T U12548 ( .A(n21687), .B(n21686), .CI(n21685), .CO(n21579), .S(
        n21688) );
  FA1D0BWP12T U12549 ( .A(n21693), .B(n21692), .CI(n21691), .CO(n21696), .S(
        n21694) );
  FA1D0BWP12T U12550 ( .A(n21697), .B(n21696), .CI(n21695), .CO(n21706), .S(
        n21698) );
  INVD1BWP12T U12551 ( .I(n21698), .ZN(n22409) );
  NR2D1BWP12T U12552 ( .A1(n22418), .A2(n21717), .ZN(n21702) );
  OAI22D1BWP12T U12553 ( .A1(n21944), .A2(n21711), .B1(n21716), .B2(n21700), 
        .ZN(n21699) );
  NR2D1BWP12T U12554 ( .A1(n21702), .A2(n21699), .ZN(n21704) );
  MAOI22D0BWP12T U12555 ( .A1(b[17]), .A2(n22977), .B1(n21711), .B2(n21700), 
        .ZN(n21701) );
  OAI211D1BWP12T U12556 ( .A1(n21944), .A2(n21716), .B(a[2]), .C(n21701), .ZN(
        n21703) );
  OAI22D1BWP12T U12557 ( .A1(n21704), .A2(a[2]), .B1(n21703), .B2(n21702), 
        .ZN(n22372) );
  FA1D0BWP12T U12558 ( .A(n21707), .B(n21706), .CI(n21705), .CO(n21569), .S(
        n21708) );
  INVD1BWP12T U12559 ( .I(n21708), .ZN(n22371) );
  NR2D1BWP12T U12560 ( .A1(n23498), .A2(n21717), .ZN(n21713) );
  OAI22D1BWP12T U12561 ( .A1(n22293), .A2(n21711), .B1(n21716), .B2(n21710), 
        .ZN(n21709) );
  NR2D1BWP12T U12562 ( .A1(n21713), .A2(n21709), .ZN(n21715) );
  MAOI22D0BWP12T U12563 ( .A1(b[21]), .A2(n22978), .B1(n21711), .B2(n21710), 
        .ZN(n21712) );
  OAI211D1BWP12T U12564 ( .A1(n21944), .A2(n21868), .B(a[2]), .C(n21712), .ZN(
        n21714) );
  OAI22D1BWP12T U12565 ( .A1(n21715), .A2(a[2]), .B1(n21714), .B2(n21713), 
        .ZN(n22314) );
  OAI22D1BWP12T U12566 ( .A1(n21886), .A2(n21717), .B1(n21716), .B2(n21759), 
        .ZN(n21718) );
  AOI211D1BWP12T U12567 ( .A1(b[23]), .A2(n21719), .B(a[2]), .C(n21718), .ZN(
        n21723) );
  AOI22D1BWP12T U12568 ( .A1(b[23]), .A2(n22978), .B1(b[22]), .B2(n21720), 
        .ZN(n21721) );
  OAI22D1BWP12T U12569 ( .A1(n21721), .A2(n21882), .B1(n22992), .B2(n21759), 
        .ZN(n21722) );
  AOI211D1BWP12T U12570 ( .A1(n21738), .A2(b[21]), .B(n21723), .C(n21722), 
        .ZN(n22229) );
  NR2D1BWP12T U12571 ( .A1(n22150), .A2(n21724), .ZN(n21729) );
  OAI22D1BWP12T U12572 ( .A1(n22088), .A2(n21727), .B1(n21726), .B2(n21725), 
        .ZN(n21728) );
  AOI211D1BWP12T U12573 ( .A1(b[24]), .A2(n21730), .B(n21729), .C(n21728), 
        .ZN(n21865) );
  NR2D1BWP12T U12574 ( .A1(n23375), .A2(n21731), .ZN(n21736) );
  OAI22D1BWP12T U12575 ( .A1(n21734), .A2(n22032), .B1(n21733), .B2(n21732), 
        .ZN(n21735) );
  AOI211D1BWP12T U12576 ( .A1(b[28]), .A2(n21737), .B(n21736), .C(n21735), 
        .ZN(n21863) );
  AOI22D1BWP12T U12577 ( .A1(b[31]), .A2(n21868), .B1(b[30]), .B2(n21738), 
        .ZN(n21741) );
  AOI21D1BWP12T U12578 ( .A1(n21741), .A2(n21740), .B(n21739), .ZN(n21861) );
  NR2D1BWP12T U12579 ( .A1(n21944), .A2(n21742), .ZN(n21747) );
  OAI22D1BWP12T U12580 ( .A1(n22418), .A2(n21745), .B1(n21744), .B2(n21743), 
        .ZN(n21746) );
  AOI211D1BWP12T U12581 ( .A1(b[20]), .A2(n21748), .B(n21747), .C(n21746), 
        .ZN(n21859) );
  NR2D1BWP12T U12582 ( .A1(n21750), .A2(n21749), .ZN(n21755) );
  OAI22D1BWP12T U12583 ( .A1(n21753), .A2(n22477), .B1(n21752), .B2(n21751), 
        .ZN(n21754) );
  AOI211D1BWP12T U12584 ( .A1(b[15]), .A2(n21756), .B(n21755), .C(n21754), 
        .ZN(n21857) );
  NR2D1BWP12T U12585 ( .A1(n21886), .A2(n21757), .ZN(n21762) );
  OAI22D1BWP12T U12586 ( .A1(n21932), .A2(n21760), .B1(n21759), .B2(n21758), 
        .ZN(n21761) );
  AOI211D1BWP12T U12587 ( .A1(b[21]), .A2(n21763), .B(n21762), .C(n21761), 
        .ZN(n21855) );
  NR2D1BWP12T U12588 ( .A1(n22547), .A2(n21764), .ZN(n21769) );
  OAI22D1BWP12T U12589 ( .A1(n21934), .A2(n21767), .B1(n21766), .B2(n21765), 
        .ZN(n21768) );
  AOI211D1BWP12T U12590 ( .A1(n21770), .A2(b[12]), .B(n21769), .C(n21768), 
        .ZN(n21853) );
  AOI22D1BWP12T U12591 ( .A1(b[9]), .A2(n21772), .B1(b[11]), .B2(n21771), .ZN(
        n21776) );
  ND2D1BWP12T U12592 ( .A1(n21774), .A2(n21773), .ZN(n21775) );
  OAI211D1BWP12T U12593 ( .A1(n22675), .A2(n21777), .B(n21776), .C(n21775), 
        .ZN(n21786) );
  AOI22D1BWP12T U12594 ( .A1(b[8]), .A2(n21779), .B1(b[7]), .B2(n21778), .ZN(
        n21783) );
  ND2D1BWP12T U12595 ( .A1(n21781), .A2(n21780), .ZN(n21782) );
  OAI211D1BWP12T U12596 ( .A1(n23370), .A2(n21784), .B(n21783), .C(n21782), 
        .ZN(n21785) );
  MAOI22D0BWP12T U12597 ( .A1(n21786), .A2(n21785), .B1(n21786), .B2(n21785), 
        .ZN(n21851) );
  NR2D1BWP12T U12598 ( .A1(n21787), .A2(n23642), .ZN(n21795) );
  MAOI22D0BWP12T U12599 ( .A1(b[2]), .A2(n21789), .B1(n22485), .B2(n21788), 
        .ZN(n21793) );
  AOI22D1BWP12T U12600 ( .A1(a[8]), .A2(n22642), .B1(a[11]), .B2(n21966), .ZN(
        n21791) );
  AOI22D1BWP12T U12601 ( .A1(a[23]), .A2(a[20]), .B1(n22404), .B2(n22267), 
        .ZN(n21790) );
  MAOI22D0BWP12T U12602 ( .A1(n21791), .A2(n21790), .B1(n21791), .B2(n21790), 
        .ZN(n21792) );
  MAOI22D0BWP12T U12603 ( .A1(n21793), .A2(n21792), .B1(n21793), .B2(n21792), 
        .ZN(n21794) );
  MAOI22D0BWP12T U12604 ( .A1(n21795), .A2(n21794), .B1(n21795), .B2(n21794), 
        .ZN(n21849) );
  NR2D1BWP12T U12605 ( .A1(n21885), .A2(n21796), .ZN(n21801) );
  OAI22D1BWP12T U12606 ( .A1(n23017), .A2(n21799), .B1(n21798), .B2(n21797), 
        .ZN(n21800) );
  AOI211D1BWP12T U12607 ( .A1(b[3]), .A2(n21802), .B(n21801), .C(n21800), .ZN(
        n21847) );
  AOI22D1BWP12T U12608 ( .A1(a[5]), .A2(a[2]), .B1(n21882), .B2(n21803), .ZN(
        n21805) );
  ND2D1BWP12T U12609 ( .A1(n23376), .A2(n22087), .ZN(n23543) );
  OAI21D1BWP12T U12610 ( .A1(n22087), .A2(n23376), .B(n23543), .ZN(n21804) );
  MAOI22D0BWP12T U12611 ( .A1(n21805), .A2(n21804), .B1(n21805), .B2(n21804), 
        .ZN(n21845) );
  FA1D0BWP12T U12612 ( .A(n21808), .B(n21807), .CI(n21806), .CO(n21811), .S(
        n23657) );
  MOAI22D0BWP12T U12613 ( .A1(n21811), .A2(n21810), .B1(n21811), .B2(n21810), 
        .ZN(n21812) );
  MAOI22D0BWP12T U12614 ( .A1(n21813), .A2(n21812), .B1(n21813), .B2(n21812), 
        .ZN(n21843) );
  FA1D0BWP12T U12615 ( .A(n21817), .B(n21816), .CI(n21815), .CO(n21818), .S(
        n21232) );
  MAOI22D0BWP12T U12616 ( .A1(n21819), .A2(n21818), .B1(n21819), .B2(n21818), 
        .ZN(n21841) );
  FA1D0BWP12T U12617 ( .A(n21823), .B(n21822), .CI(n21821), .CO(n21824), .S(
        n21248) );
  MAOI22D0BWP12T U12618 ( .A1(n21825), .A2(n21824), .B1(n21825), .B2(n21824), 
        .ZN(n21839) );
  FA1D0BWP12T U12619 ( .A(n21828), .B(n21827), .CI(n21826), .CO(n21831), .S(
        n21823) );
  MAOI22D0BWP12T U12620 ( .A1(n21831), .A2(n21830), .B1(n21831), .B2(n21830), 
        .ZN(n21837) );
  MOAI22D0BWP12T U12621 ( .A1(n21835), .A2(n21834), .B1(n21835), .B2(n21834), 
        .ZN(n21836) );
  MAOI22D0BWP12T U12622 ( .A1(n21837), .A2(n21836), .B1(n21837), .B2(n21836), 
        .ZN(n21838) );
  MAOI22D0BWP12T U12623 ( .A1(n21839), .A2(n21838), .B1(n21839), .B2(n21838), 
        .ZN(n21840) );
  MAOI22D0BWP12T U12624 ( .A1(n21841), .A2(n21840), .B1(n21841), .B2(n21840), 
        .ZN(n21842) );
  MAOI22D0BWP12T U12625 ( .A1(n21843), .A2(n21842), .B1(n21843), .B2(n21842), 
        .ZN(n21844) );
  MAOI22D0BWP12T U12626 ( .A1(n21845), .A2(n21844), .B1(n21845), .B2(n21844), 
        .ZN(n21846) );
  MAOI22D0BWP12T U12627 ( .A1(n21847), .A2(n21846), .B1(n21847), .B2(n21846), 
        .ZN(n21848) );
  MAOI22D0BWP12T U12628 ( .A1(n21849), .A2(n21848), .B1(n21849), .B2(n21848), 
        .ZN(n21850) );
  MAOI22D0BWP12T U12629 ( .A1(n21851), .A2(n21850), .B1(n21851), .B2(n21850), 
        .ZN(n21852) );
  MAOI22D0BWP12T U12630 ( .A1(n21853), .A2(n21852), .B1(n21853), .B2(n21852), 
        .ZN(n21854) );
  MAOI22D0BWP12T U12631 ( .A1(n21855), .A2(n21854), .B1(n21855), .B2(n21854), 
        .ZN(n21856) );
  MAOI22D0BWP12T U12632 ( .A1(n21857), .A2(n21856), .B1(n21857), .B2(n21856), 
        .ZN(n21858) );
  MAOI22D0BWP12T U12633 ( .A1(n21859), .A2(n21858), .B1(n21859), .B2(n21858), 
        .ZN(n21860) );
  MAOI22D0BWP12T U12634 ( .A1(n21861), .A2(n21860), .B1(n21861), .B2(n21860), 
        .ZN(n21862) );
  MAOI22D0BWP12T U12635 ( .A1(n21863), .A2(n21862), .B1(n21863), .B2(n21862), 
        .ZN(n21864) );
  MAOI22D0BWP12T U12636 ( .A1(n21865), .A2(n21864), .B1(n21865), .B2(n21864), 
        .ZN(n21867) );
  INVD1BWP12T U12637 ( .I(n23658), .ZN(n23031) );
  NR2D1BWP12T U12638 ( .A1(n23031), .A2(n21867), .ZN(n23059) );
  INVD1BWP12T U12639 ( .I(n23657), .ZN(n21866) );
  AOI32D1BWP12T U12640 ( .A1(n23658), .A2(n23657), .A3(n21867), .B1(n23059), 
        .B2(n21866), .ZN(n21871) );
  INVD1BWP12T U12641 ( .I(n21896), .ZN(n22012) );
  INVD1BWP12T U12642 ( .I(n23046), .ZN(n21902) );
  IND2D1BWP12T U12643 ( .A1(n22339), .B1(n22404), .ZN(n21898) );
  ND2D1BWP12T U12644 ( .A1(n22776), .A2(n22775), .ZN(n22728) );
  NR2D1BWP12T U12645 ( .A1(n22728), .A2(a[8]), .ZN(n23049) );
  NR2D1BWP12T U12646 ( .A1(n23021), .A2(n21918), .ZN(n23033) );
  INVD1BWP12T U12647 ( .I(n23033), .ZN(n23054) );
  NR2D1BWP12T U12648 ( .A1(a[2]), .A2(n21868), .ZN(n22942) );
  ND2D1BWP12T U12649 ( .A1(n22942), .A2(n22911), .ZN(n22910) );
  NR2D1BWP12T U12650 ( .A1(n23054), .A2(n22910), .ZN(n22874) );
  ND2D1BWP12T U12651 ( .A1(n22874), .A2(n22873), .ZN(n22856) );
  INVD1BWP12T U12652 ( .I(n22856), .ZN(n22767) );
  ND2D1BWP12T U12653 ( .A1(n23049), .A2(n22767), .ZN(n22701) );
  INVD1BWP12T U12654 ( .I(n22701), .ZN(n22670) );
  NR2D1BWP12T U12655 ( .A1(n22634), .A2(n21869), .ZN(n22587) );
  ND2D1BWP12T U12656 ( .A1(n22587), .A2(n22588), .ZN(n22490) );
  NR2D1BWP12T U12657 ( .A1(a[14]), .A2(n22490), .ZN(n21870) );
  ND2D1BWP12T U12658 ( .A1(n22670), .A2(n21870), .ZN(n22510) );
  NR2D1BWP12T U12659 ( .A1(n21897), .A2(n22510), .ZN(n22434) );
  ND2D1BWP12T U12660 ( .A1(n22434), .A2(n22441), .ZN(n22417) );
  NR2D1BWP12T U12661 ( .A1(n21898), .A2(n22417), .ZN(n22328) );
  ND2D1BWP12T U12662 ( .A1(n21902), .A2(n22328), .ZN(n22266) );
  NR2D1BWP12T U12663 ( .A1(n23047), .A2(n22266), .ZN(n22157) );
  ND2D1BWP12T U12664 ( .A1(n22012), .A2(n22157), .ZN(n22031) );
  NR2D1BWP12T U12665 ( .A1(n21895), .A2(n22031), .ZN(n21978) );
  ND3D1BWP12T U12666 ( .A1(a[31]), .A2(n23050), .A3(n21978), .ZN(n23675) );
  OAI211D1BWP12T U12667 ( .A1(n21873), .A2(n21872), .B(n21871), .C(n23675), 
        .ZN(n21874) );
  AO21D1BWP12T U12668 ( .A1(n21875), .A2(n23058), .B(n21874), .Z(v) );
  NR2D1BWP12T U12669 ( .A1(b[30]), .A2(a[30]), .ZN(n23541) );
  INVD1BWP12T U12670 ( .I(n23541), .ZN(n21925) );
  ND2D1BWP12T U12671 ( .A1(b[30]), .A2(a[30]), .ZN(n23367) );
  ND2D1BWP12T U12672 ( .A1(n21925), .A2(n23367), .ZN(n23044) );
  INVD1BWP12T U12673 ( .I(n23044), .ZN(n21938) );
  NR2D1BWP12T U12674 ( .A1(n21909), .A2(n21876), .ZN(n21877) );
  MAOI22D0BWP12T U12675 ( .A1(n21938), .A2(n21877), .B1(n21938), .B2(n21877), 
        .ZN(n23160) );
  ND2D1BWP12T U12676 ( .A1(n22342), .A2(n22757), .ZN(n23663) );
  INR2D1BWP12T U12677 ( .A1(n23663), .B1(n22806), .ZN(n22219) );
  NR2D1BWP12T U12678 ( .A1(n23663), .A2(b[3]), .ZN(n21881) );
  OR2XD1BWP12T U12679 ( .A1(n21881), .A2(n23017), .Z(n22504) );
  NR2D1BWP12T U12680 ( .A1(n22219), .A2(n22504), .ZN(n22488) );
  INVD1BWP12T U12681 ( .I(n22757), .ZN(n22640) );
  ND2D1BWP12T U12682 ( .A1(b[2]), .A2(n22640), .ZN(n22365) );
  NR2D1BWP12T U12683 ( .A1(n22867), .A2(n22365), .ZN(n22227) );
  INVD1BWP12T U12684 ( .I(b[0]), .ZN(n22605) );
  AOI22D1BWP12T U12685 ( .A1(b[0]), .A2(n22383), .B1(n22404), .B2(n22605), 
        .ZN(n22178) );
  INVD1BWP12T U12686 ( .I(n22178), .ZN(n22105) );
  AOI22D1BWP12T U12687 ( .A1(b[0]), .A2(a[21]), .B1(a[22]), .B2(n22605), .ZN(
        n21998) );
  INVD1BWP12T U12688 ( .I(n21998), .ZN(n22346) );
  ND2D1BWP12T U12689 ( .A1(n23663), .A2(n22365), .ZN(n22099) );
  INVD1BWP12T U12690 ( .I(n22099), .ZN(n22226) );
  NR2D1BWP12T U12691 ( .A1(n22864), .A2(n22226), .ZN(n22447) );
  INVD1BWP12T U12692 ( .I(n22447), .ZN(n22223) );
  NR2D1BWP12T U12693 ( .A1(n22346), .A2(n22223), .ZN(n21880) );
  AOI22D1BWP12T U12694 ( .A1(b[0]), .A2(a[15]), .B1(a[16]), .B2(n22605), .ZN(
        n22533) );
  ND2D1BWP12T U12695 ( .A1(n22864), .A2(n22533), .ZN(n21878) );
  NR2D1BWP12T U12696 ( .A1(n22864), .A2(n22099), .ZN(n22174) );
  INVD1BWP12T U12697 ( .I(n22174), .ZN(n22224) );
  OAI22D1BWP12T U12698 ( .A1(b[2]), .A2(n21878), .B1(n22224), .B2(n22196), 
        .ZN(n21879) );
  AOI211D1BWP12T U12699 ( .A1(n22227), .A2(n22105), .B(n21880), .C(n21879), 
        .ZN(n23458) );
  AOI22D1BWP12T U12700 ( .A1(b[0]), .A2(a[29]), .B1(a[30]), .B2(n22605), .ZN(
        n22011) );
  ND2D1BWP12T U12701 ( .A1(b[2]), .A2(n22842), .ZN(n22692) );
  INVD1BWP12T U12702 ( .I(n22692), .ZN(n22137) );
  ND2D1BWP12T U12703 ( .A1(b[4]), .A2(b[3]), .ZN(n23265) );
  INVD1BWP12T U12704 ( .I(n23265), .ZN(n21973) );
  ND2D1BWP12T U12705 ( .A1(n22137), .A2(n21973), .ZN(n22988) );
  ND2D1BWP12T U12706 ( .A1(n23663), .A2(n21973), .ZN(n22400) );
  INVD1BWP12T U12707 ( .I(n22400), .ZN(n22766) );
  AN2D1BWP12T U12708 ( .A1(n22365), .A2(n22766), .Z(n23445) );
  AOI22D1BWP12T U12709 ( .A1(b[0]), .A2(n22267), .B1(n23560), .B2(n22605), 
        .ZN(n22268) );
  INVD1BWP12T U12710 ( .I(n22268), .ZN(n21993) );
  ND2D1BWP12T U12711 ( .A1(n22009), .A2(n22087), .ZN(n22194) );
  INVD1BWP12T U12712 ( .I(n22194), .ZN(n22092) );
  NR2D1BWP12T U12713 ( .A1(a[25]), .A2(n22009), .ZN(n22271) );
  NR2D1BWP12T U12714 ( .A1(n22092), .A2(n22271), .ZN(n21996) );
  INVD1BWP12T U12715 ( .I(n21996), .ZN(n21997) );
  OAI22D1BWP12T U12716 ( .A1(n22867), .A2(n21993), .B1(n21997), .B2(n22864), 
        .ZN(n22102) );
  MOAI22D0BWP12T U12717 ( .A1(n22011), .A2(n22988), .B1(n23445), .B2(n22102), 
        .ZN(n21884) );
  NR2D1BWP12T U12718 ( .A1(n21881), .A2(n22219), .ZN(n22506) );
  AOI22D1BWP12T U12719 ( .A1(b[0]), .A2(a[5]), .B1(a[6]), .B2(n22009), .ZN(
        n22865) );
  INVD1BWP12T U12720 ( .I(n22865), .ZN(n22199) );
  AOI22D1BWP12T U12721 ( .A1(b[0]), .A2(a[3]), .B1(a[4]), .B2(n22605), .ZN(
        n22100) );
  INVD1BWP12T U12722 ( .I(n22100), .ZN(n22173) );
  INVD1BWP12T U12723 ( .I(n22227), .ZN(n22168) );
  AOI22D1BWP12T U12724 ( .A1(b[0]), .A2(n23011), .B1(n21882), .B2(n22605), 
        .ZN(n22001) );
  INVD1BWP12T U12725 ( .I(n22001), .ZN(n22177) );
  MOAI22D0BWP12T U12726 ( .A1(n22864), .A2(n22177), .B1(a[0]), .B2(n22843), 
        .ZN(n22933) );
  OAI222D1BWP12T U12727 ( .A1(n22199), .A2(n22223), .B1(n22173), .B2(n22168), 
        .C1(n22099), .C2(n22933), .ZN(n22288) );
  INVD1BWP12T U12728 ( .I(n22288), .ZN(n23457) );
  OAI22D1BWP12T U12729 ( .A1(n22605), .A2(a[9]), .B1(a[10]), .B2(b[0]), .ZN(
        n22721) );
  AOI22D1BWP12T U12730 ( .A1(b[0]), .A2(a[13]), .B1(a[14]), .B2(n22605), .ZN(
        n22200) );
  AOI22D1BWP12T U12731 ( .A1(b[0]), .A2(n22642), .B1(n22689), .B2(n22009), 
        .ZN(n22081) );
  ND2D1BWP12T U12732 ( .A1(b[0]), .A2(a[7]), .ZN(n22866) );
  ND2D1BWP12T U12733 ( .A1(n22009), .A2(a[8]), .ZN(n22723) );
  ND2D1BWP12T U12734 ( .A1(n22866), .A2(n22723), .ZN(n22198) );
  ND2D1BWP12T U12735 ( .A1(n22864), .A2(n22365), .ZN(n22220) );
  INVD1BWP12T U12736 ( .I(n22506), .ZN(n22505) );
  AOI22D1BWP12T U12737 ( .A1(n22506), .A2(n23457), .B1(n23437), .B2(n22505), 
        .ZN(n22542) );
  NR2D1BWP12T U12738 ( .A1(b[4]), .A2(b[3]), .ZN(n23258) );
  INVD1BWP12T U12739 ( .I(n23258), .ZN(n22691) );
  NR2D1BWP12T U12740 ( .A1(b[2]), .A2(n22691), .ZN(n22663) );
  ND2D1BWP12T U12741 ( .A1(n22757), .A2(n22663), .ZN(n23544) );
  ND2D1BWP12T U12742 ( .A1(n22504), .A2(n23544), .ZN(n23443) );
  AOI22D1BWP12T U12743 ( .A1(b[0]), .A2(a[27]), .B1(a[28]), .B2(n22605), .ZN(
        n22091) );
  IND2D1BWP12T U12744 ( .A1(n22365), .B1(n21973), .ZN(n22926) );
  NR2D1BWP12T U12745 ( .A1(n22926), .A2(n22842), .ZN(n23440) );
  INVD1BWP12T U12746 ( .I(n23440), .ZN(n22172) );
  OAI22D1BWP12T U12747 ( .A1(n22542), .A2(n23443), .B1(n22091), .B2(n22172), 
        .ZN(n21883) );
  AOI211D1BWP12T U12748 ( .A1(n22488), .A2(n23458), .B(n21884), .C(n21883), 
        .ZN(n23419) );
  ND2D1BWP12T U12749 ( .A1(op[0]), .A2(op[1]), .ZN(n21939) );
  INVD1BWP12T U12750 ( .I(n21931), .ZN(n22018) );
  NR2D1BWP12T U12751 ( .A1(n21939), .A2(n22018), .ZN(n23667) );
  INVD1BWP12T U12752 ( .I(n23667), .ZN(n22987) );
  ND4D1BWP12T U12753 ( .A1(n22699), .A2(n22741), .A3(n21935), .A4(n23370), 
        .ZN(n21893) );
  ND4D1BWP12T U12754 ( .A1(n22032), .A2(n21932), .A3(n23498), .A4(n21885), 
        .ZN(n21892) );
  ND4D1BWP12T U12755 ( .A1(n23375), .A2(n22150), .A3(n21886), .A4(n22293), 
        .ZN(n21891) );
  NR2D1BWP12T U12756 ( .A1(b[15]), .A2(b[14]), .ZN(n21889) );
  NR4D0BWP12T U12757 ( .A1(b[19]), .A2(b[18]), .A3(b[17]), .A4(b[12]), .ZN(
        n21888) );
  ND4D1BWP12T U12758 ( .A1(n21889), .A2(n21888), .A3(n22675), .A4(n21887), 
        .ZN(n21890) );
  NR4D0BWP12T U12759 ( .A1(n21893), .A2(n21892), .A3(n21891), .A4(n21890), 
        .ZN(n23538) );
  NR2D1BWP12T U12760 ( .A1(b[26]), .A2(b[16]), .ZN(n23539) );
  NR4D0BWP12T U12761 ( .A1(b[31]), .A2(b[30]), .A3(b[24]), .A4(b[13]), .ZN(
        n21894) );
  ND4D1BWP12T U12762 ( .A1(n23538), .A2(n23539), .A3(n21894), .A4(n23490), 
        .ZN(n23294) );
  NR2D1BWP12T U12763 ( .A1(op[0]), .A2(op[1]), .ZN(n22019) );
  ND2D1BWP12T U12764 ( .A1(n21931), .A2(n22019), .ZN(n22706) );
  NR2D1BWP12T U12765 ( .A1(n23294), .A2(n22706), .ZN(n22925) );
  INVD1BWP12T U12766 ( .I(n21939), .ZN(n21900) );
  NR2D1BWP12T U12767 ( .A1(op[2]), .A2(op[3]), .ZN(n21919) );
  ND2D1BWP12T U12768 ( .A1(n21900), .A2(n21919), .ZN(n23589) );
  OAI21D1BWP12T U12769 ( .A1(n23294), .A2(n23589), .B(n22987), .ZN(n22964) );
  NR2D1BWP12T U12770 ( .A1(n22925), .A2(n22964), .ZN(n23041) );
  NR2D1BWP12T U12771 ( .A1(b[4]), .A2(n23041), .ZN(n22489) );
  ND2D1BWP12T U12772 ( .A1(n22342), .A2(n22485), .ZN(n22274) );
  INVD1BWP12T U12773 ( .I(n22274), .ZN(n22607) );
  ND2D1BWP12T U12774 ( .A1(n22806), .A2(n22607), .ZN(n23012) );
  AOI22D1BWP12T U12775 ( .A1(b[0]), .A2(a[31]), .B1(a[30]), .B2(n22605), .ZN(
        n22273) );
  NR2D1BWP12T U12776 ( .A1(n23012), .A2(n22273), .ZN(n23223) );
  NR2D1BWP12T U12777 ( .A1(n21896), .A2(n21895), .ZN(n23051) );
  OR4XD1BWP12T U12778 ( .A1(a[17]), .A2(a[14]), .A3(n21897), .A4(n22490), .Z(
        n22367) );
  NR2D1BWP12T U12779 ( .A1(n22367), .A2(n21898), .ZN(n23052) );
  INVD1BWP12T U12780 ( .I(n23052), .ZN(n23572) );
  INVD1BWP12T U12781 ( .I(n21899), .ZN(n21922) );
  ND2D1BWP12T U12782 ( .A1(n21900), .A2(n21922), .ZN(n23558) );
  INVD1BWP12T U12783 ( .I(n23558), .ZN(n22905) );
  ND2D1BWP12T U12784 ( .A1(n22942), .A2(n21901), .ZN(n23048) );
  NR2D1BWP12T U12785 ( .A1(n22905), .A2(n23048), .ZN(n22857) );
  ND2D1BWP12T U12786 ( .A1(n23049), .A2(n22857), .ZN(n22585) );
  NR2D1BWP12T U12787 ( .A1(n23572), .A2(n22585), .ZN(n22344) );
  ND2D1BWP12T U12788 ( .A1(n21902), .A2(n22344), .ZN(n22228) );
  ND2D1BWP12T U12789 ( .A1(n23054), .A2(n23558), .ZN(n22586) );
  OAI21D1BWP12T U12790 ( .A1(n23047), .A2(n22228), .B(n22586), .ZN(n22209) );
  INVD1BWP12T U12791 ( .I(n22586), .ZN(n22858) );
  AOI31D1BWP12T U12792 ( .A1(n23051), .A2(n23376), .A3(n22209), .B(n22858), 
        .ZN(n23641) );
  AOI22D1BWP12T U12793 ( .A1(n22489), .A2(n23223), .B1(n21903), .B2(n23641), 
        .ZN(n21928) );
  NR2D1BWP12T U12794 ( .A1(b[4]), .A2(n23294), .ZN(n23409) );
  INVD1BWP12T U12795 ( .I(n22706), .ZN(n23585) );
  ND2D1BWP12T U12796 ( .A1(a[31]), .A2(n23585), .ZN(n23646) );
  NR2D1BWP12T U12797 ( .A1(n23409), .A2(n23646), .ZN(n22513) );
  ND2D1BWP12T U12798 ( .A1(a[31]), .A2(n23012), .ZN(n22576) );
  INVD1BWP12T U12799 ( .I(n22925), .ZN(n22986) );
  NR2D1BWP12T U12800 ( .A1(n22576), .A2(n22986), .ZN(n22539) );
  NR2D1BWP12T U12801 ( .A1(n22513), .A2(n22539), .ZN(n21982) );
  FA1D0BWP12T U12802 ( .A(n21906), .B(n21905), .CI(n21904), .CO(n21806), .S(
        n23325) );
  OAI21D1BWP12T U12803 ( .A1(n21909), .A2(n21908), .B(n21907), .ZN(n21910) );
  MAOI22D0BWP12T U12804 ( .A1(n23044), .A2(n21910), .B1(n23044), .B2(n21910), 
        .ZN(n23597) );
  MAOI22D0BWP12T U12805 ( .A1(n23658), .A2(n23325), .B1(n23597), .B2(n23653), 
        .ZN(n21927) );
  ND2D1BWP12T U12806 ( .A1(n21920), .A2(n21919), .ZN(n23298) );
  NR2D1BWP12T U12807 ( .A1(n23294), .A2(n23298), .ZN(n23644) );
  ND2D1BWP12T U12808 ( .A1(b[4]), .A2(n22806), .ZN(n22665) );
  INVD1BWP12T U12809 ( .I(n22665), .ZN(n23263) );
  NR2D1BWP12T U12810 ( .A1(b[1]), .A2(n22342), .ZN(n23259) );
  AOI22D1BWP12T U12811 ( .A1(n22607), .A2(n22200), .B1(n22721), .B2(n23259), 
        .ZN(n21912) );
  INVD1BWP12T U12812 ( .I(n22245), .ZN(n22606) );
  INVD1BWP12T U12813 ( .I(n22081), .ZN(n22201) );
  ND2D1BWP12T U12814 ( .A1(n22606), .A2(n22201), .ZN(n21911) );
  OAI211D1BWP12T U12815 ( .A1(n22198), .A2(n22244), .B(n21912), .C(n21911), 
        .ZN(n23245) );
  NR2D1BWP12T U12816 ( .A1(n22342), .A2(n22691), .ZN(n22662) );
  AOI22D1BWP12T U12817 ( .A1(n22662), .A2(n21993), .B1(n22663), .B2(n22091), 
        .ZN(n22005) );
  AOI22D1BWP12T U12818 ( .A1(n22662), .A2(n21997), .B1(n22663), .B2(n22011), 
        .ZN(n21913) );
  AOI22D1BWP12T U12819 ( .A1(b[1]), .A2(n22005), .B1(n21913), .B2(n22485), 
        .ZN(n21917) );
  AOI22D1BWP12T U12820 ( .A1(a[0]), .A2(n22843), .B1(n22485), .B2(n22001), 
        .ZN(n22077) );
  OAI222D1BWP12T U12821 ( .A1(n22274), .A2(n22865), .B1(n22245), .B2(n22100), 
        .C1(n22342), .C2(n22077), .ZN(n23271) );
  INVD1BWP12T U12822 ( .I(n22196), .ZN(n22096) );
  AOI22D1BWP12T U12823 ( .A1(n22606), .A2(n22105), .B1(n23259), .B2(n22096), 
        .ZN(n21915) );
  AOI22D1BWP12T U12824 ( .A1(n22607), .A2(n21998), .B1(n22533), .B2(n22951), 
        .ZN(n21914) );
  ND2D1BWP12T U12825 ( .A1(n21915), .A2(n21914), .ZN(n22277) );
  NR2D1BWP12T U12826 ( .A1(b[4]), .A2(n22806), .ZN(n23270) );
  MOAI22D0BWP12T U12827 ( .A1(n23265), .A2(n23271), .B1(n22277), .B2(n23270), 
        .ZN(n21916) );
  AOI211D1BWP12T U12828 ( .A1(n23263), .A2(n23245), .B(n21917), .C(n21916), 
        .ZN(n23285) );
  ND2D1BWP12T U12829 ( .A1(n22019), .A2(n22812), .ZN(n23372) );
  INVD1BWP12T U12830 ( .I(n21918), .ZN(n21930) );
  ND2D1BWP12T U12831 ( .A1(n21930), .A2(n21919), .ZN(n23499) );
  INVD1BWP12T U12832 ( .I(n23499), .ZN(n23650) );
  ND2D1BWP12T U12833 ( .A1(n21920), .A2(n21922), .ZN(n23022) );
  INVD1BWP12T U12834 ( .I(n23022), .ZN(n23509) );
  AOI22D1BWP12T U12835 ( .A1(n23650), .A2(n23367), .B1(n23509), .B2(n21921), 
        .ZN(n21923) );
  ND2D1BWP12T U12836 ( .A1(n22019), .A2(n21922), .ZN(n23645) );
  OAI211D1BWP12T U12837 ( .A1(n23372), .A2(n23367), .B(n21923), .C(n23645), 
        .ZN(n21924) );
  AOI22D1BWP12T U12838 ( .A1(n23644), .A2(n23285), .B1(n21925), .B2(n21924), 
        .ZN(n21926) );
  ND4D1BWP12T U12839 ( .A1(n21928), .A2(n21982), .A3(n21927), .A4(n21926), 
        .ZN(n21929) );
  AOI31D1BWP12T U12840 ( .A1(a[30]), .A2(n21978), .A3(n23376), .B(n21929), 
        .ZN(n21949) );
  AN2D1BWP12T U12841 ( .A1(n21931), .A2(n21930), .Z(n23027) );
  NR2D1BWP12T U12842 ( .A1(b[29]), .A2(a[29]), .ZN(n21947) );
  NR2D1BWP12T U12843 ( .A1(b[28]), .A2(a[28]), .ZN(n23540) );
  NR2D1BWP12T U12844 ( .A1(b[27]), .A2(a[27]), .ZN(n23170) );
  NR2D1BWP12T U12845 ( .A1(b[25]), .A2(a[25]), .ZN(n23174) );
  ND2D1BWP12T U12846 ( .A1(n21932), .A2(n22267), .ZN(n23093) );
  NR2D1BWP12T U12847 ( .A1(n21932), .A2(n22267), .ZN(n23352) );
  INR2D1BWP12T U12848 ( .A1(n23093), .B1(n23352), .ZN(n23065) );
  INVD1BWP12T U12849 ( .I(n23066), .ZN(n21945) );
  INVD1BWP12T U12850 ( .I(n22385), .ZN(n23099) );
  INVD1BWP12T U12851 ( .I(n23083), .ZN(n22465) );
  ND2D1BWP12T U12852 ( .A1(n21933), .A2(n22547), .ZN(n22549) );
  ND2D1BWP12T U12853 ( .A1(a[14]), .A2(b[14]), .ZN(n23341) );
  ND2D1BWP12T U12854 ( .A1(n22549), .A2(n23341), .ZN(n23178) );
  INVD1BWP12T U12855 ( .I(n23178), .ZN(n22560) );
  ND2D1BWP12T U12856 ( .A1(n21934), .A2(n22588), .ZN(n23179) );
  OAI21D1BWP12T U12857 ( .A1(n22588), .A2(n21934), .B(n23179), .ZN(n22584) );
  INVD1BWP12T U12858 ( .I(n22584), .ZN(n23180) );
  ND2D1BWP12T U12859 ( .A1(n22699), .A2(n22700), .ZN(n22694) );
  ND2D1BWP12T U12860 ( .A1(n21935), .A2(n22776), .ZN(n22772) );
  NR2D1BWP12T U12861 ( .A1(a[6]), .A2(b[6]), .ZN(n22783) );
  ND2D1BWP12T U12862 ( .A1(n23017), .A2(n22873), .ZN(n23166) );
  INVD1BWP12T U12863 ( .I(n23166), .ZN(n22828) );
  ND2D1BWP12T U12864 ( .A1(a[3]), .A2(b[3]), .ZN(n23350) );
  ND2D1BWP12T U12865 ( .A1(a[2]), .A2(b[2]), .ZN(n23349) );
  INVD1BWP12T U12866 ( .I(n22971), .ZN(n22990) );
  INVD1BWP12T U12867 ( .I(n23025), .ZN(n23639) );
  NR2D1BWP12T U12868 ( .A1(n22886), .A2(n22885), .ZN(n21936) );
  NR2D1BWP12T U12869 ( .A1(b[5]), .A2(a[5]), .ZN(n22822) );
  INVD1BWP12T U12870 ( .I(n22822), .ZN(n23087) );
  ND2D1BWP12T U12871 ( .A1(b[5]), .A2(a[5]), .ZN(n23346) );
  ND2D1BWP12T U12872 ( .A1(n23087), .A2(n23346), .ZN(n23165) );
  INVD1BWP12T U12873 ( .I(n23165), .ZN(n22832) );
  OA21D1BWP12T U12874 ( .A1(n22828), .A2(n21936), .B(n22832), .Z(n22853) );
  OAI21D1BWP12T U12875 ( .A1(n22853), .A2(n22822), .B(n22823), .ZN(n22821) );
  INVD1BWP12T U12876 ( .I(n22821), .ZN(n22784) );
  ND2D1BWP12T U12877 ( .A1(b[7]), .A2(a[7]), .ZN(n23345) );
  ND2D1BWP12T U12878 ( .A1(n22772), .A2(n23345), .ZN(n22787) );
  INVD1BWP12T U12879 ( .I(n22787), .ZN(n22782) );
  OAI21D1BWP12T U12880 ( .A1(n22783), .A2(n22784), .B(n22782), .ZN(n22794) );
  ND2D1BWP12T U12881 ( .A1(n22772), .A2(n22794), .ZN(n22743) );
  ND2D1BWP12T U12882 ( .A1(b[9]), .A2(a[9]), .ZN(n23364) );
  ND2D1BWP12T U12883 ( .A1(n22694), .A2(n23364), .ZN(n22682) );
  NR2D1BWP12T U12884 ( .A1(n21937), .A2(n22682), .ZN(n21941) );
  OAI21D1BWP12T U12885 ( .A1(n22740), .A2(n22743), .B(n21941), .ZN(n22686) );
  INVD1BWP12T U12886 ( .I(n23063), .ZN(n22668) );
  AOI21D1BWP12T U12887 ( .A1(n22694), .A2(n22686), .B(n22668), .ZN(n22681) );
  OAI21D1BWP12T U12888 ( .A1(n22629), .A2(n22681), .B(n22655), .ZN(n22624) );
  AN2D1BWP12T U12889 ( .A1(n22645), .A2(n22626), .Z(n23095) );
  NR2D1BWP12T U12890 ( .A1(n23181), .A2(n23095), .ZN(n21942) );
  OAI21D1BWP12T U12891 ( .A1(n23351), .A2(n22624), .B(n21942), .ZN(n22570) );
  ND2D1BWP12T U12892 ( .A1(n23180), .A2(n22570), .ZN(n22569) );
  ND2D1BWP12T U12893 ( .A1(n23179), .A2(n22569), .ZN(n22556) );
  ND2D1BWP12T U12894 ( .A1(n22560), .A2(n22556), .ZN(n22555) );
  ND2D1BWP12T U12895 ( .A1(n22549), .A2(n22555), .ZN(n22524) );
  ND2D1BWP12T U12896 ( .A1(n23167), .A2(n22524), .ZN(n22523) );
  INVD1BWP12T U12897 ( .I(n22523), .ZN(n23197) );
  AOI21D1BWP12T U12898 ( .A1(n23484), .A2(n22514), .B(n23197), .ZN(n22469) );
  INVD1BWP12T U12899 ( .I(n23354), .ZN(n22320) );
  OAI211D1BWP12T U12900 ( .A1(n23078), .A2(n22329), .B(n23077), .C(n22320), 
        .ZN(n22295) );
  ND2D1BWP12T U12901 ( .A1(n21945), .A2(n22295), .ZN(n22261) );
  ND2D1BWP12T U12902 ( .A1(n23065), .A2(n22261), .ZN(n22260) );
  AOI21D1BWP12T U12903 ( .A1(n23093), .A2(n22260), .B(n23092), .ZN(n22214) );
  NR2D1BWP12T U12904 ( .A1(n21946), .A2(n22214), .ZN(n22163) );
  INVD1BWP12T U12905 ( .I(n23174), .ZN(n22154) );
  ND2D1BWP12T U12906 ( .A1(b[25]), .A2(a[25]), .ZN(n23357) );
  ND2D1BWP12T U12907 ( .A1(n22154), .A2(n23357), .ZN(n23182) );
  NR2D1BWP12T U12908 ( .A1(n22163), .A2(n23182), .ZN(n22162) );
  NR2D1BWP12T U12909 ( .A1(n23174), .A2(n22162), .ZN(n22115) );
  INVD1BWP12T U12910 ( .I(n23173), .ZN(n22114) );
  NR2D1BWP12T U12911 ( .A1(n22115), .A2(n22114), .ZN(n22113) );
  NR2D1BWP12T U12912 ( .A1(n23185), .A2(n22113), .ZN(n22071) );
  ND2D1BWP12T U12913 ( .A1(b[27]), .A2(a[27]), .ZN(n23373) );
  INR2D1BWP12T U12914 ( .A1(n23373), .B1(n23170), .ZN(n23184) );
  INVD1BWP12T U12915 ( .I(n23184), .ZN(n22070) );
  NR2D1BWP12T U12916 ( .A1(n22071), .A2(n22070), .ZN(n22069) );
  NR2D1BWP12T U12917 ( .A1(n23170), .A2(n22069), .ZN(n22027) );
  NR2D1BWP12T U12918 ( .A1(n22028), .A2(n22027), .ZN(n23205) );
  NR2D1BWP12T U12919 ( .A1(n23540), .A2(n23205), .ZN(n21983) );
  MAOI22D0BWP12T U12920 ( .A1(n21938), .A2(n23045), .B1(n21938), .B2(n23045), 
        .ZN(n23204) );
  NR2D1BWP12T U12921 ( .A1(n23021), .A2(n21939), .ZN(n22945) );
  INVD1BWP12T U12922 ( .I(n22497), .ZN(n22499) );
  INVD1BWP12T U12923 ( .I(n22886), .ZN(n22882) );
  INVD1BWP12T U12924 ( .I(n21940), .ZN(n22989) );
  ND2D1BWP12T U12925 ( .A1(n23347), .A2(n22989), .ZN(n22936) );
  ND2D1BWP12T U12926 ( .A1(n22882), .A2(n22871), .ZN(n22836) );
  AOI21D1BWP12T U12927 ( .A1(n23166), .A2(n22836), .B(n23165), .ZN(n22838) );
  NR2D1BWP12T U12928 ( .A1(n22822), .A2(n22838), .ZN(n22796) );
  NR2D1BWP12T U12929 ( .A1(n23088), .A2(n22796), .ZN(n22795) );
  OAI21D1BWP12T U12930 ( .A1(n22783), .A2(n22795), .B(n22782), .ZN(n22789) );
  ND2D1BWP12T U12931 ( .A1(n22772), .A2(n22789), .ZN(n22742) );
  OAI21D1BWP12T U12932 ( .A1(n22740), .A2(n22742), .B(n21941), .ZN(n22712) );
  AOI21D1BWP12T U12933 ( .A1(n22694), .A2(n22712), .B(n22668), .ZN(n22678) );
  OAI21D1BWP12T U12934 ( .A1(n22629), .A2(n22678), .B(n22655), .ZN(n23105) );
  OAI21D1BWP12T U12935 ( .A1(n23351), .A2(n23105), .B(n21942), .ZN(n22568) );
  ND2D1BWP12T U12936 ( .A1(n22465), .A2(n22463), .ZN(n22462) );
  ND2D1BWP12T U12937 ( .A1(n23086), .A2(n22462), .ZN(n22396) );
  ND2D1BWP12T U12938 ( .A1(n22425), .A2(n22396), .ZN(n22395) );
  ND2D1BWP12T U12939 ( .A1(n21943), .A2(n22395), .ZN(n22359) );
  ND2D1BWP12T U12940 ( .A1(n23099), .A2(n22359), .ZN(n22358) );
  INVD1BWP12T U12941 ( .I(n22358), .ZN(n23111) );
  AOI21D1BWP12T U12942 ( .A1(n21944), .A2(n22383), .B(n23111), .ZN(n22334) );
  OAI211D1BWP12T U12943 ( .A1(n23078), .A2(n22304), .B(n23077), .C(n22320), 
        .ZN(n22301) );
  ND2D1BWP12T U12944 ( .A1(n21945), .A2(n22301), .ZN(n22259) );
  ND2D1BWP12T U12945 ( .A1(n23065), .A2(n22259), .ZN(n23112) );
  AOI21D1BWP12T U12946 ( .A1(n23093), .A2(n23112), .B(n23092), .ZN(n22212) );
  NR2D1BWP12T U12947 ( .A1(n21946), .A2(n22212), .ZN(n22118) );
  MOAI22D0BWP12T U12948 ( .A1(n23042), .A2(n23044), .B1(n23042), .B2(n23044), 
        .ZN(n23120) );
  AOI22D1BWP12T U12949 ( .A1(n23027), .A2(n23204), .B1(n22945), .B2(n23120), 
        .ZN(n21948) );
  OAI211D1BWP12T U12950 ( .A1(n23419), .A2(n22987), .B(n21949), .C(n21948), 
        .ZN(n21950) );
  AO21D1BWP12T U12951 ( .A1(n23160), .A2(n23674), .B(n21950), .Z(result[30])
         );
  MOAI22D0BWP12T U12952 ( .A1(n21951), .A2(n21984), .B1(n21951), .B2(n21984), 
        .ZN(n23161) );
  AOI22D1BWP12T U12953 ( .A1(b[0]), .A2(a[30]), .B1(a[29]), .B2(n22605), .ZN(
        n22309) );
  ND2D1BWP12T U12954 ( .A1(n22806), .A2(a[31]), .ZN(n23662) );
  ND2D1BWP12T U12955 ( .A1(n22009), .A2(n22606), .ZN(n22308) );
  OAI22D1BWP12T U12956 ( .A1(n22309), .A2(n23012), .B1(n23662), .B2(n22308), 
        .ZN(n23213) );
  AOI22D1BWP12T U12957 ( .A1(n22489), .A2(n23213), .B1(n23376), .B2(n23641), 
        .ZN(n21981) );
  ND2D1BWP12T U12958 ( .A1(n23645), .A2(n23499), .ZN(n22974) );
  NR2D1BWP12T U12959 ( .A1(n23509), .A2(n23650), .ZN(n23647) );
  FA1D0BWP12T U12960 ( .A(n21984), .B(n23517), .CI(n21952), .CO(n21908), .S(
        n23604) );
  FA1D0BWP12T U12961 ( .A(n21955), .B(n21954), .CI(n21953), .CO(n21904), .S(
        n23309) );
  AOI22D1BWP12T U12962 ( .A1(n23601), .A2(n23604), .B1(n23658), .B2(n23309), 
        .ZN(n21957) );
  INVD1BWP12T U12963 ( .I(n23372), .ZN(n23652) );
  INVD1BWP12T U12964 ( .I(n23645), .ZN(n22904) );
  AOI32D1BWP12T U12965 ( .A1(b[29]), .A2(a[29]), .A3(n23652), .B1(n22904), 
        .B2(a[29]), .ZN(n21956) );
  OAI211D1BWP12T U12966 ( .A1(n23647), .A2(n21958), .B(n21957), .C(n21956), 
        .ZN(n21972) );
  AOI22D1BWP12T U12967 ( .A1(b[0]), .A2(n22404), .B1(n22406), .B2(n22605), 
        .ZN(n21963) );
  AOI22D1BWP12T U12968 ( .A1(b[0]), .A2(a[14]), .B1(a[15]), .B2(n22009), .ZN(
        n22574) );
  NR3D1BWP12T U12969 ( .A1(b[2]), .A2(n22574), .A3(n22867), .ZN(n21960) );
  AOI22D1BWP12T U12970 ( .A1(b[0]), .A2(a[16]), .B1(a[17]), .B2(n22605), .ZN(
        n22243) );
  AOI22D1BWP12T U12971 ( .A1(b[0]), .A2(a[18]), .B1(a[19]), .B2(n22009), .ZN(
        n22241) );
  OAI22D1BWP12T U12972 ( .A1(n22243), .A2(n22224), .B1(n22241), .B2(n22168), 
        .ZN(n21959) );
  AOI211D1BWP12T U12973 ( .A1(n22447), .A2(n21963), .B(n21960), .C(n21959), 
        .ZN(n22325) );
  ND2D1BWP12T U12974 ( .A1(n22488), .A2(n23667), .ZN(n22377) );
  AOI22D1BWP12T U12975 ( .A1(b[0]), .A2(a[2]), .B1(a[3]), .B2(n22605), .ZN(
        n22141) );
  AOI22D1BWP12T U12976 ( .A1(b[0]), .A2(a[4]), .B1(a[5]), .B2(n22009), .ZN(
        n22045) );
  INVD1BWP12T U12977 ( .I(n22045), .ZN(n22240) );
  INVD1BWP12T U12978 ( .I(n23382), .ZN(n22991) );
  AOI21D1BWP12T U12979 ( .A1(a[1]), .A2(n22009), .B(n22991), .ZN(n23423) );
  INVD1BWP12T U12980 ( .I(n23423), .ZN(n22446) );
  OAI22D1BWP12T U12981 ( .A1(n22240), .A2(n22274), .B1(n22342), .B2(n22446), 
        .ZN(n21961) );
  AOI211D1BWP12T U12982 ( .A1(b[1]), .A2(n22141), .B(n22951), .C(n21961), .ZN(
        n23279) );
  AOI22D1BWP12T U12983 ( .A1(b[0]), .A2(a[24]), .B1(a[25]), .B2(n22605), .ZN(
        n22218) );
  INVD1BWP12T U12984 ( .I(n22218), .ZN(n21974) );
  INVD1BWP12T U12985 ( .I(n22662), .ZN(n22195) );
  AOI22D1BWP12T U12986 ( .A1(b[0]), .A2(n21962), .B1(n23376), .B2(n22009), 
        .ZN(n23441) );
  INVD1BWP12T U12987 ( .I(n22663), .ZN(n23261) );
  OAI22D1BWP12T U12988 ( .A1(n21974), .A2(n22195), .B1(n23441), .B2(n23261), 
        .ZN(n23255) );
  AOI22D1BWP12T U12989 ( .A1(b[0]), .A2(a[22]), .B1(a[23]), .B2(n22605), .ZN(
        n22306) );
  AOI22D1BWP12T U12990 ( .A1(b[0]), .A2(a[26]), .B1(a[27]), .B2(n22009), .ZN(
        n23257) );
  AOI22D1BWP12T U12991 ( .A1(n22306), .A2(n22662), .B1(n23257), .B2(n22663), 
        .ZN(n22039) );
  MAOI22D0BWP12T U12992 ( .A1(n23255), .A2(n22485), .B1(n22485), .B2(n22039), 
        .ZN(n21970) );
  AOI22D1BWP12T U12993 ( .A1(n22606), .A2(n22241), .B1(n22951), .B2(n22574), 
        .ZN(n21965) );
  INVD1BWP12T U12994 ( .I(n21963), .ZN(n22246) );
  AOI22D1BWP12T U12995 ( .A1(n23259), .A2(n22243), .B1(n22607), .B2(n22246), 
        .ZN(n21964) );
  ND2D1BWP12T U12996 ( .A1(n21965), .A2(n21964), .ZN(n22311) );
  AOI22D1BWP12T U12997 ( .A1(b[0]), .A2(a[10]), .B1(a[11]), .B2(n22605), .ZN(
        n22687) );
  AOI22D1BWP12T U12998 ( .A1(b[0]), .A2(a[12]), .B1(a[13]), .B2(n22605), .ZN(
        n22236) );
  AOI22D1BWP12T U12999 ( .A1(n22606), .A2(n22687), .B1(n22607), .B2(n22236), 
        .ZN(n21968) );
  AOI22D1BWP12T U13000 ( .A1(b[0]), .A2(n21966), .B1(n22700), .B2(n22009), 
        .ZN(n22138) );
  INVD1BWP12T U13001 ( .I(n22138), .ZN(n22235) );
  AOI22D1BWP12T U13002 ( .A1(b[0]), .A2(a[6]), .B1(a[7]), .B2(n22605), .ZN(
        n22046) );
  AOI22D1BWP12T U13003 ( .A1(n22235), .A2(n23259), .B1(n22951), .B2(n22046), 
        .ZN(n21967) );
  ND2D1BWP12T U13004 ( .A1(n21968), .A2(n21967), .ZN(n23244) );
  AOI22D1BWP12T U13005 ( .A1(n23270), .A2(n22311), .B1(n23263), .B2(n23244), 
        .ZN(n21969) );
  OAI211D1BWP12T U13006 ( .A1(n23279), .A2(n23265), .B(n21970), .C(n21969), 
        .ZN(n23247) );
  INVD1BWP12T U13007 ( .I(n23644), .ZN(n22493) );
  OAI22D1BWP12T U13008 ( .A1(n22325), .A2(n22377), .B1(n23247), .B2(n22493), 
        .ZN(n21971) );
  AOI211D1BWP12T U13009 ( .A1(n23492), .A2(n22974), .B(n21972), .C(n21971), 
        .ZN(n21980) );
  OAI22D1BWP12T U13010 ( .A1(n22141), .A2(n22168), .B1(n22223), .B2(n22045), 
        .ZN(n23414) );
  AO21D1BWP12T U13011 ( .A1(n22174), .A2(n22446), .B(n23414), .Z(n22833) );
  INVD1BWP12T U13012 ( .I(n22046), .ZN(n22239) );
  AOI22D1BWP12T U13013 ( .A1(n22506), .A2(n22833), .B1(n23456), .B2(n22505), 
        .ZN(n22580) );
  INVD1BWP12T U13014 ( .I(n22988), .ZN(n23442) );
  MAOI22D0BWP12T U13015 ( .A1(n23441), .A2(n23442), .B1(n23257), .B2(n22172), 
        .ZN(n21976) );
  ND2D1BWP12T U13016 ( .A1(n21973), .A2(n22174), .ZN(n22179) );
  INVD1BWP12T U13017 ( .I(n22179), .ZN(n22125) );
  INVD1BWP12T U13018 ( .I(n22306), .ZN(n22041) );
  NR2D1BWP12T U13019 ( .A1(n22220), .A2(n22400), .ZN(n22124) );
  AOI22D1BWP12T U13020 ( .A1(n21974), .A2(n22125), .B1(n22041), .B2(n22124), 
        .ZN(n21975) );
  OAI211D1BWP12T U13021 ( .A1(n23443), .A2(n22580), .B(n21976), .C(n21975), 
        .ZN(n21977) );
  AOI22D1BWP12T U13022 ( .A1(a[29]), .A2(n21978), .B1(n23667), .B2(n21977), 
        .ZN(n21979) );
  ND4D1BWP12T U13023 ( .A1(n21982), .A2(n21981), .A3(n21980), .A4(n21979), 
        .ZN(n21987) );
  MAOI22D0BWP12T U13024 ( .A1(n21983), .A2(n21984), .B1(n21983), .B2(n21984), 
        .ZN(n23592) );
  MAOI22D0BWP12T U13025 ( .A1(n21985), .A2(n21984), .B1(n21985), .B2(n21984), 
        .ZN(n23164) );
  INVD1BWP12T U13026 ( .I(n22945), .ZN(n23670) );
  OAI22D1BWP12T U13027 ( .A1(n23592), .A2(n23669), .B1(n23164), .B2(n23670), 
        .ZN(n21986) );
  AO211D1BWP12T U13028 ( .A1(n23161), .A2(n23674), .B(n21987), .C(n21986), .Z(
        result[29]) );
  MAOI22D0BWP12T U13029 ( .A1(n22028), .A2(n21988), .B1(n22028), .B2(n21988), 
        .ZN(n23155) );
  MOAI22D0BWP12T U13030 ( .A1(n22028), .A2(n21989), .B1(n22028), .B2(n21989), 
        .ZN(n23119) );
  INVD1BWP12T U13031 ( .I(n22124), .ZN(n22171) );
  OAI22D1BWP12T U13032 ( .A1(n21998), .A2(n22171), .B1(n22091), .B2(n22988), 
        .ZN(n21995) );
  INR2D1BWP12T U13033 ( .A1(n22721), .B1(n22867), .ZN(n21992) );
  NR2D1BWP12T U13034 ( .A1(n22867), .A2(n22199), .ZN(n21991) );
  OAI22D1BWP12T U13035 ( .A1(n22081), .A2(n22223), .B1(n22198), .B2(n22224), 
        .ZN(n21990) );
  AOI221D1BWP12T U13036 ( .A1(n21992), .A2(b[2]), .B1(n21991), .B2(n22342), 
        .C(n21990), .ZN(n23438) );
  INVD1BWP12T U13037 ( .I(n23259), .ZN(n22242) );
  MAOI22D0BWP12T U13038 ( .A1(n23438), .A2(n22505), .B1(n22505), .B2(n23424), 
        .ZN(n22609) );
  OAI22D1BWP12T U13039 ( .A1(n21993), .A2(n22179), .B1(n23443), .B2(n22609), 
        .ZN(n21994) );
  AOI211D1BWP12T U13040 ( .A1(n21996), .A2(n23440), .B(n21995), .C(n21994), 
        .ZN(n22006) );
  AOI22D1BWP12T U13041 ( .A1(n21998), .A2(n22662), .B1(n21997), .B2(n22663), 
        .ZN(n22078) );
  NR2D1BWP12T U13042 ( .A1(n22274), .A2(n22081), .ZN(n22000) );
  OAI22D1BWP12T U13043 ( .A1(n22199), .A2(n22244), .B1(n22242), .B2(n22198), 
        .ZN(n21999) );
  AOI211D1BWP12T U13044 ( .A1(n22721), .A2(n22606), .B(n22000), .C(n21999), 
        .ZN(n22336) );
  OAI22D1BWP12T U13045 ( .A1(n22485), .A2(n22001), .B1(n22173), .B2(b[1]), 
        .ZN(n22479) );
  OAI22D1BWP12T U13046 ( .A1(n23516), .A2(n22242), .B1(n22479), .B2(b[2]), 
        .ZN(n22335) );
  INVD1BWP12T U13047 ( .I(n22335), .ZN(n23278) );
  ND2D1BWP12T U13048 ( .A1(b[3]), .A2(n23278), .ZN(n23254) );
  OAI21D1BWP12T U13049 ( .A1(b[3]), .A2(n22336), .B(n23254), .ZN(n23250) );
  OAI22D1BWP12T U13050 ( .A1(n22096), .A2(n22245), .B1(n22200), .B2(n22244), 
        .ZN(n22003) );
  OAI22D1BWP12T U13051 ( .A1(n22533), .A2(n22242), .B1(n22105), .B2(n22274), 
        .ZN(n22002) );
  NR2D1BWP12T U13052 ( .A1(n22003), .A2(n22002), .ZN(n22338) );
  AOI22D1BWP12T U13053 ( .A1(b[4]), .A2(n23250), .B1(n23270), .B2(n22338), 
        .ZN(n22004) );
  OAI221D1BWP12T U13054 ( .A1(b[1]), .A2(n22005), .B1(n22485), .B2(n22078), 
        .C(n22004), .ZN(n23287) );
  OAI22D1BWP12T U13055 ( .A1(n22006), .A2(n22987), .B1(n23287), .B2(n22493), 
        .ZN(n22026) );
  INVD1BWP12T U13056 ( .I(n22220), .ZN(n22126) );
  AOI22D1BWP12T U13057 ( .A1(n22096), .A2(n22227), .B1(n22200), .B2(n22126), 
        .ZN(n22008) );
  AOI22D1BWP12T U13058 ( .A1(n22533), .A2(n22174), .B1(n22105), .B2(n22447), 
        .ZN(n22007) );
  ND2D1BWP12T U13059 ( .A1(n22008), .A2(n22007), .ZN(n22345) );
  ND2D1BWP12T U13060 ( .A1(b[0]), .A2(n22485), .ZN(n23262) );
  OAI22D1BWP12T U13061 ( .A1(a[31]), .A2(n22009), .B1(a[28]), .B2(b[1]), .ZN(
        n22010) );
  AOI22D1BWP12T U13062 ( .A1(n22864), .A2(n22011), .B1(n23262), .B2(n22010), 
        .ZN(n22348) );
  NR2D1BWP12T U13063 ( .A1(b[3]), .A2(b[2]), .ZN(n22920) );
  INVD1BWP12T U13064 ( .I(n22920), .ZN(n22844) );
  INR2D1BWP12T U13065 ( .A1(n22348), .B1(n22844), .ZN(n23221) );
  OAI21D1BWP12T U13066 ( .A1(n22012), .A2(n22858), .B(n22209), .ZN(n22076) );
  INVD1BWP12T U13067 ( .I(n22076), .ZN(n22054) );
  AOI22D1BWP12T U13068 ( .A1(b[28]), .A2(n22974), .B1(a[27]), .B2(n22586), 
        .ZN(n22013) );
  AOI21D1BWP12T U13069 ( .A1(n22054), .A2(n22013), .B(a[28]), .ZN(n22017) );
  INVD1BWP12T U13070 ( .I(n23647), .ZN(n22998) );
  AOI22D1BWP12T U13071 ( .A1(n23517), .A2(n22998), .B1(n23658), .B2(n23324), 
        .ZN(n22015) );
  INVD1BWP12T U13072 ( .I(n23646), .ZN(n22674) );
  ND2D1BWP12T U13073 ( .A1(n22674), .A2(n23294), .ZN(n22913) );
  OAI211D1BWP12T U13074 ( .A1(n22663), .A2(n23646), .B(n22015), .C(n22913), 
        .ZN(n22016) );
  AOI211D1BWP12T U13075 ( .A1(n22489), .A2(n23221), .B(n22017), .C(n22016), 
        .ZN(n22024) );
  NR2D1BWP12T U13076 ( .A1(b[28]), .A2(op[2]), .ZN(n22020) );
  ND2D1BWP12T U13077 ( .A1(n22019), .A2(n22018), .ZN(n23030) );
  OAI22D1BWP12T U13078 ( .A1(a[27]), .A2(n22031), .B1(n22020), .B2(n23030), 
        .ZN(n22022) );
  MOAI22D0BWP12T U13079 ( .A1(n22028), .A2(n22021), .B1(n22028), .B2(n22021), 
        .ZN(n23621) );
  AOI22D1BWP12T U13080 ( .A1(a[28]), .A2(n22022), .B1(n23621), .B2(n23601), 
        .ZN(n22023) );
  OAI211D1BWP12T U13081 ( .A1(n22377), .A2(n22345), .B(n22024), .C(n22023), 
        .ZN(n22025) );
  AOI211D1BWP12T U13082 ( .A1(n22945), .A2(n23119), .B(n22026), .C(n22025), 
        .ZN(n22030) );
  AOI32D1BWP12T U13083 ( .A1(n22028), .A2(n23027), .A3(n22027), .B1(n23205), 
        .B2(n23027), .ZN(n22029) );
  OAI211D1BWP12T U13084 ( .A1(n22948), .A2(n23155), .B(n22030), .C(n22029), 
        .ZN(result[28]) );
  AOI32D1BWP12T U13085 ( .A1(n22032), .A2(n22031), .A3(n22812), .B1(n23030), 
        .B2(n22031), .ZN(n22068) );
  NR2D1BWP12T U13086 ( .A1(b[0]), .A2(a[27]), .ZN(n22033) );
  NR2D1BWP12T U13087 ( .A1(a[28]), .A2(n22605), .ZN(n22134) );
  OAI32D1BWP12T U13088 ( .A1(b[1]), .A2(n22033), .A3(n22134), .B1(n22485), 
        .B2(n22309), .ZN(n22364) );
  MAOI22D0BWP12T U13089 ( .A1(n22364), .A2(n22920), .B1(n22342), .B2(n23662), 
        .ZN(n23407) );
  INVD1BWP12T U13090 ( .I(n23407), .ZN(n22641) );
  ND2D1BWP12T U13091 ( .A1(n22365), .A2(n22641), .ZN(n23230) );
  ND2D1BWP12T U13092 ( .A1(n23017), .A2(n22964), .ZN(n23661) );
  AOI22D1BWP12T U13093 ( .A1(n22662), .A2(n22246), .B1(n22663), .B2(n22218), 
        .ZN(n22146) );
  AOI22D1BWP12T U13094 ( .A1(b[1]), .A2(n23423), .B1(n22141), .B2(n22485), 
        .ZN(n22368) );
  NR2D1BWP12T U13095 ( .A1(b[2]), .A2(n22806), .ZN(n22363) );
  AOI22D1BWP12T U13096 ( .A1(n22606), .A2(n22235), .B1(n22607), .B2(n22687), 
        .ZN(n22035) );
  AOI22D1BWP12T U13097 ( .A1(n23259), .A2(n22046), .B1(n22951), .B2(n22045), 
        .ZN(n22034) );
  ND2D1BWP12T U13098 ( .A1(n22035), .A2(n22034), .ZN(n22370) );
  MAOI22D0BWP12T U13099 ( .A1(n22368), .A2(n22363), .B1(n22370), .B2(b[3]), 
        .ZN(n23290) );
  AOI22D1BWP12T U13100 ( .A1(n22607), .A2(n22241), .B1(n23259), .B2(n22574), 
        .ZN(n22037) );
  AOI22D1BWP12T U13101 ( .A1(n22606), .A2(n22243), .B1(n22951), .B2(n22236), 
        .ZN(n22036) );
  ND2D1BWP12T U13102 ( .A1(n22037), .A2(n22036), .ZN(n22369) );
  AOI22D1BWP12T U13103 ( .A1(b[4]), .A2(n23290), .B1(n23270), .B2(n22369), 
        .ZN(n22038) );
  OAI221D1BWP12T U13104 ( .A1(b[1]), .A2(n22039), .B1(n22485), .B2(n22146), 
        .C(n22038), .ZN(n22040) );
  NR2D1BWP12T U13105 ( .A1(n23294), .A2(n22040), .ZN(n23286) );
  INVD1BWP12T U13106 ( .I(n23298), .ZN(n22403) );
  ND2D1BWP12T U13107 ( .A1(n23667), .A2(n23544), .ZN(n22181) );
  AOI22D1BWP12T U13108 ( .A1(n22864), .A2(n22218), .B1(n23257), .B2(n22867), 
        .ZN(n23444) );
  OAI22D1BWP12T U13109 ( .A1(n22041), .A2(n22179), .B1(n23444), .B2(n22926), 
        .ZN(n22042) );
  AOI211D1BWP12T U13110 ( .A1(n22124), .A2(n22246), .B(n22181), .C(n22042), 
        .ZN(n22050) );
  NR2D1BWP12T U13111 ( .A1(n22867), .A2(n22236), .ZN(n22638) );
  NR2D1BWP12T U13112 ( .A1(n22574), .A2(n22224), .ZN(n22044) );
  OAI22D1BWP12T U13113 ( .A1(n22243), .A2(n22168), .B1(n22241), .B2(n22223), 
        .ZN(n22043) );
  AOI211D1BWP12T U13114 ( .A1(n22638), .A2(n22342), .B(n22044), .C(n22043), 
        .ZN(n22381) );
  AOI22D1BWP12T U13115 ( .A1(n22141), .A2(n22867), .B1(n23500), .B2(n22993), 
        .ZN(n22902) );
  ND2D1BWP12T U13116 ( .A1(n22902), .A2(n22099), .ZN(n23422) );
  OAI22D1BWP12T U13117 ( .A1(n22235), .A2(n22168), .B1(n22220), .B2(n22045), 
        .ZN(n22048) );
  OAI22D1BWP12T U13118 ( .A1(n22687), .A2(n22223), .B1(n22224), .B2(n22046), 
        .ZN(n22047) );
  NR2D1BWP12T U13119 ( .A1(n22048), .A2(n22047), .ZN(n23435) );
  OA22D1BWP12T U13120 ( .A1(n22505), .A2(n23422), .B1(n22506), .B2(n23435), 
        .Z(n22636) );
  AOI22D1BWP12T U13121 ( .A1(n22381), .A2(n22488), .B1(n22504), .B2(n22636), 
        .ZN(n22049) );
  AOI22D1BWP12T U13122 ( .A1(n23286), .A2(n22403), .B1(n22050), .B2(n22049), 
        .ZN(n22062) );
  INR2D1BWP12T U13123 ( .A1(n22052), .B1(n22051), .ZN(n22053) );
  MOAI22D0BWP12T U13124 ( .A1(n23184), .A2(n22053), .B1(n23184), .B2(n22053), 
        .ZN(n23619) );
  ND2D1BWP12T U13125 ( .A1(n23409), .A2(n23585), .ZN(n22343) );
  OAI22D1BWP12T U13126 ( .A1(n23407), .A2(n22343), .B1(a[27]), .B2(n22054), 
        .ZN(n22060) );
  FA1D0BWP12T U13127 ( .A(n22057), .B(n22056), .CI(n22055), .CO(n22014), .S(
        n23310) );
  AOI22D1BWP12T U13128 ( .A1(n23491), .A2(n22974), .B1(n23658), .B2(n23310), 
        .ZN(n22058) );
  OAI21D1BWP12T U13129 ( .A1(n23294), .A2(n22691), .B(n22674), .ZN(n22185) );
  OAI211D1BWP12T U13130 ( .A1(n23647), .A2(n23514), .B(n22058), .C(n22185), 
        .ZN(n22059) );
  AOI211D1BWP12T U13131 ( .A1(n23601), .A2(n23619), .B(n22060), .C(n22059), 
        .ZN(n22061) );
  OAI211D1BWP12T U13132 ( .A1(n23230), .A2(n23661), .B(n22062), .C(n22061), 
        .ZN(n22067) );
  MOAI22D0BWP12T U13133 ( .A1(n22063), .A2(n23184), .B1(n22063), .B2(n23184), 
        .ZN(n23116) );
  AOI22D1BWP12T U13134 ( .A1(n23184), .A2(n22065), .B1(n22070), .B2(n22064), 
        .ZN(n23156) );
  OAI22D1BWP12T U13135 ( .A1(n23116), .A2(n23670), .B1(n22948), .B2(n23156), 
        .ZN(n22066) );
  AOI211D1BWP12T U13136 ( .A1(a[27]), .A2(n22068), .B(n22067), .C(n22066), 
        .ZN(n22073) );
  AOI32D1BWP12T U13137 ( .A1(n22071), .A2(n23027), .A3(n22070), .B1(n22069), 
        .B2(n23027), .ZN(n22072) );
  ND2D1BWP12T U13138 ( .A1(n22073), .A2(n22072), .ZN(result[27]) );
  MOAI22D0BWP12T U13139 ( .A1(n23173), .A2(n22074), .B1(n23173), .B2(n22074), 
        .ZN(n23158) );
  MAOI22D0BWP12T U13140 ( .A1(n22075), .A2(n23173), .B1(n22075), .B2(n23173), 
        .ZN(n23118) );
  OA211D1BWP12T U13141 ( .A1(n22087), .A2(n22157), .B(n23553), .C(n22076), .Z(
        n22112) );
  NR2D1BWP12T U13142 ( .A1(b[2]), .A2(n22077), .ZN(n23281) );
  OAI22D1BWP12T U13143 ( .A1(n22268), .A2(n23261), .B1(n22178), .B2(n22195), 
        .ZN(n22205) );
  MAOI22D0BWP12T U13144 ( .A1(b[1]), .A2(n22205), .B1(n22078), .B2(b[1]), .ZN(
        n22085) );
  AOI22D1BWP12T U13145 ( .A1(n22865), .A2(n23259), .B1(n22951), .B2(n22100), 
        .ZN(n22080) );
  ND2D1BWP12T U13146 ( .A1(n22607), .A2(n22721), .ZN(n22079) );
  OAI211D1BWP12T U13147 ( .A1(n22245), .A2(n22198), .B(n22080), .C(n22079), 
        .ZN(n23246) );
  INVD1BWP12T U13148 ( .I(n23270), .ZN(n22727) );
  NR2D1BWP12T U13149 ( .A1(n22274), .A2(n22196), .ZN(n22083) );
  MOAI22D0BWP12T U13150 ( .A1(n22244), .A2(n22081), .B1(n22606), .B2(n22533), 
        .ZN(n22082) );
  AOI211D1BWP12T U13151 ( .A1(n23259), .A2(n22200), .B(n22083), .C(n22082), 
        .ZN(n22397) );
  MAOI22D0BWP12T U13152 ( .A1(n23263), .A2(n23246), .B1(n22727), .B2(n22397), 
        .ZN(n22084) );
  OAI211D1BWP12T U13153 ( .A1(n23281), .A2(n23265), .B(n22085), .C(n22084), 
        .ZN(n23248) );
  NR2D1BWP12T U13154 ( .A1(a[26]), .A2(n22088), .ZN(n23503) );
  AOI211D1BWP12T U13155 ( .A1(n22088), .A2(n22812), .B(n22087), .C(n23030), 
        .ZN(n22090) );
  OAI22D1BWP12T U13156 ( .A1(n23647), .A2(n23512), .B1(n22244), .B2(n23646), 
        .ZN(n22089) );
  AO211D1BWP12T U13157 ( .A1(n23326), .A2(n23658), .B(n22090), .C(n22089), .Z(
        n22095) );
  NR2D1BWP12T U13158 ( .A1(a[29]), .A2(n22009), .ZN(n22093) );
  OAI32D1BWP12T U13159 ( .A1(n22864), .A2(n22093), .A3(n22092), .B1(n22091), 
        .B2(n22867), .ZN(n22272) );
  MAOI22D0BWP12T U13160 ( .A1(n22342), .A2(n22272), .B1(n22273), .B2(n22242), 
        .ZN(n22666) );
  OAI31D1BWP12T U13161 ( .A1(n22666), .A2(n23041), .A3(n22691), .B(n22185), 
        .ZN(n22094) );
  AOI211D1BWP12T U13162 ( .A1(n23503), .A2(n22974), .B(n22095), .C(n22094), 
        .ZN(n22110) );
  NR2D1BWP12T U13163 ( .A1(n22346), .A2(n22179), .ZN(n22104) );
  OAI22D1BWP12T U13164 ( .A1(n22201), .A2(n22220), .B1(n22533), .B2(n22168), 
        .ZN(n22098) );
  OAI22D1BWP12T U13165 ( .A1(n22200), .A2(n22224), .B1(n22096), .B2(n22223), 
        .ZN(n22097) );
  NR2D1BWP12T U13166 ( .A1(n22098), .A2(n22097), .ZN(n22401) );
  ND2D1BWP12T U13167 ( .A1(n22099), .A2(n22933), .ZN(n23460) );
  INVD1BWP12T U13168 ( .I(n23460), .ZN(n22413) );
  MAOI22D0BWP12T U13169 ( .A1(n22506), .A2(n22413), .B1(n22402), .B2(n22506), 
        .ZN(n23426) );
  AOI22D1BWP12T U13170 ( .A1(n22401), .A2(n22488), .B1(n23426), .B2(n22504), 
        .ZN(n22101) );
  OAI211D1BWP12T U13171 ( .A1(n22102), .A2(n22926), .B(n22101), .C(n23544), 
        .ZN(n22103) );
  AOI211D1BWP12T U13172 ( .A1(n22124), .A2(n22105), .B(n22104), .C(n22103), 
        .ZN(n23466) );
  INR2D1BWP12T U13173 ( .A1(n22107), .B1(n22106), .ZN(n22108) );
  MOAI22D0BWP12T U13174 ( .A1(n23173), .A2(n22108), .B1(n23173), .B2(n22108), 
        .ZN(n23612) );
  AOI22D1BWP12T U13175 ( .A1(n23466), .A2(n23667), .B1(n23601), .B2(n23612), 
        .ZN(n22109) );
  OAI211D1BWP12T U13176 ( .A1(n23248), .A2(n22493), .B(n22110), .C(n22109), 
        .ZN(n22111) );
  AOI211D1BWP12T U13177 ( .A1(n22945), .A2(n23118), .B(n22112), .C(n22111), 
        .ZN(n22117) );
  AOI32D1BWP12T U13178 ( .A1(n22115), .A2(n23027), .A3(n22114), .B1(n22113), 
        .B2(n23027), .ZN(n22116) );
  OAI211D1BWP12T U13179 ( .A1(n23158), .A2(n22948), .B(n22117), .C(n22116), 
        .ZN(result[26]) );
  MAOI22D0BWP12T U13180 ( .A1(n22118), .A2(n23182), .B1(n22118), .B2(n23182), 
        .ZN(n23115) );
  IND2D1BWP12T U13181 ( .A1(n22119), .B1(n22187), .ZN(n22120) );
  MAOI22D0BWP12T U13182 ( .A1(n23182), .A2(n22120), .B1(n23182), .B2(n22120), 
        .ZN(n23154) );
  IND2D1BWP12T U13183 ( .A1(n22122), .B1(n22121), .ZN(n22123) );
  MAOI22D0BWP12T U13184 ( .A1(n23182), .A2(n22123), .B1(n23182), .B2(n22123), 
        .ZN(n23615) );
  OAI22D1BWP12T U13185 ( .A1(n23615), .A2(n23653), .B1(a[25]), .B2(n22209), 
        .ZN(n22161) );
  AOI22D1BWP12T U13186 ( .A1(n22124), .A2(n22241), .B1(n23440), .B2(n22306), 
        .ZN(n22133) );
  AOI22D1BWP12T U13187 ( .A1(n22125), .A2(n22246), .B1(n23442), .B2(n22218), 
        .ZN(n22132) );
  AOI22D1BWP12T U13188 ( .A1(n22574), .A2(n22227), .B1(n22687), .B2(n22126), 
        .ZN(n22128) );
  AOI22D1BWP12T U13189 ( .A1(n22447), .A2(n22243), .B1(n22174), .B2(n22236), 
        .ZN(n22127) );
  ND2D1BWP12T U13190 ( .A1(n22128), .A2(n22127), .ZN(n22435) );
  AOI22D1BWP12T U13191 ( .A1(n22240), .A2(n22174), .B1(n22239), .B2(n22227), 
        .ZN(n22130) );
  ND2D1BWP12T U13192 ( .A1(n22447), .A2(n22138), .ZN(n22129) );
  OAI211D1BWP12T U13193 ( .A1(n22141), .A2(n22220), .B(n22130), .C(n22129), 
        .ZN(n22460) );
  AOI32D1BWP12T U13194 ( .A1(n22447), .A2(n22506), .A3(n22446), .B1(n22505), 
        .B2(n22460), .ZN(n23427) );
  AOI22D1BWP12T U13195 ( .A1(n22488), .A2(n22435), .B1(n23427), .B2(n22504), 
        .ZN(n22131) );
  ND4D1BWP12T U13196 ( .A1(n22133), .A2(n22132), .A3(n22131), .A4(n23544), 
        .ZN(n23467) );
  NR2D1BWP12T U13197 ( .A1(b[0]), .A2(a[25]), .ZN(n22135) );
  OAI32D1BWP12T U13198 ( .A1(n22864), .A2(n22135), .A3(n22134), .B1(n23257), 
        .B2(n22867), .ZN(n22307) );
  INVD1BWP12T U13199 ( .I(n22309), .ZN(n22136) );
  OAI222D1BWP12T U13200 ( .A1(n22244), .A2(a[31]), .B1(n22307), .B2(b[2]), 
        .C1(n22242), .C2(n22136), .ZN(n23225) );
  NR2D1BWP12T U13201 ( .A1(b[3]), .A2(n23225), .ZN(n22705) );
  ND2D1BWP12T U13202 ( .A1(n22137), .A2(n22343), .ZN(n22455) );
  AOI22D1BWP12T U13203 ( .A1(n22662), .A2(n22241), .B1(n22663), .B2(n22306), 
        .ZN(n22145) );
  NR2D1BWP12T U13204 ( .A1(n23423), .A2(n22274), .ZN(n23272) );
  NR2D1BWP12T U13205 ( .A1(n22274), .A2(n22138), .ZN(n22140) );
  OAI22D1BWP12T U13206 ( .A1(n22240), .A2(n22242), .B1(n22239), .B2(n22245), 
        .ZN(n22139) );
  AOI211D1BWP12T U13207 ( .A1(n22951), .A2(n22141), .B(n22140), .C(n22139), 
        .ZN(n22437) );
  AOI22D1BWP12T U13208 ( .A1(b[3]), .A2(n23272), .B1(n22437), .B2(n22806), 
        .ZN(n23282) );
  AOI22D1BWP12T U13209 ( .A1(n22606), .A2(n22574), .B1(n22607), .B2(n22243), 
        .ZN(n22143) );
  AOI22D1BWP12T U13210 ( .A1(n22687), .A2(n22951), .B1(n23259), .B2(n22236), 
        .ZN(n22142) );
  ND2D1BWP12T U13211 ( .A1(n22143), .A2(n22142), .ZN(n22438) );
  AOI22D1BWP12T U13212 ( .A1(b[4]), .A2(n23282), .B1(n23270), .B2(n22438), 
        .ZN(n22144) );
  OAI221D1BWP12T U13213 ( .A1(b[1]), .A2(n22146), .B1(n22485), .B2(n22145), 
        .C(n22144), .ZN(n23276) );
  FA1D0BWP12T U13214 ( .A(n22149), .B(n22148), .CI(n22147), .CO(n22086), .S(
        n23313) );
  AOI22D1BWP12T U13215 ( .A1(n23650), .A2(n22151), .B1(n22150), .B2(n22998), 
        .ZN(n22152) );
  OAI211D1BWP12T U13216 ( .A1(n23372), .A2(n23357), .B(n22152), .C(n23645), 
        .ZN(n22153) );
  AOI22D1BWP12T U13217 ( .A1(n23313), .A2(n23658), .B1(n22154), .B2(n22153), 
        .ZN(n22155) );
  OAI211D1BWP12T U13218 ( .A1(n22493), .A2(n23276), .B(n22155), .C(n22185), 
        .ZN(n22156) );
  AOI31D1BWP12T U13219 ( .A1(n22705), .A2(n22489), .A3(n22455), .B(n22156), 
        .ZN(n22159) );
  ND2D1BWP12T U13220 ( .A1(a[25]), .A2(n22157), .ZN(n22158) );
  OAI211D1BWP12T U13221 ( .A1(n23467), .A2(n22987), .B(n22159), .C(n22158), 
        .ZN(n22160) );
  AOI211D1BWP12T U13222 ( .A1(n23154), .A2(n23674), .B(n22161), .C(n22160), 
        .ZN(n22165) );
  AOI32D1BWP12T U13223 ( .A1(n22163), .A2(n23027), .A3(n23182), .B1(n22162), 
        .B2(n23027), .ZN(n22164) );
  OAI211D1BWP12T U13224 ( .A1(n23115), .A2(n23670), .B(n22165), .C(n22164), 
        .ZN(result[25]) );
  AOI22D1BWP12T U13225 ( .A1(n23027), .A2(n22260), .B1(n22945), .B2(n23112), 
        .ZN(n22217) );
  ND2D1BWP12T U13226 ( .A1(n23093), .A2(n23092), .ZN(n23074) );
  INVD1BWP12T U13227 ( .I(n23030), .ZN(n23000) );
  OAI21D1BWP12T U13228 ( .A1(b[24]), .A2(op[2]), .B(n23000), .ZN(n22166) );
  OAI32D1BWP12T U13229 ( .A1(n23560), .A2(a[23]), .A3(n22266), .B1(n22166), 
        .B2(n23560), .ZN(n22211) );
  MAOI22D0BWP12T U13230 ( .A1(n23092), .A2(n22167), .B1(n23092), .B2(n22167), 
        .ZN(n23613) );
  OAI22D1BWP12T U13231 ( .A1(n22200), .A2(n22168), .B1(n22721), .B2(n22220), 
        .ZN(n22170) );
  OAI22D1BWP12T U13232 ( .A1(n22201), .A2(n22224), .B1(n22533), .B2(n22223), 
        .ZN(n22169) );
  NR2D1BWP12T U13233 ( .A1(n22170), .A2(n22169), .ZN(n23462) );
  OAI22D1BWP12T U13234 ( .A1(n22346), .A2(n22172), .B1(n22171), .B2(n22196), 
        .ZN(n22183) );
  AOI22D1BWP12T U13235 ( .A1(n22174), .A2(n22173), .B1(n22227), .B2(n22199), 
        .ZN(n22176) );
  ND2D1BWP12T U13236 ( .A1(n22447), .A2(n22198), .ZN(n22175) );
  OAI211D1BWP12T U13237 ( .A1(n22177), .A2(n22220), .B(n22176), .C(n22175), 
        .ZN(n22487) );
  ND2D1BWP12T U13238 ( .A1(b[3]), .A2(n22607), .ZN(n22310) );
  NR2D1BWP12T U13239 ( .A1(n23516), .A2(n22310), .ZN(n22197) );
  AOI21D1BWP12T U13240 ( .A1(n22487), .A2(n22505), .B(n22197), .ZN(n23425) );
  OAI22D1BWP12T U13241 ( .A1(n22268), .A2(n22988), .B1(n22179), .B2(n22178), 
        .ZN(n22180) );
  AO211D1BWP12T U13242 ( .A1(n23425), .A2(n22504), .B(n22181), .C(n22180), .Z(
        n22182) );
  AOI211D1BWP12T U13243 ( .A1(n22488), .A2(n23462), .B(n22183), .C(n22182), 
        .ZN(n22189) );
  AOI22D1BWP12T U13244 ( .A1(n23502), .A2(n22974), .B1(n23658), .B2(n23312), 
        .ZN(n22186) );
  OAI211D1BWP12T U13245 ( .A1(n23647), .A2(n22187), .B(n22186), .C(n22185), 
        .ZN(n22188) );
  AOI211D1BWP12T U13246 ( .A1(n23601), .A2(n23613), .B(n22189), .C(n22188), 
        .ZN(n22208) );
  ND2D1BWP12T U13247 ( .A1(b[0]), .A2(n22190), .ZN(n22193) );
  NR2D1BWP12T U13248 ( .A1(b[0]), .A2(a[24]), .ZN(n22191) );
  NR2D1BWP12T U13249 ( .A1(n22191), .A2(n22271), .ZN(n22192) );
  AOI32D1BWP12T U13250 ( .A1(n22194), .A2(b[1]), .A3(n22193), .B1(n22192), 
        .B2(n22485), .ZN(n22347) );
  MAOI22D0BWP12T U13251 ( .A1(b[2]), .A2(n22348), .B1(n22347), .B2(b[2]), .ZN(
        n23226) );
  NR2D1BWP12T U13252 ( .A1(b[3]), .A2(n23226), .ZN(n22736) );
  OAI22D1BWP12T U13253 ( .A1(n22346), .A2(n23261), .B1(n22196), .B2(n22195), 
        .ZN(n22206) );
  NR2D1BWP12T U13254 ( .A1(b[3]), .A2(n22342), .ZN(n23008) );
  OAI22D1BWP12T U13255 ( .A1(n22199), .A2(n22245), .B1(n22274), .B2(n22198), 
        .ZN(n22478) );
  OAI22D1BWP12T U13256 ( .A1(n22201), .A2(n22242), .B1(n22200), .B2(n22245), 
        .ZN(n22203) );
  OAI22D1BWP12T U13257 ( .A1(n22721), .A2(n22244), .B1(n22533), .B2(n22274), 
        .ZN(n22202) );
  NR2D1BWP12T U13258 ( .A1(n22203), .A2(n22202), .ZN(n22480) );
  MOAI22D0BWP12T U13259 ( .A1(n23280), .A2(n23017), .B1(n23270), .B2(n22480), 
        .ZN(n22204) );
  AOI221D1BWP12T U13260 ( .A1(b[1]), .A2(n22206), .B1(n22485), .B2(n22205), 
        .C(n22204), .ZN(n23283) );
  AOI22D1BWP12T U13261 ( .A1(n22736), .A2(n22489), .B1(n23283), .B2(n23644), 
        .ZN(n22207) );
  OAI211D1BWP12T U13262 ( .A1(a[24]), .A2(n22209), .B(n22208), .C(n22207), 
        .ZN(n22210) );
  AOI211D1BWP12T U13263 ( .A1(n22945), .A2(n22212), .B(n22211), .C(n22210), 
        .ZN(n22216) );
  MOAI22D0BWP12T U13264 ( .A1(n23092), .A2(n22213), .B1(n23092), .B2(n22213), 
        .ZN(n23153) );
  AOI22D1BWP12T U13265 ( .A1(n23153), .A2(n23674), .B1(n23027), .B2(n22214), 
        .ZN(n22215) );
  OAI211D1BWP12T U13266 ( .A1(n22217), .A2(n23074), .B(n22216), .C(n22215), 
        .ZN(result[24]) );
  ND2D1BWP12T U13267 ( .A1(a[31]), .A2(b[3]), .ZN(n22637) );
  INVD1BWP12T U13268 ( .I(n22637), .ZN(n22275) );
  AOI22D1BWP12T U13269 ( .A1(b[2]), .A2(n22364), .B1(n22362), .B2(n22342), 
        .ZN(n23406) );
  NR2D1BWP12T U13270 ( .A1(b[3]), .A2(n23406), .ZN(n22765) );
  NR2D1BWP12T U13271 ( .A1(n22275), .A2(n22765), .ZN(n23218) );
  INVD1BWP12T U13272 ( .I(n22489), .ZN(n22350) );
  AOI211D1BWP12T U13273 ( .A1(n22219), .A2(n22343), .B(n23218), .C(n22350), 
        .ZN(n22257) );
  NR2D1BWP12T U13274 ( .A1(n22867), .A2(n22246), .ZN(n22361) );
  NR2D1BWP12T U13275 ( .A1(n22241), .A2(n22224), .ZN(n22222) );
  OAI22D1BWP12T U13276 ( .A1(n22306), .A2(n22223), .B1(n22243), .B2(n22220), 
        .ZN(n22221) );
  AOI211D1BWP12T U13277 ( .A1(n22361), .A2(b[2]), .B(n22222), .C(n22221), .ZN(
        n23451) );
  ND2D1BWP12T U13278 ( .A1(n22766), .A2(n23667), .ZN(n22888) );
  NR2D1BWP12T U13279 ( .A1(n22867), .A2(n22235), .ZN(n22759) );
  OAI22D1BWP12T U13280 ( .A1(n22687), .A2(n22224), .B1(n22574), .B2(n22223), 
        .ZN(n22225) );
  AOI221D1BWP12T U13281 ( .A1(n22638), .A2(b[2]), .B1(n22759), .B2(n22342), 
        .C(n22225), .ZN(n23434) );
  OAI22D1BWP12T U13282 ( .A1(n23451), .A2(n22888), .B1(n23434), .B2(n22377), 
        .ZN(n22256) );
  AOI222D1BWP12T U13283 ( .A1(n22240), .A2(n22227), .B1(n22239), .B2(n22447), 
        .C1(n22226), .C2(n22902), .ZN(n23433) );
  ND2D1BWP12T U13284 ( .A1(n22691), .A2(n22504), .ZN(n22517) );
  NR3D1BWP12T U13285 ( .A1(n22517), .A2(n22987), .A3(n22506), .ZN(n22412) );
  INVD1BWP12T U13286 ( .I(n22412), .ZN(n22449) );
  INVD1BWP12T U13287 ( .I(n22513), .ZN(n22426) );
  OAI21D1BWP12T U13288 ( .A1(n23433), .A2(n22449), .B(n22426), .ZN(n22255) );
  ND2D1BWP12T U13289 ( .A1(n22586), .A2(n22228), .ZN(n22283) );
  FA1D0BWP12T U13290 ( .A(n22231), .B(n22230), .CI(n22229), .CO(n22184), .S(
        n23315) );
  AOI21D1BWP12T U13291 ( .A1(n22233), .A2(n23511), .B(n22232), .ZN(n22234) );
  MAOI22D0BWP12T U13292 ( .A1(n23065), .A2(n22234), .B1(n23065), .B2(n22234), 
        .ZN(n23596) );
  MAOI22D0BWP12T U13293 ( .A1(n23658), .A2(n23315), .B1(n23596), .B2(n23653), 
        .ZN(n22253) );
  AOI22D1BWP12T U13294 ( .A1(n22235), .A2(n22951), .B1(n23259), .B2(n22687), 
        .ZN(n22238) );
  AOI22D1BWP12T U13295 ( .A1(n22606), .A2(n22236), .B1(n22607), .B2(n22574), 
        .ZN(n22237) );
  ND2D1BWP12T U13296 ( .A1(n22238), .A2(n22237), .ZN(n23264) );
  INVD1BWP12T U13297 ( .I(n23294), .ZN(n23397) );
  ND2D1BWP12T U13298 ( .A1(n23397), .A2(n23265), .ZN(n22399) );
  OAI222D1BWP12T U13299 ( .A1(n22368), .A2(n22342), .B1(n22240), .B2(n22245), 
        .C1(n22239), .C2(n22274), .ZN(n23275) );
  INVD1BWP12T U13300 ( .I(n23275), .ZN(n23266) );
  OAI22D1BWP12T U13301 ( .A1(n22274), .A2(n22306), .B1(n22242), .B2(n22241), 
        .ZN(n22248) );
  OAI22D1BWP12T U13302 ( .A1(n22246), .A2(n22245), .B1(n22244), .B2(n22243), 
        .ZN(n22247) );
  NR2D1BWP12T U13303 ( .A1(n22248), .A2(n22247), .ZN(n23269) );
  MOAI22D0BWP12T U13304 ( .A1(n23266), .A2(n23017), .B1(n23258), .B2(n23269), 
        .ZN(n22249) );
  AOI211D1BWP12T U13305 ( .A1(b[3]), .A2(n23264), .B(n22399), .C(n22249), .ZN(
        n23284) );
  AOI22D1BWP12T U13306 ( .A1(n23652), .A2(n23352), .B1(n23650), .B2(n22267), 
        .ZN(n22250) );
  OAI211D1BWP12T U13307 ( .A1(b[23]), .A2(n23647), .B(n22250), .C(n23645), 
        .ZN(n22251) );
  AOI22D1BWP12T U13308 ( .A1(n22403), .A2(n23284), .B1(n23093), .B2(n22251), 
        .ZN(n22252) );
  OAI211D1BWP12T U13309 ( .A1(a[23]), .A2(n22283), .B(n22253), .C(n22252), 
        .ZN(n22254) );
  NR4D0BWP12T U13310 ( .A1(n22257), .A2(n22256), .A3(n22255), .A4(n22254), 
        .ZN(n22265) );
  MOAI22D0BWP12T U13311 ( .A1(n22258), .A2(n23065), .B1(n22258), .B2(n23065), 
        .ZN(n23152) );
  OAI32D1BWP12T U13312 ( .A1(n23670), .A2(n23065), .A3(n22259), .B1(n23112), 
        .B2(n23670), .ZN(n22263) );
  INVD1BWP12T U13313 ( .I(n23027), .ZN(n23669) );
  OAI32D1BWP12T U13314 ( .A1(n23669), .A2(n23065), .A3(n22261), .B1(n22260), 
        .B2(n23669), .ZN(n22262) );
  AOI211D1BWP12T U13315 ( .A1(n23674), .A2(n23152), .B(n22263), .C(n22262), 
        .ZN(n22264) );
  OAI211D1BWP12T U13316 ( .A1(n22267), .A2(n22266), .B(n22265), .C(n22264), 
        .ZN(result[23]) );
  NR2D1BWP12T U13317 ( .A1(b[0]), .A2(a[22]), .ZN(n22270) );
  NR2D1BWP12T U13318 ( .A1(n22268), .A2(n22867), .ZN(n22269) );
  AOI221D1BWP12T U13319 ( .A1(n22271), .A2(b[1]), .B1(n22270), .B2(n22485), 
        .C(n22269), .ZN(n22407) );
  AOI22D1BWP12T U13320 ( .A1(b[2]), .A2(n22272), .B1(n22407), .B2(n22342), 
        .ZN(n22537) );
  OAI32D1BWP12T U13321 ( .A1(n22806), .A2(n22273), .A3(n22274), .B1(b[3]), 
        .B2(n22537), .ZN(n23239) );
  INVD1BWP12T U13322 ( .I(n23239), .ZN(n22810) );
  ND2D1BWP12T U13323 ( .A1(n22275), .A2(n22274), .ZN(n22847) );
  ND2D1BWP12T U13324 ( .A1(n22810), .A2(n22847), .ZN(n22808) );
  INVD1BWP12T U13325 ( .I(n22808), .ZN(n23402) );
  NR2D1BWP12T U13326 ( .A1(a[31]), .A2(n23409), .ZN(n23401) );
  AOI211D1BWP12T U13327 ( .A1(n23409), .A2(n23402), .B(n23401), .C(n22706), 
        .ZN(n22290) );
  MOAI22D0BWP12T U13328 ( .A1(n23017), .A2(n23271), .B1(n23245), .B2(b[3]), 
        .ZN(n22276) );
  AOI211D1BWP12T U13329 ( .A1(n23258), .A2(n22277), .B(n22399), .C(n22276), 
        .ZN(n23293) );
  INVD1BWP12T U13330 ( .I(n22888), .ZN(n22834) );
  AOI22D1BWP12T U13331 ( .A1(n23293), .A2(n22403), .B1(n23458), .B2(n22834), 
        .ZN(n22287) );
  INVD1BWP12T U13332 ( .I(n22377), .ZN(n22461) );
  FA1D0BWP12T U13333 ( .A(n23077), .B(n23510), .CI(n22278), .CO(n22233), .S(
        n23598) );
  MOAI22D0BWP12T U13334 ( .A1(n23598), .A2(n23653), .B1(n23658), .B2(n23311), 
        .ZN(n22281) );
  MOAI22D0BWP12T U13335 ( .A1(n23511), .A2(n23022), .B1(n23077), .B2(n23650), 
        .ZN(n22280) );
  AOI211D1BWP12T U13336 ( .A1(n23353), .A2(n23652), .B(n22281), .C(n22280), 
        .ZN(n22282) );
  OAI21D1BWP12T U13337 ( .A1(n23066), .A2(n23645), .B(n22282), .ZN(n22285) );
  OAI22D1BWP12T U13338 ( .A1(n22810), .A2(n23661), .B1(a[22]), .B2(n22283), 
        .ZN(n22284) );
  AOI211D1BWP12T U13339 ( .A1(n23437), .A2(n22461), .B(n22285), .C(n22284), 
        .ZN(n22286) );
  OAI211D1BWP12T U13340 ( .A1(n22288), .A2(n22449), .B(n22287), .C(n22286), 
        .ZN(n22289) );
  AOI211D1BWP12T U13341 ( .A1(n22291), .A2(n22328), .B(n22290), .C(n22289), 
        .ZN(n22300) );
  NR2D1BWP12T U13342 ( .A1(n23078), .A2(n23077), .ZN(n22298) );
  ND2D1BWP12T U13343 ( .A1(n23670), .A2(n23669), .ZN(n23055) );
  OAI211D1BWP12T U13344 ( .A1(n22329), .A2(n23669), .B(n23069), .C(n22304), 
        .ZN(n22297) );
  OAI21D1BWP12T U13345 ( .A1(a[21]), .A2(n22293), .B(n22292), .ZN(n22294) );
  MOAI22D0BWP12T U13346 ( .A1(n23077), .A2(n22294), .B1(n23077), .B2(n22294), 
        .ZN(n23150) );
  OAI22D1BWP12T U13347 ( .A1(n23150), .A2(n22948), .B1(n23669), .B2(n22295), 
        .ZN(n22296) );
  AOI31D1BWP12T U13348 ( .A1(n22298), .A2(n23055), .A3(n22297), .B(n22296), 
        .ZN(n22299) );
  OAI211D1BWP12T U13349 ( .A1(n22301), .A2(n23670), .B(n22300), .C(n22299), 
        .ZN(result[22]) );
  MAOI22D0BWP12T U13350 ( .A1(n23069), .A2(n22302), .B1(n23069), .B2(n22302), 
        .ZN(n23149) );
  ND2D1BWP12T U13351 ( .A1(n23069), .A2(n22304), .ZN(n22303) );
  OAI32D1BWP12T U13352 ( .A1(n23670), .A2(n23069), .A3(n22304), .B1(n22303), 
        .B2(n23670), .ZN(n22327) );
  AOI22D1BWP12T U13353 ( .A1(n23456), .A2(n22461), .B1(n22412), .B2(n22833), 
        .ZN(n22305) );
  OA31D1BWP12T U13354 ( .A1(a[21]), .A2(n22858), .A3(n22344), .B(n22305), .Z(
        n22324) );
  OAI222D1BWP12T U13355 ( .A1(n22640), .A2(n22406), .B1(n22993), .B2(n23560), 
        .C1(n22867), .C2(n22306), .ZN(n22454) );
  AOI22D1BWP12T U13356 ( .A1(b[2]), .A2(n22307), .B1(n22454), .B2(n22342), 
        .ZN(n23452) );
  OAI222D1BWP12T U13357 ( .A1(n22310), .A2(n22309), .B1(n23452), .B2(b[3]), 
        .C1(n22308), .C2(n22637), .ZN(n23408) );
  INVD1BWP12T U13358 ( .I(n22399), .ZN(n22440) );
  AOI22D1BWP12T U13359 ( .A1(b[3]), .A2(n23244), .B1(n23258), .B2(n22311), 
        .ZN(n22312) );
  OAI211D1BWP12T U13360 ( .A1(n23279), .A2(n23017), .B(n22440), .C(n22312), 
        .ZN(n23295) );
  OAI22D1BWP12T U13361 ( .A1(n22847), .A2(n22343), .B1(n23295), .B2(n23298), 
        .ZN(n22322) );
  FA1D0BWP12T U13362 ( .A(n22313), .B(n23069), .CI(n23530), .CO(n22278), .S(
        n23599) );
  FA1D0BWP12T U13363 ( .A(n22316), .B(n22315), .CI(n22314), .CO(n22279), .S(
        n23316) );
  MOAI22D0BWP12T U13364 ( .A1(n23599), .A2(n23653), .B1(n23658), .B2(n23316), 
        .ZN(n22318) );
  OAI22D1BWP12T U13365 ( .A1(n23078), .A2(n23645), .B1(n23022), .B2(n23510), 
        .ZN(n22317) );
  AOI211D1BWP12T U13366 ( .A1(n23069), .A2(n23650), .B(n22318), .C(n22317), 
        .ZN(n22319) );
  OAI211D1BWP12T U13367 ( .A1(n23372), .A2(n22320), .B(n22319), .C(n22426), 
        .ZN(n22321) );
  AOI211D1BWP12T U13368 ( .A1(n22489), .A2(n23408), .B(n22322), .C(n22321), 
        .ZN(n22323) );
  OAI211D1BWP12T U13369 ( .A1(n22325), .A2(n22888), .B(n22324), .C(n22323), 
        .ZN(n22326) );
  AOI211D1BWP12T U13370 ( .A1(n22328), .A2(a[21]), .B(n22327), .C(n22326), 
        .ZN(n22333) );
  INVD1BWP12T U13371 ( .I(n22329), .ZN(n22331) );
  INVD1BWP12T U13372 ( .I(n23069), .ZN(n22330) );
  OAI221D1BWP12T U13373 ( .A1(n23069), .A2(n22331), .B1(n22330), .B2(n22329), 
        .C(n23027), .ZN(n22332) );
  OAI211D1BWP12T U13374 ( .A1(n23149), .A2(n22948), .B(n22333), .C(n22332), 
        .ZN(result[21]) );
  MAOI22D0BWP12T U13375 ( .A1(n22334), .A2(n22352), .B1(n22334), .B2(n22352), 
        .ZN(n23114) );
  OAI22D1BWP12T U13376 ( .A1(n22336), .A2(n22806), .B1(n23017), .B2(n22335), 
        .ZN(n22337) );
  AOI211D1BWP12T U13377 ( .A1(n23258), .A2(n22338), .B(n22399), .C(n22337), 
        .ZN(n23299) );
  NR2D1BWP12T U13378 ( .A1(n22342), .A2(n22637), .ZN(n22870) );
  AOI222D1BWP12T U13379 ( .A1(n22757), .A2(a[20]), .B1(n22842), .B2(a[23]), 
        .C1(n22864), .C2(n22346), .ZN(n22486) );
  AOI22D1BWP12T U13380 ( .A1(b[2]), .A2(n22347), .B1(n22486), .B2(n22342), 
        .ZN(n23416) );
  AOI22D1BWP12T U13381 ( .A1(n22348), .A2(n22363), .B1(n23416), .B2(n22806), 
        .ZN(n23211) );
  MAOI22D0BWP12T U13382 ( .A1(n22352), .A2(n22349), .B1(n22352), .B2(n22349), 
        .ZN(n23147) );
  MAOI22D0BWP12T U13383 ( .A1(n22352), .A2(n22351), .B1(n22352), .B2(n22351), 
        .ZN(n23636) );
  MAOI22D0BWP12T U13384 ( .A1(n22354), .A2(n22353), .B1(n22354), .B2(n22353), 
        .ZN(n23201) );
  MAOI22D0BWP12T U13385 ( .A1(n22385), .A2(n22355), .B1(n22385), .B2(n22355), 
        .ZN(n22356) );
  MAOI22D0BWP12T U13386 ( .A1(n22356), .A2(n22408), .B1(n22356), .B2(n22408), 
        .ZN(n23634) );
  MAOI22D0BWP12T U13387 ( .A1(n22357), .A2(n22385), .B1(n22357), .B2(n22385), 
        .ZN(n23203) );
  OAI32D1BWP12T U13388 ( .A1(n23670), .A2(n23099), .A3(n22359), .B1(n22358), 
        .B2(n23670), .ZN(n22391) );
  NR2D1BWP12T U13389 ( .A1(n22383), .A2(n22640), .ZN(n22360) );
  AO211D1BWP12T U13390 ( .A1(n22842), .A2(a[22]), .B(n22361), .C(n22360), .Z(
        n22755) );
  AOI22D1BWP12T U13391 ( .A1(b[2]), .A2(n22362), .B1(n22755), .B2(n22342), 
        .ZN(n23463) );
  NR2D1BWP12T U13392 ( .A1(b[3]), .A2(n23463), .ZN(n22366) );
  AOI211D1BWP12T U13393 ( .A1(n22364), .A2(n22363), .B(n22366), .C(n22870), 
        .ZN(n23212) );
  OAI31D1BWP12T U13394 ( .A1(n22366), .A2(n22925), .A3(n22365), .B(n22489), 
        .ZN(n22389) );
  OAI21D1BWP12T U13395 ( .A1(n22367), .A2(n22585), .B(n22586), .ZN(n22450) );
  ND2D1BWP12T U13396 ( .A1(n22450), .A2(n22421), .ZN(n22419) );
  ND2D1BWP12T U13397 ( .A1(n22920), .A2(n22368), .ZN(n23274) );
  AOI222D1BWP12T U13398 ( .A1(n23274), .A2(b[4]), .B1(n22370), .B2(b[3]), .C1(
        n22369), .C2(n23258), .ZN(n23252) );
  FA1D0BWP12T U13399 ( .A(n22373), .B(n22372), .CI(n22371), .CO(n22340), .S(
        n23322) );
  AOI22D1BWP12T U13400 ( .A1(n23322), .A2(n23658), .B1(n23650), .B2(n23099), 
        .ZN(n22375) );
  OAI211D1BWP12T U13401 ( .A1(a[19]), .A2(op[2]), .B(b[19]), .C(n23000), .ZN(
        n22374) );
  OAI211D1BWP12T U13402 ( .A1(n23022), .A2(n22376), .B(n22375), .C(n22374), 
        .ZN(n22379) );
  OAI22D1BWP12T U13403 ( .A1(n23435), .A2(n22377), .B1(n23422), .B2(n22449), 
        .ZN(n22378) );
  AOI211D1BWP12T U13404 ( .A1(n23252), .A2(n23644), .B(n22379), .C(n22378), 
        .ZN(n22380) );
  OAI211D1BWP12T U13405 ( .A1(n22381), .A2(n22888), .B(n22380), .C(n22426), 
        .ZN(n22382) );
  AOI31D1BWP12T U13406 ( .A1(n22383), .A2(n22586), .A3(n22419), .B(n22382), 
        .ZN(n22388) );
  OAI21D1BWP12T U13407 ( .A1(a[18]), .A2(n22417), .B(n23645), .ZN(n22386) );
  MAOI22D0BWP12T U13408 ( .A1(n22385), .A2(n22384), .B1(n22385), .B2(n22384), 
        .ZN(n23144) );
  AOI22D1BWP12T U13409 ( .A1(a[19]), .A2(n22386), .B1(n23674), .B2(n23144), 
        .ZN(n22387) );
  OAI211D1BWP12T U13410 ( .A1(n23212), .A2(n22389), .B(n22388), .C(n22387), 
        .ZN(n22390) );
  AOI211D1BWP12T U13411 ( .A1(n23027), .A2(n23203), .B(n22391), .C(n22390), 
        .ZN(n22392) );
  OAI21D1BWP12T U13412 ( .A1(n23634), .A2(n23653), .B(n22392), .ZN(result[19])
         );
  MAOI22D0BWP12T U13413 ( .A1(n22425), .A2(n22393), .B1(n22425), .B2(n22393), 
        .ZN(n23633) );
  MOAI22D0BWP12T U13414 ( .A1(n22425), .A2(n22394), .B1(n22425), .B2(n22394), 
        .ZN(n23196) );
  OAI32D1BWP12T U13415 ( .A1(n23670), .A2(n22425), .A3(n22396), .B1(n22395), 
        .B2(n23670), .ZN(n22431) );
  OAI22D1BWP12T U13416 ( .A1(n22397), .A2(n22691), .B1(n23281), .B2(n23017), 
        .ZN(n22398) );
  AOI211D1BWP12T U13417 ( .A1(n23270), .A2(n23246), .B(n22399), .C(n22398), 
        .ZN(n23301) );
  INVD1BWP12T U13418 ( .I(n22488), .ZN(n23450) );
  OAI22D1BWP12T U13419 ( .A1(n22402), .A2(n23450), .B1(n22401), .B2(n22400), 
        .ZN(n23431) );
  AOI22D1BWP12T U13420 ( .A1(n23301), .A2(n22403), .B1(n23667), .B2(n23431), 
        .ZN(n22429) );
  AOI22D1BWP12T U13421 ( .A1(b[0]), .A2(a[19]), .B1(a[18]), .B2(n22605), .ZN(
        n22483) );
  AO22D1BWP12T U13422 ( .A1(n22485), .A2(n22483), .B1(n22404), .B2(n22843), 
        .Z(n22405) );
  AOI31D1BWP12T U13423 ( .A1(b[0]), .A2(b[1]), .A3(n22406), .B(n22405), .ZN(
        n22536) );
  AOI22D1BWP12T U13424 ( .A1(b[2]), .A2(n22407), .B1(n22536), .B2(n22342), 
        .ZN(n22660) );
  ND2D1BWP12T U13425 ( .A1(n22660), .A2(n22806), .ZN(n22950) );
  INVD1BWP12T U13426 ( .I(n22950), .ZN(n22423) );
  ND2D1BWP12T U13427 ( .A1(n22951), .A2(n22674), .ZN(n22416) );
  INVD1BWP12T U13428 ( .I(n22408), .ZN(n23528) );
  FA1D0BWP12T U13429 ( .A(n22411), .B(n22410), .CI(n22409), .CO(n22373), .S(
        n23303) );
  AOI22D1BWP12T U13430 ( .A1(n23528), .A2(n22998), .B1(n23658), .B2(n23303), 
        .ZN(n22415) );
  AOI22D1BWP12T U13431 ( .A1(n23506), .A2(n22974), .B1(n22413), .B2(n22412), 
        .ZN(n22414) );
  OAI211D1BWP12T U13432 ( .A1(n22423), .A2(n22416), .B(n22415), .C(n22414), 
        .ZN(n22422) );
  AOI32D1BWP12T U13433 ( .A1(n22418), .A2(n22417), .A3(n22812), .B1(n23030), 
        .B2(n22417), .ZN(n22420) );
  OAI32D1BWP12T U13434 ( .A1(n22422), .A2(n22421), .A3(n22420), .B1(n22419), 
        .B2(n22422), .ZN(n22428) );
  OAI21D1BWP12T U13435 ( .A1(b[3]), .A2(n22660), .B(n22666), .ZN(n23216) );
  INR2D1BWP12T U13436 ( .A1(n23216), .B1(n22423), .ZN(n22965) );
  MAOI22D0BWP12T U13437 ( .A1(n22425), .A2(n22424), .B1(n22425), .B2(n22424), 
        .ZN(n23145) );
  AOI22D1BWP12T U13438 ( .A1(n22489), .A2(n22965), .B1(n23674), .B2(n23145), 
        .ZN(n22427) );
  ND4D1BWP12T U13439 ( .A1(n22429), .A2(n22428), .A3(n22427), .A4(n22426), 
        .ZN(n22430) );
  AOI211D1BWP12T U13440 ( .A1(n23027), .A2(n23196), .B(n22431), .C(n22430), 
        .ZN(n22432) );
  OAI21D1BWP12T U13441 ( .A1(n23633), .A2(n23653), .B(n22432), .ZN(result[18])
         );
  MAOI22D0BWP12T U13442 ( .A1(n22465), .A2(n22433), .B1(n22465), .B2(n22433), 
        .ZN(n23200) );
  OAI32D1BWP12T U13443 ( .A1(n22434), .A2(b[17]), .A3(op[2]), .B1(n23000), 
        .B2(n22434), .ZN(n22436) );
  OAI22D1BWP12T U13444 ( .A1(n22436), .A2(n22441), .B1(n22435), .B2(n22888), 
        .ZN(n22459) );
  MAOI22D0BWP12T U13445 ( .A1(n23258), .A2(n22438), .B1(n22806), .B2(n22437), 
        .ZN(n22439) );
  OAI211D1BWP12T U13446 ( .A1(n23272), .A2(n23017), .B(n22440), .C(n22439), 
        .ZN(n23383) );
  INVD1BWP12T U13447 ( .I(n22974), .ZN(n22907) );
  ND2D1BWP12T U13448 ( .A1(b[17]), .A2(n22441), .ZN(n23487) );
  OAI22D1BWP12T U13449 ( .A1(n23647), .A2(n22442), .B1(n22907), .B2(n23487), 
        .ZN(n22453) );
  MAOI22D0BWP12T U13450 ( .A1(n22465), .A2(n22443), .B1(n22465), .B2(n22443), 
        .ZN(n22444) );
  MAOI22D0BWP12T U13451 ( .A1(n23519), .A2(n22444), .B1(n23519), .B2(n22444), 
        .ZN(n23595) );
  MOAI22D0BWP12T U13452 ( .A1(n23653), .A2(n23595), .B1(n23658), .B2(n23331), 
        .ZN(n22452) );
  ND2D1BWP12T U13453 ( .A1(n22447), .A2(n22446), .ZN(n22448) );
  OAI22D1BWP12T U13454 ( .A1(a[17]), .A2(n22450), .B1(n22449), .B2(n22448), 
        .ZN(n22451) );
  NR4D0BWP12T U13455 ( .A1(n22513), .A2(n22453), .A3(n22452), .A4(n22451), 
        .ZN(n22457) );
  AOI22D1BWP12T U13456 ( .A1(b[0]), .A2(a[18]), .B1(a[17]), .B2(n22605), .ZN(
        n22516) );
  AOI22D1BWP12T U13457 ( .A1(b[2]), .A2(n22454), .B1(n22575), .B2(n22342), 
        .ZN(n22703) );
  NR2D1BWP12T U13458 ( .A1(b[3]), .A2(n22703), .ZN(n23222) );
  INVD1BWP12T U13459 ( .I(n23225), .ZN(n22693) );
  AO21D1BWP12T U13460 ( .A1(b[3]), .A2(n22693), .B(n23222), .Z(n22985) );
  OAI211D1BWP12T U13461 ( .A1(n23222), .A2(n22455), .B(n22489), .C(n22985), 
        .ZN(n22456) );
  OAI211D1BWP12T U13462 ( .A1(n23298), .A2(n23383), .B(n22457), .C(n22456), 
        .ZN(n22458) );
  AOI211D1BWP12T U13463 ( .A1(n22461), .A2(n22460), .B(n22459), .C(n22458), 
        .ZN(n22468) );
  OAI21D1BWP12T U13464 ( .A1(n22465), .A2(n22463), .B(n22462), .ZN(n22466) );
  MOAI22D0BWP12T U13465 ( .A1(n22465), .A2(n22464), .B1(n22465), .B2(n22464), 
        .ZN(n23146) );
  AOI22D1BWP12T U13466 ( .A1(n22945), .A2(n22466), .B1(n23146), .B2(n23674), 
        .ZN(n22467) );
  OAI211D1BWP12T U13467 ( .A1(n23200), .A2(n23669), .B(n22468), .C(n22467), 
        .ZN(result[17]) );
  MAOI22D0BWP12T U13468 ( .A1(n22469), .A2(n22497), .B1(n22469), .B2(n22497), 
        .ZN(n23199) );
  ND2D1BWP12T U13469 ( .A1(b[16]), .A2(n22515), .ZN(n23486) );
  FA1D0BWP12T U13470 ( .A(n23521), .B(n22470), .CI(n22497), .CO(n22443), .S(
        n23603) );
  FA1D0BWP12T U13471 ( .A(n22473), .B(n22472), .CI(n22471), .CO(n22445), .S(
        n23317) );
  AOI22D1BWP12T U13472 ( .A1(n23601), .A2(n23603), .B1(n23658), .B2(n23317), 
        .ZN(n22476) );
  OAI21D1BWP12T U13473 ( .A1(n23372), .A2(n23340), .B(n23645), .ZN(n22474) );
  AOI22D1BWP12T U13474 ( .A1(n23519), .A2(n22998), .B1(n23084), .B2(n22474), 
        .ZN(n22475) );
  OAI211D1BWP12T U13475 ( .A1(n23486), .A2(n23499), .B(n22476), .C(n22475), 
        .ZN(n22496) );
  OAI22D1BWP12T U13476 ( .A1(n23462), .A2(n22888), .B1(n22477), .B2(n22510), 
        .ZN(n22495) );
  NR2D1BWP12T U13477 ( .A1(n23516), .A2(n23012), .ZN(n23273) );
  AOI32D1BWP12T U13478 ( .A1(b[2]), .A2(b[3]), .A3(n22479), .B1(n22478), .B2(
        b[3]), .ZN(n22482) );
  ND2D1BWP12T U13479 ( .A1(n23258), .A2(n22480), .ZN(n22481) );
  OAI211D1BWP12T U13480 ( .A1(n23273), .A2(n23017), .B(n22482), .C(n22481), 
        .ZN(n23249) );
  ND2D1BWP12T U13481 ( .A1(a[16]), .A2(n22009), .ZN(n22484) );
  AO32D1BWP12T U13482 ( .A1(n22535), .A2(n22485), .A3(n22484), .B1(n22483), 
        .B2(b[1]), .Z(n22608) );
  OAI22D1BWP12T U13483 ( .A1(n22342), .A2(n22486), .B1(n22608), .B2(b[2]), 
        .ZN(n23455) );
  ND2D1BWP12T U13484 ( .A1(n23455), .A2(n22806), .ZN(n23224) );
  OAI21D1BWP12T U13485 ( .A1(n23226), .A2(n22806), .B(n23224), .ZN(n23018) );
  AOI22D1BWP12T U13486 ( .A1(b[4]), .A2(n23273), .B1(n22488), .B2(n22487), 
        .ZN(n23420) );
  MAOI22D0BWP12T U13487 ( .A1(n22489), .A2(n23018), .B1(n23420), .B2(n22987), 
        .ZN(n22492) );
  OAI31D1BWP12T U13488 ( .A1(a[14]), .A2(n22490), .A3(n22585), .B(n22586), 
        .ZN(n22541) );
  ND2D1BWP12T U13489 ( .A1(n22514), .A2(n22541), .ZN(n22507) );
  ND3D1BWP12T U13490 ( .A1(n22515), .A2(n22586), .A3(n22507), .ZN(n22491) );
  OAI211D1BWP12T U13491 ( .A1(n22493), .A2(n23249), .B(n22492), .C(n22491), 
        .ZN(n22494) );
  NR4D0BWP12T U13492 ( .A1(n22513), .A2(n22496), .A3(n22495), .A4(n22494), 
        .ZN(n22502) );
  MOAI22D0BWP12T U13493 ( .A1(n22498), .A2(n22497), .B1(n22498), .B2(n22497), 
        .ZN(n23138) );
  MOAI22D0BWP12T U13494 ( .A1(n22500), .A2(n22499), .B1(n22500), .B2(n22499), 
        .ZN(n23110) );
  AOI22D1BWP12T U13495 ( .A1(n23674), .A2(n23138), .B1(n22945), .B2(n23110), 
        .ZN(n22501) );
  OAI211D1BWP12T U13496 ( .A1(n23199), .A2(n23669), .B(n22502), .C(n22501), 
        .ZN(result[16]) );
  MAOI22D0BWP12T U13497 ( .A1(n22528), .A2(n22503), .B1(n22528), .B2(n22503), 
        .ZN(n23139) );
  NR2D1BWP12T U13498 ( .A1(n22504), .A2(n22987), .ZN(n22540) );
  AOI22D1BWP12T U13499 ( .A1(n22506), .A2(n23433), .B1(n23434), .B2(n22505), 
        .ZN(n23446) );
  AOI221D1BWP12T U13500 ( .A1(b[15]), .A2(n23652), .B1(n23484), .B2(n22998), 
        .C(n22514), .ZN(n22509) );
  AOI21D1BWP12T U13501 ( .A1(b[15]), .A2(n22904), .B(n22507), .ZN(n22508) );
  AOI31D1BWP12T U13502 ( .A1(n23645), .A2(n22510), .A3(n22509), .B(n22508), 
        .ZN(n22522) );
  ND2D1BWP12T U13503 ( .A1(n23270), .A2(n23644), .ZN(n22538) );
  ND2D1BWP12T U13504 ( .A1(n23258), .A2(n23644), .ZN(n22887) );
  OAI22D1BWP12T U13505 ( .A1(n22528), .A2(n23499), .B1(n22887), .B2(n23264), 
        .ZN(n22512) );
  AOI211D1BWP12T U13506 ( .A1(n23304), .A2(n23658), .B(n22513), .C(n22512), 
        .ZN(n22520) );
  OAI222D1BWP12T U13507 ( .A1(n22516), .A2(n22485), .B1(n23262), .B2(n22515), 
        .C1(n22640), .C2(n22514), .ZN(n22754) );
  AOI22D1BWP12T U13508 ( .A1(n22663), .A2(n22754), .B1(n22662), .B2(n22755), 
        .ZN(n23388) );
  AOI222D1BWP12T U13509 ( .A1(n22517), .A2(n23388), .B1(n23642), .B2(b[4]), 
        .C1(n23406), .C2(n23270), .ZN(n23227) );
  OAI21D1BWP12T U13510 ( .A1(n23406), .A2(n22727), .B(n23388), .ZN(n22518) );
  AOI22D1BWP12T U13511 ( .A1(n23227), .A2(n22964), .B1(n22925), .B2(n22518), 
        .ZN(n22519) );
  OAI211D1BWP12T U13512 ( .A1(n23275), .A2(n22538), .B(n22520), .C(n22519), 
        .ZN(n22521) );
  AOI211D1BWP12T U13513 ( .A1(n22540), .A2(n23446), .B(n22522), .C(n22521), 
        .ZN(n22532) );
  OAI32D1BWP12T U13514 ( .A1(n23669), .A2(n23167), .A3(n22524), .B1(n22523), 
        .B2(n23669), .ZN(n22530) );
  MAOI22D0BWP12T U13515 ( .A1(n23167), .A2(n22525), .B1(n23167), .B2(n22525), 
        .ZN(n23108) );
  OAI21D1BWP12T U13516 ( .A1(n22528), .A2(n22527), .B(n22526), .ZN(n23626) );
  OAI22D1BWP12T U13517 ( .A1(n23108), .A2(n23670), .B1(n23653), .B2(n23626), 
        .ZN(n22529) );
  NR2D1BWP12T U13518 ( .A1(n22530), .A2(n22529), .ZN(n22531) );
  OAI211D1BWP12T U13519 ( .A1(n23139), .A2(n22948), .B(n22532), .C(n22531), 
        .ZN(result[15]) );
  ND2D1BWP12T U13520 ( .A1(a[14]), .A2(n22009), .ZN(n22534) );
  AOI32D1BWP12T U13521 ( .A1(n22535), .A2(n22867), .A3(n22534), .B1(n22533), 
        .B2(n22864), .ZN(n22958) );
  AOI22D1BWP12T U13522 ( .A1(b[2]), .A2(n22536), .B1(n22958), .B2(n22342), 
        .ZN(n22807) );
  AOI22D1BWP12T U13523 ( .A1(n23270), .A2(n22537), .B1(n23258), .B2(n22807), 
        .ZN(n22546) );
  INVD1BWP12T U13524 ( .I(n22538), .ZN(n22671) );
  AOI22D1BWP12T U13525 ( .A1(n22546), .A2(n22539), .B1(n22671), .B2(n23271), 
        .ZN(n22567) );
  INVD1BWP12T U13526 ( .I(n22540), .ZN(n22737) );
  OAI22D1BWP12T U13527 ( .A1(n22542), .A2(n22737), .B1(a[14]), .B2(n22541), 
        .ZN(n22543) );
  AOI31D1BWP12T U13528 ( .A1(n22587), .A2(n22670), .A3(n22544), .B(n22543), 
        .ZN(n22566) );
  MAOI22D0BWP12T U13529 ( .A1(n23178), .A2(n22545), .B1(n23178), .B2(n22545), 
        .ZN(n23137) );
  OAI21D1BWP12T U13530 ( .A1(n23223), .A2(n23017), .B(n22546), .ZN(n23214) );
  OAI22D1BWP12T U13531 ( .A1(n23041), .A2(n23214), .B1(n23245), .B2(n22887), 
        .ZN(n22554) );
  AOI21D1BWP12T U13532 ( .A1(n23509), .A2(n22547), .B(n23650), .ZN(n22552) );
  INVD1BWP12T U13533 ( .I(n22549), .ZN(n23168) );
  OAI21D1BWP12T U13534 ( .A1(n23168), .A2(n22812), .B(n23341), .ZN(n22550) );
  AOI22D1BWP12T U13535 ( .A1(n23658), .A2(n23302), .B1(n23000), .B2(n22550), 
        .ZN(n22551) );
  OAI211D1BWP12T U13536 ( .A1(n22552), .A2(n23178), .B(n22551), .C(n22913), 
        .ZN(n22553) );
  AOI211D1BWP12T U13537 ( .A1(n23137), .A2(n23674), .B(n22554), .C(n22553), 
        .ZN(n22565) );
  OAI32D1BWP12T U13538 ( .A1(n23669), .A2(n22560), .A3(n22556), .B1(n22555), 
        .B2(n23669), .ZN(n22563) );
  IND2D1BWP12T U13539 ( .A1(n22558), .B1(n22557), .ZN(n22559) );
  MAOI22D0BWP12T U13540 ( .A1(n23178), .A2(n22559), .B1(n23178), .B2(n22559), 
        .ZN(n23627) );
  MAOI22D0BWP12T U13541 ( .A1(n22561), .A2(n22560), .B1(n22561), .B2(n22560), 
        .ZN(n23107) );
  OAI22D1BWP12T U13542 ( .A1(n23627), .A2(n23653), .B1(n23107), .B2(n23670), 
        .ZN(n22562) );
  NR2D1BWP12T U13543 ( .A1(n22563), .A2(n22562), .ZN(n22564) );
  ND4D1BWP12T U13544 ( .A1(n22567), .A2(n22566), .A3(n22565), .A4(n22564), 
        .ZN(result[14]) );
  MAOI22D0BWP12T U13545 ( .A1(n22568), .A2(n22584), .B1(n22568), .B2(n22584), 
        .ZN(n23104) );
  OAI32D1BWP12T U13546 ( .A1(n23669), .A2(n23180), .A3(n22570), .B1(n22569), 
        .B2(n23669), .ZN(n22600) );
  INR2D1BWP12T U13547 ( .A1(n22572), .B1(n22571), .ZN(n22573) );
  MAOI22D0BWP12T U13548 ( .A1(n23180), .A2(n22573), .B1(n23180), .B2(n22573), 
        .ZN(n23628) );
  NR2D1BWP12T U13549 ( .A1(n23017), .A2(n23213), .ZN(n22579) );
  INVD1BWP12T U13550 ( .I(n22964), .ZN(n22809) );
  AOI22D1BWP12T U13551 ( .A1(b[2]), .A2(n22575), .B1(n22690), .B2(n22342), 
        .ZN(n23417) );
  AOI22D1BWP12T U13552 ( .A1(n23270), .A2(n23452), .B1(n23258), .B2(n23417), 
        .ZN(n23208) );
  INVD1BWP12T U13553 ( .I(n23208), .ZN(n22578) );
  AOI21D1BWP12T U13554 ( .A1(n22579), .A2(n22576), .B(n22578), .ZN(n23391) );
  ND2D1BWP12T U13555 ( .A1(n23391), .A2(n22925), .ZN(n22577) );
  OAI31D1BWP12T U13556 ( .A1(n22579), .A2(n22809), .A3(n22578), .B(n22577), 
        .ZN(n22582) );
  OAI22D1BWP12T U13557 ( .A1(n23244), .A2(n22887), .B1(n22580), .B2(n22737), 
        .ZN(n22581) );
  AOI211D1BWP12T U13558 ( .A1(n23279), .A2(n22671), .B(n22582), .C(n22581), 
        .ZN(n22598) );
  MOAI22D0BWP12T U13559 ( .A1(n22584), .A2(n22583), .B1(n22584), .B2(n22583), 
        .ZN(n23136) );
  ND2D1BWP12T U13560 ( .A1(n22587), .A2(n22670), .ZN(n22590) );
  OAI21D1BWP12T U13561 ( .A1(b[13]), .A2(op[2]), .B(n23000), .ZN(n22589) );
  ND2D1BWP12T U13562 ( .A1(n22586), .A2(n22585), .ZN(n22729) );
  OA21D1BWP12T U13563 ( .A1(n22587), .A2(n23054), .B(n22729), .Z(n22617) );
  AOI32D1BWP12T U13564 ( .A1(n22590), .A2(a[13]), .A3(n22589), .B1(n22617), 
        .B2(n22588), .ZN(n22596) );
  FA1D0BWP12T U13565 ( .A(n22593), .B(n22592), .CI(n22591), .CO(n22548), .S(
        n23330) );
  AOI22D1BWP12T U13566 ( .A1(n23481), .A2(n22974), .B1(n23658), .B2(n23330), 
        .ZN(n22594) );
  OAI211D1BWP12T U13567 ( .A1(n23647), .A2(n23524), .B(n22594), .C(n22913), 
        .ZN(n22595) );
  AOI211D1BWP12T U13568 ( .A1(n23136), .A2(n23674), .B(n22596), .C(n22595), 
        .ZN(n22597) );
  OAI211D1BWP12T U13569 ( .A1(n23628), .A2(n23653), .B(n22598), .C(n22597), 
        .ZN(n22599) );
  AO211D1BWP12T U13570 ( .A1(n22945), .A2(n23104), .B(n22600), .C(n22599), .Z(
        result[13]) );
  AOI21D1BWP12T U13571 ( .A1(n22611), .A2(n22602), .B(n22601), .ZN(n23625) );
  OAI31D1BWP12T U13572 ( .A1(a[11]), .A2(n22634), .A3(n22701), .B(n23645), 
        .ZN(n22603) );
  AOI21D1BWP12T U13573 ( .A1(b[12]), .A2(n23652), .B(n22603), .ZN(n22604) );
  ND2D1BWP12T U13574 ( .A1(n23644), .A2(n23017), .ZN(n23028) );
  OAI22D1BWP12T U13575 ( .A1(n22604), .A2(n22689), .B1(n23250), .B2(n23028), 
        .ZN(n22623) );
  AOI22D1BWP12T U13576 ( .A1(b[0]), .A2(a[13]), .B1(a[12]), .B2(n22605), .ZN(
        n22724) );
  AOI22D1BWP12T U13577 ( .A1(b[0]), .A2(a[15]), .B1(a[14]), .B2(n22009), .ZN(
        n22725) );
  AOI222D1BWP12T U13578 ( .A1(n22608), .A2(b[2]), .B1(n22607), .B2(n22724), 
        .C1(n22725), .C2(n22606), .ZN(n22869) );
  INVD1BWP12T U13579 ( .I(n22869), .ZN(n23454) );
  MAOI22D0BWP12T U13580 ( .A1(n23258), .A2(n23454), .B1(n22727), .B2(n23416), 
        .ZN(n22619) );
  OAI21D1BWP12T U13581 ( .A1(n23221), .A2(n23017), .B(n22619), .ZN(n23233) );
  OAI22D1BWP12T U13582 ( .A1(n23041), .A2(n23233), .B1(n22609), .B2(n22737), 
        .ZN(n22622) );
  NR2D1BWP12T U13583 ( .A1(a[12]), .A2(n22612), .ZN(n22613) );
  AOI22D1BWP12T U13584 ( .A1(n23525), .A2(n22998), .B1(n22613), .B2(n22974), 
        .ZN(n22616) );
  AOI22D1BWP12T U13585 ( .A1(n23095), .A2(n23055), .B1(n23658), .B2(n23323), 
        .ZN(n22615) );
  OAI211D1BWP12T U13586 ( .A1(a[12]), .A2(n22617), .B(n22616), .C(n22615), 
        .ZN(n22618) );
  AOI31D1BWP12T U13587 ( .A1(n22619), .A2(n22674), .A3(n22844), .B(n22618), 
        .ZN(n22620) );
  OAI211D1BWP12T U13588 ( .A1(n23142), .A2(n22948), .B(n22620), .C(n22913), 
        .ZN(n22621) );
  NR3D1BWP12T U13589 ( .A1(n22623), .A2(n22622), .A3(n22621), .ZN(n22628) );
  OAI22D1BWP12T U13590 ( .A1(n23105), .A2(n23670), .B1(n22624), .B2(n23669), 
        .ZN(n22656) );
  NR2D1BWP12T U13591 ( .A1(n22645), .A2(n22626), .ZN(n23073) );
  AO22D1BWP12T U13592 ( .A1(n23105), .A2(n22945), .B1(n23027), .B2(n22624), 
        .Z(n22625) );
  AOI22D1BWP12T U13593 ( .A1(n22626), .A2(n22656), .B1(n23073), .B2(n22625), 
        .ZN(n22627) );
  OAI211D1BWP12T U13594 ( .A1(n23625), .A2(n23653), .B(n22628), .C(n22627), 
        .ZN(result[12]) );
  OA22D1BWP12T U13595 ( .A1(n22681), .A2(n23669), .B1(n22678), .B2(n23670), 
        .Z(n22659) );
  OR2XD1BWP12T U13596 ( .A1(n22655), .A2(n22629), .Z(n23075) );
  MAOI22D0BWP12T U13597 ( .A1(n22655), .A2(n22630), .B1(n22655), .B2(n22630), 
        .ZN(n23135) );
  FA1D0BWP12T U13598 ( .A(n22633), .B(n22632), .CI(n22631), .CO(n22614), .S(
        n23306) );
  IOA21D1BWP12T U13599 ( .A1(n22634), .A2(n23033), .B(n22729), .ZN(n22676) );
  AOI22D1BWP12T U13600 ( .A1(n23306), .A2(n23658), .B1(n22642), .B2(n22676), 
        .ZN(n22635) );
  OAI211D1BWP12T U13601 ( .A1(n22636), .A2(n22737), .B(n22635), .C(n22913), 
        .ZN(n22652) );
  ND2D1BWP12T U13602 ( .A1(n23661), .A2(n22986), .ZN(n22963) );
  INVD1BWP12T U13603 ( .I(n22963), .ZN(n22650) );
  ND2D1BWP12T U13604 ( .A1(b[4]), .A2(n22637), .ZN(n22764) );
  AOI31D1BWP12T U13605 ( .A1(a[14]), .A2(b[0]), .A3(b[1]), .B(n22638), .ZN(
        n22639) );
  OAI21D1BWP12T U13606 ( .A1(n22642), .A2(n22640), .B(n22639), .ZN(n22756) );
  AOI22D1BWP12T U13607 ( .A1(b[2]), .A2(n22754), .B1(n22756), .B2(n22342), 
        .ZN(n23453) );
  AOI22D1BWP12T U13608 ( .A1(n23463), .A2(n23270), .B1(n23258), .B2(n23453), 
        .ZN(n23209) );
  OAI21D1BWP12T U13609 ( .A1(n22764), .A2(n22641), .B(n23209), .ZN(n23385) );
  INVD1BWP12T U13610 ( .I(n23230), .ZN(n22647) );
  OAI32D1BWP12T U13611 ( .A1(n23343), .A2(n22642), .A3(n23022), .B1(n23499), 
        .B2(n23343), .ZN(n22643) );
  AOI211D1BWP12T U13612 ( .A1(n23652), .A2(n23343), .B(n22904), .C(n22643), 
        .ZN(n22644) );
  OAI22D1BWP12T U13613 ( .A1(n23290), .A2(n23028), .B1(n22645), .B2(n22644), 
        .ZN(n22646) );
  AOI31D1BWP12T U13614 ( .A1(n22647), .A2(n23209), .A3(n22964), .B(n22646), 
        .ZN(n22649) );
  ND4D1BWP12T U13615 ( .A1(a[11]), .A2(n22670), .A3(n22677), .A4(n22700), .ZN(
        n22648) );
  OAI211D1BWP12T U13616 ( .A1(n22650), .A2(n23385), .B(n22649), .C(n22648), 
        .ZN(n22651) );
  AOI211D1BWP12T U13617 ( .A1(n23135), .A2(n23674), .B(n22652), .C(n22651), 
        .ZN(n22658) );
  AOI21D1BWP12T U13618 ( .A1(n22655), .A2(n22654), .B(n22653), .ZN(n23632) );
  AOI21D1BWP12T U13619 ( .A1(n23632), .A2(n23601), .B(n22656), .ZN(n22657) );
  OAI211D1BWP12T U13620 ( .A1(n22659), .A2(n23075), .B(n22658), .C(n22657), 
        .ZN(result[11]) );
  INVD1BWP12T U13621 ( .I(n22660), .ZN(n22664) );
  ND2D1BWP12T U13622 ( .A1(a[10]), .A2(n22009), .ZN(n22661) );
  ND2D1BWP12T U13623 ( .A1(b[0]), .A2(a[11]), .ZN(n22722) );
  AOI32D1BWP12T U13624 ( .A1(n22661), .A2(n22485), .A3(n22722), .B1(n22724), 
        .B2(b[1]), .ZN(n22957) );
  AOI222D1BWP12T U13625 ( .A1(n22664), .A2(n23270), .B1(n22957), .B2(n22663), 
        .C1(n22958), .C2(n22662), .ZN(n23439) );
  OAI21D1BWP12T U13626 ( .A1(n22666), .A2(n22665), .B(n23439), .ZN(n23238) );
  INVD1BWP12T U13627 ( .I(n23041), .ZN(n22848) );
  OAI22D1BWP12T U13628 ( .A1(n23063), .A2(n22669), .B1(n22668), .B2(n22667), 
        .ZN(n23129) );
  INVD1BWP12T U13629 ( .I(n22913), .ZN(n23037) );
  NR2D1BWP12T U13630 ( .A1(a[10]), .A2(n22675), .ZN(n23480) );
  OAI21D1BWP12T U13631 ( .A1(n23063), .A2(n22680), .B(n22679), .ZN(n23631) );
  INVD1BWP12T U13632 ( .I(n22682), .ZN(n22716) );
  INR2D1BWP12T U13633 ( .A1(n22684), .B1(n22683), .ZN(n22685) );
  MAOI22D0BWP12T U13634 ( .A1(n22716), .A2(n22685), .B1(n22716), .B2(n22685), 
        .ZN(n23624) );
  INVD1BWP12T U13635 ( .I(n22686), .ZN(n22715) );
  ND2D1BWP12T U13636 ( .A1(a[9]), .A2(n22605), .ZN(n22688) );
  OAI222D1BWP12T U13637 ( .A1(n22993), .A2(n22689), .B1(n22688), .B2(n22843), 
        .C1(n22867), .C2(n22687), .ZN(n22846) );
  AOI22D1BWP12T U13638 ( .A1(b[2]), .A2(n22690), .B1(n22846), .B2(n22342), 
        .ZN(n22980) );
  OAI22D1BWP12T U13639 ( .A1(n22727), .A2(n22703), .B1(n22691), .B2(n22980), 
        .ZN(n23432) );
  AOI31D1BWP12T U13640 ( .A1(n22693), .A2(n23263), .A3(n22692), .B(n23432), 
        .ZN(n23240) );
  OAI22D1BWP12T U13641 ( .A1(n23282), .A2(n23028), .B1(n23240), .B2(n22809), 
        .ZN(n22710) );
  INVD1BWP12T U13642 ( .I(n22694), .ZN(n23064) );
  FA1D0BWP12T U13643 ( .A(n22697), .B(n22696), .CI(n22695), .CO(n22672), .S(
        n23329) );
  AOI22D1BWP12T U13644 ( .A1(n22716), .A2(n23650), .B1(n23658), .B2(n23329), 
        .ZN(n22698) );
  OAI211D1BWP12T U13645 ( .A1(n23064), .A2(n23645), .B(n22698), .C(n22913), 
        .ZN(n22709) );
  AOI22D1BWP12T U13646 ( .A1(b[9]), .A2(n23000), .B1(n23509), .B2(n22699), 
        .ZN(n22702) );
  AOI32D1BWP12T U13647 ( .A1(n22702), .A2(a[9]), .A3(n22701), .B1(n22729), 
        .B2(n22700), .ZN(n22708) );
  AOI22D1BWP12T U13648 ( .A1(n23270), .A2(n22703), .B1(n23258), .B2(n22980), 
        .ZN(n22704) );
  OAI211D1BWP12T U13649 ( .A1(n22705), .A2(n22764), .B(n23397), .C(n22704), 
        .ZN(n23583) );
  OAI22D1BWP12T U13650 ( .A1(n23427), .A2(n22737), .B1(n22706), .B2(n23583), 
        .ZN(n22707) );
  OR4XD1BWP12T U13651 ( .A1(n22710), .A2(n22709), .A3(n22708), .A4(n22707), 
        .Z(n22714) );
  MAOI22D0BWP12T U13652 ( .A1(n22716), .A2(n22711), .B1(n22716), .B2(n22711), 
        .ZN(n23132) );
  OAI22D1BWP12T U13653 ( .A1(n23132), .A2(n22948), .B1(n22712), .B2(n23670), 
        .ZN(n22713) );
  AOI211D1BWP12T U13654 ( .A1(n22715), .A2(n23027), .B(n22714), .C(n22713), 
        .ZN(n22718) );
  NR2D1BWP12T U13655 ( .A1(n22740), .A2(n22716), .ZN(n23080) );
  OAI22D1BWP12T U13656 ( .A1(n22742), .A2(n23670), .B1(n22743), .B2(n23669), 
        .ZN(n22749) );
  AOI32D1BWP12T U13657 ( .A1(n23122), .A2(n23080), .A3(n23055), .B1(n22749), 
        .B2(n23080), .ZN(n22717) );
  OAI211D1BWP12T U13658 ( .A1(n23624), .A2(n23653), .B(n22718), .C(n22717), 
        .ZN(result[9]) );
  AOI21D1BWP12T U13659 ( .A1(n23122), .A2(n22720), .B(n22719), .ZN(n23623) );
  AOI32D1BWP12T U13660 ( .A1(n22867), .A2(n22723), .A3(n22722), .B1(n22721), 
        .B2(n22864), .ZN(n22868) );
  INVD1BWP12T U13661 ( .I(n22868), .ZN(n22726) );
  AOI222D1BWP12T U13662 ( .A1(n22726), .A2(n22342), .B1(n22725), .B2(n22951), 
        .C1(n23259), .C2(n22724), .ZN(n23010) );
  IND2D1BWP12T U13663 ( .A1(n23010), .B1(n23258), .ZN(n22735) );
  OAI21D1BWP12T U13664 ( .A1(n22727), .A2(n23455), .B(n22735), .ZN(n23210) );
  INR2D1BWP12T U13665 ( .A1(n22764), .B1(n23210), .ZN(n23390) );
  OAI32D1BWP12T U13666 ( .A1(n22729), .A2(n22728), .A3(n22856), .B1(a[8]), 
        .B2(n22729), .ZN(n22734) );
  INVD1BWP12T U13667 ( .I(n23280), .ZN(n22732) );
  MAOI22D0BWP12T U13668 ( .A1(n23328), .A2(n23658), .B1(n23645), .B2(n22740), 
        .ZN(n22731) );
  OAI211D1BWP12T U13669 ( .A1(n22732), .A2(n23028), .B(n22731), .C(n22913), 
        .ZN(n22733) );
  AOI211D1BWP12T U13670 ( .A1(n23390), .A2(n22963), .B(n22734), .C(n22733), 
        .ZN(n22752) );
  ND2D1BWP12T U13671 ( .A1(n22736), .A2(n22735), .ZN(n23387) );
  OAI22D1BWP12T U13672 ( .A1(n23425), .A2(n22737), .B1(n23041), .B2(n23387), 
        .ZN(n22750) );
  NR2D1BWP12T U13673 ( .A1(n23652), .A2(n23344), .ZN(n22739) );
  OAI22D1BWP12T U13674 ( .A1(n22740), .A2(n22739), .B1(n22948), .B2(n22738), 
        .ZN(n22748) );
  AOI211D1BWP12T U13675 ( .A1(n23509), .A2(n22741), .B(n23650), .C(n23122), 
        .ZN(n22745) );
  AOI22D1BWP12T U13676 ( .A1(n23027), .A2(n22743), .B1(n22945), .B2(n22742), 
        .ZN(n22744) );
  OAI211D1BWP12T U13677 ( .A1(n22746), .A2(n22948), .B(n22745), .C(n22744), 
        .ZN(n22747) );
  OAI32D1BWP12T U13678 ( .A1(n22750), .A2(n22749), .A3(n22748), .B1(n22747), 
        .B2(n22750), .ZN(n22751) );
  OAI211D1BWP12T U13679 ( .A1(n23623), .A2(n23653), .B(n22752), .C(n22751), 
        .ZN(result[8]) );
  MAOI22D0BWP12T U13680 ( .A1(n22753), .A2(n22782), .B1(n22753), .B2(n22782), 
        .ZN(n23134) );
  OA221D1BWP12T U13681 ( .A1(n22342), .A2(n22755), .B1(b[2]), .B2(n22754), .C(
        b[3]), .Z(n22763) );
  INVD1BWP12T U13682 ( .I(n22756), .ZN(n22761) );
  INVD1BWP12T U13683 ( .I(n23008), .ZN(n22982) );
  AOI22D1BWP12T U13684 ( .A1(a[10]), .A2(n22842), .B1(a[7]), .B2(n22757), .ZN(
        n22758) );
  IND2D1BWP12T U13685 ( .A1(n22759), .B1(n22758), .ZN(n22924) );
  ND2D1BWP12T U13686 ( .A1(n22920), .A2(n22924), .ZN(n22760) );
  OAI211D1BWP12T U13687 ( .A1(n22761), .A2(n22982), .B(n23017), .C(n22760), 
        .ZN(n22762) );
  OAI22D1BWP12T U13688 ( .A1(n22765), .A2(n22764), .B1(n22763), .B2(n22762), 
        .ZN(n23386) );
  AOI211D1BWP12T U13689 ( .A1(n22766), .A2(n22986), .B(n23041), .C(n23386), 
        .ZN(n22781) );
  MAOI22D0BWP12T U13690 ( .A1(n22768), .A2(n22767), .B1(n22888), .B2(n23433), 
        .ZN(n22779) );
  FA1D0BWP12T U13691 ( .A(n22771), .B(n22770), .CI(n22769), .CO(n22730), .S(
        n23327) );
  INVD1BWP12T U13692 ( .I(n22772), .ZN(n23068) );
  AOI211D1BWP12T U13693 ( .A1(a[7]), .A2(n23645), .B(n23068), .C(n22907), .ZN(
        n22774) );
  OAI22D1BWP12T U13694 ( .A1(n23647), .A2(n23471), .B1(n23345), .B2(n23372), 
        .ZN(n22773) );
  AOI211D1BWP12T U13695 ( .A1(n23327), .A2(n23658), .B(n22774), .C(n22773), 
        .ZN(n22778) );
  INVD1BWP12T U13696 ( .I(n22887), .ZN(n23005) );
  AOI21D1BWP12T U13697 ( .A1(n22775), .A2(n22857), .B(n22858), .ZN(n22814) );
  AOI22D1BWP12T U13698 ( .A1(n23005), .A2(n23266), .B1(n22814), .B2(n22776), 
        .ZN(n22777) );
  ND4D1BWP12T U13699 ( .A1(n22779), .A2(n22778), .A3(n22777), .A4(n22913), 
        .ZN(n22780) );
  AOI211D1BWP12T U13700 ( .A1(n23674), .A2(n23134), .B(n22781), .C(n22780), 
        .ZN(n22793) );
  NR2D1BWP12T U13701 ( .A1(n22783), .A2(n22782), .ZN(n23081) );
  OAI22D1BWP12T U13702 ( .A1(n22784), .A2(n23669), .B1(n22795), .B2(n23670), 
        .ZN(n22791) );
  INR2D1BWP12T U13703 ( .A1(n22786), .B1(n22785), .ZN(n22788) );
  MOAI22D0BWP12T U13704 ( .A1(n22788), .A2(n22787), .B1(n22788), .B2(n22787), 
        .ZN(n23617) );
  OAI22D1BWP12T U13705 ( .A1(n23617), .A2(n23653), .B1(n22789), .B2(n23670), 
        .ZN(n22790) );
  AOI21D1BWP12T U13706 ( .A1(n23081), .A2(n22791), .B(n22790), .ZN(n22792) );
  OAI211D1BWP12T U13707 ( .A1(n22794), .A2(n23669), .B(n22793), .C(n22792), 
        .ZN(result[7]) );
  AOI21D1BWP12T U13708 ( .A1(n22796), .A2(n23088), .B(n22795), .ZN(n22827) );
  AOI21D1BWP12T U13709 ( .A1(n22823), .A2(n22798), .B(n22797), .ZN(n23620) );
  FA1D0BWP12T U13710 ( .A(n22801), .B(n22800), .CI(n22799), .CO(n22769), .S(
        n23308) );
  AOI22D1BWP12T U13711 ( .A1(n23658), .A2(n23308), .B1(n23005), .B2(n23271), 
        .ZN(n22802) );
  OAI211D1BWP12T U13712 ( .A1(n22907), .A2(n23482), .B(n22802), .C(n22913), 
        .ZN(n22820) );
  ND2D1BWP12T U13713 ( .A1(a[6]), .A2(n22605), .ZN(n22804) );
  AOI22D1BWP12T U13714 ( .A1(b[0]), .A2(a[9]), .B1(a[8]), .B2(n22605), .ZN(
        n22803) );
  AOI32D1BWP12T U13715 ( .A1(n22804), .A2(n22485), .A3(n22866), .B1(n22803), 
        .B2(b[1]), .ZN(n22961) );
  AOI22D1BWP12T U13716 ( .A1(n22920), .A2(n22961), .B1(n23008), .B2(n22957), 
        .ZN(n22805) );
  OAI211D1BWP12T U13717 ( .A1(n22807), .A2(n22806), .B(n22805), .C(n23017), 
        .ZN(n23207) );
  OAI21D1BWP12T U13718 ( .A1(n23017), .A2(n22808), .B(n23207), .ZN(n23393) );
  AOI21D1BWP12T U13719 ( .A1(n22810), .A2(b[4]), .B(n22809), .ZN(n22811) );
  AOI22D1BWP12T U13720 ( .A1(n22834), .A2(n23457), .B1(n22811), .B2(n23207), 
        .ZN(n22818) );
  AOI22D1BWP12T U13721 ( .A1(a[6]), .A2(n23030), .B1(n22813), .B2(n22812), 
        .ZN(n22816) );
  OAI22D1BWP12T U13722 ( .A1(a[5]), .A2(n22856), .B1(b[6]), .B2(n23647), .ZN(
        n22815) );
  OAI22D1BWP12T U13723 ( .A1(n22816), .A2(n22815), .B1(a[6]), .B2(n22814), 
        .ZN(n22817) );
  OAI211D1BWP12T U13724 ( .A1(n22986), .A2(n23393), .B(n22818), .C(n22817), 
        .ZN(n22819) );
  AOI211D1BWP12T U13725 ( .A1(n23620), .A2(n23601), .B(n22820), .C(n22819), 
        .ZN(n22826) );
  OAI31D1BWP12T U13726 ( .A1(n22822), .A2(n22823), .A3(n22853), .B(n22821), 
        .ZN(n23195) );
  MAOI22D0BWP12T U13727 ( .A1(n22824), .A2(n22823), .B1(n22824), .B2(n22823), 
        .ZN(n23126) );
  AOI22D1BWP12T U13728 ( .A1(n23027), .A2(n23195), .B1(n23674), .B2(n23126), 
        .ZN(n22825) );
  OAI211D1BWP12T U13729 ( .A1(n22827), .A2(n23670), .B(n22826), .C(n22825), 
        .ZN(result[6]) );
  NR2D1BWP12T U13730 ( .A1(n22828), .A2(n22832), .ZN(n23082) );
  INR2D1BWP12T U13731 ( .A1(n22830), .B1(n22829), .ZN(n22831) );
  MAOI22D0BWP12T U13732 ( .A1(n22832), .A2(n22831), .B1(n22832), .B2(n22831), 
        .ZN(n23616) );
  MOAI22D0BWP12T U13733 ( .A1(n23616), .A2(n23653), .B1(n22834), .B2(n22833), 
        .ZN(n22835) );
  AOI31D1BWP12T U13734 ( .A1(n23082), .A2(n22836), .A3(n23055), .B(n22835), 
        .ZN(n22863) );
  MAOI22D0BWP12T U13735 ( .A1(n23165), .A2(n22837), .B1(n23165), .B2(n22837), 
        .ZN(n23127) );
  AOI22D1BWP12T U13736 ( .A1(n22838), .A2(n22945), .B1(n23127), .B2(n23674), 
        .ZN(n22852) );
  FA1D0BWP12T U13737 ( .A(n22841), .B(n22840), .CI(n22839), .CO(n22800), .S(
        n23307) );
  AOI22D1BWP12T U13738 ( .A1(n23494), .A2(n22974), .B1(n23658), .B2(n23307), 
        .ZN(n22851) );
  OAI22D1BWP12T U13739 ( .A1(n22009), .A2(n23369), .B1(n21803), .B2(b[0]), 
        .ZN(n22921) );
  AOI222D1BWP12T U13740 ( .A1(n22485), .A2(n22921), .B1(a[7]), .B2(n22843), 
        .C1(a[8]), .C2(n22842), .ZN(n22981) );
  OAI22D1BWP12T U13741 ( .A1(n22981), .A2(n22844), .B1(n22806), .B2(n23417), 
        .ZN(n22845) );
  AOI211D1BWP12T U13742 ( .A1(n23008), .A2(n22846), .B(b[4]), .C(n22845), .ZN(
        n23236) );
  NR2D1BWP12T U13743 ( .A1(n23017), .A2(n23408), .ZN(n23235) );
  OAI32D1BWP12T U13744 ( .A1(n23236), .A2(n22847), .A3(n22986), .B1(n23235), 
        .B2(n23236), .ZN(n22849) );
  AOI22D1BWP12T U13745 ( .A1(n23279), .A2(n23005), .B1(n22849), .B2(n22848), 
        .ZN(n22850) );
  AN4XD1BWP12T U13746 ( .A1(n22852), .A2(n22851), .A3(n22850), .A4(n22913), 
        .Z(n22862) );
  AOI32D1BWP12T U13747 ( .A1(n23082), .A2(n23027), .A3(n22885), .B1(n22853), 
        .B2(n23027), .ZN(n22861) );
  OAI22D1BWP12T U13748 ( .A1(n23652), .A2(n23346), .B1(n22854), .B2(n22998), 
        .ZN(n22855) );
  ND2D1BWP12T U13749 ( .A1(n22856), .A2(n22855), .ZN(n22859) );
  NR2D1BWP12T U13750 ( .A1(n22858), .A2(n22857), .ZN(n22872) );
  OAI22D1BWP12T U13751 ( .A1(n22904), .A2(n22859), .B1(a[5]), .B2(n22872), 
        .ZN(n22860) );
  ND4D1BWP12T U13752 ( .A1(n22863), .A2(n22862), .A3(n22861), .A4(n22860), 
        .ZN(result[5]) );
  ND2D1BWP12T U13753 ( .A1(b[4]), .A2(n23211), .ZN(n22890) );
  ND2D1BWP12T U13754 ( .A1(a[4]), .A2(n22009), .ZN(n22952) );
  AOI32D1BWP12T U13755 ( .A1(n22952), .A2(n22867), .A3(n22866), .B1(n22865), 
        .B2(n22864), .ZN(n23009) );
  AOI222D1BWP12T U13756 ( .A1(b[3]), .A2(n22869), .B1(n22920), .B2(n23009), 
        .C1(n23008), .C2(n22868), .ZN(n23220) );
  ND2D1BWP12T U13757 ( .A1(n23220), .A2(n23017), .ZN(n22891) );
  OAI21D1BWP12T U13758 ( .A1(n22870), .A2(n22890), .B(n22891), .ZN(n23394) );
  MOAI22D0BWP12T U13759 ( .A1(n22882), .A2(n22871), .B1(n22882), .B2(n22871), 
        .ZN(n23103) );
  AOI22D1BWP12T U13760 ( .A1(n23477), .A2(n22998), .B1(n23497), .B2(n22974), 
        .ZN(n22878) );
  OAI21D1BWP12T U13761 ( .A1(n22874), .A2(n22873), .B(n22872), .ZN(n22877) );
  OAI211D1BWP12T U13762 ( .A1(b[4]), .A2(op[2]), .B(a[4]), .C(n23000), .ZN(
        n22876) );
  ND2D1BWP12T U13763 ( .A1(n23658), .A2(n23305), .ZN(n22875) );
  ND4D1BWP12T U13764 ( .A1(n22878), .A2(n22877), .A3(n22876), .A4(n22875), 
        .ZN(n22884) );
  AOI21D1BWP12T U13765 ( .A1(n22886), .A2(n22880), .B(n22879), .ZN(n23609) );
  MAOI22D0BWP12T U13766 ( .A1(n22882), .A2(n22881), .B1(n22882), .B2(n22881), 
        .ZN(n23130) );
  OAI22D1BWP12T U13767 ( .A1(n23609), .A2(n23653), .B1(n23130), .B2(n22948), 
        .ZN(n22883) );
  AOI211D1BWP12T U13768 ( .A1(n22945), .A2(n23103), .B(n22884), .C(n22883), 
        .ZN(n22894) );
  MAOI22D0BWP12T U13769 ( .A1(n22886), .A2(n22885), .B1(n22886), .B2(n22885), 
        .ZN(n23193) );
  OAI22D1BWP12T U13770 ( .A1(n23424), .A2(n22888), .B1(n23278), .B2(n22887), 
        .ZN(n22889) );
  AOI31D1BWP12T U13771 ( .A1(n22891), .A2(n22890), .A3(n22964), .B(n22889), 
        .ZN(n22892) );
  OA211D1BWP12T U13772 ( .A1(n23193), .A2(n23669), .B(n22892), .C(n22913), .Z(
        n22893) );
  OAI211D1BWP12T U13773 ( .A1(n23394), .A2(n22986), .B(n22894), .C(n22893), 
        .ZN(result[4]) );
  MAOI22D0BWP12T U13774 ( .A1(n22901), .A2(n22895), .B1(n22901), .B2(n22895), 
        .ZN(n23190) );
  MAOI22D0BWP12T U13775 ( .A1(n22897), .A2(n22896), .B1(n22897), .B2(n22896), 
        .ZN(n23338) );
  NR2D1BWP12T U13776 ( .A1(n22899), .A2(n22898), .ZN(n22900) );
  MAOI22D0BWP12T U13777 ( .A1(n22901), .A2(n22900), .B1(n22901), .B2(n22900), 
        .ZN(n23605) );
  NR2D1BWP12T U13778 ( .A1(n22926), .A2(n22987), .ZN(n22934) );
  AOI22D1BWP12T U13779 ( .A1(n23605), .A2(n23601), .B1(n22902), .B2(n22934), 
        .ZN(n22915) );
  MAOI22D0BWP12T U13780 ( .A1(n22917), .A2(n22903), .B1(n22917), .B2(n22903), 
        .ZN(n23123) );
  OAI22D1BWP12T U13781 ( .A1(n23123), .A2(n22948), .B1(n23647), .B2(n23515), 
        .ZN(n22909) );
  OAI22D1BWP12T U13782 ( .A1(a[3]), .A2(n22905), .B1(n22904), .B2(n23515), 
        .ZN(n22906) );
  OAI21D1BWP12T U13783 ( .A1(n22907), .A2(n22806), .B(n22906), .ZN(n22908) );
  OAI32D1BWP12T U13784 ( .A1(n22909), .A2(n23000), .A3(n22911), .B1(n22908), 
        .B2(n22909), .ZN(n22914) );
  OAI211D1BWP12T U13785 ( .A1(n22942), .A2(n22911), .B(n23033), .C(n22910), 
        .ZN(n22912) );
  ND4D1BWP12T U13786 ( .A1(n22915), .A2(n22914), .A3(n22913), .A4(n22912), 
        .ZN(n22919) );
  MAOI22D0BWP12T U13787 ( .A1(n22917), .A2(n22916), .B1(n22917), .B2(n22916), 
        .ZN(n23097) );
  OAI22D1BWP12T U13788 ( .A1(n23097), .A2(n23670), .B1(n23274), .B2(n23028), 
        .ZN(n22918) );
  AOI211D1BWP12T U13789 ( .A1(n23338), .A2(n23658), .B(n22919), .C(n22918), 
        .ZN(n22928) );
  ND2D1BWP12T U13790 ( .A1(b[4]), .A2(n23212), .ZN(n23229) );
  AOI22D1BWP12T U13791 ( .A1(b[0]), .A2(a[4]), .B1(a[3]), .B2(n22605), .ZN(
        n22984) );
  OAI21D1BWP12T U13792 ( .A1(n23012), .A2(n22984), .B(n23017), .ZN(n22923) );
  ND2D1BWP12T U13793 ( .A1(b[1]), .A2(n22920), .ZN(n23015) );
  INVD1BWP12T U13794 ( .I(n23015), .ZN(n22953) );
  MOAI22D0BWP12T U13795 ( .A1(n22806), .A2(n23453), .B1(n22953), .B2(n22921), 
        .ZN(n22922) );
  AOI211D1BWP12T U13796 ( .A1(n23008), .A2(n22924), .B(n22923), .C(n22922), 
        .ZN(n23217) );
  INR2D1BWP12T U13797 ( .A1(n23229), .B1(n23217), .ZN(n23392) );
  AOI32D1BWP12T U13798 ( .A1(n22964), .A2(n23392), .A3(n22926), .B1(n22925), 
        .B2(n23392), .ZN(n22927) );
  OAI211D1BWP12T U13799 ( .A1(n23669), .A2(n23190), .B(n22928), .C(n22927), 
        .ZN(result[3]) );
  MAOI22D0BWP12T U13800 ( .A1(n22937), .A2(n22929), .B1(n22937), .B2(n22929), 
        .ZN(n23189) );
  AOI22D1BWP12T U13801 ( .A1(n23189), .A2(n23027), .B1(n23281), .B2(n23005), 
        .ZN(n22968) );
  MAOI22D0BWP12T U13802 ( .A1(n22931), .A2(n22930), .B1(n22931), .B2(n22930), 
        .ZN(n23380) );
  MAOI22D0BWP12T U13803 ( .A1(n22937), .A2(n22932), .B1(n22937), .B2(n22932), 
        .ZN(n23124) );
  OAI21D1BWP12T U13804 ( .A1(n23372), .A2(n22342), .B(n23645), .ZN(n22935) );
  AOI22D1BWP12T U13805 ( .A1(a[2]), .A2(n22935), .B1(n22934), .B2(n22933), 
        .ZN(n22947) );
  MAOI22D0BWP12T U13806 ( .A1(n22937), .A2(n22936), .B1(n22937), .B2(n22936), 
        .ZN(n23094) );
  FA1D0BWP12T U13807 ( .A(b[1]), .B(n22938), .CI(n22937), .CO(n20753), .S(
        n23600) );
  OAI22D1BWP12T U13808 ( .A1(a[2]), .A2(n23558), .B1(n23600), .B2(n23653), 
        .ZN(n22944) );
  AOI22D1BWP12T U13809 ( .A1(n23495), .A2(n22974), .B1(n22939), .B2(n22998), 
        .ZN(n22940) );
  OAI31D1BWP12T U13810 ( .A1(n22942), .A2(n22941), .A3(n23054), .B(n22940), 
        .ZN(n22943) );
  AOI211D1BWP12T U13811 ( .A1(n23094), .A2(n22945), .B(n22944), .C(n22943), 
        .ZN(n22946) );
  OAI211D1BWP12T U13812 ( .A1(n23124), .A2(n22948), .B(n22947), .C(n22946), 
        .ZN(n22949) );
  AOI211D1BWP12T U13813 ( .A1(n23658), .A2(n23380), .B(n23037), .C(n22949), 
        .ZN(n22967) );
  AOI31D1BWP12T U13814 ( .A1(n22951), .A2(a[31]), .A3(n22950), .B(n22965), 
        .ZN(n22962) );
  AOI22D1BWP12T U13815 ( .A1(b[0]), .A2(a[3]), .B1(a[2]), .B2(n22009), .ZN(
        n23016) );
  INVD1BWP12T U13816 ( .I(n22952), .ZN(n22954) );
  OAI21D1BWP12T U13817 ( .A1(n22955), .A2(n22954), .B(n22953), .ZN(n22956) );
  OAI211D1BWP12T U13818 ( .A1(n23016), .A2(n23012), .B(n23017), .C(n22956), 
        .ZN(n22960) );
  OA221D1BWP12T U13819 ( .A1(n22342), .A2(n22958), .B1(b[2]), .B2(n22957), .C(
        b[3]), .Z(n22959) );
  AOI211D1BWP12T U13820 ( .A1(n23008), .A2(n22961), .B(n22960), .C(n22959), 
        .ZN(n23219) );
  AOI21D1BWP12T U13821 ( .A1(b[4]), .A2(n22962), .B(n23219), .ZN(n23400) );
  AOI32D1BWP12T U13822 ( .A1(n22965), .A2(n23400), .A3(n22964), .B1(n22963), 
        .B2(n23400), .ZN(n22966) );
  ND3D1BWP12T U13823 ( .A1(n22968), .A2(n22967), .A3(n22966), .ZN(result[2])
         );
  MOAI22D0BWP12T U13824 ( .A1(n22971), .A2(n22969), .B1(n22971), .B2(n22969), 
        .ZN(n23606) );
  MOAI22D0BWP12T U13825 ( .A1(n22971), .A2(n22970), .B1(n22971), .B2(n22970), 
        .ZN(n23188) );
  AOI22D1BWP12T U13826 ( .A1(n22973), .A2(n22990), .B1(n22972), .B2(n23472), 
        .ZN(n23128) );
  AOI22D1BWP12T U13827 ( .A1(n22975), .A2(n22974), .B1(n23128), .B2(n23674), 
        .ZN(n22976) );
  OAI31D1BWP12T U13828 ( .A1(n22978), .A2(n22977), .A3(n23054), .B(n22976), 
        .ZN(n22979) );
  AOI211D1BWP12T U13829 ( .A1(n23027), .A2(n23188), .B(n23037), .C(n22979), 
        .ZN(n23007) );
  NR2D1BWP12T U13830 ( .A1(n22806), .A2(n22980), .ZN(n23459) );
  AOI22D1BWP12T U13831 ( .A1(b[0]), .A2(a[2]), .B1(a[1]), .B2(n22009), .ZN(
        n22983) );
  OAI222D1BWP12T U13832 ( .A1(n22984), .A2(n23015), .B1(n23012), .B2(n22983), 
        .C1(n22982), .C2(n22981), .ZN(n23415) );
  OAI32D1BWP12T U13833 ( .A1(b[4]), .A2(n23459), .A3(n23415), .B1(n22985), 
        .B2(n23017), .ZN(n23234) );
  AOI211D1BWP12T U13834 ( .A1(n23442), .A2(n22986), .B(n23041), .C(n23234), 
        .ZN(n23004) );
  NR3D1BWP12T U13835 ( .A1(n23423), .A2(n22988), .A3(n22987), .ZN(n22997) );
  OAI21D1BWP12T U13836 ( .A1(n22991), .A2(n22990), .B(n22989), .ZN(n23090) );
  OAI22D1BWP12T U13837 ( .A1(n22993), .A2(n23559), .B1(n23262), .B2(n22992), 
        .ZN(n22994) );
  NR2D1BWP12T U13838 ( .A1(n22995), .A2(n22994), .ZN(n23339) );
  MOAI22D0BWP12T U13839 ( .A1(n23670), .A2(n23090), .B1(n23339), .B2(n23658), 
        .ZN(n22996) );
  AOI211D1BWP12T U13840 ( .A1(n22999), .A2(n22998), .B(n22997), .C(n22996), 
        .ZN(n23002) );
  OAI211D1BWP12T U13841 ( .A1(b[1]), .A2(op[2]), .B(a[1]), .C(n23000), .ZN(
        n23001) );
  OAI211D1BWP12T U13842 ( .A1(a[1]), .A2(n23558), .B(n23002), .C(n23001), .ZN(
        n23003) );
  AOI211D1BWP12T U13843 ( .A1(n23005), .A2(n23272), .B(n23004), .C(n23003), 
        .ZN(n23006) );
  OAI211D1BWP12T U13844 ( .A1(n23606), .A2(n23653), .B(n23007), .C(n23006), 
        .ZN(result[1]) );
  AOI22D1BWP12T U13845 ( .A1(b[3]), .A2(n23010), .B1(n23009), .B2(n23008), 
        .ZN(n23014) );
  OR3XD1BWP12T U13846 ( .A1(n23012), .A2(n22605), .A3(n23011), .Z(n23013) );
  OAI211D1BWP12T U13847 ( .A1(n23016), .A2(n23015), .B(n23014), .C(n23013), 
        .ZN(n23019) );
  OAI32D1BWP12T U13848 ( .A1(b[4]), .A2(n23273), .A3(n23019), .B1(n23018), 
        .B2(n23017), .ZN(n23215) );
  MAOI22D0BWP12T U13849 ( .A1(n23025), .A2(c_in), .B1(n23025), .B2(c_in), .ZN(
        n23171) );
  INVD1BWP12T U13850 ( .I(n23171), .ZN(n23608) );
  OAI22D1BWP12T U13851 ( .A1(n23034), .A2(n23022), .B1(n23021), .B2(n23020), 
        .ZN(n23023) );
  NR2D1BWP12T U13852 ( .A1(n23650), .A2(n23023), .ZN(n23024) );
  OAI22D1BWP12T U13853 ( .A1(n23025), .A2(n23024), .B1(n22605), .B2(n23645), 
        .ZN(n23026) );
  AOI221D1BWP12T U13854 ( .A1(n23027), .A2(n23608), .B1(n23601), .B2(n23171), 
        .C(n23026), .ZN(n23040) );
  INVD1BWP12T U13855 ( .I(n23028), .ZN(n23038) );
  AOI31D1BWP12T U13856 ( .A1(a[0]), .A2(n23031), .A3(n23030), .B(n23029), .ZN(
        n23032) );
  NR2D1BWP12T U13857 ( .A1(n23033), .A2(n23032), .ZN(n23035) );
  AOI22D1BWP12T U13858 ( .A1(n23035), .A2(n23645), .B1(n23034), .B2(n23558), 
        .ZN(n23036) );
  AOI211D1BWP12T U13859 ( .A1(n23273), .A2(n23038), .B(n23037), .C(n23036), 
        .ZN(n23039) );
  OAI211D1BWP12T U13860 ( .A1(n23041), .A2(n23215), .B(n23040), .C(n23039), 
        .ZN(result[0]) );
  NR2D1BWP12T U13861 ( .A1(b[31]), .A2(a[31]), .ZN(n23656) );
  NR2D1BWP12T U13862 ( .A1(n23043), .A2(n23642), .ZN(n23651) );
  NR2D1BWP12T U13863 ( .A1(n23656), .A2(n23651), .ZN(n23594) );
  INVD1BWP12T U13864 ( .I(n23594), .ZN(n23488) );
  INR3D0BWP12T U13865 ( .A1(n23206), .B1(n23656), .B2(n23669), .ZN(n23060) );
  NR2D1BWP12T U13866 ( .A1(n23047), .A2(n23046), .ZN(n23548) );
  INR2D1BWP12T U13867 ( .A1(n23049), .B1(n23048), .ZN(n23546) );
  ND4D1BWP12T U13868 ( .A1(n23052), .A2(n23546), .A3(n23051), .A4(n23050), 
        .ZN(n23053) );
  INR2D1BWP12T U13869 ( .A1(n23548), .B1(n23053), .ZN(n23569) );
  NR2D1BWP12T U13870 ( .A1(a[31]), .A2(n23054), .ZN(n23659) );
  INVD1BWP12T U13871 ( .I(n23659), .ZN(n23056) );
  MOAI22D0BWP12T U13872 ( .A1(n23569), .A2(n23056), .B1(n23055), .B2(n23651), 
        .ZN(n23057) );
  NR4D0BWP12T U13873 ( .A1(n23060), .A2(n23059), .A3(n23058), .A4(n23057), 
        .ZN(n23061) );
  OAI31D1BWP12T U13874 ( .A1(n23062), .A2(n23488), .A3(n23670), .B(n23061), 
        .ZN(c_out) );
  MOAI22D0BWP12T U13875 ( .A1(n23594), .A2(n23062), .B1(n23594), .B2(n23062), 
        .ZN(n23671) );
  OAI22D1BWP12T U13876 ( .A1(n23066), .A2(n23065), .B1(n23064), .B2(n23063), 
        .ZN(n23072) );
  OAI22D1BWP12T U13877 ( .A1(n23070), .A2(n23069), .B1(n23068), .B2(n23067), 
        .ZN(n23071) );
  INR4D0BWP12T U13878 ( .A1(n23074), .B1(n23073), .B2(n23072), .B3(n23071), 
        .ZN(n23076) );
  OAI211D1BWP12T U13879 ( .A1(n23078), .A2(n23077), .B(n23076), .C(n23075), 
        .ZN(n23079) );
  NR4D0BWP12T U13880 ( .A1(n23082), .A2(n23081), .A3(n23080), .A4(n23079), 
        .ZN(n23172) );
  AOI22D1BWP12T U13881 ( .A1(n23086), .A2(n23085), .B1(n23084), .B2(n23083), 
        .ZN(n23091) );
  ND2D1BWP12T U13882 ( .A1(n23088), .A2(n23087), .ZN(n23089) );
  ND4D1BWP12T U13883 ( .A1(n23172), .A2(n23091), .A3(n23090), .A4(n23089), 
        .ZN(n23102) );
  NR2D1BWP12T U13884 ( .A1(n23093), .A2(n23092), .ZN(n23096) );
  NR4D0BWP12T U13885 ( .A1(n23096), .A2(n23095), .A3(n23094), .A4(n23670), 
        .ZN(n23098) );
  OAI211D1BWP12T U13886 ( .A1(n23100), .A2(n23099), .B(n23098), .C(n23097), 
        .ZN(n23101) );
  NR4D0BWP12T U13887 ( .A1(n23104), .A2(n23103), .A3(n23102), .A4(n23101), 
        .ZN(n23106) );
  ND4D1BWP12T U13888 ( .A1(n23108), .A2(n23107), .A3(n23106), .A4(n23105), 
        .ZN(n23109) );
  INR4D0BWP12T U13889 ( .A1(n23112), .B1(n23111), .B2(n23110), .B3(n23109), 
        .ZN(n23113) );
  ND4D1BWP12T U13890 ( .A1(n23116), .A2(n23115), .A3(n23114), .A4(n23113), 
        .ZN(n23117) );
  NR4D0BWP12T U13891 ( .A1(n23120), .A2(n23119), .A3(n23118), .A4(n23117), 
        .ZN(n23163) );
  MAOI22D0BWP12T U13892 ( .A1(n23594), .A2(n23121), .B1(n23594), .B2(n23121), 
        .ZN(n23673) );
  ND4D1BWP12T U13893 ( .A1(n23124), .A2(n23123), .A3(n23674), .A4(n23122), 
        .ZN(n23125) );
  NR4D0BWP12T U13894 ( .A1(n23128), .A2(n23127), .A3(n23126), .A4(n23125), 
        .ZN(n23131) );
  ND4D1BWP12T U13895 ( .A1(n23132), .A2(n23131), .A3(n23130), .A4(n23129), 
        .ZN(n23133) );
  NR4D0BWP12T U13896 ( .A1(n23136), .A2(n23135), .A3(n23134), .A4(n23133), 
        .ZN(n23141) );
  NR2D1BWP12T U13897 ( .A1(n23138), .A2(n23137), .ZN(n23140) );
  ND4D1BWP12T U13898 ( .A1(n23142), .A2(n23141), .A3(n23140), .A4(n23139), 
        .ZN(n23143) );
  NR4D0BWP12T U13899 ( .A1(n23146), .A2(n23145), .A3(n23144), .A4(n23143), 
        .ZN(n23148) );
  ND4D1BWP12T U13900 ( .A1(n23150), .A2(n23149), .A3(n23148), .A4(n23147), 
        .ZN(n23151) );
  NR4D0BWP12T U13901 ( .A1(n23154), .A2(n23153), .A3(n23152), .A4(n23151), 
        .ZN(n23157) );
  ND4D1BWP12T U13902 ( .A1(n23158), .A2(n23157), .A3(n23156), .A4(n23155), 
        .ZN(n23159) );
  NR4D0BWP12T U13903 ( .A1(n23161), .A2(n23160), .A3(n23673), .A4(n23159), 
        .ZN(n23162) );
  AOI31D1BWP12T U13904 ( .A1(n23164), .A2(n23671), .A3(n23163), .B(n23162), 
        .ZN(n23640) );
  NR2D1BWP12T U13905 ( .A1(n23166), .A2(n23165), .ZN(n23177) );
  OAI22D1BWP12T U13906 ( .A1(n23170), .A2(n23169), .B1(n23168), .B2(n23167), 
        .ZN(n23176) );
  OAI211D1BWP12T U13907 ( .A1(n23174), .A2(n23173), .B(n23172), .C(n23171), 
        .ZN(n23175) );
  NR4D0BWP12T U13908 ( .A1(n23177), .A2(n23669), .A3(n23176), .A4(n23175), 
        .ZN(n23192) );
  MOAI22D0BWP12T U13909 ( .A1(n23181), .A2(n23180), .B1(n23179), .B2(n23178), 
        .ZN(n23187) );
  MOAI22D0BWP12T U13910 ( .A1(n23185), .A2(n23184), .B1(n23183), .B2(n23182), 
        .ZN(n23186) );
  NR4D0BWP12T U13911 ( .A1(n23189), .A2(n23188), .A3(n23187), .A4(n23186), 
        .ZN(n23191) );
  ND4D1BWP12T U13912 ( .A1(n23193), .A2(n23192), .A3(n23191), .A4(n23190), 
        .ZN(n23194) );
  NR4D0BWP12T U13913 ( .A1(n23197), .A2(n23196), .A3(n23195), .A4(n23194), 
        .ZN(n23198) );
  ND4D1BWP12T U13914 ( .A1(n23201), .A2(n23200), .A3(n23199), .A4(n23198), 
        .ZN(n23202) );
  NR4D0BWP12T U13915 ( .A1(n23205), .A2(n23204), .A3(n23203), .A4(n23202), 
        .ZN(n23591) );
  MOAI22D0BWP12T U13916 ( .A1(n23594), .A2(n23206), .B1(n23594), .B2(n23206), 
        .ZN(n23668) );
  INR4D0BWP12T U13917 ( .A1(n23210), .B1(n23209), .B2(n23208), .B3(n23207), 
        .ZN(n23243) );
  IND3D1BWP12T U13918 ( .A1(n23213), .B1(n23212), .B2(n23211), .ZN(n23405) );
  ND2D1BWP12T U13919 ( .A1(n23215), .A2(n23214), .ZN(n23398) );
  NR2D1BWP12T U13920 ( .A1(a[31]), .A2(n23216), .ZN(n23404) );
  ND4D1BWP12T U13921 ( .A1(n23220), .A2(n23219), .A3(n23218), .A4(n23217), 
        .ZN(n23228) );
  AOI211D1BWP12T U13922 ( .A1(n23229), .A2(n23228), .B(n23227), .C(n23411), 
        .ZN(n23231) );
  ND4D1BWP12T U13923 ( .A1(n23404), .A2(n23231), .A3(n23386), .A4(n23230), 
        .ZN(n23232) );
  NR2D1BWP12T U13924 ( .A1(n23398), .A2(n23232), .ZN(n23413) );
  OAI211D1BWP12T U13925 ( .A1(n23236), .A2(n23235), .B(n23234), .C(n23233), 
        .ZN(n23237) );
  NR2D1BWP12T U13926 ( .A1(n23238), .A2(n23237), .ZN(n23396) );
  NR2D1BWP12T U13927 ( .A1(n23408), .A2(n23239), .ZN(n23428) );
  ND4D1BWP12T U13928 ( .A1(n23413), .A2(n23396), .A3(n23428), .A4(n23240), 
        .ZN(n23241) );
  NR2D1BWP12T U13929 ( .A1(n23405), .A2(n23241), .ZN(n23242) );
  OAI32D1BWP12T U13930 ( .A1(n23294), .A2(b[4]), .A3(n23243), .B1(n23242), 
        .B2(n23294), .ZN(n23588) );
  ND4D1BWP12T U13931 ( .A1(n23246), .A2(n23264), .A3(n23245), .A4(n23244), 
        .ZN(n23253) );
  ND4D1BWP12T U13932 ( .A1(n23250), .A2(n23249), .A3(n23248), .A4(n23247), 
        .ZN(n23251) );
  AOI211D1BWP12T U13933 ( .A1(n23254), .A2(n23253), .B(n23252), .C(n23251), 
        .ZN(n23297) );
  MOAI22D0BWP12T U13934 ( .A1(a[31]), .A2(n23544), .B1(n23255), .B2(b[1]), 
        .ZN(n23256) );
  AOI31D1BWP12T U13935 ( .A1(n23259), .A2(n23258), .A3(n23257), .B(n23256), 
        .ZN(n23260) );
  OAI31D1BWP12T U13936 ( .A1(a[30]), .A2(n23262), .A3(n23261), .B(n23260), 
        .ZN(n23268) );
  MOAI22D0BWP12T U13937 ( .A1(n23266), .A2(n23265), .B1(n23264), .B2(n23263), 
        .ZN(n23267) );
  AOI211D1BWP12T U13938 ( .A1(n23270), .A2(n23269), .B(n23268), .C(n23267), 
        .ZN(n23643) );
  INR4D0BWP12T U13939 ( .A1(n23274), .B1(n23273), .B2(n23272), .B3(n23271), 
        .ZN(n23277) );
  ND4D1BWP12T U13940 ( .A1(n23278), .A2(n23277), .A3(n23276), .A4(n23275), 
        .ZN(n23292) );
  INR4D0BWP12T U13941 ( .A1(n23282), .B1(n23281), .B2(n23280), .B3(n23279), 
        .ZN(n23289) );
  NR4D0BWP12T U13942 ( .A1(n23286), .A2(n23285), .A3(n23284), .A4(n23283), 
        .ZN(n23288) );
  ND4D1BWP12T U13943 ( .A1(n23290), .A2(n23289), .A3(n23288), .A4(n23287), 
        .ZN(n23291) );
  NR4D0BWP12T U13944 ( .A1(n23643), .A2(n23293), .A3(n23292), .A4(n23291), 
        .ZN(n23296) );
  AOI31D1BWP12T U13945 ( .A1(n23297), .A2(n23296), .A3(n23295), .B(n23294), 
        .ZN(n23300) );
  NR4D0BWP12T U13946 ( .A1(n23301), .A2(n23300), .A3(n23299), .A4(n23298), 
        .ZN(n23384) );
  NR4D0BWP12T U13947 ( .A1(n23305), .A2(n23304), .A3(n23303), .A4(n23302), 
        .ZN(n23321) );
  NR4D0BWP12T U13948 ( .A1(n23309), .A2(n23308), .A3(n23307), .A4(n23306), 
        .ZN(n23320) );
  NR4D0BWP12T U13949 ( .A1(n23313), .A2(n23312), .A3(n23311), .A4(n23310), 
        .ZN(n23319) );
  NR4D0BWP12T U13950 ( .A1(n23317), .A2(n23316), .A3(n23315), .A4(n23314), 
        .ZN(n23318) );
  ND4D1BWP12T U13951 ( .A1(n23321), .A2(n23320), .A3(n23319), .A4(n23318), 
        .ZN(n23337) );
  NR4D0BWP12T U13952 ( .A1(n23324), .A2(n23323), .A3(n23322), .A4(n23657), 
        .ZN(n23335) );
  NR4D0BWP12T U13953 ( .A1(n23328), .A2(n23327), .A3(n23326), .A4(n23325), 
        .ZN(n23334) );
  NR4D0BWP12T U13954 ( .A1(n23332), .A2(n23331), .A3(n23330), .A4(n23329), 
        .ZN(n23333) );
  ND4D1BWP12T U13955 ( .A1(n23658), .A2(n23335), .A3(n23334), .A4(n23333), 
        .ZN(n23336) );
  OR4XD1BWP12T U13956 ( .A1(n23339), .A2(n23338), .A3(n23337), .A4(n23336), 
        .Z(n23379) );
  AOI211D1BWP12T U13957 ( .A1(a[13]), .A2(b[13]), .B(n23343), .C(n23342), .ZN(
        n23366) );
  ND4D1BWP12T U13958 ( .A1(n23347), .A2(n23346), .A3(n23345), .A4(n23344), 
        .ZN(n23362) );
  ND2D1BWP12T U13959 ( .A1(b[19]), .A2(a[19]), .ZN(n23348) );
  IND4D1BWP12T U13960 ( .A1(n23351), .B1(n23350), .B2(n23349), .B3(n23348), 
        .ZN(n23361) );
  OR4XD1BWP12T U13961 ( .A1(n23355), .A2(n23354), .A3(n23353), .A4(n23352), 
        .Z(n23360) );
  INVD1BWP12T U13962 ( .I(n23651), .ZN(n23649) );
  ND4D1BWP12T U13963 ( .A1(n23649), .A2(n23358), .A3(n23357), .A4(n23356), 
        .ZN(n23359) );
  NR4D0BWP12T U13964 ( .A1(n23362), .A2(n23361), .A3(n23360), .A4(n23359), 
        .ZN(n23365) );
  ND2D1BWP12T U13965 ( .A1(b[10]), .A2(a[10]), .ZN(n23363) );
  ND4D1BWP12T U13966 ( .A1(n23366), .A2(n23365), .A3(n23364), .A4(n23363), 
        .ZN(n23378) );
  AOI22D1BWP12T U13967 ( .A1(b[15]), .A2(a[15]), .B1(b[4]), .B2(a[4]), .ZN(
        n23368) );
  OAI211D1BWP12T U13968 ( .A1(n23370), .A2(n23369), .B(n23368), .C(n23367), 
        .ZN(n23371) );
  AOI211D1BWP12T U13969 ( .A1(b[28]), .A2(a[28]), .B(n23372), .C(n23371), .ZN(
        n23374) );
  OAI211D1BWP12T U13970 ( .A1(n23376), .A2(n23375), .B(n23374), .C(n23373), 
        .ZN(n23377) );
  OAI22D1BWP12T U13971 ( .A1(n23380), .A2(n23379), .B1(n23378), .B2(n23377), 
        .ZN(n23381) );
  AOI22D1BWP12T U13972 ( .A1(n23384), .A2(n23383), .B1(n23382), .B2(n23381), 
        .ZN(n23587) );
  ND4D1BWP12T U13973 ( .A1(n23388), .A2(n23387), .A3(n23386), .A4(n23385), 
        .ZN(n23389) );
  NR4D0BWP12T U13974 ( .A1(n23392), .A2(n23391), .A3(n23390), .A4(n23389), 
        .ZN(n23395) );
  ND4D1BWP12T U13975 ( .A1(n23396), .A2(n23395), .A3(n23394), .A4(n23393), 
        .ZN(n23399) );
  OAI31D1BWP12T U13976 ( .A1(n23400), .A2(n23399), .A3(n23398), .B(n23397), 
        .ZN(n23403) );
  AOI32D1BWP12T U13977 ( .A1(n23404), .A2(n23403), .A3(n23402), .B1(n23401), 
        .B2(n23403), .ZN(n23412) );
  INVD1BWP12T U13978 ( .I(n23405), .ZN(n23421) );
  IND4D1BWP12T U13979 ( .A1(n23408), .B1(n23407), .B2(n23421), .B3(n23406), 
        .ZN(n23410) );
  OAI32D1BWP12T U13980 ( .A1(n23412), .A2(n23411), .A3(n23410), .B1(n23409), 
        .B2(n23412), .ZN(n23584) );
  INVD1BWP12T U13981 ( .I(n23413), .ZN(n23581) );
  INR4D0BWP12T U13982 ( .A1(n23417), .B1(n23416), .B2(n23415), .B3(n23414), 
        .ZN(n23418) );
  ND4D1BWP12T U13983 ( .A1(n23421), .A2(n23420), .A3(n23419), .A4(n23418), 
        .ZN(n23580) );
  ND4D1BWP12T U13984 ( .A1(n23424), .A2(n23423), .A3(n23667), .A4(n23422), 
        .ZN(n23430) );
  ND4D1BWP12T U13985 ( .A1(n23428), .A2(n23427), .A3(n23426), .A4(n23425), 
        .ZN(n23429) );
  NR4D0BWP12T U13986 ( .A1(n23432), .A2(n23431), .A3(n23430), .A4(n23429), 
        .ZN(n23470) );
  ND4D1BWP12T U13987 ( .A1(n23435), .A2(n23434), .A3(n23433), .A4(n23451), 
        .ZN(n23436) );
  INR4D0BWP12T U13988 ( .A1(n23439), .B1(n23438), .B2(n23437), .B3(n23436), 
        .ZN(n23469) );
  AOI22D1BWP12T U13989 ( .A1(a[30]), .A2(n23442), .B1(n23441), .B2(n23440), 
        .ZN(n23449) );
  INVD1BWP12T U13990 ( .I(n23443), .ZN(n23447) );
  AOI22D1BWP12T U13991 ( .A1(n23447), .A2(n23446), .B1(n23445), .B2(n23444), 
        .ZN(n23448) );
  OAI211D1BWP12T U13992 ( .A1(n23451), .A2(n23450), .B(n23449), .C(n23448), 
        .ZN(n23666) );
  IND4D1BWP12T U13993 ( .A1(n23455), .B1(n23454), .B2(n23453), .B3(n23452), 
        .ZN(n23465) );
  NR4D0BWP12T U13994 ( .A1(n23459), .A2(n23458), .A3(n23457), .A4(n23456), 
        .ZN(n23461) );
  ND4D1BWP12T U13995 ( .A1(n23463), .A2(n23462), .A3(n23461), .A4(n23460), 
        .ZN(n23464) );
  NR4D0BWP12T U13996 ( .A1(n23466), .A2(n23666), .A3(n23465), .A4(n23464), 
        .ZN(n23468) );
  ND4D1BWP12T U13997 ( .A1(n23470), .A2(n23469), .A3(n23468), .A4(n23467), 
        .ZN(n23579) );
  AN4XD1BWP12T U13998 ( .A1(n23474), .A2(n23473), .A3(n23472), .A4(n23471), 
        .Z(n23577) );
  INR4D0BWP12T U13999 ( .A1(n23478), .B1(n23477), .B2(n23476), .B3(n23475), 
        .ZN(n23576) );
  IND4D1BWP12T U14000 ( .A1(n23513), .B1(n23512), .B2(n23511), .B3(n23510), 
        .ZN(n23536) );
  IND4D1BWP12T U14001 ( .A1(n23517), .B1(n23516), .B2(n23515), .B3(n23514), 
        .ZN(n23535) );
  NR4D0BWP12T U14002 ( .A1(n23521), .A2(n23520), .A3(n23519), .A4(n23518), 
        .ZN(n23532) );
  IND4D1BWP12T U14003 ( .A1(n23525), .B1(n23524), .B2(n23523), .B3(n23522), 
        .ZN(n23526) );
  NR4D0BWP12T U14004 ( .A1(n23529), .A2(n23528), .A3(n23527), .A4(n23526), 
        .ZN(n23531) );
  IND4D1BWP12T U14005 ( .A1(n23533), .B1(n23532), .B2(n23531), .B3(n23530), 
        .ZN(n23534) );
  NR4D0BWP12T U14006 ( .A1(n23537), .A2(n23536), .A3(n23535), .A4(n23534), 
        .ZN(n23575) );
  INVD1BWP12T U14007 ( .I(n23538), .ZN(n23573) );
  ND4D1BWP12T U14008 ( .A1(n23656), .A2(n23541), .A3(n23540), .A4(n23539), 
        .ZN(n23542) );
  NR4D0BWP12T U14009 ( .A1(b[24]), .A2(b[13]), .A3(n23543), .A4(n23542), .ZN(
        n23547) );
  NR4D0BWP12T U14010 ( .A1(a[27]), .A2(a[25]), .A3(n23544), .A4(n23645), .ZN(
        n23545) );
  ND4D1BWP12T U14011 ( .A1(n23548), .A2(n23547), .A3(n23546), .A4(n23545), 
        .ZN(n23571) );
  INR4D0BWP12T U14012 ( .A1(n23552), .B1(n23551), .B2(n23550), .B3(n23549), 
        .ZN(n23568) );
  ND4D1BWP12T U14013 ( .A1(a[23]), .A2(a[20]), .A3(a[13]), .A4(a[8]), .ZN(
        n23564) );
  INR4D0BWP12T U14014 ( .A1(n23556), .B1(n23555), .B2(n23554), .B3(n23553), 
        .ZN(n23562) );
  NR4D0BWP12T U14015 ( .A1(n23560), .A2(n23559), .A3(n23558), .A4(n23557), 
        .ZN(n23561) );
  ND4D1BWP12T U14016 ( .A1(a[31]), .A2(a[5]), .A3(n23562), .A4(n23561), .ZN(
        n23563) );
  NR4D0BWP12T U14017 ( .A1(n23566), .A2(n23565), .A3(n23564), .A4(n23563), 
        .ZN(n23567) );
  AOI22D1BWP12T U14018 ( .A1(n23659), .A2(n23569), .B1(n23568), .B2(n23567), 
        .ZN(n23570) );
  OAI31D1BWP12T U14019 ( .A1(n23573), .A2(n23572), .A3(n23571), .B(n23570), 
        .ZN(n23574) );
  AOI31D1BWP12T U14020 ( .A1(n23577), .A2(n23576), .A3(n23575), .B(n23574), 
        .ZN(n23578) );
  OAI31D1BWP12T U14021 ( .A1(n23581), .A2(n23580), .A3(n23579), .B(n23578), 
        .ZN(n23582) );
  AOI31D1BWP12T U14022 ( .A1(n23585), .A2(n23584), .A3(n23583), .B(n23582), 
        .ZN(n23586) );
  OAI211D1BWP12T U14023 ( .A1(n23589), .A2(n23588), .B(n23587), .C(n23586), 
        .ZN(n23590) );
  AOI31D1BWP12T U14024 ( .A1(n23592), .A2(n23591), .A3(n23668), .B(n23590), 
        .ZN(n23638) );
  MAOI22D0BWP12T U14025 ( .A1(n23594), .A2(n23593), .B1(n23594), .B2(n23593), 
        .ZN(n23654) );
  ND4D1BWP12T U14026 ( .A1(n23597), .A2(n23654), .A3(n23596), .A4(n23595), 
        .ZN(n23611) );
  ND4D1BWP12T U14027 ( .A1(n23601), .A2(n23600), .A3(n23599), .A4(n23598), 
        .ZN(n23602) );
  NR4D0BWP12T U14028 ( .A1(n23605), .A2(n23604), .A3(n23603), .A4(n23602), 
        .ZN(n23607) );
  ND4D1BWP12T U14029 ( .A1(n23609), .A2(n23608), .A3(n23607), .A4(n23606), 
        .ZN(n23610) );
  NR4D0BWP12T U14030 ( .A1(n23613), .A2(n23612), .A3(n23611), .A4(n23610), 
        .ZN(n23614) );
  ND4D1BWP12T U14031 ( .A1(n23617), .A2(n23616), .A3(n23615), .A4(n23614), 
        .ZN(n23618) );
  NR4D0BWP12T U14032 ( .A1(n23621), .A2(n23620), .A3(n23619), .A4(n23618), 
        .ZN(n23622) );
  ND4D1BWP12T U14033 ( .A1(n23625), .A2(n23624), .A3(n23623), .A4(n23622), 
        .ZN(n23630) );
  ND3D1BWP12T U14034 ( .A1(n23628), .A2(n23627), .A3(n23626), .ZN(n23629) );
  NR4D0BWP12T U14035 ( .A1(n23632), .A2(n23631), .A3(n23630), .A4(n23629), 
        .ZN(n23635) );
  ND4D1BWP12T U14036 ( .A1(n23636), .A2(n23635), .A3(n23634), .A4(n23633), 
        .ZN(n23637) );
  OAI211D1BWP12T U14037 ( .A1(n23640), .A2(n23639), .B(n23638), .C(n23637), 
        .ZN(z) );
  AOI22D1BWP12T U14038 ( .A1(n23644), .A2(n23643), .B1(n23642), .B2(n23641), 
        .ZN(n23678) );
  OAI211D1BWP12T U14039 ( .A1(b[31]), .A2(n23647), .B(n23646), .C(n23645), 
        .ZN(n23648) );
  AOI221D1BWP12T U14040 ( .A1(n23652), .A2(n23651), .B1(n23650), .B2(n23649), 
        .C(n23648), .ZN(n23655) );
  OAI22D1BWP12T U14041 ( .A1(n23656), .A2(n23655), .B1(n23654), .B2(n23653), 
        .ZN(n23665) );
  AOI22D1BWP12T U14042 ( .A1(a[30]), .A2(n23659), .B1(n23658), .B2(n23657), 
        .ZN(n23660) );
  OAI31D1BWP12T U14043 ( .A1(n23663), .A2(n23662), .A3(n23661), .B(n23660), 
        .ZN(n23664) );
  AOI211D1BWP12T U14044 ( .A1(n23667), .A2(n23666), .B(n23665), .C(n23664), 
        .ZN(n23677) );
  OAI22D1BWP12T U14045 ( .A1(n23671), .A2(n23670), .B1(n23669), .B2(n23668), 
        .ZN(n23672) );
  AOI21D1BWP12T U14046 ( .A1(n23674), .A2(n23673), .B(n23672), .ZN(n23676) );
  ND4D1BWP12T U14047 ( .A1(n23678), .A2(n23677), .A3(n23676), .A4(n23675), 
        .ZN(result[31]) );
  CKBD1BWP12T U14048 ( .I(result[31]), .Z(n) );
endmodule

