
module register_file ( readA_sel, readB_sel, readC_sel, readD_sel, write1_sel, 
        write2_sel, write1_en, write2_en, write1_in, write2_in, immediate1_in, 
        immediate2_in, next_pc_in, next_cpsr_in, next_sp_in, clk, reset, 
        regA_out, regB_out, regC_out, regD_out, pc_out, cpsr_out, sp_out, 
        next_pc_en_BAR );
  input [4:0] readA_sel;
  input [4:0] readB_sel;
  input [4:0] readC_sel;
  input [4:0] readD_sel;
  input [4:0] write1_sel;
  input [4:0] write2_sel;
  input [31:0] write1_in;
  input [31:0] write2_in;
  input [31:0] immediate1_in;
  input [31:0] immediate2_in;
  input [31:0] next_pc_in;
  input [3:0] next_cpsr_in;
  input [31:0] next_sp_in;
  output [31:0] regA_out;
  output [31:0] regB_out;
  output [31:0] regC_out;
  output [31:0] regD_out;
  output [31:0] pc_out;
  output [3:0] cpsr_out;
  output [31:0] sp_out;
  input write1_en, write2_en, clk, reset, next_pc_en_BAR;
  wire   n2136, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009;
  wire   [2010:2041] n;
  wire   [31:0] r0;
  wire   [31:0] r1;
  wire   [31:0] r2;
  wire   [31:0] r3;
  wire   [31:0] r4;
  wire   [31:0] r5;
  wire   [31:0] r6;
  wire   [31:0] r7;
  wire   [31:0] r8;
  wire   [31:0] r9;
  wire   [31:0] r10;
  wire   [31:0] r11;
  wire   [31:0] r12;
  wire   [31:0] lr;
  wire   [31:0] tmp1;
  wire   [31:0] spin;
  wire   [3:0] cpsrin;

  DFQD1BWP12T r0_reg_31_ ( .D(n2648), .CP(clk), .Q(r0[31]) );
  DFQD1BWP12T r0_reg_30_ ( .D(n2647), .CP(clk), .Q(r0[30]) );
  DFQD1BWP12T r0_reg_29_ ( .D(n2646), .CP(clk), .Q(r0[29]) );
  DFQD1BWP12T r0_reg_28_ ( .D(n2645), .CP(clk), .Q(r0[28]) );
  DFQD1BWP12T r0_reg_27_ ( .D(n2644), .CP(clk), .Q(r0[27]) );
  DFQD1BWP12T r0_reg_26_ ( .D(n2643), .CP(clk), .Q(r0[26]) );
  DFQD1BWP12T r0_reg_25_ ( .D(n2642), .CP(clk), .Q(r0[25]) );
  DFQD1BWP12T r0_reg_24_ ( .D(n2641), .CP(clk), .Q(r0[24]) );
  DFQD1BWP12T r0_reg_23_ ( .D(n2640), .CP(clk), .Q(r0[23]) );
  DFQD1BWP12T r0_reg_22_ ( .D(n2639), .CP(clk), .Q(r0[22]) );
  DFQD1BWP12T r0_reg_21_ ( .D(n2638), .CP(clk), .Q(r0[21]) );
  DFQD1BWP12T r0_reg_20_ ( .D(n2637), .CP(clk), .Q(r0[20]) );
  DFQD1BWP12T r0_reg_19_ ( .D(n2636), .CP(clk), .Q(r0[19]) );
  DFQD1BWP12T r0_reg_18_ ( .D(n2635), .CP(clk), .Q(r0[18]) );
  DFQD1BWP12T r0_reg_17_ ( .D(n2634), .CP(clk), .Q(r0[17]) );
  DFQD1BWP12T r0_reg_16_ ( .D(n2633), .CP(clk), .Q(r0[16]) );
  DFQD1BWP12T r0_reg_15_ ( .D(n2632), .CP(clk), .Q(r0[15]) );
  DFQD1BWP12T r0_reg_14_ ( .D(n2631), .CP(clk), .Q(r0[14]) );
  DFQD1BWP12T r0_reg_13_ ( .D(n2630), .CP(clk), .Q(r0[13]) );
  DFQD1BWP12T r0_reg_12_ ( .D(n2629), .CP(clk), .Q(r0[12]) );
  DFQD1BWP12T r0_reg_11_ ( .D(n2628), .CP(clk), .Q(r0[11]) );
  DFQD1BWP12T r0_reg_10_ ( .D(n2627), .CP(clk), .Q(r0[10]) );
  DFQD1BWP12T r0_reg_9_ ( .D(n2626), .CP(clk), .Q(r0[9]) );
  DFQD1BWP12T r0_reg_8_ ( .D(n2625), .CP(clk), .Q(r0[8]) );
  DFQD1BWP12T r0_reg_7_ ( .D(n2624), .CP(clk), .Q(r0[7]) );
  DFQD1BWP12T r0_reg_6_ ( .D(n2623), .CP(clk), .Q(r0[6]) );
  DFQD1BWP12T r0_reg_5_ ( .D(n2622), .CP(clk), .Q(r0[5]) );
  DFQD1BWP12T r0_reg_4_ ( .D(n2621), .CP(clk), .Q(r0[4]) );
  DFQD1BWP12T r0_reg_3_ ( .D(n2620), .CP(clk), .Q(r0[3]) );
  DFQD1BWP12T r0_reg_2_ ( .D(n2619), .CP(clk), .Q(r0[2]) );
  DFQD1BWP12T r0_reg_1_ ( .D(n2618), .CP(clk), .Q(r0[1]) );
  DFQD1BWP12T r0_reg_0_ ( .D(n2617), .CP(clk), .Q(r0[0]) );
  DFQD1BWP12T r1_reg_31_ ( .D(n2616), .CP(clk), .Q(r1[31]) );
  DFQD1BWP12T r1_reg_30_ ( .D(n2615), .CP(clk), .Q(r1[30]) );
  DFQD1BWP12T r1_reg_29_ ( .D(n2614), .CP(clk), .Q(r1[29]) );
  DFQD1BWP12T r1_reg_28_ ( .D(n2613), .CP(clk), .Q(r1[28]) );
  DFQD1BWP12T r1_reg_27_ ( .D(n2612), .CP(clk), .Q(r1[27]) );
  DFQD1BWP12T r1_reg_26_ ( .D(n2611), .CP(clk), .Q(r1[26]) );
  DFQD1BWP12T r1_reg_25_ ( .D(n2610), .CP(clk), .Q(r1[25]) );
  DFQD1BWP12T r1_reg_24_ ( .D(n2609), .CP(clk), .Q(r1[24]) );
  DFQD1BWP12T r1_reg_23_ ( .D(n2608), .CP(clk), .Q(r1[23]) );
  DFQD1BWP12T r1_reg_22_ ( .D(n2607), .CP(clk), .Q(r1[22]) );
  DFQD1BWP12T r1_reg_21_ ( .D(n2606), .CP(clk), .Q(r1[21]) );
  DFQD1BWP12T r1_reg_20_ ( .D(n2605), .CP(clk), .Q(r1[20]) );
  DFQD1BWP12T r1_reg_19_ ( .D(n2604), .CP(clk), .Q(r1[19]) );
  DFQD1BWP12T r1_reg_18_ ( .D(n2603), .CP(clk), .Q(r1[18]) );
  DFQD1BWP12T r1_reg_17_ ( .D(n2602), .CP(clk), .Q(r1[17]) );
  DFQD1BWP12T r1_reg_16_ ( .D(n2601), .CP(clk), .Q(r1[16]) );
  DFQD1BWP12T r1_reg_15_ ( .D(n2600), .CP(clk), .Q(r1[15]) );
  DFQD1BWP12T r1_reg_14_ ( .D(n2599), .CP(clk), .Q(r1[14]) );
  DFQD1BWP12T r1_reg_13_ ( .D(n2598), .CP(clk), .Q(r1[13]) );
  DFQD1BWP12T r1_reg_12_ ( .D(n2597), .CP(clk), .Q(r1[12]) );
  DFQD1BWP12T r1_reg_11_ ( .D(n2596), .CP(clk), .Q(r1[11]) );
  DFQD1BWP12T r1_reg_10_ ( .D(n2595), .CP(clk), .Q(r1[10]) );
  DFQD1BWP12T r1_reg_9_ ( .D(n2594), .CP(clk), .Q(r1[9]) );
  DFQD1BWP12T r1_reg_8_ ( .D(n2593), .CP(clk), .Q(r1[8]) );
  DFQD1BWP12T r1_reg_7_ ( .D(n2592), .CP(clk), .Q(r1[7]) );
  DFQD1BWP12T r1_reg_6_ ( .D(n2591), .CP(clk), .Q(r1[6]) );
  DFQD1BWP12T r1_reg_5_ ( .D(n2590), .CP(clk), .Q(r1[5]) );
  DFQD1BWP12T r1_reg_4_ ( .D(n2589), .CP(clk), .Q(r1[4]) );
  DFQD1BWP12T r1_reg_3_ ( .D(n2588), .CP(clk), .Q(r1[3]) );
  DFQD1BWP12T r1_reg_2_ ( .D(n2587), .CP(clk), .Q(r1[2]) );
  DFQD1BWP12T r1_reg_1_ ( .D(n2586), .CP(clk), .Q(r1[1]) );
  DFQD1BWP12T r1_reg_0_ ( .D(n2585), .CP(clk), .Q(r1[0]) );
  DFQD1BWP12T r2_reg_31_ ( .D(n2584), .CP(clk), .Q(r2[31]) );
  DFQD1BWP12T r2_reg_30_ ( .D(n2583), .CP(clk), .Q(r2[30]) );
  DFQD1BWP12T r2_reg_29_ ( .D(n2582), .CP(clk), .Q(r2[29]) );
  DFQD1BWP12T r2_reg_28_ ( .D(n2581), .CP(clk), .Q(r2[28]) );
  DFQD1BWP12T r2_reg_27_ ( .D(n2580), .CP(clk), .Q(r2[27]) );
  DFQD1BWP12T r2_reg_26_ ( .D(n2579), .CP(clk), .Q(r2[26]) );
  DFQD1BWP12T r2_reg_25_ ( .D(n2578), .CP(clk), .Q(r2[25]) );
  DFQD1BWP12T r2_reg_24_ ( .D(n2577), .CP(clk), .Q(r2[24]) );
  DFQD1BWP12T r2_reg_23_ ( .D(n2576), .CP(clk), .Q(r2[23]) );
  DFQD1BWP12T r2_reg_22_ ( .D(n2575), .CP(clk), .Q(r2[22]) );
  DFQD1BWP12T r2_reg_21_ ( .D(n2574), .CP(clk), .Q(r2[21]) );
  DFQD1BWP12T r2_reg_20_ ( .D(n2573), .CP(clk), .Q(r2[20]) );
  DFQD1BWP12T r2_reg_19_ ( .D(n2572), .CP(clk), .Q(r2[19]) );
  DFQD1BWP12T r2_reg_18_ ( .D(n2571), .CP(clk), .Q(r2[18]) );
  DFQD1BWP12T r2_reg_17_ ( .D(n2570), .CP(clk), .Q(r2[17]) );
  DFQD1BWP12T r2_reg_16_ ( .D(n2569), .CP(clk), .Q(r2[16]) );
  DFQD1BWP12T r2_reg_15_ ( .D(n2568), .CP(clk), .Q(r2[15]) );
  DFQD1BWP12T r2_reg_14_ ( .D(n2567), .CP(clk), .Q(r2[14]) );
  DFQD1BWP12T r2_reg_13_ ( .D(n2566), .CP(clk), .Q(r2[13]) );
  DFQD1BWP12T r2_reg_12_ ( .D(n2565), .CP(clk), .Q(r2[12]) );
  DFQD1BWP12T r2_reg_11_ ( .D(n2564), .CP(clk), .Q(r2[11]) );
  DFQD1BWP12T r2_reg_10_ ( .D(n2563), .CP(clk), .Q(r2[10]) );
  DFQD1BWP12T r2_reg_9_ ( .D(n2562), .CP(clk), .Q(r2[9]) );
  DFQD1BWP12T r2_reg_8_ ( .D(n2561), .CP(clk), .Q(r2[8]) );
  DFQD1BWP12T r2_reg_7_ ( .D(n2560), .CP(clk), .Q(r2[7]) );
  DFQD1BWP12T r2_reg_6_ ( .D(n2559), .CP(clk), .Q(r2[6]) );
  DFQD1BWP12T r2_reg_5_ ( .D(n2558), .CP(clk), .Q(r2[5]) );
  DFQD1BWP12T r2_reg_4_ ( .D(n2557), .CP(clk), .Q(r2[4]) );
  DFQD1BWP12T r2_reg_3_ ( .D(n2556), .CP(clk), .Q(r2[3]) );
  DFQD1BWP12T r2_reg_2_ ( .D(n2555), .CP(clk), .Q(r2[2]) );
  DFQD1BWP12T r2_reg_1_ ( .D(n2554), .CP(clk), .Q(r2[1]) );
  DFQD1BWP12T r2_reg_0_ ( .D(n2553), .CP(clk), .Q(r2[0]) );
  DFQD1BWP12T r3_reg_31_ ( .D(n2552), .CP(clk), .Q(r3[31]) );
  DFQD1BWP12T r3_reg_30_ ( .D(n2551), .CP(clk), .Q(r3[30]) );
  DFQD1BWP12T r3_reg_29_ ( .D(n2550), .CP(clk), .Q(r3[29]) );
  DFQD1BWP12T r3_reg_28_ ( .D(n2549), .CP(clk), .Q(r3[28]) );
  DFQD1BWP12T r3_reg_27_ ( .D(n2548), .CP(clk), .Q(r3[27]) );
  DFQD1BWP12T r3_reg_26_ ( .D(n2547), .CP(clk), .Q(r3[26]) );
  DFQD1BWP12T r3_reg_25_ ( .D(n2546), .CP(clk), .Q(r3[25]) );
  DFQD1BWP12T r3_reg_24_ ( .D(n2545), .CP(clk), .Q(r3[24]) );
  DFQD1BWP12T r3_reg_23_ ( .D(n2544), .CP(clk), .Q(r3[23]) );
  DFQD1BWP12T r3_reg_22_ ( .D(n2543), .CP(clk), .Q(r3[22]) );
  DFQD1BWP12T r3_reg_21_ ( .D(n2542), .CP(clk), .Q(r3[21]) );
  DFQD1BWP12T r3_reg_20_ ( .D(n2541), .CP(clk), .Q(r3[20]) );
  DFQD1BWP12T r3_reg_19_ ( .D(n2540), .CP(clk), .Q(r3[19]) );
  DFQD1BWP12T r3_reg_18_ ( .D(n2539), .CP(clk), .Q(r3[18]) );
  DFQD1BWP12T r3_reg_17_ ( .D(n2538), .CP(clk), .Q(r3[17]) );
  DFQD1BWP12T r3_reg_16_ ( .D(n2537), .CP(clk), .Q(r3[16]) );
  DFQD1BWP12T r3_reg_15_ ( .D(n2536), .CP(clk), .Q(r3[15]) );
  DFQD1BWP12T r3_reg_14_ ( .D(n2535), .CP(clk), .Q(r3[14]) );
  DFQD1BWP12T r3_reg_13_ ( .D(n2534), .CP(clk), .Q(r3[13]) );
  DFQD1BWP12T r3_reg_12_ ( .D(n2533), .CP(clk), .Q(r3[12]) );
  DFQD1BWP12T r3_reg_11_ ( .D(n2532), .CP(clk), .Q(r3[11]) );
  DFQD1BWP12T r3_reg_10_ ( .D(n2531), .CP(clk), .Q(r3[10]) );
  DFQD1BWP12T r3_reg_9_ ( .D(n2530), .CP(clk), .Q(r3[9]) );
  DFQD1BWP12T r3_reg_8_ ( .D(n2529), .CP(clk), .Q(r3[8]) );
  DFQD1BWP12T r3_reg_7_ ( .D(n2528), .CP(clk), .Q(r3[7]) );
  DFQD1BWP12T r3_reg_6_ ( .D(n2527), .CP(clk), .Q(r3[6]) );
  DFQD1BWP12T r3_reg_5_ ( .D(n2526), .CP(clk), .Q(r3[5]) );
  DFQD1BWP12T r3_reg_4_ ( .D(n2525), .CP(clk), .Q(r3[4]) );
  DFQD1BWP12T r3_reg_3_ ( .D(n2524), .CP(clk), .Q(r3[3]) );
  DFQD1BWP12T r3_reg_2_ ( .D(n2523), .CP(clk), .Q(r3[2]) );
  DFQD1BWP12T r3_reg_1_ ( .D(n2522), .CP(clk), .Q(r3[1]) );
  DFQD1BWP12T r3_reg_0_ ( .D(n2521), .CP(clk), .Q(r3[0]) );
  DFQD1BWP12T r4_reg_31_ ( .D(n2520), .CP(clk), .Q(r4[31]) );
  DFQD1BWP12T r4_reg_30_ ( .D(n2519), .CP(clk), .Q(r4[30]) );
  DFQD1BWP12T r4_reg_29_ ( .D(n2518), .CP(clk), .Q(r4[29]) );
  DFQD1BWP12T r4_reg_28_ ( .D(n2517), .CP(clk), .Q(r4[28]) );
  DFQD1BWP12T r4_reg_27_ ( .D(n2516), .CP(clk), .Q(r4[27]) );
  DFQD1BWP12T r4_reg_26_ ( .D(n2515), .CP(clk), .Q(r4[26]) );
  DFQD1BWP12T r4_reg_25_ ( .D(n2514), .CP(clk), .Q(r4[25]) );
  DFQD1BWP12T r4_reg_24_ ( .D(n2513), .CP(clk), .Q(r4[24]) );
  DFQD1BWP12T r4_reg_23_ ( .D(n2512), .CP(clk), .Q(r4[23]) );
  DFQD1BWP12T r4_reg_22_ ( .D(n2511), .CP(clk), .Q(r4[22]) );
  DFQD1BWP12T r4_reg_21_ ( .D(n2510), .CP(clk), .Q(r4[21]) );
  DFQD1BWP12T r4_reg_20_ ( .D(n2509), .CP(clk), .Q(r4[20]) );
  DFQD1BWP12T r4_reg_19_ ( .D(n2508), .CP(clk), .Q(r4[19]) );
  DFQD1BWP12T r4_reg_18_ ( .D(n2507), .CP(clk), .Q(r4[18]) );
  DFQD1BWP12T r4_reg_17_ ( .D(n2506), .CP(clk), .Q(r4[17]) );
  DFQD1BWP12T r4_reg_16_ ( .D(n2505), .CP(clk), .Q(r4[16]) );
  DFQD1BWP12T r4_reg_15_ ( .D(n2504), .CP(clk), .Q(r4[15]) );
  DFQD1BWP12T r4_reg_14_ ( .D(n2503), .CP(clk), .Q(r4[14]) );
  DFQD1BWP12T r4_reg_13_ ( .D(n2502), .CP(clk), .Q(r4[13]) );
  DFQD1BWP12T r4_reg_12_ ( .D(n2501), .CP(clk), .Q(r4[12]) );
  DFQD1BWP12T r4_reg_11_ ( .D(n2500), .CP(clk), .Q(r4[11]) );
  DFQD1BWP12T r4_reg_10_ ( .D(n2499), .CP(clk), .Q(r4[10]) );
  DFQD1BWP12T r4_reg_9_ ( .D(n2498), .CP(clk), .Q(r4[9]) );
  DFQD1BWP12T r4_reg_8_ ( .D(n2497), .CP(clk), .Q(r4[8]) );
  DFQD1BWP12T r4_reg_7_ ( .D(n2496), .CP(clk), .Q(r4[7]) );
  DFQD1BWP12T r4_reg_6_ ( .D(n2495), .CP(clk), .Q(r4[6]) );
  DFQD1BWP12T r4_reg_5_ ( .D(n2494), .CP(clk), .Q(r4[5]) );
  DFQD1BWP12T r4_reg_4_ ( .D(n2493), .CP(clk), .Q(r4[4]) );
  DFQD1BWP12T r4_reg_3_ ( .D(n2492), .CP(clk), .Q(r4[3]) );
  DFQD1BWP12T r4_reg_2_ ( .D(n2491), .CP(clk), .Q(r4[2]) );
  DFQD1BWP12T r4_reg_1_ ( .D(n2490), .CP(clk), .Q(r4[1]) );
  DFQD1BWP12T r4_reg_0_ ( .D(n2489), .CP(clk), .Q(r4[0]) );
  DFQD1BWP12T r5_reg_31_ ( .D(n2488), .CP(clk), .Q(r5[31]) );
  DFQD1BWP12T r5_reg_30_ ( .D(n2487), .CP(clk), .Q(r5[30]) );
  DFQD1BWP12T r5_reg_29_ ( .D(n2486), .CP(clk), .Q(r5[29]) );
  DFQD1BWP12T r5_reg_28_ ( .D(n2485), .CP(clk), .Q(r5[28]) );
  DFQD1BWP12T r5_reg_27_ ( .D(n2484), .CP(clk), .Q(r5[27]) );
  DFQD1BWP12T r5_reg_26_ ( .D(n2483), .CP(clk), .Q(r5[26]) );
  DFQD1BWP12T r5_reg_25_ ( .D(n2482), .CP(clk), .Q(r5[25]) );
  DFQD1BWP12T r5_reg_24_ ( .D(n2481), .CP(clk), .Q(r5[24]) );
  DFQD1BWP12T r5_reg_23_ ( .D(n2480), .CP(clk), .Q(r5[23]) );
  DFQD1BWP12T r5_reg_22_ ( .D(n2479), .CP(clk), .Q(r5[22]) );
  DFQD1BWP12T r5_reg_21_ ( .D(n2478), .CP(clk), .Q(r5[21]) );
  DFQD1BWP12T r5_reg_20_ ( .D(n2477), .CP(clk), .Q(r5[20]) );
  DFQD1BWP12T r5_reg_19_ ( .D(n2476), .CP(clk), .Q(r5[19]) );
  DFQD1BWP12T r5_reg_18_ ( .D(n2475), .CP(clk), .Q(r5[18]) );
  DFQD1BWP12T r5_reg_17_ ( .D(n2474), .CP(clk), .Q(r5[17]) );
  DFQD1BWP12T r5_reg_16_ ( .D(n2473), .CP(clk), .Q(r5[16]) );
  DFQD1BWP12T r5_reg_15_ ( .D(n2472), .CP(clk), .Q(r5[15]) );
  DFQD1BWP12T r5_reg_14_ ( .D(n2471), .CP(clk), .Q(r5[14]) );
  DFQD1BWP12T r5_reg_13_ ( .D(n2470), .CP(clk), .Q(r5[13]) );
  DFQD1BWP12T r5_reg_12_ ( .D(n2469), .CP(clk), .Q(r5[12]) );
  DFQD1BWP12T r5_reg_11_ ( .D(n2468), .CP(clk), .Q(r5[11]) );
  DFQD1BWP12T r5_reg_10_ ( .D(n2467), .CP(clk), .Q(r5[10]) );
  DFQD1BWP12T r5_reg_9_ ( .D(n2466), .CP(clk), .Q(r5[9]) );
  DFQD1BWP12T r5_reg_8_ ( .D(n2465), .CP(clk), .Q(r5[8]) );
  DFQD1BWP12T r5_reg_7_ ( .D(n2464), .CP(clk), .Q(r5[7]) );
  DFQD1BWP12T r5_reg_6_ ( .D(n2463), .CP(clk), .Q(r5[6]) );
  DFQD1BWP12T r5_reg_5_ ( .D(n2462), .CP(clk), .Q(r5[5]) );
  DFQD1BWP12T r5_reg_4_ ( .D(n2461), .CP(clk), .Q(r5[4]) );
  DFQD1BWP12T r5_reg_3_ ( .D(n2460), .CP(clk), .Q(r5[3]) );
  DFQD1BWP12T r5_reg_2_ ( .D(n2459), .CP(clk), .Q(r5[2]) );
  DFQD1BWP12T r5_reg_1_ ( .D(n2458), .CP(clk), .Q(r5[1]) );
  DFQD1BWP12T r5_reg_0_ ( .D(n2457), .CP(clk), .Q(r5[0]) );
  DFQD1BWP12T r6_reg_31_ ( .D(n2456), .CP(clk), .Q(r6[31]) );
  DFQD1BWP12T r6_reg_30_ ( .D(n2455), .CP(clk), .Q(r6[30]) );
  DFQD1BWP12T r6_reg_29_ ( .D(n2454), .CP(clk), .Q(r6[29]) );
  DFQD1BWP12T r6_reg_28_ ( .D(n2453), .CP(clk), .Q(r6[28]) );
  DFQD1BWP12T r6_reg_27_ ( .D(n2452), .CP(clk), .Q(r6[27]) );
  DFQD1BWP12T r6_reg_26_ ( .D(n2451), .CP(clk), .Q(r6[26]) );
  DFQD1BWP12T r6_reg_25_ ( .D(n2450), .CP(clk), .Q(r6[25]) );
  DFQD1BWP12T r6_reg_24_ ( .D(n2449), .CP(clk), .Q(r6[24]) );
  DFQD1BWP12T r6_reg_23_ ( .D(n2448), .CP(clk), .Q(r6[23]) );
  DFQD1BWP12T r6_reg_22_ ( .D(n2447), .CP(clk), .Q(r6[22]) );
  DFQD1BWP12T r6_reg_21_ ( .D(n2446), .CP(clk), .Q(r6[21]) );
  DFQD1BWP12T r6_reg_20_ ( .D(n2445), .CP(clk), .Q(r6[20]) );
  DFQD1BWP12T r6_reg_19_ ( .D(n2444), .CP(clk), .Q(r6[19]) );
  DFQD1BWP12T r6_reg_18_ ( .D(n2443), .CP(clk), .Q(r6[18]) );
  DFQD1BWP12T r6_reg_17_ ( .D(n2442), .CP(clk), .Q(r6[17]) );
  DFQD1BWP12T r6_reg_16_ ( .D(n2441), .CP(clk), .Q(r6[16]) );
  DFQD1BWP12T r6_reg_15_ ( .D(n2440), .CP(clk), .Q(r6[15]) );
  DFQD1BWP12T r6_reg_14_ ( .D(n2439), .CP(clk), .Q(r6[14]) );
  DFQD1BWP12T r6_reg_13_ ( .D(n2438), .CP(clk), .Q(r6[13]) );
  DFQD1BWP12T r6_reg_12_ ( .D(n2437), .CP(clk), .Q(r6[12]) );
  DFQD1BWP12T r6_reg_11_ ( .D(n2436), .CP(clk), .Q(r6[11]) );
  DFQD1BWP12T r6_reg_10_ ( .D(n2435), .CP(clk), .Q(r6[10]) );
  DFQD1BWP12T r6_reg_9_ ( .D(n2434), .CP(clk), .Q(r6[9]) );
  DFQD1BWP12T r6_reg_8_ ( .D(n2433), .CP(clk), .Q(r6[8]) );
  DFQD1BWP12T r6_reg_7_ ( .D(n2432), .CP(clk), .Q(r6[7]) );
  DFQD1BWP12T r6_reg_6_ ( .D(n2431), .CP(clk), .Q(r6[6]) );
  DFQD1BWP12T r6_reg_5_ ( .D(n2430), .CP(clk), .Q(r6[5]) );
  DFQD1BWP12T r6_reg_4_ ( .D(n2429), .CP(clk), .Q(r6[4]) );
  DFQD1BWP12T r6_reg_3_ ( .D(n2428), .CP(clk), .Q(r6[3]) );
  DFQD1BWP12T r6_reg_2_ ( .D(n2427), .CP(clk), .Q(r6[2]) );
  DFQD1BWP12T r6_reg_1_ ( .D(n2426), .CP(clk), .Q(r6[1]) );
  DFQD1BWP12T r6_reg_0_ ( .D(n2425), .CP(clk), .Q(r6[0]) );
  DFQD1BWP12T r7_reg_31_ ( .D(n2424), .CP(clk), .Q(r7[31]) );
  DFQD1BWP12T r7_reg_30_ ( .D(n2423), .CP(clk), .Q(r7[30]) );
  DFQD1BWP12T r7_reg_29_ ( .D(n2422), .CP(clk), .Q(r7[29]) );
  DFQD1BWP12T r7_reg_28_ ( .D(n2421), .CP(clk), .Q(r7[28]) );
  DFQD1BWP12T r7_reg_27_ ( .D(n2420), .CP(clk), .Q(r7[27]) );
  DFQD1BWP12T r7_reg_26_ ( .D(n2419), .CP(clk), .Q(r7[26]) );
  DFQD1BWP12T r7_reg_25_ ( .D(n2418), .CP(clk), .Q(r7[25]) );
  DFQD1BWP12T r7_reg_24_ ( .D(n2417), .CP(clk), .Q(r7[24]) );
  DFQD1BWP12T r7_reg_23_ ( .D(n2416), .CP(clk), .Q(r7[23]) );
  DFQD1BWP12T r7_reg_22_ ( .D(n2415), .CP(clk), .Q(r7[22]) );
  DFQD1BWP12T r7_reg_21_ ( .D(n2414), .CP(clk), .Q(r7[21]) );
  DFQD1BWP12T r7_reg_20_ ( .D(n2413), .CP(clk), .Q(r7[20]) );
  DFQD1BWP12T r7_reg_19_ ( .D(n2412), .CP(clk), .Q(r7[19]) );
  DFQD1BWP12T r7_reg_18_ ( .D(n2411), .CP(clk), .Q(r7[18]) );
  DFQD1BWP12T r7_reg_17_ ( .D(n2410), .CP(clk), .Q(r7[17]) );
  DFQD1BWP12T r7_reg_16_ ( .D(n2409), .CP(clk), .Q(r7[16]) );
  DFQD1BWP12T r7_reg_15_ ( .D(n2408), .CP(clk), .Q(r7[15]) );
  DFQD1BWP12T r7_reg_14_ ( .D(n2407), .CP(clk), .Q(r7[14]) );
  DFQD1BWP12T r7_reg_13_ ( .D(n2406), .CP(clk), .Q(r7[13]) );
  DFQD1BWP12T r7_reg_12_ ( .D(n2405), .CP(clk), .Q(r7[12]) );
  DFQD1BWP12T r7_reg_11_ ( .D(n2404), .CP(clk), .Q(r7[11]) );
  DFQD1BWP12T r7_reg_10_ ( .D(n2403), .CP(clk), .Q(r7[10]) );
  DFQD1BWP12T r7_reg_9_ ( .D(n2402), .CP(clk), .Q(r7[9]) );
  DFQD1BWP12T r7_reg_8_ ( .D(n2401), .CP(clk), .Q(r7[8]) );
  DFQD1BWP12T r7_reg_7_ ( .D(n2400), .CP(clk), .Q(r7[7]) );
  DFQD1BWP12T r7_reg_6_ ( .D(n2399), .CP(clk), .Q(r7[6]) );
  DFQD1BWP12T r7_reg_5_ ( .D(n2398), .CP(clk), .Q(r7[5]) );
  DFQD1BWP12T r7_reg_4_ ( .D(n2397), .CP(clk), .Q(r7[4]) );
  DFQD1BWP12T r7_reg_3_ ( .D(n2396), .CP(clk), .Q(r7[3]) );
  DFQD1BWP12T r7_reg_2_ ( .D(n2395), .CP(clk), .Q(r7[2]) );
  DFQD1BWP12T r7_reg_1_ ( .D(n2394), .CP(clk), .Q(r7[1]) );
  DFQD1BWP12T r7_reg_0_ ( .D(n2393), .CP(clk), .Q(r7[0]) );
  DFQD1BWP12T r8_reg_31_ ( .D(n2392), .CP(clk), .Q(r8[31]) );
  DFQD1BWP12T r8_reg_30_ ( .D(n2391), .CP(clk), .Q(r8[30]) );
  DFQD1BWP12T r8_reg_29_ ( .D(n2390), .CP(clk), .Q(r8[29]) );
  DFQD1BWP12T r8_reg_28_ ( .D(n2389), .CP(clk), .Q(r8[28]) );
  DFQD1BWP12T r8_reg_27_ ( .D(n2388), .CP(clk), .Q(r8[27]) );
  DFQD1BWP12T r8_reg_26_ ( .D(n2387), .CP(clk), .Q(r8[26]) );
  DFQD1BWP12T r8_reg_25_ ( .D(n2386), .CP(clk), .Q(r8[25]) );
  DFQD1BWP12T r8_reg_24_ ( .D(n2385), .CP(clk), .Q(r8[24]) );
  DFQD1BWP12T r8_reg_23_ ( .D(n2384), .CP(clk), .Q(r8[23]) );
  DFQD1BWP12T r8_reg_22_ ( .D(n2383), .CP(clk), .Q(r8[22]) );
  DFQD1BWP12T r8_reg_21_ ( .D(n2382), .CP(clk), .Q(r8[21]) );
  DFQD1BWP12T r8_reg_20_ ( .D(n2381), .CP(clk), .Q(r8[20]) );
  DFQD1BWP12T r8_reg_19_ ( .D(n2380), .CP(clk), .Q(r8[19]) );
  DFQD1BWP12T r8_reg_18_ ( .D(n2379), .CP(clk), .Q(r8[18]) );
  DFQD1BWP12T r8_reg_17_ ( .D(n2378), .CP(clk), .Q(r8[17]) );
  DFQD1BWP12T r8_reg_16_ ( .D(n2377), .CP(clk), .Q(r8[16]) );
  DFQD1BWP12T r8_reg_15_ ( .D(n2376), .CP(clk), .Q(r8[15]) );
  DFQD1BWP12T r8_reg_14_ ( .D(n2375), .CP(clk), .Q(r8[14]) );
  DFQD1BWP12T r8_reg_13_ ( .D(n2374), .CP(clk), .Q(r8[13]) );
  DFQD1BWP12T r8_reg_12_ ( .D(n2373), .CP(clk), .Q(r8[12]) );
  DFQD1BWP12T r8_reg_11_ ( .D(n2372), .CP(clk), .Q(r8[11]) );
  DFQD1BWP12T r8_reg_10_ ( .D(n2371), .CP(clk), .Q(r8[10]) );
  DFQD1BWP12T r8_reg_9_ ( .D(n2370), .CP(clk), .Q(r8[9]) );
  DFQD1BWP12T r8_reg_8_ ( .D(n2369), .CP(clk), .Q(r8[8]) );
  DFQD1BWP12T r8_reg_7_ ( .D(n2368), .CP(clk), .Q(r8[7]) );
  DFQD1BWP12T r8_reg_6_ ( .D(n2367), .CP(clk), .Q(r8[6]) );
  DFQD1BWP12T r8_reg_5_ ( .D(n2366), .CP(clk), .Q(r8[5]) );
  DFQD1BWP12T r8_reg_4_ ( .D(n2365), .CP(clk), .Q(r8[4]) );
  DFQD1BWP12T r8_reg_3_ ( .D(n2364), .CP(clk), .Q(r8[3]) );
  DFQD1BWP12T r8_reg_2_ ( .D(n2363), .CP(clk), .Q(r8[2]) );
  DFQD1BWP12T r8_reg_1_ ( .D(n2362), .CP(clk), .Q(r8[1]) );
  DFQD1BWP12T r8_reg_0_ ( .D(n2361), .CP(clk), .Q(r8[0]) );
  DFQD1BWP12T r9_reg_31_ ( .D(n2360), .CP(clk), .Q(r9[31]) );
  DFQD1BWP12T r9_reg_30_ ( .D(n2359), .CP(clk), .Q(r9[30]) );
  DFQD1BWP12T r9_reg_29_ ( .D(n2358), .CP(clk), .Q(r9[29]) );
  DFQD1BWP12T r9_reg_28_ ( .D(n2357), .CP(clk), .Q(r9[28]) );
  DFQD1BWP12T r9_reg_27_ ( .D(n2356), .CP(clk), .Q(r9[27]) );
  DFQD1BWP12T r9_reg_26_ ( .D(n2355), .CP(clk), .Q(r9[26]) );
  DFQD1BWP12T r9_reg_25_ ( .D(n2354), .CP(clk), .Q(r9[25]) );
  DFQD1BWP12T r9_reg_24_ ( .D(n2353), .CP(clk), .Q(r9[24]) );
  DFQD1BWP12T r9_reg_23_ ( .D(n2352), .CP(clk), .Q(r9[23]) );
  DFQD1BWP12T r9_reg_22_ ( .D(n2351), .CP(clk), .Q(r9[22]) );
  DFQD1BWP12T r9_reg_21_ ( .D(n2350), .CP(clk), .Q(r9[21]) );
  DFQD1BWP12T r9_reg_20_ ( .D(n2349), .CP(clk), .Q(r9[20]) );
  DFQD1BWP12T r9_reg_19_ ( .D(n2348), .CP(clk), .Q(r9[19]) );
  DFQD1BWP12T r9_reg_18_ ( .D(n2347), .CP(clk), .Q(r9[18]) );
  DFQD1BWP12T r9_reg_17_ ( .D(n2346), .CP(clk), .Q(r9[17]) );
  DFQD1BWP12T r9_reg_16_ ( .D(n2345), .CP(clk), .Q(r9[16]) );
  DFQD1BWP12T r9_reg_15_ ( .D(n2344), .CP(clk), .Q(r9[15]) );
  DFQD1BWP12T r9_reg_14_ ( .D(n2343), .CP(clk), .Q(r9[14]) );
  DFQD1BWP12T r9_reg_13_ ( .D(n2342), .CP(clk), .Q(r9[13]) );
  DFQD1BWP12T r9_reg_12_ ( .D(n2341), .CP(clk), .Q(r9[12]) );
  DFQD1BWP12T r9_reg_11_ ( .D(n2340), .CP(clk), .Q(r9[11]) );
  DFQD1BWP12T r9_reg_10_ ( .D(n2339), .CP(clk), .Q(r9[10]) );
  DFQD1BWP12T r9_reg_9_ ( .D(n2338), .CP(clk), .Q(r9[9]) );
  DFQD1BWP12T r9_reg_8_ ( .D(n2337), .CP(clk), .Q(r9[8]) );
  DFQD1BWP12T r9_reg_7_ ( .D(n2336), .CP(clk), .Q(r9[7]) );
  DFQD1BWP12T r9_reg_6_ ( .D(n2335), .CP(clk), .Q(r9[6]) );
  DFQD1BWP12T r9_reg_5_ ( .D(n2334), .CP(clk), .Q(r9[5]) );
  DFQD1BWP12T r9_reg_4_ ( .D(n2333), .CP(clk), .Q(r9[4]) );
  DFQD1BWP12T r9_reg_3_ ( .D(n2332), .CP(clk), .Q(r9[3]) );
  DFQD1BWP12T r9_reg_2_ ( .D(n2331), .CP(clk), .Q(r9[2]) );
  DFQD1BWP12T r9_reg_1_ ( .D(n2330), .CP(clk), .Q(r9[1]) );
  DFQD1BWP12T r9_reg_0_ ( .D(n2329), .CP(clk), .Q(r9[0]) );
  DFQD1BWP12T r10_reg_31_ ( .D(n2328), .CP(clk), .Q(r10[31]) );
  DFQD1BWP12T r10_reg_30_ ( .D(n2327), .CP(clk), .Q(r10[30]) );
  DFQD1BWP12T r10_reg_29_ ( .D(n2326), .CP(clk), .Q(r10[29]) );
  DFQD1BWP12T r10_reg_28_ ( .D(n2325), .CP(clk), .Q(r10[28]) );
  DFQD1BWP12T r10_reg_27_ ( .D(n2324), .CP(clk), .Q(r10[27]) );
  DFQD1BWP12T r10_reg_26_ ( .D(n2323), .CP(clk), .Q(r10[26]) );
  DFQD1BWP12T r10_reg_25_ ( .D(n2322), .CP(clk), .Q(r10[25]) );
  DFQD1BWP12T r10_reg_24_ ( .D(n2321), .CP(clk), .Q(r10[24]) );
  DFQD1BWP12T r10_reg_23_ ( .D(n2320), .CP(clk), .Q(r10[23]) );
  DFQD1BWP12T r10_reg_22_ ( .D(n2319), .CP(clk), .Q(r10[22]) );
  DFQD1BWP12T r10_reg_21_ ( .D(n2318), .CP(clk), .Q(r10[21]) );
  DFQD1BWP12T r10_reg_20_ ( .D(n2317), .CP(clk), .Q(r10[20]) );
  DFQD1BWP12T r10_reg_19_ ( .D(n2316), .CP(clk), .Q(r10[19]) );
  DFQD1BWP12T r10_reg_18_ ( .D(n2315), .CP(clk), .Q(r10[18]) );
  DFQD1BWP12T r10_reg_17_ ( .D(n2314), .CP(clk), .Q(r10[17]) );
  DFQD1BWP12T r10_reg_16_ ( .D(n2313), .CP(clk), .Q(r10[16]) );
  DFQD1BWP12T r10_reg_15_ ( .D(n2312), .CP(clk), .Q(r10[15]) );
  DFQD1BWP12T r10_reg_14_ ( .D(n2311), .CP(clk), .Q(r10[14]) );
  DFQD1BWP12T r10_reg_13_ ( .D(n2310), .CP(clk), .Q(r10[13]) );
  DFQD1BWP12T r10_reg_12_ ( .D(n2309), .CP(clk), .Q(r10[12]) );
  DFQD1BWP12T r10_reg_11_ ( .D(n2308), .CP(clk), .Q(r10[11]) );
  DFQD1BWP12T r10_reg_10_ ( .D(n2307), .CP(clk), .Q(r10[10]) );
  DFQD1BWP12T r10_reg_9_ ( .D(n2306), .CP(clk), .Q(r10[9]) );
  DFQD1BWP12T r10_reg_8_ ( .D(n2305), .CP(clk), .Q(r10[8]) );
  DFQD1BWP12T r10_reg_7_ ( .D(n2304), .CP(clk), .Q(r10[7]) );
  DFQD1BWP12T r10_reg_6_ ( .D(n2303), .CP(clk), .Q(r10[6]) );
  DFQD1BWP12T r10_reg_5_ ( .D(n2302), .CP(clk), .Q(r10[5]) );
  DFQD1BWP12T r10_reg_4_ ( .D(n2301), .CP(clk), .Q(r10[4]) );
  DFQD1BWP12T r10_reg_3_ ( .D(n2300), .CP(clk), .Q(r10[3]) );
  DFQD1BWP12T r10_reg_2_ ( .D(n2299), .CP(clk), .Q(r10[2]) );
  DFQD1BWP12T r10_reg_1_ ( .D(n2298), .CP(clk), .Q(r10[1]) );
  DFQD1BWP12T r10_reg_0_ ( .D(n2297), .CP(clk), .Q(r10[0]) );
  DFQD1BWP12T r11_reg_31_ ( .D(n2296), .CP(clk), .Q(r11[31]) );
  DFQD1BWP12T r11_reg_30_ ( .D(n2295), .CP(clk), .Q(r11[30]) );
  DFQD1BWP12T r11_reg_29_ ( .D(n2294), .CP(clk), .Q(r11[29]) );
  DFQD1BWP12T r11_reg_28_ ( .D(n2293), .CP(clk), .Q(r11[28]) );
  DFQD1BWP12T r11_reg_27_ ( .D(n2292), .CP(clk), .Q(r11[27]) );
  DFQD1BWP12T r11_reg_26_ ( .D(n2291), .CP(clk), .Q(r11[26]) );
  DFQD1BWP12T r11_reg_25_ ( .D(n2290), .CP(clk), .Q(r11[25]) );
  DFQD1BWP12T r11_reg_24_ ( .D(n2289), .CP(clk), .Q(r11[24]) );
  DFQD1BWP12T r11_reg_23_ ( .D(n2288), .CP(clk), .Q(r11[23]) );
  DFQD1BWP12T r11_reg_22_ ( .D(n2287), .CP(clk), .Q(r11[22]) );
  DFQD1BWP12T r11_reg_21_ ( .D(n2286), .CP(clk), .Q(r11[21]) );
  DFQD1BWP12T r11_reg_20_ ( .D(n2285), .CP(clk), .Q(r11[20]) );
  DFQD1BWP12T r11_reg_19_ ( .D(n2284), .CP(clk), .Q(r11[19]) );
  DFQD1BWP12T r11_reg_18_ ( .D(n2283), .CP(clk), .Q(r11[18]) );
  DFQD1BWP12T r11_reg_17_ ( .D(n2282), .CP(clk), .Q(r11[17]) );
  DFQD1BWP12T r11_reg_16_ ( .D(n2281), .CP(clk), .Q(r11[16]) );
  DFQD1BWP12T r11_reg_15_ ( .D(n2280), .CP(clk), .Q(r11[15]) );
  DFQD1BWP12T r11_reg_14_ ( .D(n2279), .CP(clk), .Q(r11[14]) );
  DFQD1BWP12T r11_reg_13_ ( .D(n2278), .CP(clk), .Q(r11[13]) );
  DFQD1BWP12T r11_reg_12_ ( .D(n2277), .CP(clk), .Q(r11[12]) );
  DFQD1BWP12T r11_reg_11_ ( .D(n2276), .CP(clk), .Q(r11[11]) );
  DFQD1BWP12T r11_reg_10_ ( .D(n2275), .CP(clk), .Q(r11[10]) );
  DFQD1BWP12T r11_reg_9_ ( .D(n2274), .CP(clk), .Q(r11[9]) );
  DFQD1BWP12T r11_reg_8_ ( .D(n2273), .CP(clk), .Q(r11[8]) );
  DFQD1BWP12T r11_reg_7_ ( .D(n2272), .CP(clk), .Q(r11[7]) );
  DFQD1BWP12T r11_reg_6_ ( .D(n2271), .CP(clk), .Q(r11[6]) );
  DFQD1BWP12T r11_reg_5_ ( .D(n2270), .CP(clk), .Q(r11[5]) );
  DFQD1BWP12T r11_reg_4_ ( .D(n2269), .CP(clk), .Q(r11[4]) );
  DFQD1BWP12T r11_reg_3_ ( .D(n2268), .CP(clk), .Q(r11[3]) );
  DFQD1BWP12T r11_reg_2_ ( .D(n2267), .CP(clk), .Q(r11[2]) );
  DFQD1BWP12T r11_reg_1_ ( .D(n2266), .CP(clk), .Q(r11[1]) );
  DFQD1BWP12T r11_reg_0_ ( .D(n2265), .CP(clk), .Q(r11[0]) );
  DFQD1BWP12T r12_reg_31_ ( .D(n2264), .CP(clk), .Q(r12[31]) );
  DFQD1BWP12T r12_reg_30_ ( .D(n2263), .CP(clk), .Q(r12[30]) );
  DFQD1BWP12T r12_reg_29_ ( .D(n2262), .CP(clk), .Q(r12[29]) );
  DFQD1BWP12T r12_reg_28_ ( .D(n2261), .CP(clk), .Q(r12[28]) );
  DFQD1BWP12T r12_reg_27_ ( .D(n2260), .CP(clk), .Q(r12[27]) );
  DFQD1BWP12T r12_reg_26_ ( .D(n2259), .CP(clk), .Q(r12[26]) );
  DFQD1BWP12T r12_reg_25_ ( .D(n2258), .CP(clk), .Q(r12[25]) );
  DFQD1BWP12T r12_reg_24_ ( .D(n2257), .CP(clk), .Q(r12[24]) );
  DFQD1BWP12T r12_reg_23_ ( .D(n2256), .CP(clk), .Q(r12[23]) );
  DFQD1BWP12T r12_reg_22_ ( .D(n2255), .CP(clk), .Q(r12[22]) );
  DFQD1BWP12T r12_reg_21_ ( .D(n2254), .CP(clk), .Q(r12[21]) );
  DFQD1BWP12T r12_reg_20_ ( .D(n2253), .CP(clk), .Q(r12[20]) );
  DFQD1BWP12T r12_reg_19_ ( .D(n2252), .CP(clk), .Q(r12[19]) );
  DFQD1BWP12T r12_reg_18_ ( .D(n2251), .CP(clk), .Q(r12[18]) );
  DFQD1BWP12T r12_reg_17_ ( .D(n2250), .CP(clk), .Q(r12[17]) );
  DFQD1BWP12T r12_reg_16_ ( .D(n2249), .CP(clk), .Q(r12[16]) );
  DFQD1BWP12T r12_reg_15_ ( .D(n2248), .CP(clk), .Q(r12[15]) );
  DFQD1BWP12T r12_reg_14_ ( .D(n2247), .CP(clk), .Q(r12[14]) );
  DFQD1BWP12T r12_reg_13_ ( .D(n2246), .CP(clk), .Q(r12[13]) );
  DFQD1BWP12T r12_reg_12_ ( .D(n2245), .CP(clk), .Q(r12[12]) );
  DFQD1BWP12T r12_reg_11_ ( .D(n2244), .CP(clk), .Q(r12[11]) );
  DFQD1BWP12T r12_reg_10_ ( .D(n2243), .CP(clk), .Q(r12[10]) );
  DFQD1BWP12T r12_reg_9_ ( .D(n2242), .CP(clk), .Q(r12[9]) );
  DFQD1BWP12T r12_reg_8_ ( .D(n2241), .CP(clk), .Q(r12[8]) );
  DFQD1BWP12T r12_reg_7_ ( .D(n2240), .CP(clk), .Q(r12[7]) );
  DFQD1BWP12T r12_reg_6_ ( .D(n2239), .CP(clk), .Q(r12[6]) );
  DFQD1BWP12T r12_reg_5_ ( .D(n2238), .CP(clk), .Q(r12[5]) );
  DFQD1BWP12T r12_reg_4_ ( .D(n2237), .CP(clk), .Q(r12[4]) );
  DFQD1BWP12T r12_reg_3_ ( .D(n2236), .CP(clk), .Q(r12[3]) );
  DFQD1BWP12T r12_reg_2_ ( .D(n2235), .CP(clk), .Q(r12[2]) );
  DFQD1BWP12T r12_reg_1_ ( .D(n2234), .CP(clk), .Q(r12[1]) );
  DFQD1BWP12T r12_reg_0_ ( .D(n2233), .CP(clk), .Q(r12[0]) );
  DFQD1BWP12T lr_reg_31_ ( .D(n2232), .CP(clk), .Q(lr[31]) );
  DFQD1BWP12T lr_reg_30_ ( .D(n2231), .CP(clk), .Q(lr[30]) );
  DFQD1BWP12T lr_reg_29_ ( .D(n2230), .CP(clk), .Q(lr[29]) );
  DFQD1BWP12T lr_reg_28_ ( .D(n2229), .CP(clk), .Q(lr[28]) );
  DFQD1BWP12T lr_reg_27_ ( .D(n2228), .CP(clk), .Q(lr[27]) );
  DFQD1BWP12T lr_reg_26_ ( .D(n2227), .CP(clk), .Q(lr[26]) );
  DFQD1BWP12T lr_reg_25_ ( .D(n2226), .CP(clk), .Q(lr[25]) );
  DFQD1BWP12T lr_reg_24_ ( .D(n2225), .CP(clk), .Q(lr[24]) );
  DFQD1BWP12T lr_reg_23_ ( .D(n2224), .CP(clk), .Q(lr[23]) );
  DFQD1BWP12T lr_reg_22_ ( .D(n2223), .CP(clk), .Q(lr[22]) );
  DFQD1BWP12T lr_reg_21_ ( .D(n2222), .CP(clk), .Q(lr[21]) );
  DFQD1BWP12T lr_reg_20_ ( .D(n2221), .CP(clk), .Q(lr[20]) );
  DFQD1BWP12T lr_reg_19_ ( .D(n2220), .CP(clk), .Q(lr[19]) );
  DFQD1BWP12T lr_reg_18_ ( .D(n2219), .CP(clk), .Q(lr[18]) );
  DFQD1BWP12T lr_reg_17_ ( .D(n2218), .CP(clk), .Q(lr[17]) );
  DFQD1BWP12T lr_reg_16_ ( .D(n2217), .CP(clk), .Q(lr[16]) );
  DFQD1BWP12T lr_reg_15_ ( .D(n2216), .CP(clk), .Q(lr[15]) );
  DFQD1BWP12T lr_reg_14_ ( .D(n2215), .CP(clk), .Q(lr[14]) );
  DFQD1BWP12T lr_reg_13_ ( .D(n2214), .CP(clk), .Q(lr[13]) );
  DFQD1BWP12T lr_reg_12_ ( .D(n2213), .CP(clk), .Q(lr[12]) );
  DFQD1BWP12T lr_reg_11_ ( .D(n2212), .CP(clk), .Q(lr[11]) );
  DFQD1BWP12T lr_reg_10_ ( .D(n2211), .CP(clk), .Q(lr[10]) );
  DFQD1BWP12T lr_reg_9_ ( .D(n2210), .CP(clk), .Q(lr[9]) );
  DFQD1BWP12T lr_reg_8_ ( .D(n2209), .CP(clk), .Q(lr[8]) );
  DFQD1BWP12T lr_reg_7_ ( .D(n2208), .CP(clk), .Q(lr[7]) );
  DFQD1BWP12T lr_reg_6_ ( .D(n2207), .CP(clk), .Q(lr[6]) );
  DFQD1BWP12T lr_reg_5_ ( .D(n2206), .CP(clk), .Q(lr[5]) );
  DFQD1BWP12T lr_reg_4_ ( .D(n2205), .CP(clk), .Q(lr[4]) );
  DFQD1BWP12T lr_reg_3_ ( .D(n2204), .CP(clk), .Q(lr[3]) );
  DFQD1BWP12T lr_reg_2_ ( .D(n2203), .CP(clk), .Q(lr[2]) );
  DFQD1BWP12T lr_reg_1_ ( .D(n2202), .CP(clk), .Q(lr[1]) );
  DFQD1BWP12T lr_reg_0_ ( .D(n2201), .CP(clk), .Q(lr[0]) );
  DFQD1BWP12T sp_reg_31_ ( .D(spin[31]), .CP(clk), .Q(n[2010]) );
  DFQD1BWP12T sp_reg_30_ ( .D(spin[30]), .CP(clk), .Q(n[2011]) );
  DFQD1BWP12T sp_reg_29_ ( .D(spin[29]), .CP(clk), .Q(n[2012]) );
  DFQD1BWP12T sp_reg_28_ ( .D(spin[28]), .CP(clk), .Q(n[2013]) );
  DFQD1BWP12T sp_reg_27_ ( .D(spin[27]), .CP(clk), .Q(n[2014]) );
  DFQD1BWP12T sp_reg_26_ ( .D(spin[26]), .CP(clk), .Q(n[2015]) );
  DFQD1BWP12T sp_reg_25_ ( .D(spin[25]), .CP(clk), .Q(n[2016]) );
  DFQD1BWP12T sp_reg_24_ ( .D(spin[24]), .CP(clk), .Q(n[2017]) );
  DFQD1BWP12T sp_reg_23_ ( .D(spin[23]), .CP(clk), .Q(n[2018]) );
  DFQD1BWP12T sp_reg_22_ ( .D(spin[22]), .CP(clk), .Q(n[2019]) );
  DFQD1BWP12T sp_reg_21_ ( .D(spin[21]), .CP(clk), .Q(n[2020]) );
  DFQD1BWP12T sp_reg_20_ ( .D(spin[20]), .CP(clk), .Q(n[2021]) );
  DFQD1BWP12T sp_reg_19_ ( .D(spin[19]), .CP(clk), .Q(n[2022]) );
  DFQD1BWP12T sp_reg_18_ ( .D(spin[18]), .CP(clk), .Q(n[2023]) );
  DFQD1BWP12T sp_reg_17_ ( .D(spin[17]), .CP(clk), .Q(n[2024]) );
  DFQD1BWP12T sp_reg_16_ ( .D(spin[16]), .CP(clk), .Q(n[2025]) );
  DFQD1BWP12T sp_reg_15_ ( .D(spin[15]), .CP(clk), .Q(n[2026]) );
  DFQD1BWP12T sp_reg_14_ ( .D(spin[14]), .CP(clk), .Q(n[2027]) );
  DFQD1BWP12T sp_reg_13_ ( .D(spin[13]), .CP(clk), .Q(n[2028]) );
  DFQD1BWP12T sp_reg_12_ ( .D(spin[12]), .CP(clk), .Q(n[2029]) );
  DFQD1BWP12T sp_reg_11_ ( .D(spin[11]), .CP(clk), .Q(n[2030]) );
  DFQD1BWP12T sp_reg_10_ ( .D(spin[10]), .CP(clk), .Q(n[2031]) );
  DFQD1BWP12T sp_reg_9_ ( .D(spin[9]), .CP(clk), .Q(n[2032]) );
  DFQD1BWP12T sp_reg_8_ ( .D(spin[8]), .CP(clk), .Q(n[2033]) );
  DFQD1BWP12T sp_reg_7_ ( .D(spin[7]), .CP(clk), .Q(n[2034]) );
  DFQD1BWP12T sp_reg_6_ ( .D(spin[6]), .CP(clk), .Q(n[2035]) );
  DFQD1BWP12T sp_reg_5_ ( .D(spin[5]), .CP(clk), .Q(n[2036]) );
  DFQD1BWP12T sp_reg_4_ ( .D(spin[4]), .CP(clk), .Q(n[2037]) );
  DFQD1BWP12T sp_reg_3_ ( .D(spin[3]), .CP(clk), .Q(n[2038]) );
  DFQD1BWP12T sp_reg_2_ ( .D(spin[2]), .CP(clk), .Q(n[2039]) );
  DFQD1BWP12T sp_reg_1_ ( .D(spin[1]), .CP(clk), .Q(n[2040]) );
  DFQD1BWP12T sp_reg_0_ ( .D(spin[0]), .CP(clk), .Q(n[2041]) );
  DFQD1BWP12T pc_reg_30_ ( .D(n2199), .CP(clk), .Q(pc_out[30]) );
  DFQD1BWP12T pc_reg_29_ ( .D(n2198), .CP(clk), .Q(pc_out[29]) );
  DFQD1BWP12T pc_reg_28_ ( .D(n2197), .CP(clk), .Q(pc_out[28]) );
  DFQD1BWP12T pc_reg_27_ ( .D(n2196), .CP(clk), .Q(pc_out[27]) );
  DFQD1BWP12T pc_reg_26_ ( .D(n2195), .CP(clk), .Q(pc_out[26]) );
  DFQD1BWP12T pc_reg_25_ ( .D(n2194), .CP(clk), .Q(pc_out[25]) );
  DFQD1BWP12T pc_reg_24_ ( .D(n2193), .CP(clk), .Q(pc_out[24]) );
  DFQD1BWP12T pc_reg_23_ ( .D(n2192), .CP(clk), .Q(pc_out[23]) );
  DFQD1BWP12T pc_reg_22_ ( .D(n2191), .CP(clk), .Q(pc_out[22]) );
  DFQD1BWP12T pc_reg_21_ ( .D(n2190), .CP(clk), .Q(pc_out[21]) );
  DFQD1BWP12T pc_reg_20_ ( .D(n2189), .CP(clk), .Q(pc_out[20]) );
  DFQD1BWP12T pc_reg_19_ ( .D(n2188), .CP(clk), .Q(pc_out[19]) );
  DFQD1BWP12T pc_reg_18_ ( .D(n2187), .CP(clk), .Q(pc_out[18]) );
  DFQD1BWP12T pc_reg_17_ ( .D(n2186), .CP(clk), .Q(pc_out[17]) );
  DFQD1BWP12T pc_reg_16_ ( .D(n2185), .CP(clk), .Q(pc_out[16]) );
  DFQD1BWP12T pc_reg_15_ ( .D(n2184), .CP(clk), .Q(pc_out[15]) );
  DFQD1BWP12T pc_reg_14_ ( .D(n2183), .CP(clk), .Q(pc_out[14]) );
  DFQD1BWP12T pc_reg_13_ ( .D(n2182), .CP(clk), .Q(pc_out[13]) );
  DFQD1BWP12T pc_reg_12_ ( .D(n2181), .CP(clk), .Q(pc_out[12]) );
  DFQD1BWP12T pc_reg_11_ ( .D(n2180), .CP(clk), .Q(pc_out[11]) );
  DFQD1BWP12T pc_reg_10_ ( .D(n2179), .CP(clk), .Q(pc_out[10]) );
  DFQD1BWP12T pc_reg_9_ ( .D(n2178), .CP(clk), .Q(pc_out[9]) );
  DFQD1BWP12T pc_reg_8_ ( .D(n2177), .CP(clk), .Q(pc_out[8]) );
  DFQD1BWP12T pc_reg_7_ ( .D(n2176), .CP(clk), .Q(pc_out[7]) );
  DFQD1BWP12T pc_reg_6_ ( .D(n2175), .CP(clk), .Q(pc_out[6]) );
  DFQD1BWP12T pc_reg_5_ ( .D(n2174), .CP(clk), .Q(pc_out[5]) );
  DFQD1BWP12T pc_reg_4_ ( .D(n2173), .CP(clk), .Q(pc_out[4]) );
  DFQD1BWP12T pc_reg_3_ ( .D(n2172), .CP(clk), .Q(pc_out[3]) );
  DFQD1BWP12T pc_reg_2_ ( .D(n2171), .CP(clk), .Q(pc_out[2]) );
  DFQD1BWP12T pc_reg_1_ ( .D(n2170), .CP(clk), .Q(pc_out[1]) );
  DFQD1BWP12T pc_reg_0_ ( .D(n2169), .CP(clk), .Q(pc_out[0]) );
  DFQD1BWP12T cpsr_reg_3_ ( .D(cpsrin[3]), .CP(clk), .Q(cpsr_out[3]) );
  DFQD1BWP12T cpsr_reg_2_ ( .D(cpsrin[2]), .CP(clk), .Q(cpsr_out[2]) );
  DFQD1BWP12T cpsr_reg_1_ ( .D(cpsrin[1]), .CP(clk), .Q(cpsr_out[1]) );
  DFQD1BWP12T cpsr_reg_0_ ( .D(cpsrin[0]), .CP(clk), .Q(cpsr_out[0]) );
  DFQD1BWP12T tmp1_reg_31_ ( .D(n2168), .CP(clk), .Q(tmp1[31]) );
  DFQD1BWP12T tmp1_reg_30_ ( .D(n2167), .CP(clk), .Q(tmp1[30]) );
  DFQD1BWP12T tmp1_reg_29_ ( .D(n2166), .CP(clk), .Q(tmp1[29]) );
  DFQD1BWP12T tmp1_reg_28_ ( .D(n2165), .CP(clk), .Q(tmp1[28]) );
  DFQD1BWP12T tmp1_reg_27_ ( .D(n2164), .CP(clk), .Q(tmp1[27]) );
  DFQD1BWP12T tmp1_reg_26_ ( .D(n2163), .CP(clk), .Q(tmp1[26]) );
  DFQD1BWP12T tmp1_reg_25_ ( .D(n2162), .CP(clk), .Q(tmp1[25]) );
  DFQD1BWP12T tmp1_reg_24_ ( .D(n2161), .CP(clk), .Q(tmp1[24]) );
  DFQD1BWP12T tmp1_reg_23_ ( .D(n2160), .CP(clk), .Q(tmp1[23]) );
  DFQD1BWP12T tmp1_reg_22_ ( .D(n2159), .CP(clk), .Q(tmp1[22]) );
  DFQD1BWP12T tmp1_reg_21_ ( .D(n2158), .CP(clk), .Q(tmp1[21]) );
  DFQD1BWP12T tmp1_reg_20_ ( .D(n2157), .CP(clk), .Q(tmp1[20]) );
  DFQD1BWP12T tmp1_reg_19_ ( .D(n2156), .CP(clk), .Q(tmp1[19]) );
  DFQD1BWP12T tmp1_reg_18_ ( .D(n2155), .CP(clk), .Q(tmp1[18]) );
  DFQD1BWP12T tmp1_reg_17_ ( .D(n2154), .CP(clk), .Q(tmp1[17]) );
  DFQD1BWP12T tmp1_reg_16_ ( .D(n2153), .CP(clk), .Q(tmp1[16]) );
  DFQD1BWP12T tmp1_reg_15_ ( .D(n2152), .CP(clk), .Q(tmp1[15]) );
  DFQD1BWP12T tmp1_reg_14_ ( .D(n2151), .CP(clk), .Q(tmp1[14]) );
  DFQD1BWP12T tmp1_reg_13_ ( .D(n2150), .CP(clk), .Q(tmp1[13]) );
  DFQD1BWP12T tmp1_reg_12_ ( .D(n2149), .CP(clk), .Q(tmp1[12]) );
  DFQD1BWP12T tmp1_reg_11_ ( .D(n2148), .CP(clk), .Q(tmp1[11]) );
  DFQD1BWP12T tmp1_reg_10_ ( .D(n2147), .CP(clk), .Q(tmp1[10]) );
  DFQD1BWP12T tmp1_reg_9_ ( .D(n2146), .CP(clk), .Q(tmp1[9]) );
  DFQD1BWP12T tmp1_reg_8_ ( .D(n2145), .CP(clk), .Q(tmp1[8]) );
  DFQD1BWP12T tmp1_reg_7_ ( .D(n2144), .CP(clk), .Q(tmp1[7]) );
  DFQD1BWP12T tmp1_reg_6_ ( .D(n2143), .CP(clk), .Q(tmp1[6]) );
  DFQD1BWP12T tmp1_reg_5_ ( .D(n2142), .CP(clk), .Q(tmp1[5]) );
  DFQD1BWP12T tmp1_reg_4_ ( .D(n2141), .CP(clk), .Q(tmp1[4]) );
  DFQD1BWP12T tmp1_reg_3_ ( .D(n2140), .CP(clk), .Q(tmp1[3]) );
  DFQD1BWP12T tmp1_reg_2_ ( .D(n2139), .CP(clk), .Q(tmp1[2]) );
  DFQD1BWP12T tmp1_reg_1_ ( .D(n2138), .CP(clk), .Q(tmp1[1]) );
  DFQD1BWP12T tmp1_reg_0_ ( .D(n2136), .CP(clk), .Q(tmp1[0]) );
  DFQD1BWP12T pc_reg_31_ ( .D(n2200), .CP(clk), .Q(pc_out[31]) );
  AOI22D1BWP12T U3 ( .A1(pc_out[26]), .A2(n174), .B1(n1996), .B2(r6[26]), .ZN(
        n793) );
  AOI22D1BWP12T U4 ( .A1(r3[26]), .A2(n1994), .B1(n168), .B2(lr[26]), .ZN(n795) );
  NR2D2BWP12T U5 ( .A1(readA_sel[2]), .A2(readA_sel[1]), .ZN(n128) );
  ND2D3BWP12T U6 ( .A1(n113), .A2(n119), .ZN(n139) );
  INR2D2BWP12T U7 ( .A1(readB_sel[2]), .B1(readB_sel[1]), .ZN(n172) );
  INVD1BWP12T U8 ( .I(n1370), .ZN(n1363) );
  AN2D1BWP12T U9 ( .A1(next_cpsr_in[0]), .A2(n804), .Z(cpsrin[0]) );
  OAI22D1BWP12T U10 ( .A1(n1923), .A2(n1910), .B1(n1909), .B2(n1936), .ZN(n609) );
  OAI22D1BWP12T U11 ( .A1(n1907), .A2(n1862), .B1(n1905), .B2(n1861), .ZN(n501) );
  OAI22D1BWP12T U12 ( .A1(n1915), .A2(n1852), .B1(n1913), .B2(n498), .ZN(n499)
         );
  AOI22D1BWP12T U13 ( .A1(n112), .A2(r12[5]), .B1(n273), .B2(tmp1[5]), .ZN(
        n549) );
  NR4D0BWP12T U14 ( .A1(n558), .A2(n557), .A3(n556), .A4(n555), .ZN(n559) );
  OAI22D1BWP12T U15 ( .A1(n1907), .A2(n1837), .B1(n1905), .B2(n1836), .ZN(n557) );
  INVD1BWP12T U16 ( .I(n1366), .ZN(n70) );
  INVD1BWP12T U17 ( .I(write2_in[30]), .ZN(n69) );
  ND2D1BWP12T U18 ( .A1(n745), .A2(n744), .ZN(regA_out[6]) );
  INVD3BWP12T U19 ( .I(readA_sel[4]), .ZN(n119) );
  IND2XD2BWP12T U20 ( .A1(readA_sel[2]), .B1(readA_sel[1]), .ZN(n135) );
  INVD1BWP12T U21 ( .I(n135), .ZN(n140) );
  INVD1BWP12T U22 ( .I(n97), .ZN(n1303) );
  INVD1BWP12T U23 ( .I(reset), .ZN(n804) );
  IOA21D1BWP12T U24 ( .A1(n1247), .A2(n1350), .B(n1246), .ZN(n1251) );
  AOI21D1BWP12T U25 ( .A1(n1322), .A2(n1350), .B(n1321), .ZN(n1333) );
  NR2D1BWP12T U26 ( .A1(n1355), .A2(n1377), .ZN(n1359) );
  NR2D1BWP12T U27 ( .A1(n101), .A2(n100), .ZN(n1299) );
  AN3XD1BWP12T U28 ( .A1(n348), .A2(n225), .A3(n86), .Z(n1288) );
  AN3XD1BWP12T U29 ( .A1(n228), .A2(n804), .A3(n227), .Z(n1293) );
  BUFFD2BWP12T U30 ( .I(write1_in[15]), .Z(n1245) );
  BUFFD2BWP12T U31 ( .I(write1_in[27]), .Z(n1337) );
  INVD1BWP12T U32 ( .I(readC_sel[4]), .ZN(n1208) );
  AN3XD1BWP12T U33 ( .A1(n239), .A2(n238), .A3(n237), .Z(n242) );
  AN3XD1BWP12T U34 ( .A1(n799), .A2(n798), .A3(n797), .Z(n802) );
  NR2D1BWP12T U35 ( .A1(readB_sel[1]), .A2(readB_sel[2]), .ZN(n170) );
  ND3D2BWP12T U36 ( .A1(n119), .A2(readA_sel[0]), .A3(readA_sel[3]), .ZN(n136)
         );
  INR2D2BWP12T U37 ( .A1(readB_sel[1]), .B1(readB_sel[2]), .ZN(n166) );
  NR2D2BWP12T U38 ( .A1(n127), .A2(n135), .ZN(n1803) );
  INR2XD2BWP12T U39 ( .A1(n128), .B1(n127), .ZN(n1812) );
  INVD2BWP12T U40 ( .I(n1819), .ZN(n1888) );
  INR2D4BWP12T U41 ( .A1(n121), .B1(n139), .ZN(n112) );
  INVD2BWP12T U42 ( .I(n1802), .ZN(n1893) );
  INVD2BWP12T U43 ( .I(n1989), .ZN(n1959) );
  INR2XD2BWP12T U44 ( .A1(n172), .B1(n169), .ZN(n1993) );
  INR2XD2BWP12T U45 ( .A1(n172), .B1(n173), .ZN(n1995) );
  INR2XD2BWP12T U46 ( .A1(n170), .B1(n173), .ZN(n152) );
  NR2D1BWP12T U47 ( .A1(n1339), .A2(n1338), .ZN(n1341) );
  INR2D1BWP12T U48 ( .A1(n166), .B1(n165), .ZN(n167) );
  OAI22D1BWP12T U49 ( .A1(n1911), .A2(n1949), .B1(n1948), .B2(n1886), .ZN(n216) );
  OAI22D1BWP12T U50 ( .A1(n1977), .A2(n1906), .B1(n1975), .B2(n1904), .ZN(n218) );
  OAI22D1BWP12T U51 ( .A1(n1981), .A2(n1885), .B1(n1979), .B2(n1900), .ZN(n217) );
  INVD1BWP12T U52 ( .I(n172), .ZN(n154) );
  INR2D0BWP12T U53 ( .A1(n357), .B1(n356), .ZN(n1258) );
  INR2D0BWP12T U54 ( .A1(n363), .B1(n362), .ZN(n1261) );
  MAOI22D0BWP12T U55 ( .A1(n1241), .A2(n1240), .B1(n1241), .B2(n1240), .ZN(n1)
         );
  AO222D0BWP12T U56 ( .A1(pc_out[13]), .A2(n1363), .B1(n1), .B2(n1364), .C1(
        next_pc_in[13]), .C2(n1375), .Z(n2182) );
  MAOI22D0BWP12T U57 ( .A1(n1243), .A2(n1242), .B1(n1243), .B2(n1242), .ZN(n2)
         );
  AO222D0BWP12T U58 ( .A1(pc_out[14]), .A2(n1363), .B1(n2), .B2(n1364), .C1(
        next_pc_in[14]), .C2(n1375), .Z(n2183) );
  MAOI22D0BWP12T U59 ( .A1(n1249), .A2(n1248), .B1(n1249), .B2(n1248), .ZN(n3)
         );
  AO222D0BWP12T U60 ( .A1(pc_out[15]), .A2(n1363), .B1(n3), .B2(n1364), .C1(
        next_pc_in[15]), .C2(n1375), .Z(n2184) );
  INR2D0BWP12T U61 ( .A1(n342), .B1(n341), .ZN(n1270) );
  MAOI22D0BWP12T U62 ( .A1(n1251), .A2(n1250), .B1(n1251), .B2(n1250), .ZN(n4)
         );
  AO222D0BWP12T U63 ( .A1(pc_out[16]), .A2(n1363), .B1(n4), .B2(n1364), .C1(
        next_pc_in[16]), .C2(n1375), .Z(n2185) );
  INR2D0BWP12T U64 ( .A1(n344), .B1(n343), .ZN(n1267) );
  MAOI22D0BWP12T U65 ( .A1(n1254), .A2(n1253), .B1(n1254), .B2(n1253), .ZN(n5)
         );
  AO222D0BWP12T U66 ( .A1(pc_out[17]), .A2(n1363), .B1(n5), .B2(n1364), .C1(
        next_pc_in[17]), .C2(n1375), .Z(n2186) );
  INR2D0BWP12T U67 ( .A1(n369), .B1(n368), .ZN(n1276) );
  MAOI22D0BWP12T U68 ( .A1(n1305), .A2(n1304), .B1(n1305), .B2(n1304), .ZN(n6)
         );
  AO222D0BWP12T U69 ( .A1(pc_out[18]), .A2(n1363), .B1(n6), .B2(n1364), .C1(
        next_pc_in[18]), .C2(n1375), .Z(n2187) );
  IND3D0BWP12T U70 ( .A1(write1_sel[0]), .B1(write1_sel[3]), .B2(write1_en), 
        .ZN(n96) );
  AOI22D0BWP12T U71 ( .A1(n1366), .A2(write2_in[21]), .B1(n1350), .B2(
        write1_in[21]), .ZN(n1315) );
  OA211D1BWP12T U72 ( .A1(n1806), .A2(n257), .B(n256), .C(n255), .Z(n7) );
  AN4XD1BWP12T U73 ( .A1(n258), .A2(n259), .A3(n260), .A4(n261), .Z(n8) );
  AOI22D1BWP12T U74 ( .A1(n1818), .A2(r10[26]), .B1(n1819), .B2(lr[26]), .ZN(
        n9) );
  AOI22D1BWP12T U75 ( .A1(n1817), .A2(r11[26]), .B1(n134), .B2(pc_out[26]), 
        .ZN(n10) );
  ND4D2BWP12T U76 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(regA_out[26]) );
  MAOI22D0BWP12T U77 ( .A1(n1311), .A2(n1310), .B1(n1311), .B2(n1310), .ZN(n11) );
  AO222D0BWP12T U78 ( .A1(pc_out[19]), .A2(n1363), .B1(n11), .B2(n1364), .C1(
        next_pc_in[19]), .C2(n1375), .Z(n2188) );
  INR2D1BWP12T U79 ( .A1(n98), .B1(n99), .ZN(n1302) );
  CKND0BWP12T U80 ( .I(r4[30]), .ZN(n12) );
  AOI22D0BWP12T U81 ( .A1(n1801), .A2(tmp1[30]), .B1(n112), .B2(r12[30]), .ZN(
        n13) );
  AOI22D0BWP12T U82 ( .A1(n1803), .A2(r2[30]), .B1(n1802), .B2(r1[30]), .ZN(
        n14) );
  OA211D1BWP12T U83 ( .A1(n1806), .A2(n12), .B(n13), .C(n14), .Z(n15) );
  AOI22D1BWP12T U84 ( .A1(n123), .A2(r5[30]), .B1(n1811), .B2(r3[30]), .ZN(n16) );
  AOI22D0BWP12T U85 ( .A1(n126), .A2(r7[30]), .B1(n1812), .B2(r0[30]), .ZN(n17) );
  AOI22D0BWP12T U86 ( .A1(n1809), .A2(n[2011]), .B1(n1810), .B2(r8[30]), .ZN(
        n18) );
  AOI22D0BWP12T U87 ( .A1(n120), .A2(r6[30]), .B1(n1808), .B2(r9[30]), .ZN(n19) );
  AN4XD1BWP12T U88 ( .A1(n16), .A2(n17), .A3(n18), .A4(n19), .Z(n20) );
  AOI22D1BWP12T U89 ( .A1(n1818), .A2(r10[30]), .B1(n1819), .B2(lr[30]), .ZN(
        n21) );
  AOI22D1BWP12T U90 ( .A1(n1817), .A2(r11[30]), .B1(n134), .B2(pc_out[30]), 
        .ZN(n22) );
  ND4D1BWP12T U91 ( .A1(n15), .A2(n20), .A3(n21), .A4(n22), .ZN(regA_out[30])
         );
  MAOI22D0BWP12T U92 ( .A1(n1316), .A2(n1315), .B1(n1316), .B2(n1315), .ZN(n23) );
  AO222D0BWP12T U93 ( .A1(pc_out[21]), .A2(n1363), .B1(n23), .B2(n1364), .C1(
        next_pc_in[21]), .C2(n1375), .Z(n2190) );
  AO22D0BWP12T U94 ( .A1(n1366), .A2(write2_in[10]), .B1(n1350), .B2(
        write1_in[10]), .Z(n1230) );
  INR2D1BWP12T U95 ( .A1(n101), .B1(n100), .ZN(n1300) );
  IND2D0BWP12T U96 ( .A1(n228), .B1(n227), .ZN(n467) );
  OA211D1BWP12T U97 ( .A1(n1806), .A2(n1784), .B(n1783), .C(n1782), .Z(n24) );
  AOI22D1BWP12T U98 ( .A1(n1818), .A2(r10[23]), .B1(n1819), .B2(lr[23]), .ZN(
        n25) );
  AOI22D0BWP12T U99 ( .A1(n1817), .A2(r11[23]), .B1(n134), .B2(pc_out[23]), 
        .ZN(n26) );
  ND4D1BWP12T U100 ( .A1(n24), .A2(n1789), .A3(n25), .A4(n26), .ZN(
        regA_out[23]) );
  MAOI22D0BWP12T U101 ( .A1(n1320), .A2(n1319), .B1(n1320), .B2(n1319), .ZN(
        n27) );
  AO222D0BWP12T U102 ( .A1(pc_out[22]), .A2(n1363), .B1(n27), .B2(n1364), .C1(
        next_pc_in[22]), .C2(n1375), .Z(n2191) );
  NR2D0BWP12T U103 ( .A1(write2_sel[0]), .A2(n107), .ZN(n28) );
  ND4D0BWP12T U104 ( .A1(write2_en), .A2(write2_sel[4]), .A3(write2_sel[3]), 
        .A4(n28), .ZN(n98) );
  AN2D0BWP12T U105 ( .A1(write1_sel[2]), .A2(write1_sel[1]), .Z(n102) );
  AO22D0BWP12T U106 ( .A1(n1366), .A2(write2_in[8]), .B1(n1350), .B2(
        write1_in[8]), .Z(n1226) );
  INR3D0BWP12T U107 ( .A1(n94), .B1(reset), .B2(n95), .ZN(n1290) );
  INR2D0BWP12T U108 ( .A1(n340), .B1(n339), .ZN(n1273) );
  OA211D1BWP12T U109 ( .A1(n1806), .A2(n1807), .B(n1805), .C(n1804), .Z(n29)
         );
  AOI22D1BWP12T U110 ( .A1(n1818), .A2(r10[25]), .B1(n1819), .B2(lr[25]), .ZN(
        n30) );
  AOI22D0BWP12T U111 ( .A1(n1817), .A2(r11[25]), .B1(n134), .B2(pc_out[25]), 
        .ZN(n31) );
  ND4D1BWP12T U112 ( .A1(n29), .A2(n1820), .A3(n30), .A4(n31), .ZN(
        regA_out[25]) );
  MAOI22D0BWP12T U113 ( .A1(n1331), .A2(n1333), .B1(n1331), .B2(n1333), .ZN(
        n32) );
  AO222D0BWP12T U114 ( .A1(pc_out[23]), .A2(n1363), .B1(n32), .B2(n1364), .C1(
        next_pc_in[23]), .C2(n1375), .Z(n2192) );
  NR2D0BWP12T U115 ( .A1(write1_sel[3]), .A2(n82), .ZN(n89) );
  INR3D0BWP12T U116 ( .A1(write1_sel[2]), .B1(reset), .B2(write1_sel[1]), .ZN(
        n364) );
  AO22D1BWP12T U117 ( .A1(n1366), .A2(write2_in[14]), .B1(n1350), .B2(
        write1_in[14]), .Z(n1243) );
  INR2D0BWP12T U118 ( .A1(n346), .B1(n345), .ZN(n1264) );
  AN4XD1BWP12T U119 ( .A1(n787), .A2(n788), .A3(n789), .A4(n790), .Z(n33) );
  AOI22D0BWP12T U120 ( .A1(n1989), .A2(r2[23]), .B1(n1990), .B2(r7[23]), .ZN(
        n34) );
  AOI22D0BWP12T U121 ( .A1(n152), .A2(r9[23]), .B1(n2002), .B2(r4[23]), .ZN(
        n35) );
  AOI22D1BWP12T U122 ( .A1(n1988), .A2(r5[23]), .B1(n158), .B2(r10[23]), .ZN(
        n36) );
  AN4D0BWP12T U123 ( .A1(n792), .A2(n35), .A3(n791), .A4(n36), .Z(n37) );
  ND3D1BWP12T U124 ( .A1(n33), .A2(n34), .A3(n37), .ZN(regB_out[23]) );
  IND2XD2BWP12T U125 ( .A1(n127), .B1(n121), .ZN(n1806) );
  MAOI22D0BWP12T U126 ( .A1(n1210), .A2(n1209), .B1(n1210), .B2(n1209), .ZN(
        n38) );
  AO222D0BWP12T U127 ( .A1(pc_out[2]), .A2(n1363), .B1(n1364), .B2(n38), .C1(
        next_pc_in[2]), .C2(n1375), .Z(n2171) );
  MOAI22D0BWP12T U128 ( .A1(n1326), .A2(n1332), .B1(n1326), .B2(n1332), .ZN(
        n39) );
  AO222D0BWP12T U129 ( .A1(n39), .A2(n1364), .B1(next_pc_in[24]), .B2(n1375), 
        .C1(pc_out[24]), .C2(n1363), .Z(n2193) );
  IND3D0BWP12T U130 ( .A1(n96), .B1(write1_sel[4]), .B2(n358), .ZN(n97) );
  AO222D1BWP12T U131 ( .A1(n1891), .A2(r4[20]), .B1(n112), .B2(r12[20]), .C1(
        tmp1[20]), .C2(n1801), .Z(n482) );
  INR3D0BWP12T U132 ( .A1(n79), .B1(reset), .B2(n80), .ZN(n1296) );
  AN4XD1BWP12T U133 ( .A1(n780), .A2(n781), .A3(n782), .A4(n783), .Z(n40) );
  AOI22D0BWP12T U134 ( .A1(n1989), .A2(r2[22]), .B1(n1990), .B2(r7[22]), .ZN(
        n41) );
  AOI22D1BWP12T U135 ( .A1(n158), .A2(r10[22]), .B1(n1988), .B2(r5[22]), .ZN(
        n42) );
  AN4D0BWP12T U136 ( .A1(n786), .A2(n784), .A3(n785), .A4(n42), .Z(n43) );
  ND3D1BWP12T U137 ( .A1(n40), .A2(n41), .A3(n43), .ZN(regB_out[22]) );
  AN2D0BWP12T U138 ( .A1(n804), .A2(next_cpsr_in[2]), .Z(cpsrin[2]) );
  MAOI22D0BWP12T U139 ( .A1(n230), .A2(n229), .B1(n230), .B2(n229), .ZN(n44)
         );
  AO222D0BWP12T U140 ( .A1(pc_out[3]), .A2(n1363), .B1(n44), .B2(n1364), .C1(
        next_pc_in[3]), .C2(n1375), .Z(n2172) );
  MAOI22D0BWP12T U141 ( .A1(n1223), .A2(n1222), .B1(n1223), .B2(n1222), .ZN(
        n45) );
  AO222D0BWP12T U142 ( .A1(pc_out[7]), .A2(n1363), .B1(n45), .B2(n1364), .C1(
        next_pc_in[7]), .C2(n1375), .Z(n2176) );
  MAOI22D0BWP12T U143 ( .A1(n1228), .A2(n1227), .B1(n1228), .B2(n1227), .ZN(
        n46) );
  AO222D0BWP12T U144 ( .A1(pc_out[9]), .A2(n1363), .B1(n46), .B2(n1364), .C1(
        next_pc_in[9]), .C2(n1375), .Z(n2178) );
  MAOI22D0BWP12T U145 ( .A1(n1344), .A2(n1343), .B1(n1344), .B2(n1343), .ZN(
        n47) );
  AO222D0BWP12T U146 ( .A1(pc_out[27]), .A2(n1363), .B1(n47), .B2(n1364), .C1(
        next_pc_in[27]), .C2(n1375), .Z(n2196) );
  NR2D0BWP12T U147 ( .A1(n96), .A2(write1_sel[4]), .ZN(n352) );
  AN2D0BWP12T U148 ( .A1(write1_sel[0]), .A2(n89), .Z(n359) );
  AOI22D0BWP12T U149 ( .A1(n1954), .A2(r0[0]), .B1(n1955), .B2(r11[0]), .ZN(
        n48) );
  AOI22D0BWP12T U150 ( .A1(n1953), .A2(r4[0]), .B1(n152), .B2(r9[0]), .ZN(n49)
         );
  CKND2D0BWP12T U151 ( .A1(n48), .A2(n49), .ZN(n1873) );
  OAI22D0BWP12T U152 ( .A1(write1_in[0]), .A2(n1366), .B1(write2_in[0]), .B2(
        n1350), .ZN(n50) );
  AOI22D0BWP12T U153 ( .A1(pc_out[0]), .A2(n1363), .B1(next_pc_in[0]), .B2(
        n1375), .ZN(n51) );
  OAI21D0BWP12T U154 ( .A1(n1367), .A2(n50), .B(n51), .ZN(n2169) );
  MAOI22D0BWP12T U155 ( .A1(n1213), .A2(n1212), .B1(n1213), .B2(n1212), .ZN(
        n52) );
  AO222D0BWP12T U156 ( .A1(pc_out[4]), .A2(n1363), .B1(n52), .B2(n1364), .C1(
        next_pc_in[4]), .C2(n1375), .Z(n2173) );
  MAOI22D0BWP12T U157 ( .A1(n1226), .A2(n1225), .B1(n1226), .B2(n1225), .ZN(
        n53) );
  AO222D0BWP12T U158 ( .A1(pc_out[8]), .A2(n1363), .B1(n53), .B2(n1364), .C1(
        next_pc_in[8]), .C2(n1375), .Z(n2177) );
  MAOI22D0BWP12T U159 ( .A1(n1231), .A2(n1230), .B1(n1231), .B2(n1230), .ZN(
        n54) );
  AO222D0BWP12T U160 ( .A1(pc_out[10]), .A2(n1363), .B1(n54), .B2(n1364), .C1(
        next_pc_in[10]), .C2(n1375), .Z(n2179) );
  MAOI22D0BWP12T U161 ( .A1(n1348), .A2(n1347), .B1(n1348), .B2(n1347), .ZN(
        n55) );
  AO222D0BWP12T U162 ( .A1(pc_out[28]), .A2(n1363), .B1(n55), .B2(n1364), .C1(
        next_pc_in[28]), .C2(n1375), .Z(n2197) );
  AOI22D0BWP12T U163 ( .A1(r9[30]), .A2(n1194), .B1(r10[30]), .B2(n1201), .ZN(
        n56) );
  AOI22D0BWP12T U164 ( .A1(n[2011]), .A2(n1196), .B1(lr[30]), .B2(n1197), .ZN(
        n57) );
  AOI22D0BWP12T U165 ( .A1(r4[30]), .A2(n1182), .B1(r7[30]), .B2(n1183), .ZN(
        n58) );
  AOI22D0BWP12T U166 ( .A1(r6[30]), .A2(n1184), .B1(r2[30]), .B2(n1185), .ZN(
        n59) );
  AOI22D0BWP12T U167 ( .A1(r1[30]), .A2(n1186), .B1(r5[30]), .B2(n1187), .ZN(
        n60) );
  AOI22D0BWP12T U168 ( .A1(r0[30]), .A2(n1189), .B1(r3[30]), .B2(n1188), .ZN(
        n61) );
  ND4D0BWP12T U169 ( .A1(n58), .A2(n59), .A3(n60), .A4(n61), .ZN(n62) );
  MOAI22D0BWP12T U170 ( .A1(n1356), .A2(n883), .B1(r8[30]), .B2(n1195), .ZN(
        n63) );
  CKND0BWP12T U171 ( .I(r12[30]), .ZN(n64) );
  CKND0BWP12T U172 ( .I(r11[30]), .ZN(n65) );
  OAI22D0BWP12T U173 ( .A1(n1172), .A2(n64), .B1(n1112), .B2(n65), .ZN(n66) );
  AOI211D0BWP12T U174 ( .A1(n1208), .A2(n62), .B(n63), .C(n66), .ZN(n67) );
  ND3D0BWP12T U175 ( .A1(n56), .A2(n57), .A3(n67), .ZN(regC_out[30]) );
  TPND2D2BWP12T U176 ( .A1(n1348), .A2(n1347), .ZN(n1362) );
  AOI21D4BWP12T U177 ( .A1(n1337), .A2(n1350), .B(n1336), .ZN(n1343) );
  BUFFXD8BWP12T U178 ( .I(write1_in[30]), .Z(n1352) );
  TPNR2D2BWP12T U179 ( .A1(n1344), .A2(n1343), .ZN(n1348) );
  CKND2D2BWP12T U180 ( .A1(n1335), .A2(n1334), .ZN(n1344) );
  TPNR2D2BWP12T U181 ( .A1(n1223), .A2(n1222), .ZN(n1225) );
  TPND2D2BWP12T U182 ( .A1(n1354), .A2(n1364), .ZN(n1377) );
  CKND2D2BWP12T U183 ( .A1(n600), .A2(n599), .ZN(regA_out[11]) );
  MUX2D1BWP12T U184 ( .I0(n69), .I1(n68), .S(n70), .Z(n1353) );
  INVD18BWP12T U185 ( .I(n1352), .ZN(n68) );
  INR2XD2BWP12T U186 ( .A1(n170), .B1(n165), .ZN(n164) );
  TPNR2D2BWP12T U187 ( .A1(n127), .A2(n133), .ZN(n120) );
  ND4D2BWP12T U188 ( .A1(n756), .A2(n755), .A3(n754), .A4(n753), .ZN(
        regB_out[21]) );
  ND4D2BWP12T U189 ( .A1(n243), .A2(n242), .A3(n241), .A4(n240), .ZN(
        regB_out[27]) );
  TPNR2D3BWP12T U190 ( .A1(n125), .A2(n133), .ZN(n126) );
  INR2XD2BWP12T U191 ( .A1(n170), .B1(n169), .ZN(n171) );
  INR2XD2BWP12T U192 ( .A1(n166), .B1(n169), .ZN(n158) );
  ND4D2BWP12T U193 ( .A1(n779), .A2(n778), .A3(n777), .A4(n776), .ZN(
        regB_out[25]) );
  ND4D2BWP12T U194 ( .A1(n768), .A2(n767), .A3(n766), .A4(n765), .ZN(
        regB_out[24]) );
  INR2XD2BWP12T U195 ( .A1(n138), .B1(n136), .ZN(n134) );
  NR2D3BWP12T U196 ( .A1(n125), .A2(n122), .ZN(n123) );
  INR2XD2BWP12T U197 ( .A1(n175), .B1(n169), .ZN(n168) );
  INR2XD2BWP12T U198 ( .A1(n175), .B1(n173), .ZN(n174) );
  INR2D2BWP12T U199 ( .A1(readB_sel[0]), .B1(n149), .ZN(n150) );
  INR2D2BWP12T U200 ( .A1(n170), .B1(n177), .ZN(n236) );
  BUFFD2BWP12T U201 ( .I(n236), .Z(n1954) );
  ND2D1BWP12T U202 ( .A1(n364), .A2(n352), .ZN(n460) );
  INVD1BWP12T U203 ( .I(n460), .ZN(n1286) );
  BUFFD2BWP12T U204 ( .I(write1_in[28]), .Z(n1346) );
  INR2D1BWP12T U205 ( .A1(write2_en), .B1(write2_sel[4]), .ZN(n77) );
  INR2D1BWP12T U206 ( .A1(n77), .B1(write2_sel[0]), .ZN(n91) );
  AN2XD1BWP12T U207 ( .A1(n91), .A2(write2_sel[3]), .Z(n355) );
  INR2D1BWP12T U208 ( .A1(write2_sel[2]), .B1(write2_sel[1]), .ZN(n366) );
  CKND2D1BWP12T U209 ( .A1(n355), .A2(n366), .ZN(n73) );
  INVD1BWP12T U210 ( .I(n73), .ZN(n71) );
  ND2D1BWP12T U211 ( .A1(n460), .A2(n804), .ZN(n72) );
  NR2D1BWP12T U212 ( .A1(n71), .A2(n72), .ZN(n1285) );
  NR2D1BWP12T U213 ( .A1(n73), .A2(n72), .ZN(n1284) );
  AO222D1BWP12T U214 ( .A1(n1286), .A2(n1346), .B1(n1285), .B2(r12[28]), .C1(
        write2_in[28]), .C2(n1284), .Z(n2261) );
  INR2D1BWP12T U215 ( .A1(n102), .B1(reset), .ZN(n358) );
  ND2D1BWP12T U216 ( .A1(n358), .A2(n352), .ZN(n473) );
  INVD1BWP12T U217 ( .I(n473), .ZN(n1280) );
  ND2D1BWP12T U218 ( .A1(write2_sel[2]), .A2(write2_sel[1]), .ZN(n107) );
  INVD1BWP12T U219 ( .I(n107), .ZN(n360) );
  ND2D1BWP12T U220 ( .A1(n355), .A2(n360), .ZN(n76) );
  INVD1BWP12T U221 ( .I(n76), .ZN(n74) );
  ND2D1BWP12T U222 ( .A1(n473), .A2(n804), .ZN(n75) );
  NR2D1BWP12T U223 ( .A1(n74), .A2(n75), .ZN(n1279) );
  NR2D1BWP12T U224 ( .A1(n76), .A2(n75), .ZN(n1278) );
  AO222D1BWP12T U225 ( .A1(n1280), .A2(n1346), .B1(n1279), .B2(lr[28]), .C1(
        write2_in[28]), .C2(n1278), .Z(n2229) );
  IND2XD1BWP12T U226 ( .A1(write1_sel[4]), .B1(write1_en), .ZN(n82) );
  INVD1BWP12T U227 ( .I(n359), .ZN(n78) );
  IND2D1BWP12T U228 ( .A1(write1_sel[2]), .B1(write1_sel[1]), .ZN(n92) );
  INVD1BWP12T U229 ( .I(n92), .ZN(n226) );
  ND2D1BWP12T U230 ( .A1(n226), .A2(n804), .ZN(n224) );
  NR2D1BWP12T U231 ( .A1(n78), .A2(n224), .ZN(n1298) );
  BUFFD2BWP12T U232 ( .I(write1_in[20]), .Z(n1309) );
  AN2XD1BWP12T U233 ( .A1(write2_sel[0]), .A2(n77), .Z(n84) );
  INVD1BWP12T U234 ( .I(write2_sel[3]), .ZN(n90) );
  AN2XD1BWP12T U235 ( .A1(n84), .A2(n90), .Z(n361) );
  INVD1BWP12T U236 ( .I(write2_sel[1]), .ZN(n85) );
  NR3D1BWP12T U237 ( .A1(n85), .A2(reset), .A3(write2_sel[2]), .ZN(n225) );
  CKND2D1BWP12T U238 ( .A1(n361), .A2(n225), .ZN(n79) );
  NR2D1BWP12T U239 ( .A1(n78), .A2(n92), .ZN(n80) );
  NR2D1BWP12T U240 ( .A1(n79), .A2(n80), .ZN(n1297) );
  AO222D0BWP12T U241 ( .A1(n1298), .A2(n1309), .B1(n1297), .B2(write2_in[20]), 
        .C1(n1296), .C2(r3[20]), .Z(n2541) );
  CKND2D1BWP12T U242 ( .A1(write1_sel[3]), .A2(write1_sel[0]), .ZN(n81) );
  NR2D1BWP12T U243 ( .A1(n82), .A2(n81), .ZN(n347) );
  CKND0BWP12T U244 ( .I(n347), .ZN(n83) );
  NR2D1BWP12T U245 ( .A1(n83), .A2(n224), .ZN(n1289) );
  ND2D1BWP12T U246 ( .A1(n84), .A2(write2_sel[3]), .ZN(n108) );
  INVD1BWP12T U247 ( .I(n108), .ZN(n348) );
  TPND2D0BWP12T U248 ( .A1(n347), .A2(n226), .ZN(n86) );
  NR2D0BWP12T U249 ( .A1(n85), .A2(write2_sel[2]), .ZN(n88) );
  INVD1BWP12T U250 ( .I(n86), .ZN(n87) );
  AOI211D1BWP12T U251 ( .A1(n348), .A2(n88), .B(reset), .C(n87), .ZN(n1287) );
  AO222D0BWP12T U252 ( .A1(n1289), .A2(n1309), .B1(n1288), .B2(write2_in[20]), 
        .C1(n1287), .C2(r11[20]), .Z(n2285) );
  INR2D1BWP12T U253 ( .A1(n89), .B1(write1_sel[0]), .ZN(n365) );
  INVD1BWP12T U254 ( .I(n365), .ZN(n93) );
  NR2D1BWP12T U255 ( .A1(n93), .A2(n224), .ZN(n1292) );
  AN2XD1BWP12T U256 ( .A1(n91), .A2(n90), .Z(n367) );
  CKND2D1BWP12T U257 ( .A1(n367), .A2(n225), .ZN(n94) );
  NR2D1BWP12T U258 ( .A1(n93), .A2(n92), .ZN(n95) );
  NR2D1BWP12T U259 ( .A1(n94), .A2(n95), .ZN(n1291) );
  AO222D0BWP12T U260 ( .A1(n1292), .A2(n1309), .B1(n1291), .B2(write2_in[20]), 
        .C1(n1290), .C2(r2[20]), .Z(n2573) );
  BUFFD2BWP12T U261 ( .I(write1_in[19]), .Z(n1307) );
  ND2D1BWP12T U262 ( .A1(n97), .A2(n804), .ZN(n99) );
  NR2D1BWP12T U263 ( .A1(n99), .A2(n98), .ZN(n757) );
  AO222D1BWP12T U264 ( .A1(n1303), .A2(n1307), .B1(n757), .B2(write2_in[19]), 
        .C1(n1302), .C2(tmp1[19]), .Z(n2156) );
  BUFFD2BWP12T U265 ( .I(write1_in[18]), .Z(n1256) );
  AO222D1BWP12T U266 ( .A1(n1303), .A2(n1256), .B1(n757), .B2(write2_in[18]), 
        .C1(n1302), .C2(tmp1[18]), .Z(n2155) );
  ND2D1BWP12T U267 ( .A1(n347), .A2(n364), .ZN(n470) );
  INVD1BWP12T U268 ( .I(n470), .ZN(n1301) );
  ND2D1BWP12T U269 ( .A1(n348), .A2(n366), .ZN(n101) );
  ND2D1BWP12T U270 ( .A1(n470), .A2(n804), .ZN(n100) );
  AO222D1BWP12T U271 ( .A1(n1301), .A2(n1256), .B1(n1300), .B2(n[2023]), .C1(
        write2_in[18]), .C2(n1299), .Z(spin[18]) );
  AO222D1BWP12T U272 ( .A1(n1303), .A2(write1_in[21]), .B1(n757), .B2(
        write2_in[21]), .C1(n1302), .C2(tmp1[21]), .Z(n2158) );
  CKND2D2BWP12T U273 ( .A1(n347), .A2(n102), .ZN(n1366) );
  INVD2BWP12T U274 ( .I(n1366), .ZN(n1350) );
  AN2XD0BWP12T U275 ( .A1(write2_in[3]), .A2(n1366), .Z(n103) );
  AOI21D1BWP12T U276 ( .A1(write1_in[3]), .A2(n1350), .B(n103), .ZN(n230) );
  CKND2D0BWP12T U277 ( .A1(write2_in[2]), .A2(n1366), .ZN(n104) );
  IOA21D2BWP12T U278 ( .A1(write1_in[2]), .A2(n1350), .B(n104), .ZN(n1210) );
  CKND2D0BWP12T U279 ( .A1(write2_in[1]), .A2(n1366), .ZN(n105) );
  IOA21D1BWP12T U280 ( .A1(write1_in[1]), .A2(n1350), .B(n105), .ZN(n1209) );
  TPND2D1BWP12T U281 ( .A1(n1210), .A2(n1209), .ZN(n229) );
  NR2D1BWP12T U282 ( .A1(n230), .A2(n229), .ZN(n1213) );
  CKND2D0BWP12T U283 ( .A1(write2_in[4]), .A2(n1366), .ZN(n106) );
  IOA21D1BWP12T U284 ( .A1(write1_in[4]), .A2(n1350), .B(n106), .ZN(n1212) );
  OAI21D1BWP12T U285 ( .A1(n108), .A2(n107), .B(n1366), .ZN(n1178) );
  ND2D1BWP12T U286 ( .A1(n1178), .A2(n804), .ZN(n1367) );
  INVD2BWP12T U287 ( .I(n1367), .ZN(n1364) );
  NR2D1BWP12T U288 ( .A1(n1178), .A2(reset), .ZN(n110) );
  INVD1BWP12T U289 ( .I(n110), .ZN(n109) );
  NR2D2BWP12T U290 ( .A1(next_pc_en_BAR), .A2(n109), .ZN(n1375) );
  ND2D1BWP12T U291 ( .A1(next_pc_en_BAR), .A2(n110), .ZN(n1370) );
  INVD1BWP12T U292 ( .I(r4[28]), .ZN(n118) );
  TPNR2D3BWP12T U293 ( .A1(readA_sel[0]), .A2(readA_sel[3]), .ZN(n111) );
  TPND2D2BWP12T U294 ( .A1(n111), .A2(n119), .ZN(n127) );
  INR2D4BWP12T U295 ( .A1(readA_sel[2]), .B1(readA_sel[1]), .ZN(n121) );
  INR2D4BWP12T U296 ( .A1(readA_sel[3]), .B1(readA_sel[0]), .ZN(n113) );
  ND2D3BWP12T U297 ( .A1(readA_sel[2]), .A2(readA_sel[1]), .ZN(n133) );
  INVD2BWP12T U298 ( .I(n113), .ZN(n114) );
  INR3D2BWP12T U299 ( .A1(readA_sel[4]), .B1(n133), .B2(n114), .ZN(n273) );
  BUFFD2BWP12T U300 ( .I(n273), .Z(n1801) );
  AOI22D1BWP12T U301 ( .A1(n112), .A2(r12[28]), .B1(n1801), .B2(tmp1[28]), 
        .ZN(n117) );
  TPNR2D1BWP12T U302 ( .A1(readA_sel[4]), .A2(readA_sel[3]), .ZN(n115) );
  CKND2D2BWP12T U303 ( .A1(n115), .A2(readA_sel[0]), .ZN(n125) );
  INR2D4BWP12T U304 ( .A1(n128), .B1(n125), .ZN(n1802) );
  AOI22D0BWP12T U305 ( .A1(r2[28]), .A2(n1803), .B1(n1802), .B2(r1[28]), .ZN(
        n116) );
  OA211D1BWP12T U306 ( .A1(n118), .A2(n1806), .B(n117), .C(n116), .Z(n144) );
  INR2D4BWP12T U307 ( .A1(n128), .B1(n136), .ZN(n1808) );
  AOI22D1BWP12T U308 ( .A1(r9[28]), .A2(n1808), .B1(n120), .B2(r6[28]), .ZN(
        n132) );
  INR2D8BWP12T U309 ( .A1(n128), .B1(n139), .ZN(n1810) );
  INR2D4BWP12T U310 ( .A1(n121), .B1(n136), .ZN(n1809) );
  AOI22D1BWP12T U311 ( .A1(r8[28]), .A2(n1810), .B1(n1809), .B2(n[2013]), .ZN(
        n131) );
  INVD2BWP12T U312 ( .I(n121), .ZN(n122) );
  TPNR2D1BWP12T U313 ( .A1(n125), .A2(n135), .ZN(n124) );
  BUFFXD4BWP12T U314 ( .I(n124), .Z(n1811) );
  AOI22D1BWP12T U315 ( .A1(r5[28]), .A2(n123), .B1(n1811), .B2(r3[28]), .ZN(
        n130) );
  RCAOI22D0BWP12T U316 ( .A1(r7[28]), .A2(n126), .B1(n1812), .B2(r0[28]), .ZN(
        n129) );
  AN4XD1BWP12T U317 ( .A1(n132), .A2(n131), .A3(n130), .A4(n129), .Z(n143) );
  INVD2P3BWP12T U318 ( .I(n133), .ZN(n138) );
  INR2XD2BWP12T U319 ( .A1(n140), .B1(n136), .ZN(n137) );
  BUFFXD4BWP12T U320 ( .I(n137), .Z(n1817) );
  AOI22D1BWP12T U321 ( .A1(pc_out[28]), .A2(n134), .B1(n1817), .B2(r11[28]), 
        .ZN(n142) );
  INR2D8BWP12T U322 ( .A1(n138), .B1(n139), .ZN(n1819) );
  INR2XD2BWP12T U323 ( .A1(n140), .B1(n139), .ZN(n1818) );
  AOI22D1BWP12T U324 ( .A1(lr[28]), .A2(n1819), .B1(n1818), .B2(r10[28]), .ZN(
        n141) );
  ND4D2BWP12T U325 ( .A1(n144), .A2(n143), .A3(n142), .A4(n141), .ZN(
        regA_out[28]) );
  INVD1BWP12T U326 ( .I(tmp1[8]), .ZN(n151) );
  INVD1BWP12T U327 ( .I(readB_sel[0]), .ZN(n148) );
  INVD2BWP12T U328 ( .I(readB_sel[1]), .ZN(n145) );
  INR2D4BWP12T U329 ( .A1(readB_sel[2]), .B1(n145), .ZN(n175) );
  CKND2BWP12T U330 ( .I(readB_sel[3]), .ZN(n146) );
  INR2D2BWP12T U331 ( .A1(readB_sel[4]), .B1(n146), .ZN(n147) );
  TPND2D2BWP12T U332 ( .A1(n175), .A2(n147), .ZN(n149) );
  INR2D2BWP12T U333 ( .A1(n148), .B1(n149), .ZN(n2001) );
  INVD3BWP12T U334 ( .I(n2001), .ZN(n1951) );
  MOAI22D0BWP12T U335 ( .A1(n151), .A2(n1951), .B1(n150), .B2(immediate2_in[8]), .ZN(n163) );
  INVD4BWP12T U336 ( .I(readB_sel[4]), .ZN(n157) );
  ND3D2BWP12T U337 ( .A1(n157), .A2(readB_sel[3]), .A3(readB_sel[0]), .ZN(n173) );
  NR2D1BWP12T U338 ( .A1(readB_sel[3]), .A2(readB_sel[0]), .ZN(n153) );
  TPND2D4BWP12T U339 ( .A1(n153), .A2(n157), .ZN(n177) );
  TPNR2D3BWP12T U340 ( .A1(n177), .A2(n154), .ZN(n235) );
  BUFFD2BWP12T U341 ( .I(n235), .Z(n1732) );
  AOI22D1BWP12T U342 ( .A1(r9[8]), .A2(n152), .B1(n1732), .B2(r4[8]), .ZN(n156) );
  INR2XD2BWP12T U343 ( .A1(n166), .B1(n173), .ZN(n1955) );
  BUFFD3BWP12T U344 ( .I(n236), .Z(n1733) );
  AOI22D1BWP12T U345 ( .A1(r11[8]), .A2(n1955), .B1(n1733), .B2(r0[8]), .ZN(
        n155) );
  ND2D1BWP12T U346 ( .A1(n156), .A2(n155), .ZN(n162) );
  INVD1BWP12T U347 ( .I(r5[8]), .ZN(n1697) );
  IND3D4BWP12T U348 ( .A1(readB_sel[3]), .B1(readB_sel[0]), .B2(n157), .ZN(
        n165) );
  INR2XD2BWP12T U349 ( .A1(n172), .B1(n165), .ZN(n1988) );
  CKND4BWP12T U350 ( .I(n1988), .ZN(n1949) );
  IND3D4BWP12T U351 ( .A1(readB_sel[0]), .B1(readB_sel[3]), .B2(n157), .ZN(
        n169) );
  INVD4BWP12T U352 ( .I(n158), .ZN(n1948) );
  INVD1BWP12T U353 ( .I(r10[8]), .ZN(n1682) );
  OAI22D1BWP12T U354 ( .A1(n1697), .A2(n1949), .B1(n1948), .B2(n1682), .ZN(
        n161) );
  INR2D4BWP12T U355 ( .A1(n175), .B1(n165), .ZN(n1990) );
  INVD2BWP12T U356 ( .I(n1990), .ZN(n1961) );
  INVD1BWP12T U357 ( .I(r7[8]), .ZN(n1699) );
  INVD2BWP12T U358 ( .I(n166), .ZN(n159) );
  NR2XD3BWP12T U359 ( .A1(n177), .A2(n159), .ZN(n1989) );
  INVD1BWP12T U360 ( .I(r2[8]), .ZN(n1687) );
  OAI22D1BWP12T U361 ( .A1(n1961), .A2(n1699), .B1(n1959), .B2(n1687), .ZN(
        n160) );
  NR4D0BWP12T U362 ( .A1(n163), .A2(n162), .A3(n161), .A4(n160), .ZN(n183) );
  INVD1BWP12T U363 ( .I(r1[8]), .ZN(n1686) );
  INVD3BWP12T U364 ( .I(n164), .ZN(n1968) );
  INVD2BWP12T U365 ( .I(n1993), .ZN(n1967) );
  INVD1BWP12T U366 ( .I(r12[8]), .ZN(n937) );
  OAI22D1BWP12T U367 ( .A1(n1686), .A2(n1968), .B1(n1967), .B2(n937), .ZN(n181) );
  INVD1BWP12T U368 ( .I(r3[8]), .ZN(n1696) );
  BUFFXD8BWP12T U369 ( .I(n167), .Z(n1994) );
  INVD2BWP12T U370 ( .I(n1994), .ZN(n1972) );
  INVD6BWP12T U371 ( .I(n168), .ZN(n1971) );
  INVD1BWP12T U372 ( .I(lr[8]), .ZN(n1683) );
  OAI22D1BWP12T U373 ( .A1(n1696), .A2(n1972), .B1(n1971), .B2(n1683), .ZN(
        n180) );
  INVD2BWP12T U374 ( .I(n171), .ZN(n1977) );
  INVD1BWP12T U375 ( .I(r8[8]), .ZN(n1695) );
  INVD3BWP12T U376 ( .I(n1995), .ZN(n1975) );
  INVD1BWP12T U377 ( .I(n[2033]), .ZN(n1694) );
  OAI22D1BWP12T U378 ( .A1(n1977), .A2(n1695), .B1(n1975), .B2(n1694), .ZN(
        n179) );
  INVD8BWP12T U379 ( .I(n174), .ZN(n1981) );
  INVD1BWP12T U380 ( .I(pc_out[8]), .ZN(n1681) );
  INVD3BWP12T U381 ( .I(n175), .ZN(n176) );
  TPNR2D8BWP12T U382 ( .A1(n177), .A2(n176), .ZN(n1996) );
  INVD3BWP12T U383 ( .I(n1996), .ZN(n1979) );
  INVD1BWP12T U384 ( .I(r6[8]), .ZN(n1692) );
  OAI22D1BWP12T U385 ( .A1(n1981), .A2(n1681), .B1(n1979), .B2(n1692), .ZN(
        n178) );
  NR4D0BWP12T U386 ( .A1(n181), .A2(n180), .A3(n179), .A4(n178), .ZN(n182) );
  CKND2D1BWP12T U387 ( .A1(n183), .A2(n182), .ZN(regB_out[8]) );
  INVD0BWP12T U388 ( .I(tmp1[11]), .ZN(n184) );
  MOAI22D0BWP12T U389 ( .A1(n184), .A2(n1951), .B1(n150), .B2(
        immediate2_in[11]), .ZN(n190) );
  AOI22D1BWP12T U390 ( .A1(r9[11]), .A2(n152), .B1(n1732), .B2(r4[11]), .ZN(
        n186) );
  CKBD1BWP12T U391 ( .I(n1955), .Z(n2003) );
  AOI22D1BWP12T U392 ( .A1(r11[11]), .A2(n2003), .B1(n1733), .B2(r0[11]), .ZN(
        n185) );
  ND2D1BWP12T U393 ( .A1(n186), .A2(n185), .ZN(n189) );
  INVD1BWP12T U394 ( .I(r5[11]), .ZN(n592) );
  INVD1BWP12T U395 ( .I(r10[11]), .ZN(n579) );
  OAI22D1BWP12T U396 ( .A1(n592), .A2(n1949), .B1(n1948), .B2(n579), .ZN(n188)
         );
  INVD1BWP12T U397 ( .I(r7[11]), .ZN(n594) );
  INVD1BWP12T U398 ( .I(r2[11]), .ZN(n583) );
  OAI22D1BWP12T U399 ( .A1(n1961), .A2(n594), .B1(n1959), .B2(n583), .ZN(n187)
         );
  NR4D0BWP12T U400 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(n196) );
  INVD1BWP12T U401 ( .I(r1[11]), .ZN(n582) );
  INVD1BWP12T U402 ( .I(r12[11]), .ZN(n1089) );
  OAI22D1BWP12T U403 ( .A1(n582), .A2(n1968), .B1(n1967), .B2(n1089), .ZN(n194) );
  INVD1BWP12T U404 ( .I(r3[11]), .ZN(n591) );
  INVD1BWP12T U405 ( .I(lr[11]), .ZN(n580) );
  OAI22D1BWP12T U406 ( .A1(n591), .A2(n1972), .B1(n1971), .B2(n580), .ZN(n193)
         );
  INVD1BWP12T U407 ( .I(r8[11]), .ZN(n590) );
  INVD1BWP12T U408 ( .I(n[2030]), .ZN(n1090) );
  OAI22D1BWP12T U409 ( .A1(n1977), .A2(n590), .B1(n1975), .B2(n1090), .ZN(n192) );
  INVD1BWP12T U410 ( .I(pc_out[11]), .ZN(n578) );
  INVD1BWP12T U411 ( .I(r6[11]), .ZN(n588) );
  OAI22D1BWP12T U412 ( .A1(n1981), .A2(n578), .B1(n1979), .B2(n588), .ZN(n191)
         );
  NR4D0BWP12T U413 ( .A1(n194), .A2(n193), .A3(n192), .A4(n191), .ZN(n195) );
  CKND2D1BWP12T U414 ( .A1(n196), .A2(n195), .ZN(regB_out[11]) );
  INVD1BWP12T U415 ( .I(tmp1[10]), .ZN(n197) );
  MOAI22D0BWP12T U416 ( .A1(n197), .A2(n1951), .B1(n150), .B2(
        immediate2_in[10]), .ZN(n203) );
  AOI22D1BWP12T U417 ( .A1(r9[10]), .A2(n152), .B1(n1732), .B2(r4[10]), .ZN(
        n199) );
  AOI22D1BWP12T U418 ( .A1(r11[10]), .A2(n1955), .B1(n1733), .B2(r0[10]), .ZN(
        n198) );
  ND2D1BWP12T U419 ( .A1(n199), .A2(n198), .ZN(n202) );
  INVD1BWP12T U420 ( .I(r5[10]), .ZN(n1671) );
  INVD1BWP12T U421 ( .I(r10[10]), .ZN(n1657) );
  OAI22D1BWP12T U422 ( .A1(n1671), .A2(n1949), .B1(n1948), .B2(n1657), .ZN(
        n201) );
  INVD1BWP12T U423 ( .I(r7[10]), .ZN(n1673) );
  INVD1BWP12T U424 ( .I(r2[10]), .ZN(n1661) );
  OAI22D1BWP12T U425 ( .A1(n1961), .A2(n1673), .B1(n1959), .B2(n1661), .ZN(
        n200) );
  NR4D0BWP12T U426 ( .A1(n203), .A2(n202), .A3(n201), .A4(n200), .ZN(n209) );
  INVD1BWP12T U427 ( .I(r1[10]), .ZN(n1660) );
  INVD1BWP12T U428 ( .I(r12[10]), .ZN(n397) );
  OAI22D1BWP12T U429 ( .A1(n1660), .A2(n1968), .B1(n1967), .B2(n397), .ZN(n207) );
  INVD1BWP12T U430 ( .I(r3[10]), .ZN(n1670) );
  INVD1BWP12T U431 ( .I(lr[10]), .ZN(n1658) );
  OAI22D1BWP12T U432 ( .A1(n1670), .A2(n1972), .B1(n1971), .B2(n1658), .ZN(
        n206) );
  INVD1BWP12T U433 ( .I(r8[10]), .ZN(n1669) );
  INVD1BWP12T U434 ( .I(n[2031]), .ZN(n1668) );
  OAI22D1BWP12T U435 ( .A1(n1977), .A2(n1669), .B1(n1975), .B2(n1668), .ZN(
        n205) );
  INVD1BWP12T U436 ( .I(pc_out[10]), .ZN(n1656) );
  INVD1BWP12T U437 ( .I(r6[10]), .ZN(n1666) );
  OAI22D1BWP12T U438 ( .A1(n1981), .A2(n1656), .B1(n1979), .B2(n1666), .ZN(
        n204) );
  NR4D0BWP12T U439 ( .A1(n207), .A2(n206), .A3(n205), .A4(n204), .ZN(n208) );
  CKND2D1BWP12T U440 ( .A1(n209), .A2(n208), .ZN(regB_out[10]) );
  INVD1BWP12T U441 ( .I(r5[4]), .ZN(n1911) );
  INVD1BWP12T U442 ( .I(r10[4]), .ZN(n1886) );
  INVD1BWP12T U443 ( .I(tmp1[4]), .ZN(n210) );
  MOAI22D0BWP12T U444 ( .A1(n210), .A2(n1951), .B1(n150), .B2(immediate2_in[4]), .ZN(n215) );
  BUFFD2BWP12T U445 ( .I(n235), .Z(n1953) );
  AOI22D1BWP12T U446 ( .A1(r9[4]), .A2(n152), .B1(n1953), .B2(r4[4]), .ZN(n212) );
  AOI22D1BWP12T U447 ( .A1(r11[4]), .A2(n1955), .B1(n1954), .B2(r0[4]), .ZN(
        n211) );
  ND2D1BWP12T U448 ( .A1(n212), .A2(n211), .ZN(n214) );
  INVD1BWP12T U449 ( .I(r7[4]), .ZN(n1914) );
  INVD1BWP12T U450 ( .I(r2[4]), .ZN(n1894) );
  OAI22D1BWP12T U451 ( .A1(n1961), .A2(n1914), .B1(n1959), .B2(n1894), .ZN(
        n213) );
  NR4D0BWP12T U452 ( .A1(n216), .A2(n215), .A3(n214), .A4(n213), .ZN(n222) );
  INVD1BWP12T U453 ( .I(r1[4]), .ZN(n1892) );
  INVD1BWP12T U454 ( .I(r12[4]), .ZN(n419) );
  OAI22D1BWP12T U455 ( .A1(n1892), .A2(n1968), .B1(n1967), .B2(n419), .ZN(n220) );
  INVD1BWP12T U456 ( .I(r3[4]), .ZN(n1908) );
  INVD1BWP12T U457 ( .I(lr[4]), .ZN(n1889) );
  OAI22D1BWP12T U458 ( .A1(n1908), .A2(n1972), .B1(n1971), .B2(n1889), .ZN(
        n219) );
  INVD1BWP12T U459 ( .I(r8[4]), .ZN(n1906) );
  INVD1BWP12T U460 ( .I(n[2037]), .ZN(n1904) );
  INVD1BWP12T U461 ( .I(pc_out[4]), .ZN(n1885) );
  INVD1BWP12T U462 ( .I(r6[4]), .ZN(n1900) );
  NR4D0BWP12T U463 ( .A1(n220), .A2(n219), .A3(n218), .A4(n217), .ZN(n221) );
  ND2D1BWP12T U464 ( .A1(n222), .A2(n221), .ZN(regB_out[4]) );
  AN2XD1BWP12T U465 ( .A1(next_cpsr_in[3]), .A2(n804), .Z(cpsrin[3]) );
  CKND0BWP12T U466 ( .I(n352), .ZN(n223) );
  NR2D1BWP12T U467 ( .A1(n224), .A2(n223), .ZN(n1295) );
  CKND2D1BWP12T U468 ( .A1(n355), .A2(n225), .ZN(n228) );
  TPND2D0BWP12T U469 ( .A1(n226), .A2(n352), .ZN(n227) );
  INVD1BWP12T U470 ( .I(n467), .ZN(n1294) );
  AO222D1BWP12T U471 ( .A1(n1295), .A2(write1_in[17]), .B1(n1294), .B2(
        write2_in[17]), .C1(n1293), .C2(r10[17]), .Z(n2314) );
  AO222D0BWP12T U472 ( .A1(n1303), .A2(write1_in[14]), .B1(n757), .B2(
        write2_in[14]), .C1(n1302), .C2(tmp1[14]), .Z(n2151) );
  AOI22D1BWP12T U473 ( .A1(r1[27]), .A2(n164), .B1(n1993), .B2(r12[27]), .ZN(
        n234) );
  AOI22D1BWP12T U474 ( .A1(r3[27]), .A2(n1994), .B1(n168), .B2(lr[27]), .ZN(
        n233) );
  AOI22D1BWP12T U475 ( .A1(r8[27]), .A2(n171), .B1(n1995), .B2(n[2014]), .ZN(
        n232) );
  AOI22D1BWP12T U476 ( .A1(pc_out[27]), .A2(n174), .B1(n1996), .B2(r6[27]), 
        .ZN(n231) );
  AN4XD1BWP12T U477 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .Z(n243) );
  AOI22D1BWP12T U478 ( .A1(tmp1[27]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[27]), .ZN(n239) );
  BUFFXD4BWP12T U479 ( .I(n235), .Z(n2002) );
  AOI22D1BWP12T U480 ( .A1(r9[27]), .A2(n152), .B1(n2002), .B2(r4[27]), .ZN(
        n238) );
  AOI22D1BWP12T U481 ( .A1(r11[27]), .A2(n2003), .B1(n1954), .B2(r0[27]), .ZN(
        n237) );
  AOI22D1BWP12T U482 ( .A1(r5[27]), .A2(n1988), .B1(n158), .B2(r10[27]), .ZN(
        n241) );
  AOI22D1BWP12T U483 ( .A1(r7[27]), .A2(n1990), .B1(n1989), .B2(r2[27]), .ZN(
        n240) );
  AOI22D1BWP12T U484 ( .A1(r1[31]), .A2(n164), .B1(n1993), .B2(r12[31]), .ZN(
        n247) );
  AOI22D1BWP12T U485 ( .A1(r3[31]), .A2(n1994), .B1(n168), .B2(lr[31]), .ZN(
        n246) );
  AOI22D1BWP12T U486 ( .A1(r8[31]), .A2(n171), .B1(n1995), .B2(n[2010]), .ZN(
        n245) );
  AOI22D1BWP12T U487 ( .A1(pc_out[31]), .A2(n174), .B1(n1996), .B2(r6[31]), 
        .ZN(n244) );
  AN4XD1BWP12T U488 ( .A1(n247), .A2(n246), .A3(n245), .A4(n244), .Z(n254) );
  AOI22D1BWP12T U489 ( .A1(tmp1[31]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[31]), .ZN(n250) );
  AOI22D1BWP12T U490 ( .A1(r9[31]), .A2(n152), .B1(n2002), .B2(r4[31]), .ZN(
        n249) );
  AOI22D1BWP12T U491 ( .A1(r11[31]), .A2(n2003), .B1(n1954), .B2(r0[31]), .ZN(
        n248) );
  AN3XD1BWP12T U492 ( .A1(n250), .A2(n249), .A3(n248), .Z(n253) );
  AOI22D1BWP12T U493 ( .A1(r5[31]), .A2(n1988), .B1(n158), .B2(r10[31]), .ZN(
        n252) );
  AOI22D1BWP12T U494 ( .A1(r7[31]), .A2(n1990), .B1(n1989), .B2(r2[31]), .ZN(
        n251) );
  ND4D2BWP12T U495 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(
        regB_out[31]) );
  INVD1BWP12T U496 ( .I(r4[26]), .ZN(n257) );
  AOI22D1BWP12T U497 ( .A1(n112), .A2(r12[26]), .B1(n1801), .B2(tmp1[26]), 
        .ZN(n256) );
  AOI22D1BWP12T U498 ( .A1(r2[26]), .A2(n1803), .B1(n1802), .B2(r1[26]), .ZN(
        n255) );
  AOI22D1BWP12T U499 ( .A1(r9[26]), .A2(n1808), .B1(n120), .B2(r6[26]), .ZN(
        n261) );
  AOI22D1BWP12T U500 ( .A1(r8[26]), .A2(n1810), .B1(n1809), .B2(n[2015]), .ZN(
        n260) );
  AOI22D1BWP12T U501 ( .A1(r5[26]), .A2(n123), .B1(n1811), .B2(r3[26]), .ZN(
        n259) );
  AOI22D1BWP12T U502 ( .A1(r7[26]), .A2(n126), .B1(n1812), .B2(r0[26]), .ZN(
        n258) );
  INVD1BWP12T U503 ( .I(pc_out[9]), .ZN(n631) );
  INVD6BWP12T U504 ( .I(n134), .ZN(n1884) );
  INVD6BWP12T U505 ( .I(n1817), .ZN(n1883) );
  INVD1BWP12T U506 ( .I(r11[9]), .ZN(n380) );
  OAI22D1BWP12T U507 ( .A1(n631), .A2(n1884), .B1(n1883), .B2(n380), .ZN(n266)
         );
  INVD1BWP12T U508 ( .I(lr[9]), .ZN(n627) );
  DCCKND8BWP12T U509 ( .I(n1818), .ZN(n1887) );
  INVD1BWP12T U510 ( .I(r10[9]), .ZN(n617) );
  OAI22D1BWP12T U511 ( .A1(n627), .A2(n1888), .B1(n1887), .B2(n617), .ZN(n265)
         );
  INVD3BWP12T U512 ( .I(n1806), .ZN(n1891) );
  BUFFD2BWP12T U513 ( .I(n273), .Z(n1684) );
  AOI22D1BWP12T U514 ( .A1(n112), .A2(r12[9]), .B1(n1684), .B2(tmp1[9]), .ZN(
        n262) );
  IOA21D1BWP12T U515 ( .A1(n1891), .A2(r4[9]), .B(n262), .ZN(n264) );
  INVD3BWP12T U516 ( .I(n1803), .ZN(n1895) );
  INVD1BWP12T U517 ( .I(r2[9]), .ZN(n619) );
  INVD1BWP12T U518 ( .I(r1[9]), .ZN(n626) );
  OAI22D1BWP12T U519 ( .A1(n1895), .A2(n619), .B1(n1893), .B2(n626), .ZN(n263)
         );
  NR4D0BWP12T U520 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(n272) );
  INVD3BWP12T U521 ( .I(n1808), .ZN(n1903) );
  INVD1BWP12T U522 ( .I(r9[9]), .ZN(n1053) );
  INVD4BWP12T U523 ( .I(n120), .ZN(n1901) );
  INVD1BWP12T U524 ( .I(r6[9]), .ZN(n630) );
  OAI22D1BWP12T U525 ( .A1(n1903), .A2(n1053), .B1(n1901), .B2(n630), .ZN(n270) );
  INVD3BWP12T U526 ( .I(n1810), .ZN(n1907) );
  INVD1BWP12T U527 ( .I(r8[9]), .ZN(n1054) );
  INVD3BWP12T U528 ( .I(n1809), .ZN(n1905) );
  INVD1BWP12T U529 ( .I(n[2032]), .ZN(n629) );
  OAI22D1BWP12T U530 ( .A1(n1907), .A2(n1054), .B1(n1905), .B2(n629), .ZN(n269) );
  INVD1BWP12T U531 ( .I(r5[9]), .ZN(n618) );
  INVD6BWP12T U532 ( .I(n123), .ZN(n1910) );
  INVD4BWP12T U533 ( .I(n1811), .ZN(n1909) );
  INVD1BWP12T U534 ( .I(r3[9]), .ZN(n628) );
  OAI22D1BWP12T U535 ( .A1(n618), .A2(n1910), .B1(n1909), .B2(n628), .ZN(n268)
         );
  INVD3BWP12T U536 ( .I(n126), .ZN(n1915) );
  INVD1BWP12T U537 ( .I(r7[9]), .ZN(n620) );
  INVD3BWP12T U538 ( .I(n1812), .ZN(n1913) );
  INVD1BWP12T U539 ( .I(r0[9]), .ZN(n382) );
  OAI22D1BWP12T U540 ( .A1(n1915), .A2(n620), .B1(n1913), .B2(n382), .ZN(n267)
         );
  NR4D0BWP12T U541 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(n271) );
  TPND2D1BWP12T U542 ( .A1(n272), .A2(n271), .ZN(regA_out[9]) );
  INVD1BWP12T U543 ( .I(pc_out[2]), .ZN(n1980) );
  INVD1BWP12T U544 ( .I(r11[2]), .ZN(n403) );
  OAI22D1BWP12T U545 ( .A1(n1980), .A2(n1884), .B1(n1883), .B2(n403), .ZN(n278) );
  INVD1BWP12T U546 ( .I(lr[2]), .ZN(n1970) );
  INVD1BWP12T U547 ( .I(r10[2]), .ZN(n1947) );
  OAI22D1BWP12T U548 ( .A1(n1970), .A2(n1888), .B1(n1887), .B2(n1947), .ZN(
        n277) );
  AOI22D1BWP12T U549 ( .A1(n112), .A2(r12[2]), .B1(n273), .B2(tmp1[2]), .ZN(
        n274) );
  IOA21D1BWP12T U550 ( .A1(n1891), .A2(r4[2]), .B(n274), .ZN(n276) );
  INVD1BWP12T U551 ( .I(r2[2]), .ZN(n1958) );
  INVD1BWP12T U552 ( .I(r1[2]), .ZN(n1969) );
  OAI22D1BWP12T U553 ( .A1(n1895), .A2(n1958), .B1(n1893), .B2(n1969), .ZN(
        n275) );
  NR4D0BWP12T U554 ( .A1(n278), .A2(n277), .A3(n276), .A4(n275), .ZN(n284) );
  INVD1BWP12T U555 ( .I(r9[2]), .ZN(n381) );
  INVD1BWP12T U556 ( .I(r6[2]), .ZN(n1978) );
  OAI22D1BWP12T U557 ( .A1(n1903), .A2(n381), .B1(n1901), .B2(n1978), .ZN(n282) );
  INVD1BWP12T U558 ( .I(r8[2]), .ZN(n1976) );
  INVD1BWP12T U559 ( .I(n[2039]), .ZN(n1974) );
  OAI22D1BWP12T U560 ( .A1(n1907), .A2(n1976), .B1(n1905), .B2(n1974), .ZN(
        n281) );
  INVD1BWP12T U561 ( .I(r5[2]), .ZN(n1950) );
  INVD1BWP12T U562 ( .I(r3[2]), .ZN(n1973) );
  OAI22D1BWP12T U563 ( .A1(n1950), .A2(n1910), .B1(n1909), .B2(n1973), .ZN(
        n280) );
  INVD1BWP12T U564 ( .I(r7[2]), .ZN(n1960) );
  INVD1BWP12T U565 ( .I(r0[2]), .ZN(n828) );
  OAI22D1BWP12T U566 ( .A1(n1915), .A2(n1960), .B1(n1913), .B2(n828), .ZN(n279) );
  NR4D0BWP12T U567 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(n283) );
  ND2D1BWP12T U568 ( .A1(n284), .A2(n283), .ZN(regA_out[2]) );
  NR2D1BWP12T U569 ( .A1(readD_sel[1]), .A2(readD_sel[0]), .ZN(n298) );
  INVD1BWP12T U570 ( .I(n298), .ZN(n289) );
  IND2D1BWP12T U571 ( .A1(readD_sel[2]), .B1(readD_sel[3]), .ZN(n288) );
  NR2D1BWP12T U572 ( .A1(n289), .A2(n288), .ZN(n705) );
  IND2D1BWP12T U573 ( .A1(readD_sel[3]), .B1(readD_sel[2]), .ZN(n287) );
  NR2D1BWP12T U574 ( .A1(n289), .A2(n287), .ZN(n704) );
  AOI22D0BWP12T U575 ( .A1(r8[12]), .A2(n705), .B1(n704), .B2(r4[12]), .ZN(
        n286) );
  ND2D1BWP12T U576 ( .A1(readD_sel[3]), .A2(readD_sel[2]), .ZN(n300) );
  IND2D1BWP12T U577 ( .A1(readD_sel[1]), .B1(readD_sel[0]), .ZN(n294) );
  NR2D1BWP12T U578 ( .A1(n300), .A2(n294), .ZN(n707) );
  IND2D1BWP12T U579 ( .A1(readD_sel[0]), .B1(readD_sel[1]), .ZN(n296) );
  NR2D1BWP12T U580 ( .A1(n288), .A2(n296), .ZN(n706) );
  AOI22D0BWP12T U581 ( .A1(n[2029]), .A2(n707), .B1(n706), .B2(r10[12]), .ZN(
        n285) );
  CKND2D1BWP12T U582 ( .A1(n286), .A2(n285), .ZN(n305) );
  ND2D1BWP12T U583 ( .A1(readD_sel[1]), .A2(readD_sel[0]), .ZN(n299) );
  NR2D1BWP12T U584 ( .A1(n299), .A2(n287), .ZN(n711) );
  NR2D1BWP12T U585 ( .A1(n294), .A2(n287), .ZN(n710) );
  AOI22D0BWP12T U586 ( .A1(r7[12]), .A2(n711), .B1(n710), .B2(r5[12]), .ZN(
        n293) );
  NR2D1BWP12T U587 ( .A1(n300), .A2(n296), .ZN(n713) );
  NR2D1BWP12T U588 ( .A1(n288), .A2(n294), .ZN(n712) );
  AOI22D0BWP12T U589 ( .A1(lr[12]), .A2(n713), .B1(n712), .B2(r9[12]), .ZN(
        n292) );
  NR2D1BWP12T U590 ( .A1(n296), .A2(n287), .ZN(n715) );
  NR2D1BWP12T U591 ( .A1(n288), .A2(n299), .ZN(n714) );
  AOI22D0BWP12T U592 ( .A1(r6[12]), .A2(n715), .B1(n714), .B2(r11[12]), .ZN(
        n291) );
  NR2D1BWP12T U593 ( .A1(n300), .A2(n289), .ZN(n716) );
  CKND2D0BWP12T U594 ( .A1(n716), .A2(r12[12]), .ZN(n290) );
  ND4D1BWP12T U595 ( .A1(n293), .A2(n292), .A3(n291), .A4(n290), .ZN(n304) );
  INVD1BWP12T U596 ( .I(r1[12]), .ZN(n1642) );
  NR2D1BWP12T U597 ( .A1(readD_sel[3]), .A2(readD_sel[2]), .ZN(n297) );
  INVD1BWP12T U598 ( .I(n297), .ZN(n295) );
  OR2XD1BWP12T U599 ( .A1(n294), .A2(n295), .Z(n727) );
  NR2D1BWP12T U600 ( .A1(n299), .A2(n295), .ZN(n722) );
  NR2D1BWP12T U601 ( .A1(n296), .A2(n295), .ZN(n721) );
  AOI22D0BWP12T U602 ( .A1(r3[12]), .A2(n722), .B1(n721), .B2(r2[12]), .ZN(
        n302) );
  AN2XD1BWP12T U603 ( .A1(n298), .A2(n297), .Z(n724) );
  NR2D1BWP12T U604 ( .A1(n300), .A2(n299), .ZN(n723) );
  AOI22D0BWP12T U605 ( .A1(n724), .A2(r0[12]), .B1(pc_out[12]), .B2(n723), 
        .ZN(n301) );
  OAI211D0BWP12T U606 ( .A1(n1642), .A2(n727), .B(n302), .C(n301), .ZN(n303)
         );
  INVD1BWP12T U607 ( .I(readD_sel[4]), .ZN(n728) );
  OA31D0BWP12T U608 ( .A1(n305), .A2(n304), .A3(n303), .B(n728), .Z(
        regD_out[12]) );
  AOI22D0BWP12T U609 ( .A1(r8[11]), .A2(n705), .B1(n704), .B2(r4[11]), .ZN(
        n307) );
  AOI22D0BWP12T U610 ( .A1(n[2030]), .A2(n707), .B1(n706), .B2(r10[11]), .ZN(
        n306) );
  CKND2D1BWP12T U611 ( .A1(n307), .A2(n306), .ZN(n316) );
  AOI22D0BWP12T U612 ( .A1(r7[11]), .A2(n711), .B1(n710), .B2(r5[11]), .ZN(
        n311) );
  AOI22D0BWP12T U613 ( .A1(lr[11]), .A2(n713), .B1(n712), .B2(r9[11]), .ZN(
        n310) );
  AOI22D0BWP12T U614 ( .A1(r6[11]), .A2(n715), .B1(n714), .B2(r11[11]), .ZN(
        n309) );
  CKND2D0BWP12T U615 ( .A1(n716), .A2(r12[11]), .ZN(n308) );
  ND4D1BWP12T U616 ( .A1(n311), .A2(n310), .A3(n309), .A4(n308), .ZN(n315) );
  AOI22D0BWP12T U617 ( .A1(r3[11]), .A2(n722), .B1(n721), .B2(r2[11]), .ZN(
        n313) );
  AOI22D0BWP12T U618 ( .A1(n724), .A2(r0[11]), .B1(pc_out[11]), .B2(n723), 
        .ZN(n312) );
  OAI211D0BWP12T U619 ( .A1(n582), .A2(n727), .B(n313), .C(n312), .ZN(n314) );
  OA31D0BWP12T U620 ( .A1(n316), .A2(n315), .A3(n314), .B(n728), .Z(
        regD_out[11]) );
  AOI22D0BWP12T U621 ( .A1(r8[7]), .A2(n705), .B1(n704), .B2(r4[7]), .ZN(n318)
         );
  AOI22D0BWP12T U622 ( .A1(n[2034]), .A2(n707), .B1(n706), .B2(r10[7]), .ZN(
        n317) );
  CKND2D1BWP12T U623 ( .A1(n318), .A2(n317), .ZN(n327) );
  AOI22D0BWP12T U624 ( .A1(r7[7]), .A2(n711), .B1(n710), .B2(r5[7]), .ZN(n322)
         );
  AOI22D0BWP12T U625 ( .A1(lr[7]), .A2(n713), .B1(n712), .B2(r9[7]), .ZN(n321)
         );
  AOI22D0BWP12T U626 ( .A1(r6[7]), .A2(n715), .B1(n714), .B2(r11[7]), .ZN(n320) );
  CKND2D0BWP12T U627 ( .A1(n716), .A2(r12[7]), .ZN(n319) );
  ND4D1BWP12T U628 ( .A1(n322), .A2(n321), .A3(n320), .A4(n319), .ZN(n326) );
  INVD1BWP12T U629 ( .I(r1[7]), .ZN(n1718) );
  AOI22D0BWP12T U630 ( .A1(r3[7]), .A2(n722), .B1(n721), .B2(r2[7]), .ZN(n324)
         );
  AOI22D0BWP12T U631 ( .A1(n724), .A2(r0[7]), .B1(pc_out[7]), .B2(n723), .ZN(
        n323) );
  OAI211D0BWP12T U632 ( .A1(n1718), .A2(n727), .B(n324), .C(n323), .ZN(n325)
         );
  OA31D0BWP12T U633 ( .A1(n327), .A2(n326), .A3(n325), .B(n728), .Z(
        regD_out[7]) );
  AOI22D0BWP12T U634 ( .A1(r8[9]), .A2(n705), .B1(n704), .B2(r4[9]), .ZN(n329)
         );
  AOI22D0BWP12T U635 ( .A1(n[2032]), .A2(n707), .B1(n706), .B2(r10[9]), .ZN(
        n328) );
  CKND2D1BWP12T U636 ( .A1(n329), .A2(n328), .ZN(n338) );
  AOI22D0BWP12T U637 ( .A1(r7[9]), .A2(n711), .B1(n710), .B2(r5[9]), .ZN(n333)
         );
  AOI22D0BWP12T U638 ( .A1(lr[9]), .A2(n713), .B1(n712), .B2(r9[9]), .ZN(n332)
         );
  AOI22D0BWP12T U639 ( .A1(r6[9]), .A2(n715), .B1(n714), .B2(r11[9]), .ZN(n331) );
  CKND2D0BWP12T U640 ( .A1(n716), .A2(r12[9]), .ZN(n330) );
  ND4D1BWP12T U641 ( .A1(n333), .A2(n332), .A3(n331), .A4(n330), .ZN(n337) );
  AOI22D0BWP12T U642 ( .A1(r3[9]), .A2(n722), .B1(n721), .B2(r2[9]), .ZN(n335)
         );
  AOI22D0BWP12T U643 ( .A1(n724), .A2(r0[9]), .B1(pc_out[9]), .B2(n723), .ZN(
        n334) );
  OAI211D0BWP12T U644 ( .A1(n626), .A2(n727), .B(n335), .C(n334), .ZN(n336) );
  OA31D0BWP12T U645 ( .A1(n338), .A2(n337), .A3(n336), .B(n728), .Z(
        regD_out[9]) );
  INR3D0BWP12T U646 ( .A1(n804), .B1(write1_sel[2]), .B2(write1_sel[1]), .ZN(
        n353) );
  ND2D1BWP12T U647 ( .A1(n359), .A2(n353), .ZN(n457) );
  INVD1BWP12T U648 ( .I(n457), .ZN(n1274) );
  NR2D1BWP12T U649 ( .A1(write2_sel[2]), .A2(write2_sel[1]), .ZN(n354) );
  CKND2D1BWP12T U650 ( .A1(n361), .A2(n354), .ZN(n340) );
  ND2D1BWP12T U651 ( .A1(n457), .A2(n804), .ZN(n339) );
  NR2D1BWP12T U652 ( .A1(n340), .A2(n339), .ZN(n1272) );
  AO222D1BWP12T U653 ( .A1(n1274), .A2(n1352), .B1(n1273), .B2(r1[30]), .C1(
        write2_in[30]), .C2(n1272), .Z(n2615) );
  ND2D1BWP12T U654 ( .A1(n365), .A2(n358), .ZN(n451) );
  INVD1BWP12T U655 ( .I(n451), .ZN(n1271) );
  ND2D1BWP12T U656 ( .A1(n367), .A2(n360), .ZN(n342) );
  ND2D1BWP12T U657 ( .A1(n451), .A2(n804), .ZN(n341) );
  NR2D1BWP12T U658 ( .A1(n342), .A2(n341), .ZN(n1269) );
  AO222D1BWP12T U659 ( .A1(n1271), .A2(n1352), .B1(n1270), .B2(r6[30]), .C1(
        write2_in[30]), .C2(n1269), .Z(n2455) );
  AO222D1BWP12T U660 ( .A1(n1280), .A2(n1352), .B1(n1279), .B2(lr[30]), .C1(
        write2_in[30]), .C2(n1278), .Z(n2231) );
  ND2D1BWP12T U661 ( .A1(n359), .A2(n364), .ZN(n441) );
  INVD1BWP12T U662 ( .I(n441), .ZN(n1268) );
  CKND2D1BWP12T U663 ( .A1(n361), .A2(n366), .ZN(n344) );
  ND2D1BWP12T U664 ( .A1(n441), .A2(n804), .ZN(n343) );
  NR2D1BWP12T U665 ( .A1(n344), .A2(n343), .ZN(n1266) );
  AO222D1BWP12T U666 ( .A1(n1268), .A2(n1352), .B1(n1267), .B2(r5[30]), .C1(
        write2_in[30]), .C2(n1266), .Z(n2487) );
  AO222D1BWP12T U667 ( .A1(n1289), .A2(n1352), .B1(n1288), .B2(write2_in[30]), 
        .C1(n1287), .C2(r11[30]), .Z(n2295) );
  ND2D1BWP12T U668 ( .A1(n365), .A2(n353), .ZN(n448) );
  INVD1BWP12T U669 ( .I(n448), .ZN(n1265) );
  CKND2D1BWP12T U670 ( .A1(n367), .A2(n354), .ZN(n346) );
  ND2D1BWP12T U671 ( .A1(n448), .A2(n804), .ZN(n345) );
  NR2D1BWP12T U672 ( .A1(n346), .A2(n345), .ZN(n1263) );
  AO222D1BWP12T U673 ( .A1(n1265), .A2(n1352), .B1(n1264), .B2(r0[30]), .C1(
        write2_in[30]), .C2(n1263), .Z(n2647) );
  ND2D1BWP12T U674 ( .A1(n347), .A2(n353), .ZN(n463) );
  INVD1BWP12T U675 ( .I(n463), .ZN(n1283) );
  CKND2D1BWP12T U676 ( .A1(n348), .A2(n354), .ZN(n351) );
  INVD1BWP12T U677 ( .I(n351), .ZN(n349) );
  ND2D1BWP12T U678 ( .A1(n463), .A2(n804), .ZN(n350) );
  NR2D1BWP12T U679 ( .A1(n349), .A2(n350), .ZN(n1282) );
  NR2D1BWP12T U680 ( .A1(n351), .A2(n350), .ZN(n1281) );
  AO222D1BWP12T U681 ( .A1(n1283), .A2(n1352), .B1(n1282), .B2(r9[30]), .C1(
        write2_in[30]), .C2(n1281), .Z(n2359) );
  AO222D1BWP12T U682 ( .A1(n1303), .A2(n1352), .B1(n757), .B2(write2_in[30]), 
        .C1(n1302), .C2(tmp1[30]), .Z(n2167) );
  ND2D1BWP12T U683 ( .A1(n353), .A2(n352), .ZN(n432) );
  INVD1BWP12T U684 ( .I(n432), .ZN(n1259) );
  CKND2D1BWP12T U685 ( .A1(n355), .A2(n354), .ZN(n357) );
  ND2D1BWP12T U686 ( .A1(n432), .A2(n804), .ZN(n356) );
  NR2D1BWP12T U687 ( .A1(n357), .A2(n356), .ZN(n1257) );
  AO222D1BWP12T U688 ( .A1(n1259), .A2(n1352), .B1(n1258), .B2(r8[30]), .C1(
        write2_in[30]), .C2(n1257), .Z(n2391) );
  AO222D1BWP12T U689 ( .A1(n1301), .A2(n1352), .B1(n1300), .B2(n[2011]), .C1(
        write2_in[30]), .C2(n1299), .Z(spin[30]) );
  AO222D1BWP12T U690 ( .A1(n1286), .A2(n1352), .B1(n1285), .B2(r12[30]), .C1(
        write2_in[30]), .C2(n1284), .Z(n2263) );
  AO222D1BWP12T U691 ( .A1(n1295), .A2(n1352), .B1(n1294), .B2(write2_in[30]), 
        .C1(n1293), .C2(r10[30]), .Z(n2327) );
  ND2D1BWP12T U692 ( .A1(n359), .A2(n358), .ZN(n438) );
  INVD1BWP12T U693 ( .I(n438), .ZN(n1262) );
  ND2D1BWP12T U694 ( .A1(n361), .A2(n360), .ZN(n363) );
  ND2D1BWP12T U695 ( .A1(n438), .A2(n804), .ZN(n362) );
  NR2D1BWP12T U696 ( .A1(n363), .A2(n362), .ZN(n1260) );
  AO222D1BWP12T U697 ( .A1(n1262), .A2(n1352), .B1(n1261), .B2(r7[30]), .C1(
        write2_in[30]), .C2(n1260), .Z(n2423) );
  ND2D1BWP12T U698 ( .A1(n365), .A2(n364), .ZN(n444) );
  INVD1BWP12T U699 ( .I(n444), .ZN(n1277) );
  CKND2D1BWP12T U700 ( .A1(n367), .A2(n366), .ZN(n369) );
  ND2D1BWP12T U701 ( .A1(n444), .A2(n804), .ZN(n368) );
  NR2D1BWP12T U702 ( .A1(n369), .A2(n368), .ZN(n1275) );
  AO222D1BWP12T U703 ( .A1(n1277), .A2(n1352), .B1(n1276), .B2(r4[30]), .C1(
        write2_in[30]), .C2(n1275), .Z(n2519) );
  AO222D1BWP12T U704 ( .A1(n1303), .A2(n1346), .B1(n757), .B2(write2_in[28]), 
        .C1(n1302), .C2(tmp1[28]), .Z(n2165) );
  AO222D1BWP12T U705 ( .A1(n1301), .A2(n1346), .B1(n1300), .B2(n[2013]), .C1(
        write2_in[28]), .C2(n1299), .Z(spin[28]) );
  AO222D1BWP12T U706 ( .A1(n1295), .A2(n1346), .B1(n1294), .B2(write2_in[28]), 
        .C1(n1293), .C2(r10[28]), .Z(n2325) );
  BUFFXD4BWP12T U707 ( .I(write1_in[23]), .Z(n1322) );
  AO222D1BWP12T U708 ( .A1(n1295), .A2(n1322), .B1(n1294), .B2(write2_in[23]), 
        .C1(n1293), .C2(r10[23]), .Z(n2320) );
  AO222D0BWP12T U709 ( .A1(n1271), .A2(n1309), .B1(n1270), .B2(r6[20]), .C1(
        write2_in[20]), .C2(n1269), .Z(n2445) );
  AO222D0BWP12T U710 ( .A1(n1280), .A2(n1309), .B1(n1279), .B2(lr[20]), .C1(
        write2_in[20]), .C2(n1278), .Z(n2221) );
  AO222D0BWP12T U711 ( .A1(n1262), .A2(n1309), .B1(n1261), .B2(r7[20]), .C1(
        write2_in[20]), .C2(n1260), .Z(n2413) );
  AO222D0BWP12T U712 ( .A1(n1268), .A2(n1307), .B1(n1267), .B2(r5[19]), .C1(
        write2_in[19]), .C2(n1266), .Z(n2476) );
  AO222D0BWP12T U713 ( .A1(n1271), .A2(n1256), .B1(n1270), .B2(r6[18]), .C1(
        write2_in[18]), .C2(n1269), .Z(n2443) );
  AO222D0BWP12T U714 ( .A1(n1283), .A2(write1_in[17]), .B1(n1282), .B2(r9[17]), 
        .C1(write2_in[17]), .C2(n1281), .Z(n2346) );
  AO222D0BWP12T U715 ( .A1(n1259), .A2(n1256), .B1(n1258), .B2(r8[18]), .C1(
        write2_in[18]), .C2(n1257), .Z(n2379) );
  AO222D0BWP12T U716 ( .A1(n1283), .A2(n1307), .B1(n1282), .B2(r9[19]), .C1(
        write2_in[19]), .C2(n1281), .Z(n2348) );
  AO222D0BWP12T U717 ( .A1(n1289), .A2(write1_in[17]), .B1(n1288), .B2(
        write2_in[17]), .C1(n1287), .C2(r11[17]), .Z(n2282) );
  AO222D0BWP12T U718 ( .A1(n1262), .A2(write1_in[17]), .B1(n1261), .B2(r7[17]), 
        .C1(write2_in[17]), .C2(n1260), .Z(n2410) );
  AO222D0BWP12T U719 ( .A1(n1277), .A2(n1307), .B1(n1276), .B2(r4[19]), .C1(
        write2_in[19]), .C2(n1275), .Z(n2508) );
  AO222D0BWP12T U720 ( .A1(n1277), .A2(n1256), .B1(n1276), .B2(r4[18]), .C1(
        write2_in[18]), .C2(n1275), .Z(n2507) );
  AO222D0BWP12T U721 ( .A1(n1277), .A2(write1_in[17]), .B1(n1276), .B2(r4[17]), 
        .C1(write2_in[17]), .C2(n1275), .Z(n2506) );
  AO222D0BWP12T U722 ( .A1(n1268), .A2(n1256), .B1(n1267), .B2(r5[18]), .C1(
        write2_in[18]), .C2(n1266), .Z(n2475) );
  AO222D0BWP12T U723 ( .A1(n1268), .A2(write1_in[17]), .B1(n1267), .B2(r5[17]), 
        .C1(write2_in[17]), .C2(n1266), .Z(n2474) );
  AO222D0BWP12T U724 ( .A1(n1283), .A2(n1256), .B1(n1282), .B2(r9[18]), .C1(
        write2_in[18]), .C2(n1281), .Z(n2347) );
  AO222D0BWP12T U725 ( .A1(n1259), .A2(write1_in[17]), .B1(n1258), .B2(r8[17]), 
        .C1(write2_in[17]), .C2(n1257), .Z(n2378) );
  AO222D0BWP12T U726 ( .A1(n1259), .A2(n1307), .B1(n1258), .B2(r8[19]), .C1(
        write2_in[19]), .C2(n1257), .Z(n2380) );
  AO222D0BWP12T U727 ( .A1(n1295), .A2(n1256), .B1(n1294), .B2(write2_in[18]), 
        .C1(n1293), .C2(r10[18]), .Z(n2315) );
  AO222D0BWP12T U728 ( .A1(n1274), .A2(write1_in[17]), .B1(n1273), .B2(r1[17]), 
        .C1(write2_in[17]), .C2(n1272), .Z(n2602) );
  AO222D0BWP12T U729 ( .A1(n1295), .A2(n1307), .B1(n1294), .B2(write2_in[19]), 
        .C1(n1293), .C2(r10[19]), .Z(n2316) );
  AO222D0BWP12T U730 ( .A1(n1274), .A2(n1256), .B1(n1273), .B2(r1[18]), .C1(
        write2_in[18]), .C2(n1272), .Z(n2603) );
  AO222D0BWP12T U731 ( .A1(n1298), .A2(n1307), .B1(n1297), .B2(write2_in[19]), 
        .C1(n1296), .C2(r3[19]), .Z(n2540) );
  AO222D0BWP12T U732 ( .A1(n1298), .A2(n1256), .B1(n1297), .B2(write2_in[18]), 
        .C1(n1296), .C2(r3[18]), .Z(n2539) );
  AO222D0BWP12T U733 ( .A1(n1298), .A2(write1_in[17]), .B1(n1297), .B2(
        write2_in[17]), .C1(n1296), .C2(r3[17]), .Z(n2538) );
  AO222D0BWP12T U734 ( .A1(n1265), .A2(n1307), .B1(n1264), .B2(r0[19]), .C1(
        write2_in[19]), .C2(n1263), .Z(n2636) );
  AO222D0BWP12T U735 ( .A1(n1265), .A2(write1_in[17]), .B1(n1264), .B2(r0[17]), 
        .C1(write2_in[17]), .C2(n1263), .Z(n2634) );
  AO222D0BWP12T U736 ( .A1(n1265), .A2(n1256), .B1(n1264), .B2(r0[18]), .C1(
        write2_in[18]), .C2(n1263), .Z(n2635) );
  AO222D0BWP12T U737 ( .A1(n1289), .A2(n1256), .B1(n1288), .B2(write2_in[18]), 
        .C1(n1287), .C2(r11[18]), .Z(n2283) );
  AO222D0BWP12T U738 ( .A1(n1286), .A2(n1307), .B1(n1285), .B2(r12[19]), .C1(
        write2_in[19]), .C2(n1284), .Z(n2252) );
  AO222D0BWP12T U739 ( .A1(n1274), .A2(n1307), .B1(n1273), .B2(r1[19]), .C1(
        write2_in[19]), .C2(n1272), .Z(n2604) );
  AO222D0BWP12T U740 ( .A1(n1262), .A2(n1256), .B1(n1261), .B2(r7[18]), .C1(
        write2_in[18]), .C2(n1260), .Z(n2411) );
  AO222D0BWP12T U741 ( .A1(n1262), .A2(n1307), .B1(n1261), .B2(r7[19]), .C1(
        write2_in[19]), .C2(n1260), .Z(n2412) );
  AO222D0BWP12T U742 ( .A1(n1289), .A2(n1307), .B1(n1288), .B2(write2_in[19]), 
        .C1(n1287), .C2(r11[19]), .Z(n2284) );
  AO222D0BWP12T U743 ( .A1(n1280), .A2(n1307), .B1(n1279), .B2(lr[19]), .C1(
        write2_in[19]), .C2(n1278), .Z(n2220) );
  AO222D0BWP12T U744 ( .A1(n1286), .A2(n1256), .B1(n1285), .B2(r12[18]), .C1(
        write2_in[18]), .C2(n1284), .Z(n2251) );
  AO222D0BWP12T U745 ( .A1(n1286), .A2(write1_in[17]), .B1(n1285), .B2(r12[17]), .C1(write2_in[17]), .C2(n1284), .Z(n2250) );
  AO222D0BWP12T U746 ( .A1(n1280), .A2(n1256), .B1(n1279), .B2(lr[18]), .C1(
        write2_in[18]), .C2(n1278), .Z(n2219) );
  AO222D0BWP12T U747 ( .A1(n1292), .A2(n1307), .B1(n1291), .B2(write2_in[19]), 
        .C1(n1290), .C2(r2[19]), .Z(n2572) );
  AO222D0BWP12T U748 ( .A1(n1280), .A2(write1_in[17]), .B1(n1279), .B2(lr[17]), 
        .C1(write2_in[17]), .C2(n1278), .Z(n2218) );
  AO222D0BWP12T U749 ( .A1(n1292), .A2(n1256), .B1(n1291), .B2(write2_in[18]), 
        .C1(n1290), .C2(r2[18]), .Z(n2571) );
  AO222D0BWP12T U750 ( .A1(n1271), .A2(write1_in[17]), .B1(n1270), .B2(r6[17]), 
        .C1(write2_in[17]), .C2(n1269), .Z(n2442) );
  AO222D0BWP12T U751 ( .A1(n1271), .A2(n1307), .B1(n1270), .B2(r6[19]), .C1(
        write2_in[19]), .C2(n1269), .Z(n2444) );
  AO222D0BWP12T U752 ( .A1(n1292), .A2(write1_in[17]), .B1(n1291), .B2(
        write2_in[17]), .C1(n1290), .C2(r2[17]), .Z(n2570) );
  AO222D0BWP12T U753 ( .A1(n1280), .A2(n1245), .B1(n1279), .B2(lr[15]), .C1(
        write2_in[15]), .C2(n1278), .Z(n2216) );
  AO222D0BWP12T U754 ( .A1(n1271), .A2(n1245), .B1(n1270), .B2(r6[15]), .C1(
        write2_in[15]), .C2(n1269), .Z(n2440) );
  AO222D0BWP12T U755 ( .A1(n1301), .A2(n1245), .B1(n1300), .B2(n[2026]), .C1(
        write2_in[15]), .C2(n1299), .Z(spin[15]) );
  AO222D0BWP12T U756 ( .A1(n1283), .A2(write1_in[21]), .B1(n1282), .B2(r9[21]), 
        .C1(write2_in[21]), .C2(n1281), .Z(n2350) );
  AO222D0BWP12T U757 ( .A1(n1265), .A2(write1_in[21]), .B1(n1264), .B2(r0[21]), 
        .C1(write2_in[21]), .C2(n1263), .Z(n2638) );
  AO222D0BWP12T U758 ( .A1(n1277), .A2(n1245), .B1(n1276), .B2(r4[15]), .C1(
        write2_in[15]), .C2(n1275), .Z(n2504) );
  AO222D0BWP12T U759 ( .A1(n1292), .A2(n1245), .B1(n1291), .B2(write2_in[15]), 
        .C1(n1290), .C2(r2[15]), .Z(n2568) );
  AO222D0BWP12T U760 ( .A1(n1277), .A2(write1_in[21]), .B1(n1276), .B2(r4[21]), 
        .C1(write2_in[21]), .C2(n1275), .Z(n2510) );
  AO222D0BWP12T U761 ( .A1(n1268), .A2(write1_in[21]), .B1(n1267), .B2(r5[21]), 
        .C1(write2_in[21]), .C2(n1266), .Z(n2478) );
  AO222D0BWP12T U762 ( .A1(n1298), .A2(n1245), .B1(n1297), .B2(write2_in[15]), 
        .C1(n1296), .C2(r3[15]), .Z(n2536) );
  AO222D0BWP12T U763 ( .A1(n1268), .A2(n1245), .B1(n1267), .B2(r5[15]), .C1(
        write2_in[15]), .C2(n1266), .Z(n2472) );
  AO222D0BWP12T U764 ( .A1(n1265), .A2(n1245), .B1(n1264), .B2(r0[15]), .C1(
        write2_in[15]), .C2(n1263), .Z(n2632) );
  AO222D0BWP12T U765 ( .A1(n1286), .A2(write1_in[21]), .B1(n1285), .B2(r12[21]), .C1(write2_in[21]), .C2(n1284), .Z(n2254) );
  AO222D0BWP12T U766 ( .A1(n1295), .A2(n1245), .B1(n1294), .B2(write2_in[15]), 
        .C1(n1293), .C2(r10[15]), .Z(n2312) );
  AO222D0BWP12T U767 ( .A1(n1259), .A2(n1245), .B1(n1258), .B2(r8[15]), .C1(
        write2_in[15]), .C2(n1257), .Z(n2376) );
  AO222D0BWP12T U768 ( .A1(n1295), .A2(write1_in[21]), .B1(n1294), .B2(
        write2_in[21]), .C1(n1293), .C2(r10[21]), .Z(n2318) );
  AO222D0BWP12T U769 ( .A1(n1289), .A2(n1245), .B1(n1288), .B2(write2_in[15]), 
        .C1(n1287), .C2(r11[15]), .Z(n2280) );
  AO222D0BWP12T U770 ( .A1(n1274), .A2(n1245), .B1(n1273), .B2(r1[15]), .C1(
        write2_in[15]), .C2(n1272), .Z(n2600) );
  AO222D0BWP12T U771 ( .A1(n1298), .A2(write1_in[21]), .B1(n1297), .B2(
        write2_in[21]), .C1(n1296), .C2(r3[21]), .Z(n2542) );
  AO222D0BWP12T U772 ( .A1(n1271), .A2(write1_in[21]), .B1(n1270), .B2(r6[21]), 
        .C1(write2_in[21]), .C2(n1269), .Z(n2446) );
  AO222D0BWP12T U773 ( .A1(n1303), .A2(n1245), .B1(n757), .B2(write2_in[15]), 
        .C1(n1302), .C2(tmp1[15]), .Z(n2152) );
  AO222D0BWP12T U774 ( .A1(n1262), .A2(n1245), .B1(n1261), .B2(r7[15]), .C1(
        write2_in[15]), .C2(n1260), .Z(n2408) );
  AO222D0BWP12T U775 ( .A1(n1262), .A2(write1_in[21]), .B1(n1261), .B2(r7[21]), 
        .C1(write2_in[21]), .C2(n1260), .Z(n2414) );
  AO222D0BWP12T U776 ( .A1(n1259), .A2(write1_in[21]), .B1(n1258), .B2(r8[21]), 
        .C1(write2_in[21]), .C2(n1257), .Z(n2382) );
  AO222D0BWP12T U777 ( .A1(n1286), .A2(n1245), .B1(n1285), .B2(r12[15]), .C1(
        write2_in[15]), .C2(n1284), .Z(n2248) );
  AO222D0BWP12T U778 ( .A1(n1280), .A2(write1_in[21]), .B1(n1279), .B2(lr[21]), 
        .C1(write2_in[21]), .C2(n1278), .Z(n2222) );
  AO222D0BWP12T U779 ( .A1(n1289), .A2(write1_in[21]), .B1(n1288), .B2(
        write2_in[21]), .C1(n1287), .C2(r11[21]), .Z(n2286) );
  AO222D0BWP12T U780 ( .A1(n1292), .A2(write1_in[21]), .B1(n1291), .B2(
        write2_in[21]), .C1(n1290), .C2(r2[21]), .Z(n2574) );
  AO222D0BWP12T U781 ( .A1(n1274), .A2(write1_in[21]), .B1(n1273), .B2(r1[21]), 
        .C1(write2_in[21]), .C2(n1272), .Z(n2606) );
  AO222D0BWP12T U782 ( .A1(n1283), .A2(n1245), .B1(n1282), .B2(r9[15]), .C1(
        write2_in[15]), .C2(n1281), .Z(n2344) );
  INVD1BWP12T U783 ( .I(r9[12]), .ZN(n1622) );
  INVD1BWP12T U784 ( .I(n1282), .ZN(n464) );
  INVD1BWP12T U785 ( .I(write1_in[12]), .ZN(n374) );
  INVD1BWP12T U786 ( .I(write2_in[12]), .ZN(n373) );
  INVD1BWP12T U787 ( .I(n1281), .ZN(n462) );
  OAI222D0BWP12T U788 ( .A1(n1622), .A2(n464), .B1(n374), .B2(n463), .C1(n373), 
        .C2(n462), .ZN(n2341) );
  AO222D0BWP12T U789 ( .A1(n1262), .A2(write1_in[14]), .B1(n1261), .B2(r7[14]), 
        .C1(write2_in[14]), .C2(n1260), .Z(n2407) );
  CKND0BWP12T U790 ( .I(r4[12]), .ZN(n370) );
  INVD1BWP12T U791 ( .I(n1276), .ZN(n445) );
  INVD1BWP12T U792 ( .I(n1275), .ZN(n443) );
  OAI222D0BWP12T U793 ( .A1(n370), .A2(n445), .B1(n374), .B2(n444), .C1(n373), 
        .C2(n443), .ZN(n2501) );
  AO222D0BWP12T U794 ( .A1(n1301), .A2(write1_in[14]), .B1(n1300), .B2(n[2027]), .C1(write2_in[14]), .C2(n1299), .Z(spin[14]) );
  AO222D0BWP12T U795 ( .A1(n1259), .A2(write1_in[14]), .B1(n1258), .B2(r8[14]), 
        .C1(write2_in[14]), .C2(n1257), .Z(n2375) );
  AO222D0BWP12T U796 ( .A1(n1265), .A2(write1_in[14]), .B1(n1264), .B2(r0[14]), 
        .C1(write2_in[14]), .C2(n1263), .Z(n2631) );
  AO222D0BWP12T U797 ( .A1(n1271), .A2(write1_in[14]), .B1(n1270), .B2(r6[14]), 
        .C1(write2_in[14]), .C2(n1269), .Z(n2439) );
  AO222D0BWP12T U798 ( .A1(n1286), .A2(write1_in[14]), .B1(n1285), .B2(r12[14]), .C1(write2_in[14]), .C2(n1284), .Z(n2247) );
  INVD1BWP12T U799 ( .I(r7[12]), .ZN(n1636) );
  INVD1BWP12T U800 ( .I(n1261), .ZN(n439) );
  INVD1BWP12T U801 ( .I(n1260), .ZN(n437) );
  OAI222D0BWP12T U802 ( .A1(n1636), .A2(n439), .B1(n374), .B2(n438), .C1(n373), 
        .C2(n437), .ZN(n2405) );
  AO222D0BWP12T U803 ( .A1(n1292), .A2(write1_in[14]), .B1(n1291), .B2(
        write2_in[14]), .C1(n1290), .C2(r2[14]), .Z(n2567) );
  INVD1BWP12T U804 ( .I(n1291), .ZN(n430) );
  INVD1BWP12T U805 ( .I(n1292), .ZN(n429) );
  INVD1BWP12T U806 ( .I(n1290), .ZN(n428) );
  INVD1BWP12T U807 ( .I(r2[12]), .ZN(n1635) );
  OAI222D0BWP12T U808 ( .A1(n373), .A2(n430), .B1(n374), .B2(n429), .C1(n428), 
        .C2(n1635), .ZN(n2565) );
  INVD1BWP12T U809 ( .I(n1273), .ZN(n458) );
  INVD1BWP12T U810 ( .I(n1272), .ZN(n456) );
  OAI222D0BWP12T U811 ( .A1(n1642), .A2(n458), .B1(n374), .B2(n457), .C1(n373), 
        .C2(n456), .ZN(n2597) );
  AO222D0BWP12T U812 ( .A1(n1295), .A2(write1_in[14]), .B1(n1294), .B2(
        write2_in[14]), .C1(n1293), .C2(r10[14]), .Z(n2311) );
  INVD1BWP12T U813 ( .I(r0[12]), .ZN(n1623) );
  INVD1BWP12T U814 ( .I(n1264), .ZN(n449) );
  INVD1BWP12T U815 ( .I(n1263), .ZN(n447) );
  OAI222D0BWP12T U816 ( .A1(n1623), .A2(n449), .B1(n374), .B2(n448), .C1(n373), 
        .C2(n447), .ZN(n2629) );
  INVD1BWP12T U817 ( .I(r12[12]), .ZN(n1641) );
  INVD1BWP12T U818 ( .I(n1285), .ZN(n461) );
  INVD1BWP12T U819 ( .I(n1284), .ZN(n459) );
  OAI222D0BWP12T U820 ( .A1(n1641), .A2(n461), .B1(n374), .B2(n460), .C1(n373), 
        .C2(n459), .ZN(n2245) );
  AO222D0BWP12T U821 ( .A1(n1298), .A2(write1_in[14]), .B1(n1297), .B2(
        write2_in[14]), .C1(n1296), .C2(r3[14]), .Z(n2535) );
  AO222D0BWP12T U822 ( .A1(n1289), .A2(write1_in[14]), .B1(n1288), .B2(
        write2_in[14]), .C1(n1287), .C2(r11[14]), .Z(n2279) );
  INVD1BWP12T U823 ( .I(r8[12]), .ZN(n1646) );
  INVD1BWP12T U824 ( .I(n1258), .ZN(n433) );
  INVD1BWP12T U825 ( .I(n1257), .ZN(n431) );
  OAI222D0BWP12T U826 ( .A1(n1646), .A2(n433), .B1(n374), .B2(n432), .C1(n373), 
        .C2(n431), .ZN(n2373) );
  AO222D0BWP12T U827 ( .A1(n1268), .A2(write1_in[14]), .B1(n1267), .B2(r5[14]), 
        .C1(write2_in[14]), .C2(n1266), .Z(n2471) );
  INVD1BWP12T U828 ( .I(lr[12]), .ZN(n1643) );
  INVD1BWP12T U829 ( .I(n1279), .ZN(n475) );
  INVD1BWP12T U830 ( .I(n1278), .ZN(n471) );
  OAI222D0BWP12T U831 ( .A1(n1643), .A2(n475), .B1(n374), .B2(n473), .C1(n373), 
        .C2(n471), .ZN(n2213) );
  AO222D0BWP12T U832 ( .A1(n1280), .A2(write1_in[14]), .B1(n1279), .B2(lr[14]), 
        .C1(write2_in[14]), .C2(n1278), .Z(n2215) );
  INVD1BWP12T U833 ( .I(n1295), .ZN(n466) );
  INVD1BWP12T U834 ( .I(n1293), .ZN(n465) );
  INVD1BWP12T U835 ( .I(r10[12]), .ZN(n1633) );
  OAI222D0BWP12T U836 ( .A1(n373), .A2(n467), .B1(n374), .B2(n466), .C1(n465), 
        .C2(n1633), .ZN(n2309) );
  AO222D0BWP12T U837 ( .A1(n1274), .A2(write1_in[14]), .B1(n1273), .B2(r1[14]), 
        .C1(write2_in[14]), .C2(n1272), .Z(n2599) );
  INVD1BWP12T U838 ( .I(n1297), .ZN(n436) );
  INVD1BWP12T U839 ( .I(n1298), .ZN(n435) );
  INVD1BWP12T U840 ( .I(n1296), .ZN(n434) );
  INVD1BWP12T U841 ( .I(r3[12]), .ZN(n1644) );
  OAI222D0BWP12T U842 ( .A1(n373), .A2(n436), .B1(n374), .B2(n435), .C1(n434), 
        .C2(n1644), .ZN(n2533) );
  AO222D0BWP12T U843 ( .A1(n1277), .A2(write1_in[14]), .B1(n1276), .B2(r4[14]), 
        .C1(write2_in[14]), .C2(n1275), .Z(n2503) );
  TPAOI21D0BWP12T U844 ( .A1(n1300), .A2(n[2029]), .B(reset), .ZN(n372) );
  CKND2D0BWP12T U845 ( .A1(write2_in[12]), .A2(n1299), .ZN(n371) );
  OAI211D0BWP12T U846 ( .A1(n470), .A2(n374), .B(n372), .C(n371), .ZN(spin[12]) );
  INVD1BWP12T U847 ( .I(r5[12]), .ZN(n1634) );
  INVD1BWP12T U848 ( .I(n1267), .ZN(n442) );
  INVD1BWP12T U849 ( .I(n1266), .ZN(n440) );
  OAI222D0BWP12T U850 ( .A1(n1634), .A2(n442), .B1(n374), .B2(n441), .C1(n373), 
        .C2(n440), .ZN(n2469) );
  AO222D0BWP12T U851 ( .A1(n1283), .A2(write1_in[14]), .B1(n1282), .B2(r9[14]), 
        .C1(write2_in[14]), .C2(n1281), .Z(n2343) );
  INVD1BWP12T U852 ( .I(n1288), .ZN(n455) );
  INVD1BWP12T U853 ( .I(n1289), .ZN(n454) );
  INVD1BWP12T U854 ( .I(n1287), .ZN(n453) );
  INVD1BWP12T U855 ( .I(r11[12]), .ZN(n1616) );
  OAI222D0BWP12T U856 ( .A1(n373), .A2(n455), .B1(n374), .B2(n454), .C1(n453), 
        .C2(n1616), .ZN(n2277) );
  INVD1BWP12T U857 ( .I(r6[12]), .ZN(n1647) );
  INVD1BWP12T U858 ( .I(n1270), .ZN(n452) );
  INVD1BWP12T U859 ( .I(n1269), .ZN(n450) );
  OAI222D0BWP12T U860 ( .A1(n1647), .A2(n452), .B1(n374), .B2(n451), .C1(n373), 
        .C2(n450), .ZN(n2437) );
  INVD1BWP12T U861 ( .I(write1_in[11]), .ZN(n379) );
  INVD1BWP12T U862 ( .I(write2_in[11]), .ZN(n376) );
  OAI222D0BWP12T U863 ( .A1(n594), .A2(n439), .B1(n379), .B2(n438), .C1(n376), 
        .C2(n437), .ZN(n2404) );
  AO222D0BWP12T U864 ( .A1(n1289), .A2(write1_in[13]), .B1(n1288), .B2(
        write2_in[13]), .C1(n1287), .C2(r11[13]), .Z(n2278) );
  INVD1BWP12T U865 ( .I(r0[11]), .ZN(n593) );
  OAI222D0BWP12T U866 ( .A1(n593), .A2(n449), .B1(n379), .B2(n448), .C1(n376), 
        .C2(n447), .ZN(n2628) );
  AO222D0BWP12T U867 ( .A1(n1268), .A2(write1_in[13]), .B1(n1267), .B2(r5[13]), 
        .C1(write2_in[13]), .C2(n1266), .Z(n2470) );
  OAI222D0BWP12T U868 ( .A1(n582), .A2(n458), .B1(n379), .B2(n457), .C1(n376), 
        .C2(n456), .ZN(n2596) );
  AO222D0BWP12T U869 ( .A1(n1271), .A2(write1_in[13]), .B1(n1270), .B2(r6[13]), 
        .C1(write2_in[13]), .C2(n1269), .Z(n2438) );
  AO222D0BWP12T U870 ( .A1(n1283), .A2(write1_in[13]), .B1(n1282), .B2(r9[13]), 
        .C1(write2_in[13]), .C2(n1281), .Z(n2342) );
  OAI222D0BWP12T U871 ( .A1(n376), .A2(n430), .B1(n379), .B2(n429), .C1(n428), 
        .C2(n583), .ZN(n2564) );
  OAI222D0BWP12T U872 ( .A1(n376), .A2(n436), .B1(n379), .B2(n435), .C1(n434), 
        .C2(n591), .ZN(n2532) );
  OAI222D0BWP12T U873 ( .A1(n588), .A2(n452), .B1(n379), .B2(n451), .C1(n376), 
        .C2(n450), .ZN(n2436) );
  AO222D0BWP12T U874 ( .A1(n1298), .A2(write1_in[13]), .B1(n1297), .B2(
        write2_in[13]), .C1(n1296), .C2(r3[13]), .Z(n2534) );
  AO222D0BWP12T U875 ( .A1(n1301), .A2(write1_in[13]), .B1(n1300), .B2(n[2028]), .C1(write2_in[13]), .C2(n1299), .Z(spin[13]) );
  INVD1BWP12T U876 ( .I(r9[11]), .ZN(n589) );
  OAI222D0BWP12T U877 ( .A1(n589), .A2(n464), .B1(n379), .B2(n463), .C1(n376), 
        .C2(n462), .ZN(n2340) );
  OAI222D0BWP12T U878 ( .A1(n376), .A2(n467), .B1(n379), .B2(n466), .C1(n465), 
        .C2(n579), .ZN(n2308) );
  CKND0BWP12T U879 ( .I(r4[11]), .ZN(n375) );
  OAI222D0BWP12T U880 ( .A1(n375), .A2(n445), .B1(n379), .B2(n444), .C1(n376), 
        .C2(n443), .ZN(n2500) );
  AO222D0BWP12T U881 ( .A1(n1259), .A2(write1_in[13]), .B1(n1258), .B2(r8[13]), 
        .C1(write2_in[13]), .C2(n1257), .Z(n2374) );
  AO222D0BWP12T U882 ( .A1(n1295), .A2(write1_in[13]), .B1(n1294), .B2(
        write2_in[13]), .C1(n1293), .C2(r10[13]), .Z(n2310) );
  OAI222D0BWP12T U883 ( .A1(n592), .A2(n442), .B1(n379), .B2(n441), .C1(n376), 
        .C2(n440), .ZN(n2468) );
  AO222D0BWP12T U884 ( .A1(n1303), .A2(write1_in[12]), .B1(n757), .B2(
        write2_in[12]), .C1(n1302), .C2(tmp1[12]), .Z(n2149) );
  AO222D0BWP12T U885 ( .A1(n1274), .A2(write1_in[13]), .B1(n1273), .B2(r1[13]), 
        .C1(write2_in[13]), .C2(n1272), .Z(n2598) );
  OAI222D0BWP12T U886 ( .A1(n590), .A2(n433), .B1(n379), .B2(n432), .C1(n376), 
        .C2(n431), .ZN(n2372) );
  AO222D0BWP12T U887 ( .A1(n1303), .A2(write1_in[13]), .B1(n757), .B2(
        write2_in[13]), .C1(n1302), .C2(tmp1[13]), .Z(n2150) );
  AO222D0BWP12T U888 ( .A1(n1277), .A2(write1_in[13]), .B1(n1276), .B2(r4[13]), 
        .C1(write2_in[13]), .C2(n1275), .Z(n2502) );
  AO222D0BWP12T U889 ( .A1(n1280), .A2(write1_in[13]), .B1(n1279), .B2(lr[13]), 
        .C1(write2_in[13]), .C2(n1278), .Z(n2214) );
  INVD1BWP12T U890 ( .I(r11[11]), .ZN(n577) );
  OAI222D0BWP12T U891 ( .A1(n376), .A2(n455), .B1(n379), .B2(n454), .C1(n453), 
        .C2(n577), .ZN(n2276) );
  OAI222D0BWP12T U892 ( .A1(n580), .A2(n475), .B1(n379), .B2(n473), .C1(n376), 
        .C2(n471), .ZN(n2212) );
  AO222D0BWP12T U893 ( .A1(n1262), .A2(write1_in[13]), .B1(n1261), .B2(r7[13]), 
        .C1(write2_in[13]), .C2(n1260), .Z(n2406) );
  OAI222D0BWP12T U894 ( .A1(n1089), .A2(n461), .B1(n379), .B2(n460), .C1(n376), 
        .C2(n459), .ZN(n2244) );
  AO222D0BWP12T U895 ( .A1(n1292), .A2(write1_in[13]), .B1(n1291), .B2(
        write2_in[13]), .C1(n1290), .C2(r2[13]), .Z(n2566) );
  AO222D0BWP12T U896 ( .A1(n1265), .A2(write1_in[13]), .B1(n1264), .B2(r0[13]), 
        .C1(write2_in[13]), .C2(n1263), .Z(n2630) );
  AO222D0BWP12T U897 ( .A1(n1286), .A2(write1_in[13]), .B1(n1285), .B2(r12[13]), .C1(write2_in[13]), .C2(n1284), .Z(n2246) );
  TPAOI21D0BWP12T U898 ( .A1(n1300), .A2(n[2030]), .B(reset), .ZN(n378) );
  CKND2D0BWP12T U899 ( .A1(write2_in[11]), .A2(n1299), .ZN(n377) );
  OAI211D0BWP12T U900 ( .A1(n470), .A2(n379), .B(n378), .C(n377), .ZN(spin[11]) );
  INVD1BWP12T U901 ( .I(r9[8]), .ZN(n1693) );
  INVD1BWP12T U902 ( .I(write1_in[8]), .ZN(n401) );
  INVD1BWP12T U903 ( .I(write2_in[8]), .ZN(n400) );
  OAI222D0BWP12T U904 ( .A1(n1693), .A2(n464), .B1(n401), .B2(n463), .C1(n400), 
        .C2(n462), .ZN(n2337) );
  INVD1BWP12T U905 ( .I(write2_in[9]), .ZN(n407) );
  INVD1BWP12T U906 ( .I(write1_in[9]), .ZN(n408) );
  OAI222D0BWP12T U907 ( .A1(n407), .A2(n455), .B1(n408), .B2(n454), .C1(n453), 
        .C2(n380), .ZN(n2274) );
  OAI222D0BWP12T U908 ( .A1(n627), .A2(n475), .B1(n408), .B2(n473), .C1(n407), 
        .C2(n471), .ZN(n2210) );
  INVD1BWP12T U909 ( .I(write2_in[7]), .ZN(n416) );
  INVD1BWP12T U910 ( .I(write1_in[7]), .ZN(n417) );
  INVD1BWP12T U911 ( .I(r11[7]), .ZN(n520) );
  OAI222D0BWP12T U912 ( .A1(n416), .A2(n455), .B1(n417), .B2(n454), .C1(n453), 
        .C2(n520), .ZN(n2272) );
  INVD1BWP12T U913 ( .I(write1_in[2]), .ZN(n410) );
  INVD1BWP12T U914 ( .I(write2_in[2]), .ZN(n409) );
  OAI222D0BWP12T U915 ( .A1(n381), .A2(n464), .B1(n410), .B2(n463), .C1(n409), 
        .C2(n462), .ZN(n2331) );
  OAI222D0BWP12T U916 ( .A1(n626), .A2(n458), .B1(n408), .B2(n457), .C1(n407), 
        .C2(n456), .ZN(n2594) );
  INVD1BWP12T U917 ( .I(write2_in[10]), .ZN(n414) );
  INVD1BWP12T U918 ( .I(write1_in[10]), .ZN(n415) );
  INVD1BWP12T U919 ( .I(r11[10]), .ZN(n1655) );
  OAI222D0BWP12T U920 ( .A1(n414), .A2(n455), .B1(n415), .B2(n454), .C1(n453), 
        .C2(n1655), .ZN(n2275) );
  OAI222D0BWP12T U921 ( .A1(n1683), .A2(n475), .B1(n401), .B2(n473), .C1(n400), 
        .C2(n471), .ZN(n2209) );
  INVD1BWP12T U922 ( .I(lr[7]), .ZN(n1719) );
  OAI222D0BWP12T U923 ( .A1(n1719), .A2(n475), .B1(n417), .B2(n473), .C1(n416), 
        .C2(n471), .ZN(n2208) );
  OAI222D0BWP12T U924 ( .A1(n1658), .A2(n475), .B1(n415), .B2(n473), .C1(n414), 
        .C2(n471), .ZN(n2211) );
  INVD1BWP12T U925 ( .I(write2_in[5]), .ZN(n404) );
  INVD1BWP12T U926 ( .I(write1_in[5]), .ZN(n405) );
  INVD1BWP12T U927 ( .I(r11[5]), .ZN(n548) );
  OAI222D0BWP12T U928 ( .A1(n404), .A2(n455), .B1(n405), .B2(n454), .C1(n453), 
        .C2(n548), .ZN(n2270) );
  INVD1BWP12T U929 ( .I(r2[5]), .ZN(n1826) );
  OAI222D0BWP12T U930 ( .A1(n404), .A2(n430), .B1(n405), .B2(n429), .C1(n428), 
        .C2(n1826), .ZN(n2558) );
  OAI222D0BWP12T U931 ( .A1(n1686), .A2(n458), .B1(n401), .B2(n457), .C1(n400), 
        .C2(n456), .ZN(n2593) );
  INVD1BWP12T U932 ( .I(r9[10]), .ZN(n1667) );
  OAI222D0BWP12T U933 ( .A1(n1667), .A2(n464), .B1(n415), .B2(n463), .C1(n414), 
        .C2(n462), .ZN(n2339) );
  INVD1BWP12T U934 ( .I(r9[5]), .ZN(n983) );
  OAI222D0BWP12T U935 ( .A1(n983), .A2(n464), .B1(n405), .B2(n463), .C1(n404), 
        .C2(n462), .ZN(n2334) );
  INVD1BWP12T U936 ( .I(r9[7]), .ZN(n526) );
  OAI222D0BWP12T U937 ( .A1(n526), .A2(n464), .B1(n417), .B2(n463), .C1(n416), 
        .C2(n462), .ZN(n2336) );
  INVD1BWP12T U938 ( .I(r9[1]), .ZN(n497) );
  INVD1BWP12T U939 ( .I(write1_in[1]), .ZN(n412) );
  INVD1BWP12T U940 ( .I(write2_in[1]), .ZN(n411) );
  OAI222D0BWP12T U941 ( .A1(n497), .A2(n464), .B1(n412), .B2(n463), .C1(n411), 
        .C2(n462), .ZN(n2330) );
  OAI222D0BWP12T U942 ( .A1(n1970), .A2(n475), .B1(n410), .B2(n473), .C1(n409), 
        .C2(n471), .ZN(n2203) );
  OAI222D0BWP12T U943 ( .A1(n1718), .A2(n458), .B1(n417), .B2(n457), .C1(n416), 
        .C2(n456), .ZN(n2592) );
  INVD1BWP12T U944 ( .I(lr[1]), .ZN(n1859) );
  OAI222D0BWP12T U945 ( .A1(n1859), .A2(n475), .B1(n412), .B2(n473), .C1(n411), 
        .C2(n471), .ZN(n2202) );
  INVD1BWP12T U946 ( .I(r0[7]), .ZN(n527) );
  OAI222D0BWP12T U947 ( .A1(n527), .A2(n449), .B1(n417), .B2(n448), .C1(n416), 
        .C2(n447), .ZN(n2624) );
  INVD1BWP12T U948 ( .I(lr[5]), .ZN(n1834) );
  OAI222D0BWP12T U949 ( .A1(n1834), .A2(n475), .B1(n405), .B2(n473), .C1(n404), 
        .C2(n471), .ZN(n2206) );
  OAI222D0BWP12T U950 ( .A1(n828), .A2(n449), .B1(n410), .B2(n448), .C1(n409), 
        .C2(n447), .ZN(n2619) );
  OAI222D0BWP12T U951 ( .A1(n1666), .A2(n452), .B1(n415), .B2(n451), .C1(n414), 
        .C2(n450), .ZN(n2435) );
  OAI222D0BWP12T U952 ( .A1(n630), .A2(n452), .B1(n408), .B2(n451), .C1(n407), 
        .C2(n450), .ZN(n2434) );
  OAI222D0BWP12T U953 ( .A1(n1692), .A2(n452), .B1(n401), .B2(n451), .C1(n400), 
        .C2(n450), .ZN(n2433) );
  INVD1BWP12T U954 ( .I(r11[8]), .ZN(n1680) );
  OAI222D0BWP12T U955 ( .A1(n400), .A2(n455), .B1(n401), .B2(n454), .C1(n453), 
        .C2(n1680), .ZN(n2273) );
  INVD1BWP12T U956 ( .I(r6[7]), .ZN(n1723) );
  OAI222D0BWP12T U957 ( .A1(n1723), .A2(n452), .B1(n417), .B2(n451), .C1(n416), 
        .C2(n450), .ZN(n2432) );
  INVD1BWP12T U958 ( .I(r6[5]), .ZN(n1838) );
  OAI222D0BWP12T U959 ( .A1(n1838), .A2(n452), .B1(n405), .B2(n451), .C1(n404), 
        .C2(n450), .ZN(n2430) );
  OAI222D0BWP12T U960 ( .A1(n1978), .A2(n452), .B1(n410), .B2(n451), .C1(n409), 
        .C2(n450), .ZN(n2427) );
  INVD1BWP12T U961 ( .I(r6[1]), .ZN(n1863) );
  OAI222D0BWP12T U962 ( .A1(n1863), .A2(n452), .B1(n412), .B2(n451), .C1(n411), 
        .C2(n450), .ZN(n2426) );
  INVD1BWP12T U963 ( .I(r3[1]), .ZN(n1860) );
  OAI222D0BWP12T U964 ( .A1(n411), .A2(n436), .B1(n412), .B2(n435), .C1(n434), 
        .C2(n1860), .ZN(n2522) );
  INVD1BWP12T U965 ( .I(r0[5]), .ZN(n554) );
  OAI222D0BWP12T U966 ( .A1(n554), .A2(n449), .B1(n405), .B2(n448), .C1(n404), 
        .C2(n447), .ZN(n2622) );
  OAI222D0BWP12T U967 ( .A1(n409), .A2(n436), .B1(n410), .B2(n435), .C1(n434), 
        .C2(n1973), .ZN(n2523) );
  INVD1BWP12T U968 ( .I(r0[8]), .ZN(n1698) );
  OAI222D0BWP12T U969 ( .A1(n1698), .A2(n449), .B1(n401), .B2(n448), .C1(n400), 
        .C2(n447), .ZN(n2625) );
  INVD1BWP12T U970 ( .I(r3[5]), .ZN(n1835) );
  OAI222D0BWP12T U971 ( .A1(n404), .A2(n436), .B1(n405), .B2(n435), .C1(n434), 
        .C2(n1835), .ZN(n2526) );
  INVD1BWP12T U972 ( .I(r3[7]), .ZN(n1720) );
  OAI222D0BWP12T U973 ( .A1(n416), .A2(n436), .B1(n417), .B2(n435), .C1(n434), 
        .C2(n1720), .ZN(n2528) );
  OAI222D0BWP12T U974 ( .A1(n400), .A2(n436), .B1(n401), .B2(n435), .C1(n434), 
        .C2(n1696), .ZN(n2529) );
  OAI222D0BWP12T U975 ( .A1(n407), .A2(n436), .B1(n408), .B2(n435), .C1(n434), 
        .C2(n628), .ZN(n2530) );
  OAI222D0BWP12T U976 ( .A1(n414), .A2(n436), .B1(n415), .B2(n435), .C1(n434), 
        .C2(n1670), .ZN(n2531) );
  OAI222D0BWP12T U977 ( .A1(n382), .A2(n449), .B1(n408), .B2(n448), .C1(n407), 
        .C2(n447), .ZN(n2626) );
  TPAOI21D0BWP12T U978 ( .A1(n1300), .A2(n[2031]), .B(reset), .ZN(n384) );
  CKND2D0BWP12T U979 ( .A1(write2_in[10]), .A2(n1299), .ZN(n383) );
  OAI211D0BWP12T U980 ( .A1(n470), .A2(n415), .B(n384), .C(n383), .ZN(spin[10]) );
  INVD1BWP12T U981 ( .I(r1[5]), .ZN(n1833) );
  OAI222D0BWP12T U982 ( .A1(n1833), .A2(n458), .B1(n405), .B2(n457), .C1(n404), 
        .C2(n456), .ZN(n2590) );
  INVD1BWP12T U983 ( .I(r0[10]), .ZN(n1672) );
  OAI222D0BWP12T U984 ( .A1(n1672), .A2(n449), .B1(n415), .B2(n448), .C1(n414), 
        .C2(n447), .ZN(n2627) );
  AO222D0BWP12T U985 ( .A1(n1303), .A2(write1_in[11]), .B1(n757), .B2(
        write2_in[11]), .C1(n1302), .C2(tmp1[11]), .Z(n2148) );
  OAI222D0BWP12T U986 ( .A1(n1673), .A2(n439), .B1(n415), .B2(n438), .C1(n414), 
        .C2(n437), .ZN(n2403) );
  OAI222D0BWP12T U987 ( .A1(n620), .A2(n439), .B1(n408), .B2(n438), .C1(n407), 
        .C2(n437), .ZN(n2402) );
  OAI222D0BWP12T U988 ( .A1(n1699), .A2(n439), .B1(n401), .B2(n438), .C1(n400), 
        .C2(n437), .ZN(n2401) );
  INVD1BWP12T U989 ( .I(r10[1]), .ZN(n1846) );
  OAI222D0BWP12T U990 ( .A1(n411), .A2(n467), .B1(n412), .B2(n466), .C1(n465), 
        .C2(n1846), .ZN(n2298) );
  INVD1BWP12T U991 ( .I(r7[7]), .ZN(n1712) );
  OAI222D0BWP12T U992 ( .A1(n1712), .A2(n439), .B1(n417), .B2(n438), .C1(n416), 
        .C2(n437), .ZN(n2400) );
  OAI222D0BWP12T U993 ( .A1(n409), .A2(n467), .B1(n410), .B2(n466), .C1(n465), 
        .C2(n1947), .ZN(n2299) );
  OAI222D0BWP12T U994 ( .A1(n1969), .A2(n458), .B1(n410), .B2(n457), .C1(n409), 
        .C2(n456), .ZN(n2587) );
  TPAOI21D0BWP12T U995 ( .A1(n1300), .A2(n[2032]), .B(reset), .ZN(n386) );
  CKND2D0BWP12T U996 ( .A1(write2_in[9]), .A2(n1299), .ZN(n385) );
  OAI211D0BWP12T U997 ( .A1(n470), .A2(n408), .B(n386), .C(n385), .ZN(spin[9])
         );
  INVD1BWP12T U998 ( .I(r7[5]), .ZN(n1827) );
  OAI222D0BWP12T U999 ( .A1(n1827), .A2(n439), .B1(n405), .B2(n438), .C1(n404), 
        .C2(n437), .ZN(n2398) );
  INVD1BWP12T U1000 ( .I(r10[5]), .ZN(n1824) );
  OAI222D0BWP12T U1001 ( .A1(n404), .A2(n467), .B1(n405), .B2(n466), .C1(n465), 
        .C2(n1824), .ZN(n2302) );
  INVD1BWP12T U1002 ( .I(r1[1]), .ZN(n1858) );
  OAI222D0BWP12T U1003 ( .A1(n1858), .A2(n458), .B1(n412), .B2(n457), .C1(n411), .C2(n456), .ZN(n2586) );
  OAI222D0BWP12T U1004 ( .A1(n1053), .A2(n464), .B1(n408), .B2(n463), .C1(n407), .C2(n462), .ZN(n2338) );
  OAI222D0BWP12T U1005 ( .A1(n1960), .A2(n439), .B1(n410), .B2(n438), .C1(n409), .C2(n437), .ZN(n2395) );
  INVD1BWP12T U1006 ( .I(r10[7]), .ZN(n1709) );
  OAI222D0BWP12T U1007 ( .A1(n416), .A2(n467), .B1(n417), .B2(n466), .C1(n465), 
        .C2(n1709), .ZN(n2304) );
  INVD1BWP12T U1008 ( .I(r7[1]), .ZN(n1852) );
  OAI222D0BWP12T U1009 ( .A1(n1852), .A2(n439), .B1(n412), .B2(n438), .C1(n411), .C2(n437), .ZN(n2394) );
  OAI222D0BWP12T U1010 ( .A1(n400), .A2(n467), .B1(n401), .B2(n466), .C1(n465), 
        .C2(n1682), .ZN(n2305) );
  OAI222D0BWP12T U1011 ( .A1(n407), .A2(n467), .B1(n408), .B2(n466), .C1(n465), 
        .C2(n617), .ZN(n2306) );
  TPAOI21D0BWP12T U1012 ( .A1(n1300), .A2(n[2033]), .B(reset), .ZN(n388) );
  CKND2D0BWP12T U1013 ( .A1(write2_in[8]), .A2(n1299), .ZN(n387) );
  OAI211D0BWP12T U1014 ( .A1(n470), .A2(n401), .B(n388), .C(n387), .ZN(spin[8]) );
  OAI222D0BWP12T U1015 ( .A1(n414), .A2(n430), .B1(n415), .B2(n429), .C1(n428), 
        .C2(n1661), .ZN(n2563) );
  OAI222D0BWP12T U1016 ( .A1(n414), .A2(n467), .B1(n415), .B2(n466), .C1(n465), 
        .C2(n1657), .ZN(n2307) );
  TPAOI21D0BWP12T U1017 ( .A1(n1300), .A2(n[2034]), .B(reset), .ZN(n390) );
  CKND2D0BWP12T U1018 ( .A1(write2_in[7]), .A2(n1299), .ZN(n389) );
  OAI211D0BWP12T U1019 ( .A1(n470), .A2(n417), .B(n390), .C(n389), .ZN(spin[7]) );
  OAI222D0BWP12T U1020 ( .A1(n407), .A2(n430), .B1(n408), .B2(n429), .C1(n428), 
        .C2(n619), .ZN(n2562) );
  OAI222D0BWP12T U1021 ( .A1(n400), .A2(n430), .B1(n401), .B2(n429), .C1(n428), 
        .C2(n1687), .ZN(n2561) );
  AOI21D0BWP12T U1022 ( .A1(n1300), .A2(n[2036]), .B(reset), .ZN(n392) );
  CKND2D0BWP12T U1023 ( .A1(write2_in[5]), .A2(n1299), .ZN(n391) );
  OAI211D0BWP12T U1024 ( .A1(n470), .A2(n405), .B(n392), .C(n391), .ZN(spin[5]) );
  INVD1BWP12T U1025 ( .I(r2[7]), .ZN(n1711) );
  OAI222D0BWP12T U1026 ( .A1(n416), .A2(n430), .B1(n417), .B2(n429), .C1(n428), 
        .C2(n1711), .ZN(n2560) );
  AOI21D0BWP12T U1027 ( .A1(n1300), .A2(n[2039]), .B(reset), .ZN(n394) );
  CKND2D0BWP12T U1028 ( .A1(write2_in[2]), .A2(n1299), .ZN(n393) );
  OAI211D0BWP12T U1029 ( .A1(n470), .A2(n410), .B(n394), .C(n393), .ZN(spin[2]) );
  INVD1BWP12T U1030 ( .I(r8[1]), .ZN(n1862) );
  OAI222D0BWP12T U1031 ( .A1(n1862), .A2(n433), .B1(n412), .B2(n432), .C1(n411), .C2(n431), .ZN(n2362) );
  OAI222D0BWP12T U1032 ( .A1(n1669), .A2(n433), .B1(n415), .B2(n432), .C1(n414), .C2(n431), .ZN(n2371) );
  INVD1BWP12T U1033 ( .I(r2[1]), .ZN(n1851) );
  OAI222D0BWP12T U1034 ( .A1(n411), .A2(n430), .B1(n412), .B2(n429), .C1(n428), 
        .C2(n1851), .ZN(n2554) );
  AOI21D0BWP12T U1035 ( .A1(n1300), .A2(n[2040]), .B(reset), .ZN(n396) );
  CKND2D0BWP12T U1036 ( .A1(write2_in[1]), .A2(n1299), .ZN(n395) );
  OAI211D0BWP12T U1037 ( .A1(n470), .A2(n412), .B(n396), .C(n395), .ZN(spin[1]) );
  OAI222D0BWP12T U1038 ( .A1(n1054), .A2(n433), .B1(n408), .B2(n432), .C1(n407), .C2(n431), .ZN(n2370) );
  OAI222D0BWP12T U1039 ( .A1(n1695), .A2(n433), .B1(n401), .B2(n432), .C1(n400), .C2(n431), .ZN(n2369) );
  INVD1BWP12T U1040 ( .I(r8[7]), .ZN(n1722) );
  OAI222D0BWP12T U1041 ( .A1(n1722), .A2(n433), .B1(n417), .B2(n432), .C1(n416), .C2(n431), .ZN(n2368) );
  OAI222D0BWP12T U1042 ( .A1(n409), .A2(n430), .B1(n410), .B2(n429), .C1(n428), 
        .C2(n1958), .ZN(n2555) );
  OAI222D0BWP12T U1043 ( .A1(n1976), .A2(n433), .B1(n410), .B2(n432), .C1(n409), .C2(n431), .ZN(n2363) );
  INVD1BWP12T U1044 ( .I(r0[1]), .ZN(n498) );
  OAI222D0BWP12T U1045 ( .A1(n498), .A2(n449), .B1(n412), .B2(n448), .C1(n411), 
        .C2(n447), .ZN(n2618) );
  INVD1BWP12T U1046 ( .I(r8[5]), .ZN(n1837) );
  OAI222D0BWP12T U1047 ( .A1(n1837), .A2(n433), .B1(n405), .B2(n432), .C1(n404), .C2(n431), .ZN(n2366) );
  OAI222D0BWP12T U1048 ( .A1(n1660), .A2(n458), .B1(n415), .B2(n457), .C1(n414), .C2(n456), .ZN(n2595) );
  INVD1BWP12T U1049 ( .I(r12[5]), .ZN(n1832) );
  OAI222D0BWP12T U1050 ( .A1(n1832), .A2(n461), .B1(n405), .B2(n460), .C1(n404), .C2(n459), .ZN(n2238) );
  OAI222D0BWP12T U1051 ( .A1(n397), .A2(n461), .B1(n415), .B2(n460), .C1(n414), 
        .C2(n459), .ZN(n2243) );
  OAI222D0BWP12T U1052 ( .A1(n1950), .A2(n442), .B1(n410), .B2(n441), .C1(n409), .C2(n440), .ZN(n2459) );
  INVD1BWP12T U1053 ( .I(r5[1]), .ZN(n1847) );
  OAI222D0BWP12T U1054 ( .A1(n1847), .A2(n442), .B1(n412), .B2(n441), .C1(n411), .C2(n440), .ZN(n2458) );
  CKND0BWP12T U1055 ( .I(r4[8]), .ZN(n398) );
  OAI222D0BWP12T U1056 ( .A1(n398), .A2(n445), .B1(n401), .B2(n444), .C1(n400), 
        .C2(n443), .ZN(n2497) );
  INVD1BWP12T U1057 ( .I(r11[1]), .ZN(n491) );
  OAI222D0BWP12T U1058 ( .A1(n411), .A2(n455), .B1(n412), .B2(n454), .C1(n453), 
        .C2(n491), .ZN(n2266) );
  OAI222D0BWP12T U1059 ( .A1(n618), .A2(n442), .B1(n408), .B2(n441), .C1(n407), 
        .C2(n440), .ZN(n2466) );
  OAI222D0BWP12T U1060 ( .A1(n1697), .A2(n442), .B1(n401), .B2(n441), .C1(n400), .C2(n440), .ZN(n2465) );
  OAI222D0BWP12T U1061 ( .A1(n1671), .A2(n442), .B1(n415), .B2(n441), .C1(n414), .C2(n440), .ZN(n2467) );
  INVD1BWP12T U1062 ( .I(r12[1]), .ZN(n1857) );
  OAI222D0BWP12T U1063 ( .A1(n1857), .A2(n461), .B1(n412), .B2(n460), .C1(n411), .C2(n459), .ZN(n2234) );
  INVD1BWP12T U1064 ( .I(r12[7]), .ZN(n1717) );
  OAI222D0BWP12T U1065 ( .A1(n1717), .A2(n461), .B1(n417), .B2(n460), .C1(n416), .C2(n459), .ZN(n2240) );
  CKND0BWP12T U1066 ( .I(r4[7]), .ZN(n399) );
  OAI222D0BWP12T U1067 ( .A1(n399), .A2(n445), .B1(n417), .B2(n444), .C1(n416), 
        .C2(n443), .ZN(n2496) );
  OAI222D0BWP12T U1068 ( .A1(n937), .A2(n461), .B1(n401), .B2(n460), .C1(n400), 
        .C2(n459), .ZN(n2241) );
  CKND0BWP12T U1069 ( .I(r4[9]), .ZN(n402) );
  OAI222D0BWP12T U1070 ( .A1(n402), .A2(n445), .B1(n408), .B2(n444), .C1(n407), 
        .C2(n443), .ZN(n2498) );
  OAI222D0BWP12T U1071 ( .A1(n409), .A2(n455), .B1(n410), .B2(n454), .C1(n453), 
        .C2(n403), .ZN(n2267) );
  INVD1BWP12T U1072 ( .I(r5[5]), .ZN(n1825) );
  OAI222D0BWP12T U1073 ( .A1(n1825), .A2(n442), .B1(n405), .B2(n441), .C1(n404), .C2(n440), .ZN(n2462) );
  CKND0BWP12T U1074 ( .I(r4[5]), .ZN(n406) );
  OAI222D0BWP12T U1075 ( .A1(n406), .A2(n445), .B1(n405), .B2(n444), .C1(n404), 
        .C2(n443), .ZN(n2494) );
  INVD1BWP12T U1076 ( .I(r12[9]), .ZN(n625) );
  OAI222D0BWP12T U1077 ( .A1(n625), .A2(n461), .B1(n408), .B2(n460), .C1(n407), 
        .C2(n459), .ZN(n2242) );
  CKND0BWP12T U1078 ( .I(r4[2]), .ZN(n827) );
  OAI222D0BWP12T U1079 ( .A1(n827), .A2(n445), .B1(n410), .B2(n444), .C1(n409), 
        .C2(n443), .ZN(n2491) );
  INVD1BWP12T U1080 ( .I(r12[2]), .ZN(n1966) );
  OAI222D0BWP12T U1081 ( .A1(n1966), .A2(n461), .B1(n410), .B2(n460), .C1(n409), .C2(n459), .ZN(n2235) );
  CKND0BWP12T U1082 ( .I(r4[1]), .ZN(n413) );
  OAI222D0BWP12T U1083 ( .A1(n413), .A2(n445), .B1(n412), .B2(n444), .C1(n411), 
        .C2(n443), .ZN(n2490) );
  CKND0BWP12T U1084 ( .I(r4[10]), .ZN(n1135) );
  OAI222D0BWP12T U1085 ( .A1(n1135), .A2(n445), .B1(n415), .B2(n444), .C1(n414), .C2(n443), .ZN(n2499) );
  INVD1BWP12T U1086 ( .I(r5[7]), .ZN(n1710) );
  OAI222D0BWP12T U1087 ( .A1(n1710), .A2(n442), .B1(n417), .B2(n441), .C1(n416), .C2(n440), .ZN(n2464) );
  INVD1BWP12T U1088 ( .I(r12[3]), .ZN(n1933) );
  INVD1BWP12T U1089 ( .I(write1_in[3]), .ZN(n426) );
  INVD1BWP12T U1090 ( .I(write2_in[3]), .ZN(n427) );
  OAI222D0BWP12T U1091 ( .A1(n1933), .A2(n461), .B1(n426), .B2(n460), .C1(n427), .C2(n459), .ZN(n2236) );
  INVD1BWP12T U1092 ( .I(write1_in[4]), .ZN(n425) );
  INVD1BWP12T U1093 ( .I(write2_in[4]), .ZN(n424) );
  OAI222D0BWP12T U1094 ( .A1(n1900), .A2(n452), .B1(n425), .B2(n451), .C1(n424), .C2(n450), .ZN(n2429) );
  CKND0BWP12T U1095 ( .I(r4[3]), .ZN(n839) );
  OAI222D0BWP12T U1096 ( .A1(n839), .A2(n445), .B1(n426), .B2(n444), .C1(n427), 
        .C2(n443), .ZN(n2492) );
  INVD1BWP12T U1097 ( .I(r6[3]), .ZN(n1939) );
  OAI222D0BWP12T U1098 ( .A1(n1939), .A2(n452), .B1(n426), .B2(n451), .C1(n427), .C2(n450), .ZN(n2428) );
  CKND0BWP12T U1099 ( .I(r4[4]), .ZN(n418) );
  OAI222D0BWP12T U1100 ( .A1(n418), .A2(n445), .B1(n425), .B2(n444), .C1(n424), 
        .C2(n443), .ZN(n2493) );
  OAI222D0BWP12T U1101 ( .A1(n419), .A2(n461), .B1(n425), .B2(n460), .C1(n424), 
        .C2(n459), .ZN(n2237) );
  AOI21D0BWP12T U1102 ( .A1(n1300), .A2(n[2037]), .B(reset), .ZN(n421) );
  CKND2D0BWP12T U1103 ( .A1(write2_in[4]), .A2(n1299), .ZN(n420) );
  OAI211D0BWP12T U1104 ( .A1(n470), .A2(n425), .B(n421), .C(n420), .ZN(spin[4]) );
  AOI21D0BWP12T U1105 ( .A1(n1300), .A2(n[2038]), .B(reset), .ZN(n423) );
  CKND2D0BWP12T U1106 ( .A1(write2_in[3]), .A2(n1299), .ZN(n422) );
  OAI211D0BWP12T U1107 ( .A1(n470), .A2(n426), .B(n423), .C(n422), .ZN(spin[3]) );
  OAI222D0BWP12T U1108 ( .A1(n1889), .A2(n475), .B1(n425), .B2(n473), .C1(n424), .C2(n471), .ZN(n2205) );
  INVD1BWP12T U1109 ( .I(r2[3]), .ZN(n1927) );
  OAI222D0BWP12T U1110 ( .A1(n427), .A2(n430), .B1(n426), .B2(n429), .C1(n428), 
        .C2(n1927), .ZN(n2556) );
  INVD1BWP12T U1111 ( .I(lr[3]), .ZN(n1935) );
  OAI222D0BWP12T U1112 ( .A1(n1935), .A2(n475), .B1(n426), .B2(n473), .C1(n427), .C2(n471), .ZN(n2204) );
  OAI222D0BWP12T U1113 ( .A1(n424), .A2(n430), .B1(n425), .B2(n429), .C1(n428), 
        .C2(n1894), .ZN(n2557) );
  OAI222D0BWP12T U1114 ( .A1(n1906), .A2(n433), .B1(n425), .B2(n432), .C1(n424), .C2(n431), .ZN(n2365) );
  INVD1BWP12T U1115 ( .I(r8[3]), .ZN(n1938) );
  OAI222D0BWP12T U1116 ( .A1(n1938), .A2(n433), .B1(n426), .B2(n432), .C1(n427), .C2(n431), .ZN(n2364) );
  AO222D0BWP12T U1117 ( .A1(n1303), .A2(write1_in[1]), .B1(n757), .B2(
        write2_in[1]), .C1(n1302), .C2(tmp1[1]), .Z(n2138) );
  AO222D0BWP12T U1118 ( .A1(n1303), .A2(write1_in[5]), .B1(n757), .B2(
        write2_in[5]), .C1(n1302), .C2(tmp1[5]), .Z(n2142) );
  AO222D0BWP12T U1119 ( .A1(n1303), .A2(write1_in[7]), .B1(n757), .B2(
        write2_in[7]), .C1(n1302), .C2(tmp1[7]), .Z(n2144) );
  AO222D0BWP12T U1120 ( .A1(n1303), .A2(write1_in[8]), .B1(n757), .B2(
        write2_in[8]), .C1(n1302), .C2(tmp1[8]), .Z(n2145) );
  AO222D0BWP12T U1121 ( .A1(n1303), .A2(write1_in[9]), .B1(n757), .B2(
        write2_in[9]), .C1(n1302), .C2(tmp1[9]), .Z(n2146) );
  AO222D0BWP12T U1122 ( .A1(n1303), .A2(write1_in[10]), .B1(n757), .B2(
        write2_in[10]), .C1(n1302), .C2(tmp1[10]), .Z(n2147) );
  INVD1BWP12T U1123 ( .I(r5[3]), .ZN(n1923) );
  OAI222D0BWP12T U1124 ( .A1(n1923), .A2(n442), .B1(n426), .B2(n441), .C1(n427), .C2(n440), .ZN(n2460) );
  INVD1BWP12T U1125 ( .I(r11[4]), .ZN(n1882) );
  OAI222D0BWP12T U1126 ( .A1(n424), .A2(n455), .B1(n425), .B2(n454), .C1(n453), 
        .C2(n1882), .ZN(n2269) );
  INVD1BWP12T U1127 ( .I(r0[3]), .ZN(n840) );
  OAI222D0BWP12T U1128 ( .A1(n840), .A2(n449), .B1(n426), .B2(n448), .C1(n427), 
        .C2(n447), .ZN(n2620) );
  OAI222D0BWP12T U1129 ( .A1(n1892), .A2(n458), .B1(n425), .B2(n457), .C1(n424), .C2(n456), .ZN(n2589) );
  INVD1BWP12T U1130 ( .I(r11[3]), .ZN(n601) );
  OAI222D0BWP12T U1131 ( .A1(n427), .A2(n455), .B1(n426), .B2(n454), .C1(n453), 
        .C2(n601), .ZN(n2268) );
  OAI222D0BWP12T U1132 ( .A1(n1911), .A2(n442), .B1(n425), .B2(n441), .C1(n424), .C2(n440), .ZN(n2461) );
  INVD1BWP12T U1133 ( .I(r9[4]), .ZN(n1902) );
  OAI222D0BWP12T U1134 ( .A1(n1902), .A2(n464), .B1(n425), .B2(n463), .C1(n424), .C2(n462), .ZN(n2333) );
  INVD1BWP12T U1135 ( .I(r1[3]), .ZN(n1934) );
  OAI222D0BWP12T U1136 ( .A1(n1934), .A2(n458), .B1(n426), .B2(n457), .C1(n427), .C2(n456), .ZN(n2588) );
  INVD1BWP12T U1137 ( .I(r10[3]), .ZN(n1922) );
  OAI222D0BWP12T U1138 ( .A1(n427), .A2(n467), .B1(n426), .B2(n466), .C1(n465), 
        .C2(n1922), .ZN(n2300) );
  INVD1BWP12T U1139 ( .I(r0[4]), .ZN(n1912) );
  OAI222D0BWP12T U1140 ( .A1(n1912), .A2(n449), .B1(n425), .B2(n448), .C1(n424), .C2(n447), .ZN(n2621) );
  INVD1BWP12T U1141 ( .I(r9[3]), .ZN(n607) );
  OAI222D0BWP12T U1142 ( .A1(n607), .A2(n464), .B1(n426), .B2(n463), .C1(n427), 
        .C2(n462), .ZN(n2332) );
  OAI222D0BWP12T U1143 ( .A1(n424), .A2(n436), .B1(n425), .B2(n435), .C1(n434), 
        .C2(n1908), .ZN(n2525) );
  INVD1BWP12T U1144 ( .I(r7[3]), .ZN(n1928) );
  OAI222D0BWP12T U1145 ( .A1(n1928), .A2(n439), .B1(n426), .B2(n438), .C1(n427), .C2(n437), .ZN(n2396) );
  OAI222D0BWP12T U1146 ( .A1(n424), .A2(n467), .B1(n425), .B2(n466), .C1(n465), 
        .C2(n1886), .ZN(n2301) );
  OAI222D0BWP12T U1147 ( .A1(n1914), .A2(n439), .B1(n425), .B2(n438), .C1(n424), .C2(n437), .ZN(n2397) );
  INVD1BWP12T U1148 ( .I(r3[3]), .ZN(n1936) );
  OAI222D0BWP12T U1149 ( .A1(n427), .A2(n436), .B1(n426), .B2(n435), .C1(n434), 
        .C2(n1936), .ZN(n2524) );
  AO222D0BWP12T U1150 ( .A1(n1303), .A2(write1_in[3]), .B1(n757), .B2(
        write2_in[3]), .C1(n1302), .C2(tmp1[3]), .Z(n2140) );
  INVD1BWP12T U1151 ( .I(write2_in[6]), .ZN(n472) );
  INVD1BWP12T U1152 ( .I(write1_in[6]), .ZN(n474) );
  INVD1BWP12T U1153 ( .I(r2[6]), .ZN(n1738) );
  OAI222D0BWP12T U1154 ( .A1(n472), .A2(n430), .B1(n474), .B2(n429), .C1(n428), 
        .C2(n1738), .ZN(n2559) );
  AO222D0BWP12T U1155 ( .A1(n1303), .A2(write1_in[4]), .B1(n757), .B2(
        write2_in[4]), .C1(n1302), .C2(tmp1[4]), .Z(n2141) );
  INVD1BWP12T U1156 ( .I(r8[6]), .ZN(n1749) );
  OAI222D0BWP12T U1157 ( .A1(n1749), .A2(n433), .B1(n474), .B2(n432), .C1(n472), .C2(n431), .ZN(n2367) );
  INVD1BWP12T U1158 ( .I(r3[6]), .ZN(n1747) );
  OAI222D0BWP12T U1159 ( .A1(n472), .A2(n436), .B1(n474), .B2(n435), .C1(n434), 
        .C2(n1747), .ZN(n2527) );
  INVD1BWP12T U1160 ( .I(r7[6]), .ZN(n1739) );
  OAI222D0BWP12T U1161 ( .A1(n1739), .A2(n439), .B1(n474), .B2(n438), .C1(n472), .C2(n437), .ZN(n2399) );
  INVD1BWP12T U1162 ( .I(r5[6]), .ZN(n1737) );
  OAI222D0BWP12T U1163 ( .A1(n1737), .A2(n442), .B1(n474), .B2(n441), .C1(n472), .C2(n440), .ZN(n2463) );
  CKND0BWP12T U1164 ( .I(r4[6]), .ZN(n446) );
  OAI222D0BWP12T U1165 ( .A1(n446), .A2(n445), .B1(n474), .B2(n444), .C1(n472), 
        .C2(n443), .ZN(n2495) );
  INVD1BWP12T U1166 ( .I(r0[6]), .ZN(n739) );
  OAI222D0BWP12T U1167 ( .A1(n739), .A2(n449), .B1(n474), .B2(n448), .C1(n472), 
        .C2(n447), .ZN(n2623) );
  INVD1BWP12T U1168 ( .I(r6[6]), .ZN(n1750) );
  OAI222D0BWP12T U1169 ( .A1(n1750), .A2(n452), .B1(n474), .B2(n451), .C1(n472), .C2(n450), .ZN(n2431) );
  INVD1BWP12T U1170 ( .I(r11[6]), .ZN(n732) );
  OAI222D0BWP12T U1171 ( .A1(n472), .A2(n455), .B1(n474), .B2(n454), .C1(n453), 
        .C2(n732), .ZN(n2271) );
  INVD1BWP12T U1172 ( .I(r1[6]), .ZN(n1745) );
  OAI222D0BWP12T U1173 ( .A1(n1745), .A2(n458), .B1(n474), .B2(n457), .C1(n472), .C2(n456), .ZN(n2591) );
  INVD1BWP12T U1174 ( .I(r12[6]), .ZN(n1744) );
  OAI222D0BWP12T U1175 ( .A1(n1744), .A2(n461), .B1(n474), .B2(n460), .C1(n472), .C2(n459), .ZN(n2239) );
  INVD1BWP12T U1176 ( .I(r9[6]), .ZN(n738) );
  OAI222D0BWP12T U1177 ( .A1(n738), .A2(n464), .B1(n474), .B2(n463), .C1(n472), 
        .C2(n462), .ZN(n2335) );
  INVD1BWP12T U1178 ( .I(r10[6]), .ZN(n1736) );
  OAI222D0BWP12T U1179 ( .A1(n472), .A2(n467), .B1(n474), .B2(n466), .C1(n465), 
        .C2(n1736), .ZN(n2303) );
  TPAOI21D0BWP12T U1180 ( .A1(n1300), .A2(n[2035]), .B(reset), .ZN(n469) );
  CKND2D0BWP12T U1181 ( .A1(write2_in[6]), .A2(n1299), .ZN(n468) );
  OAI211D0BWP12T U1182 ( .A1(n470), .A2(n474), .B(n469), .C(n468), .ZN(spin[6]) );
  INVD1BWP12T U1183 ( .I(lr[6]), .ZN(n1746) );
  OAI222D0BWP12T U1184 ( .A1(n1746), .A2(n475), .B1(n474), .B2(n473), .C1(n472), .C2(n471), .ZN(n2207) );
  AO222D0BWP12T U1185 ( .A1(n1303), .A2(write1_in[6]), .B1(n757), .B2(
        write2_in[6]), .C1(n1302), .C2(tmp1[6]), .Z(n2143) );
  AO222D0BWP12T U1186 ( .A1(n1280), .A2(write1_in[0]), .B1(n1279), .B2(lr[0]), 
        .C1(write2_in[0]), .C2(n1278), .Z(n2201) );
  AO222D0BWP12T U1187 ( .A1(n1295), .A2(write1_in[0]), .B1(n1294), .B2(
        write2_in[0]), .C1(n1293), .C2(r10[0]), .Z(n2297) );
  AO222D0BWP12T U1188 ( .A1(n1286), .A2(write1_in[0]), .B1(n1285), .B2(r12[0]), 
        .C1(write2_in[0]), .C2(n1284), .Z(n2233) );
  AO222D0BWP12T U1189 ( .A1(n1274), .A2(write1_in[0]), .B1(n1273), .B2(r1[0]), 
        .C1(write2_in[0]), .C2(n1272), .Z(n2585) );
  AO222D0BWP12T U1190 ( .A1(n1289), .A2(write1_in[0]), .B1(n1288), .B2(
        write2_in[0]), .C1(n1287), .C2(r11[0]), .Z(n2265) );
  AO222D0BWP12T U1191 ( .A1(n1265), .A2(write1_in[0]), .B1(n1264), .B2(r0[0]), 
        .C1(write2_in[0]), .C2(n1263), .Z(n2617) );
  AO222D0BWP12T U1192 ( .A1(n1262), .A2(write1_in[0]), .B1(n1261), .B2(r7[0]), 
        .C1(write2_in[0]), .C2(n1260), .Z(n2393) );
  AO222D0BWP12T U1193 ( .A1(n1268), .A2(write1_in[0]), .B1(n1267), .B2(r5[0]), 
        .C1(write2_in[0]), .C2(n1266), .Z(n2457) );
  AO222D0BWP12T U1194 ( .A1(n1277), .A2(write1_in[0]), .B1(n1276), .B2(r4[0]), 
        .C1(write2_in[0]), .C2(n1275), .Z(n2489) );
  AO222D0BWP12T U1195 ( .A1(n1271), .A2(write1_in[0]), .B1(n1270), .B2(r6[0]), 
        .C1(write2_in[0]), .C2(n1269), .Z(n2425) );
  AO222D0BWP12T U1196 ( .A1(n1301), .A2(write1_in[0]), .B1(n1300), .B2(n[2041]), .C1(write2_in[0]), .C2(n1299), .Z(spin[0]) );
  AO222D0BWP12T U1197 ( .A1(n1298), .A2(write1_in[0]), .B1(n1297), .B2(
        write2_in[0]), .C1(n1296), .C2(r3[0]), .Z(n2521) );
  AO222D0BWP12T U1198 ( .A1(n1292), .A2(write1_in[0]), .B1(n1291), .B2(
        write2_in[0]), .C1(n1290), .C2(r2[0]), .Z(n2553) );
  AO222D0BWP12T U1199 ( .A1(n1303), .A2(write1_in[0]), .B1(n757), .B2(
        write2_in[0]), .C1(n1302), .C2(tmp1[0]), .Z(n2136) );
  AO222D0BWP12T U1200 ( .A1(n1259), .A2(write1_in[0]), .B1(n1258), .B2(r8[0]), 
        .C1(write2_in[0]), .C2(n1257), .Z(n2361) );
  AO222D0BWP12T U1201 ( .A1(n1283), .A2(write1_in[0]), .B1(n1282), .B2(r9[0]), 
        .C1(write2_in[0]), .C2(n1281), .Z(n2329) );
  INVD1BWP12T U1202 ( .I(pc_out[20]), .ZN(n476) );
  INVD1BWP12T U1203 ( .I(r11[20]), .ZN(n994) );
  OAI22D1BWP12T U1204 ( .A1(n476), .A2(n1884), .B1(n1883), .B2(n994), .ZN(n484) );
  INVD1BWP12T U1205 ( .I(lr[20]), .ZN(n478) );
  INVD1BWP12T U1206 ( .I(r10[20]), .ZN(n477) );
  OAI22D1BWP12T U1207 ( .A1(n478), .A2(n1888), .B1(n1887), .B2(n477), .ZN(n483) );
  INVD1BWP12T U1208 ( .I(r2[20]), .ZN(n480) );
  INVD1BWP12T U1209 ( .I(r1[20]), .ZN(n479) );
  OAI22D1BWP12T U1210 ( .A1(n1895), .A2(n480), .B1(n1893), .B2(n479), .ZN(n481) );
  NR4D0BWP12T U1211 ( .A1(n484), .A2(n483), .A3(n482), .A4(n481), .ZN(n490) );
  AOI22D1BWP12T U1212 ( .A1(r9[20]), .A2(n1808), .B1(n120), .B2(r6[20]), .ZN(
        n488) );
  AOI22D1BWP12T U1213 ( .A1(r8[20]), .A2(n1810), .B1(n1809), .B2(n[2021]), 
        .ZN(n487) );
  AOI22D1BWP12T U1214 ( .A1(r5[20]), .A2(n123), .B1(n1811), .B2(r3[20]), .ZN(
        n486) );
  AOI22D1BWP12T U1215 ( .A1(r7[20]), .A2(n126), .B1(n1812), .B2(r0[20]), .ZN(
        n485) );
  AN4XD1BWP12T U1216 ( .A1(n488), .A2(n487), .A3(n486), .A4(n485), .Z(n489) );
  CKND2D1BWP12T U1217 ( .A1(n490), .A2(n489), .ZN(regA_out[20]) );
  INVD1BWP12T U1218 ( .I(pc_out[1]), .ZN(n1864) );
  OAI22D1BWP12T U1219 ( .A1(n1864), .A2(n1884), .B1(n1883), .B2(n491), .ZN(
        n496) );
  OAI22D1BWP12T U1220 ( .A1(n1859), .A2(n1888), .B1(n1887), .B2(n1846), .ZN(
        n495) );
  AOI22D1BWP12T U1221 ( .A1(n112), .A2(r12[1]), .B1(n273), .B2(tmp1[1]), .ZN(
        n492) );
  IOA21D1BWP12T U1222 ( .A1(n1891), .A2(r4[1]), .B(n492), .ZN(n494) );
  OAI22D1BWP12T U1223 ( .A1(n1895), .A2(n1851), .B1(n1893), .B2(n1858), .ZN(
        n493) );
  NR4D1BWP12T U1224 ( .A1(n496), .A2(n495), .A3(n494), .A4(n493), .ZN(n504) );
  OAI22D1BWP12T U1225 ( .A1(n1903), .A2(n497), .B1(n1901), .B2(n1863), .ZN(
        n502) );
  INVD1BWP12T U1226 ( .I(n[2040]), .ZN(n1861) );
  OAI22D1BWP12T U1227 ( .A1(n1847), .A2(n1910), .B1(n1909), .B2(n1860), .ZN(
        n500) );
  NR4D0BWP12T U1228 ( .A1(n502), .A2(n501), .A3(n500), .A4(n499), .ZN(n503) );
  TPND2D1BWP12T U1229 ( .A1(n504), .A2(n503), .ZN(regA_out[1]) );
  INVD1BWP12T U1230 ( .I(pc_out[0]), .ZN(n506) );
  INVD1BWP12T U1231 ( .I(r11[0]), .ZN(n505) );
  OAI22D1BWP12T U1232 ( .A1(n506), .A2(n1884), .B1(n1883), .B2(n505), .ZN(n513) );
  INVD1BWP12T U1233 ( .I(lr[0]), .ZN(n972) );
  INVD1BWP12T U1234 ( .I(r10[0]), .ZN(n971) );
  OAI22D1BWP12T U1235 ( .A1(n972), .A2(n1888), .B1(n1887), .B2(n971), .ZN(n512) );
  AOI22D1BWP12T U1236 ( .A1(n112), .A2(r12[0]), .B1(n273), .B2(tmp1[0]), .ZN(
        n507) );
  IOA21D1BWP12T U1237 ( .A1(n1891), .A2(r4[0]), .B(n507), .ZN(n511) );
  INVD1BWP12T U1238 ( .I(r2[0]), .ZN(n509) );
  INVD1BWP12T U1239 ( .I(r1[0]), .ZN(n508) );
  OAI22D1BWP12T U1240 ( .A1(n1895), .A2(n509), .B1(n1893), .B2(n508), .ZN(n510) );
  NR4D0BWP12T U1241 ( .A1(n513), .A2(n512), .A3(n511), .A4(n510), .ZN(n519) );
  AOI22D1BWP12T U1242 ( .A1(r9[0]), .A2(n1808), .B1(n120), .B2(r6[0]), .ZN(
        n517) );
  AOI22D1BWP12T U1243 ( .A1(r8[0]), .A2(n1810), .B1(n1809), .B2(n[2041]), .ZN(
        n516) );
  AOI22D1BWP12T U1244 ( .A1(r5[0]), .A2(n123), .B1(n1811), .B2(r3[0]), .ZN(
        n515) );
  AOI22D1BWP12T U1245 ( .A1(r7[0]), .A2(n126), .B1(n1812), .B2(r0[0]), .ZN(
        n514) );
  AN4XD1BWP12T U1246 ( .A1(n517), .A2(n516), .A3(n515), .A4(n514), .Z(n518) );
  CKND2D1BWP12T U1247 ( .A1(n519), .A2(n518), .ZN(regA_out[0]) );
  INVD1BWP12T U1248 ( .I(pc_out[7]), .ZN(n1724) );
  OAI22D1BWP12T U1249 ( .A1(n1724), .A2(n1884), .B1(n1883), .B2(n520), .ZN(
        n525) );
  OAI22D1BWP12T U1250 ( .A1(n1719), .A2(n1888), .B1(n1887), .B2(n1709), .ZN(
        n524) );
  AOI22D1BWP12T U1251 ( .A1(n112), .A2(r12[7]), .B1(n1684), .B2(tmp1[7]), .ZN(
        n521) );
  IOA21D1BWP12T U1252 ( .A1(n1891), .A2(r4[7]), .B(n521), .ZN(n523) );
  OAI22D1BWP12T U1253 ( .A1(n1895), .A2(n1711), .B1(n1893), .B2(n1718), .ZN(
        n522) );
  NR4D1BWP12T U1254 ( .A1(n525), .A2(n524), .A3(n523), .A4(n522), .ZN(n533) );
  OAI22D1BWP12T U1255 ( .A1(n1903), .A2(n526), .B1(n1901), .B2(n1723), .ZN(
        n531) );
  INVD1BWP12T U1256 ( .I(n[2034]), .ZN(n1721) );
  OAI22D1BWP12T U1257 ( .A1(n1907), .A2(n1722), .B1(n1905), .B2(n1721), .ZN(
        n530) );
  OAI22D1BWP12T U1258 ( .A1(n1710), .A2(n1910), .B1(n1909), .B2(n1720), .ZN(
        n529) );
  OAI22D1BWP12T U1259 ( .A1(n1915), .A2(n1712), .B1(n1913), .B2(n527), .ZN(
        n528) );
  NR4D0BWP12T U1260 ( .A1(n531), .A2(n530), .A3(n529), .A4(n528), .ZN(n532) );
  CKND2D2BWP12T U1261 ( .A1(n533), .A2(n532), .ZN(regA_out[7]) );
  INVD0BWP12T U1262 ( .I(pc_out[14]), .ZN(n535) );
  INVD1BWP12T U1263 ( .I(r11[14]), .ZN(n534) );
  OAI22D1BWP12T U1264 ( .A1(n535), .A2(n1884), .B1(n1883), .B2(n534), .ZN(n541) );
  INVD1BWP12T U1265 ( .I(lr[14]), .ZN(n1067) );
  INVD1BWP12T U1266 ( .I(r10[14]), .ZN(n1065) );
  OAI22D1BWP12T U1267 ( .A1(n1067), .A2(n1888), .B1(n1887), .B2(n1065), .ZN(
        n540) );
  AOI22D1BWP12T U1268 ( .A1(n112), .A2(r12[14]), .B1(n1684), .B2(tmp1[14]), 
        .ZN(n536) );
  IOA21D1BWP12T U1269 ( .A1(n1891), .A2(r4[14]), .B(n536), .ZN(n539) );
  INVD1BWP12T U1270 ( .I(r2[14]), .ZN(n565) );
  INVD1BWP12T U1271 ( .I(r1[14]), .ZN(n537) );
  OAI22D1BWP12T U1272 ( .A1(n1895), .A2(n565), .B1(n1893), .B2(n537), .ZN(n538) );
  NR4D0BWP12T U1273 ( .A1(n541), .A2(n540), .A3(n539), .A4(n538), .ZN(n547) );
  AOI22D1BWP12T U1274 ( .A1(r9[14]), .A2(n1808), .B1(n120), .B2(r6[14]), .ZN(
        n545) );
  AOI22D1BWP12T U1275 ( .A1(r8[14]), .A2(n1810), .B1(n1809), .B2(n[2027]), 
        .ZN(n544) );
  AOI22D1BWP12T U1276 ( .A1(r5[14]), .A2(n123), .B1(n1811), .B2(r3[14]), .ZN(
        n543) );
  AOI22D1BWP12T U1277 ( .A1(r7[14]), .A2(n126), .B1(n1812), .B2(r0[14]), .ZN(
        n542) );
  AN4XD1BWP12T U1278 ( .A1(n545), .A2(n544), .A3(n543), .A4(n542), .Z(n546) );
  CKND2D1BWP12T U1279 ( .A1(n547), .A2(n546), .ZN(regA_out[14]) );
  INVD1BWP12T U1280 ( .I(pc_out[5]), .ZN(n1839) );
  OAI22D1BWP12T U1281 ( .A1(n1839), .A2(n1884), .B1(n1883), .B2(n548), .ZN(
        n553) );
  OAI22D1BWP12T U1282 ( .A1(n1834), .A2(n1888), .B1(n1887), .B2(n1824), .ZN(
        n552) );
  IOA21D1BWP12T U1283 ( .A1(n1891), .A2(r4[5]), .B(n549), .ZN(n551) );
  OAI22D1BWP12T U1284 ( .A1(n1895), .A2(n1826), .B1(n1893), .B2(n1833), .ZN(
        n550) );
  NR4D1BWP12T U1285 ( .A1(n553), .A2(n552), .A3(n551), .A4(n550), .ZN(n560) );
  OAI22D1BWP12T U1286 ( .A1(n1903), .A2(n983), .B1(n1901), .B2(n1838), .ZN(
        n558) );
  INVD1BWP12T U1287 ( .I(n[2036]), .ZN(n1836) );
  OAI22D1BWP12T U1288 ( .A1(n1825), .A2(n1910), .B1(n1909), .B2(n1835), .ZN(
        n556) );
  OAI22D1BWP12T U1289 ( .A1(n1915), .A2(n1827), .B1(n1913), .B2(n554), .ZN(
        n555) );
  CKND2D2BWP12T U1290 ( .A1(n560), .A2(n559), .ZN(regA_out[5]) );
  INVD1BWP12T U1291 ( .I(tmp1[14]), .ZN(n561) );
  MOAI22D0BWP12T U1292 ( .A1(n561), .A2(n1951), .B1(n150), .B2(
        immediate2_in[14]), .ZN(n570) );
  AOI22D1BWP12T U1293 ( .A1(r9[14]), .A2(n152), .B1(n1732), .B2(r4[14]), .ZN(
        n563) );
  BUFFD3BWP12T U1294 ( .I(n1955), .Z(n1571) );
  AOI22D1BWP12T U1295 ( .A1(r11[14]), .A2(n1571), .B1(n1733), .B2(r0[14]), 
        .ZN(n562) );
  ND2D1BWP12T U1296 ( .A1(n563), .A2(n562), .ZN(n569) );
  INVD1BWP12T U1297 ( .I(r5[14]), .ZN(n564) );
  OAI22D1BWP12T U1298 ( .A1(n564), .A2(n1949), .B1(n1948), .B2(n1065), .ZN(
        n568) );
  INVD1BWP12T U1299 ( .I(r7[14]), .ZN(n566) );
  OAI22D1BWP12T U1300 ( .A1(n1961), .A2(n566), .B1(n1959), .B2(n565), .ZN(n567) );
  NR4D0BWP12T U1301 ( .A1(n570), .A2(n569), .A3(n568), .A4(n567), .ZN(n576) );
  AOI22D1BWP12T U1302 ( .A1(r1[14]), .A2(n164), .B1(n1993), .B2(r12[14]), .ZN(
        n574) );
  AOI22D1BWP12T U1303 ( .A1(r3[14]), .A2(n1994), .B1(n168), .B2(lr[14]), .ZN(
        n573) );
  AOI22D1BWP12T U1304 ( .A1(r8[14]), .A2(n171), .B1(n1995), .B2(n[2027]), .ZN(
        n572) );
  AOI22D1BWP12T U1305 ( .A1(pc_out[14]), .A2(n174), .B1(n1996), .B2(r6[14]), 
        .ZN(n571) );
  AN4XD1BWP12T U1306 ( .A1(n574), .A2(n573), .A3(n572), .A4(n571), .Z(n575) );
  CKND2D1BWP12T U1307 ( .A1(n576), .A2(n575), .ZN(regB_out[14]) );
  OAI22D1BWP12T U1308 ( .A1(n578), .A2(n1884), .B1(n1883), .B2(n577), .ZN(n587) );
  OAI22D1BWP12T U1309 ( .A1(n580), .A2(n1888), .B1(n1887), .B2(n579), .ZN(n586) );
  AOI22D1BWP12T U1310 ( .A1(n112), .A2(r12[11]), .B1(n1684), .B2(tmp1[11]), 
        .ZN(n581) );
  IOA21D1BWP12T U1311 ( .A1(n1891), .A2(r4[11]), .B(n581), .ZN(n585) );
  OAI22D1BWP12T U1312 ( .A1(n1895), .A2(n583), .B1(n1893), .B2(n582), .ZN(n584) );
  NR4D0BWP12T U1313 ( .A1(n587), .A2(n586), .A3(n585), .A4(n584), .ZN(n600) );
  OAI22D1BWP12T U1314 ( .A1(n1903), .A2(n589), .B1(n1901), .B2(n588), .ZN(n598) );
  OAI22D1BWP12T U1315 ( .A1(n1907), .A2(n590), .B1(n1905), .B2(n1090), .ZN(
        n597) );
  OAI22D1BWP12T U1316 ( .A1(n592), .A2(n1910), .B1(n1909), .B2(n591), .ZN(n596) );
  OAI22D1BWP12T U1317 ( .A1(n1915), .A2(n594), .B1(n1913), .B2(n593), .ZN(n595) );
  NR4D0BWP12T U1318 ( .A1(n598), .A2(n597), .A3(n596), .A4(n595), .ZN(n599) );
  INVD1BWP12T U1319 ( .I(pc_out[3]), .ZN(n1940) );
  OAI22D1BWP12T U1320 ( .A1(n1940), .A2(n1884), .B1(n1883), .B2(n601), .ZN(
        n606) );
  OAI22D1BWP12T U1321 ( .A1(n1935), .A2(n1888), .B1(n1887), .B2(n1922), .ZN(
        n605) );
  AOI22D1BWP12T U1322 ( .A1(n112), .A2(r12[3]), .B1(n1684), .B2(tmp1[3]), .ZN(
        n602) );
  IOA21D1BWP12T U1323 ( .A1(n1891), .A2(r4[3]), .B(n602), .ZN(n604) );
  OAI22D1BWP12T U1324 ( .A1(n1895), .A2(n1927), .B1(n1893), .B2(n1934), .ZN(
        n603) );
  NR4D0BWP12T U1325 ( .A1(n606), .A2(n605), .A3(n604), .A4(n603), .ZN(n613) );
  OAI22D1BWP12T U1326 ( .A1(n1903), .A2(n607), .B1(n1901), .B2(n1939), .ZN(
        n611) );
  INVD1BWP12T U1327 ( .I(n[2038]), .ZN(n1937) );
  OAI22D1BWP12T U1328 ( .A1(n1907), .A2(n1938), .B1(n1905), .B2(n1937), .ZN(
        n610) );
  OAI22D1BWP12T U1329 ( .A1(n1915), .A2(n1928), .B1(n1913), .B2(n840), .ZN(
        n608) );
  NR4D0BWP12T U1330 ( .A1(n611), .A2(n610), .A3(n609), .A4(n608), .ZN(n612) );
  ND2D1BWP12T U1331 ( .A1(n613), .A2(n612), .ZN(regA_out[3]) );
  INVD0BWP12T U1332 ( .I(tmp1[9]), .ZN(n614) );
  MOAI22D0BWP12T U1333 ( .A1(n614), .A2(n1951), .B1(n150), .B2(
        immediate2_in[9]), .ZN(n624) );
  AOI22D1BWP12T U1334 ( .A1(r9[9]), .A2(n152), .B1(n1732), .B2(r4[9]), .ZN(
        n616) );
  AOI22D1BWP12T U1335 ( .A1(r11[9]), .A2(n1955), .B1(n1733), .B2(r0[9]), .ZN(
        n615) );
  ND2D1BWP12T U1336 ( .A1(n616), .A2(n615), .ZN(n623) );
  OAI22D1BWP12T U1337 ( .A1(n618), .A2(n1949), .B1(n1948), .B2(n617), .ZN(n622) );
  OAI22D1BWP12T U1338 ( .A1(n1961), .A2(n620), .B1(n1959), .B2(n619), .ZN(n621) );
  NR4D0BWP12T U1339 ( .A1(n624), .A2(n623), .A3(n622), .A4(n621), .ZN(n637) );
  OAI22D1BWP12T U1340 ( .A1(n626), .A2(n1968), .B1(n1967), .B2(n625), .ZN(n635) );
  OAI22D1BWP12T U1341 ( .A1(n628), .A2(n1972), .B1(n1971), .B2(n627), .ZN(n634) );
  OAI22D1BWP12T U1342 ( .A1(n1977), .A2(n1054), .B1(n1975), .B2(n629), .ZN(
        n633) );
  OAI22D1BWP12T U1343 ( .A1(n1981), .A2(n631), .B1(n1979), .B2(n630), .ZN(n632) );
  NR4D0BWP12T U1344 ( .A1(n635), .A2(n634), .A3(n633), .A4(n632), .ZN(n636) );
  CKND2D1BWP12T U1345 ( .A1(n637), .A2(n636), .ZN(regB_out[9]) );
  AOI22D0BWP12T U1346 ( .A1(r8[3]), .A2(n705), .B1(n704), .B2(r4[3]), .ZN(n639) );
  AOI22D0BWP12T U1347 ( .A1(n[2038]), .A2(n707), .B1(n706), .B2(r10[3]), .ZN(
        n638) );
  CKND2D1BWP12T U1348 ( .A1(n639), .A2(n638), .ZN(n648) );
  AOI22D0BWP12T U1349 ( .A1(r7[3]), .A2(n711), .B1(n710), .B2(r5[3]), .ZN(n643) );
  AOI22D0BWP12T U1350 ( .A1(lr[3]), .A2(n713), .B1(n712), .B2(r9[3]), .ZN(n642) );
  AOI22D0BWP12T U1351 ( .A1(r6[3]), .A2(n715), .B1(n714), .B2(r11[3]), .ZN(
        n641) );
  CKND2D0BWP12T U1352 ( .A1(n716), .A2(r12[3]), .ZN(n640) );
  ND4D1BWP12T U1353 ( .A1(n643), .A2(n642), .A3(n641), .A4(n640), .ZN(n647) );
  AOI22D0BWP12T U1354 ( .A1(r3[3]), .A2(n722), .B1(n721), .B2(r2[3]), .ZN(n645) );
  AOI22D0BWP12T U1355 ( .A1(n724), .A2(r0[3]), .B1(pc_out[3]), .B2(n723), .ZN(
        n644) );
  OAI211D0BWP12T U1356 ( .A1(n1934), .A2(n727), .B(n645), .C(n644), .ZN(n646)
         );
  OA31D0BWP12T U1357 ( .A1(n648), .A2(n647), .A3(n646), .B(n728), .Z(
        regD_out[3]) );
  AOI22D0BWP12T U1358 ( .A1(r8[10]), .A2(n705), .B1(n704), .B2(r4[10]), .ZN(
        n650) );
  AOI22D0BWP12T U1359 ( .A1(n[2031]), .A2(n707), .B1(n706), .B2(r10[10]), .ZN(
        n649) );
  CKND2D1BWP12T U1360 ( .A1(n650), .A2(n649), .ZN(n659) );
  AOI22D0BWP12T U1361 ( .A1(r7[10]), .A2(n711), .B1(n710), .B2(r5[10]), .ZN(
        n654) );
  AOI22D0BWP12T U1362 ( .A1(lr[10]), .A2(n713), .B1(n712), .B2(r9[10]), .ZN(
        n653) );
  AOI22D0BWP12T U1363 ( .A1(r6[10]), .A2(n715), .B1(n714), .B2(r11[10]), .ZN(
        n652) );
  CKND2D0BWP12T U1364 ( .A1(n716), .A2(r12[10]), .ZN(n651) );
  ND4D1BWP12T U1365 ( .A1(n654), .A2(n653), .A3(n652), .A4(n651), .ZN(n658) );
  AOI22D0BWP12T U1366 ( .A1(r3[10]), .A2(n722), .B1(n721), .B2(r2[10]), .ZN(
        n656) );
  AOI22D0BWP12T U1367 ( .A1(n724), .A2(r0[10]), .B1(pc_out[10]), .B2(n723), 
        .ZN(n655) );
  OAI211D0BWP12T U1368 ( .A1(n1660), .A2(n727), .B(n656), .C(n655), .ZN(n657)
         );
  OA31D0BWP12T U1369 ( .A1(n659), .A2(n658), .A3(n657), .B(n728), .Z(
        regD_out[10]) );
  AOI22D0BWP12T U1370 ( .A1(r8[4]), .A2(n705), .B1(n704), .B2(r4[4]), .ZN(n661) );
  AOI22D0BWP12T U1371 ( .A1(n[2037]), .A2(n707), .B1(n706), .B2(r10[4]), .ZN(
        n660) );
  CKND2D1BWP12T U1372 ( .A1(n661), .A2(n660), .ZN(n670) );
  AOI22D0BWP12T U1373 ( .A1(r7[4]), .A2(n711), .B1(n710), .B2(r5[4]), .ZN(n665) );
  AOI22D0BWP12T U1374 ( .A1(lr[4]), .A2(n713), .B1(n712), .B2(r9[4]), .ZN(n664) );
  AOI22D0BWP12T U1375 ( .A1(r6[4]), .A2(n715), .B1(n714), .B2(r11[4]), .ZN(
        n663) );
  CKND2D0BWP12T U1376 ( .A1(n716), .A2(r12[4]), .ZN(n662) );
  ND4D1BWP12T U1377 ( .A1(n665), .A2(n664), .A3(n663), .A4(n662), .ZN(n669) );
  AOI22D0BWP12T U1378 ( .A1(r3[4]), .A2(n722), .B1(n721), .B2(r2[4]), .ZN(n667) );
  AOI22D0BWP12T U1379 ( .A1(n724), .A2(r0[4]), .B1(pc_out[4]), .B2(n723), .ZN(
        n666) );
  OAI211D0BWP12T U1380 ( .A1(n1892), .A2(n727), .B(n667), .C(n666), .ZN(n668)
         );
  OA31D0BWP12T U1381 ( .A1(n670), .A2(n669), .A3(n668), .B(n728), .Z(
        regD_out[4]) );
  AOI22D0BWP12T U1382 ( .A1(r8[5]), .A2(n705), .B1(n704), .B2(r4[5]), .ZN(n672) );
  AOI22D0BWP12T U1383 ( .A1(n[2036]), .A2(n707), .B1(n706), .B2(r10[5]), .ZN(
        n671) );
  CKND2D1BWP12T U1384 ( .A1(n672), .A2(n671), .ZN(n681) );
  AOI22D0BWP12T U1385 ( .A1(r7[5]), .A2(n711), .B1(n710), .B2(r5[5]), .ZN(n676) );
  AOI22D0BWP12T U1386 ( .A1(lr[5]), .A2(n713), .B1(n712), .B2(r9[5]), .ZN(n675) );
  AOI22D0BWP12T U1387 ( .A1(r6[5]), .A2(n715), .B1(n714), .B2(r11[5]), .ZN(
        n674) );
  CKND2D0BWP12T U1388 ( .A1(n716), .A2(r12[5]), .ZN(n673) );
  ND4D1BWP12T U1389 ( .A1(n676), .A2(n675), .A3(n674), .A4(n673), .ZN(n680) );
  AOI22D0BWP12T U1390 ( .A1(r3[5]), .A2(n722), .B1(n721), .B2(r2[5]), .ZN(n678) );
  AOI22D0BWP12T U1391 ( .A1(n724), .A2(r0[5]), .B1(pc_out[5]), .B2(n723), .ZN(
        n677) );
  OAI211D0BWP12T U1392 ( .A1(n1833), .A2(n727), .B(n678), .C(n677), .ZN(n679)
         );
  OA31D0BWP12T U1393 ( .A1(n681), .A2(n680), .A3(n679), .B(n728), .Z(
        regD_out[5]) );
  AOI22D0BWP12T U1394 ( .A1(r8[8]), .A2(n705), .B1(n704), .B2(r4[8]), .ZN(n683) );
  AOI22D0BWP12T U1395 ( .A1(n[2033]), .A2(n707), .B1(n706), .B2(r10[8]), .ZN(
        n682) );
  CKND2D1BWP12T U1396 ( .A1(n683), .A2(n682), .ZN(n692) );
  AOI22D0BWP12T U1397 ( .A1(r7[8]), .A2(n711), .B1(n710), .B2(r5[8]), .ZN(n687) );
  AOI22D0BWP12T U1398 ( .A1(lr[8]), .A2(n713), .B1(n712), .B2(r9[8]), .ZN(n686) );
  AOI22D0BWP12T U1399 ( .A1(r6[8]), .A2(n715), .B1(n714), .B2(r11[8]), .ZN(
        n685) );
  CKND2D0BWP12T U1400 ( .A1(n716), .A2(r12[8]), .ZN(n684) );
  ND4D1BWP12T U1401 ( .A1(n687), .A2(n686), .A3(n685), .A4(n684), .ZN(n691) );
  AOI22D0BWP12T U1402 ( .A1(r3[8]), .A2(n722), .B1(n721), .B2(r2[8]), .ZN(n689) );
  AOI22D0BWP12T U1403 ( .A1(n724), .A2(r0[8]), .B1(pc_out[8]), .B2(n723), .ZN(
        n688) );
  OAI211D0BWP12T U1404 ( .A1(n1686), .A2(n727), .B(n689), .C(n688), .ZN(n690)
         );
  OA31D0BWP12T U1405 ( .A1(n692), .A2(n691), .A3(n690), .B(n728), .Z(
        regD_out[8]) );
  AOI22D0BWP12T U1406 ( .A1(r8[6]), .A2(n705), .B1(n704), .B2(r4[6]), .ZN(n694) );
  AOI22D0BWP12T U1407 ( .A1(n[2035]), .A2(n707), .B1(n706), .B2(r10[6]), .ZN(
        n693) );
  CKND2D1BWP12T U1408 ( .A1(n694), .A2(n693), .ZN(n703) );
  AOI22D0BWP12T U1409 ( .A1(r7[6]), .A2(n711), .B1(n710), .B2(r5[6]), .ZN(n698) );
  AOI22D0BWP12T U1410 ( .A1(lr[6]), .A2(n713), .B1(n712), .B2(r9[6]), .ZN(n697) );
  AOI22D0BWP12T U1411 ( .A1(r6[6]), .A2(n715), .B1(n714), .B2(r11[6]), .ZN(
        n696) );
  CKND2D0BWP12T U1412 ( .A1(n716), .A2(r12[6]), .ZN(n695) );
  ND4D1BWP12T U1413 ( .A1(n698), .A2(n697), .A3(n696), .A4(n695), .ZN(n702) );
  AOI22D0BWP12T U1414 ( .A1(r3[6]), .A2(n722), .B1(n721), .B2(r2[6]), .ZN(n700) );
  AOI22D0BWP12T U1415 ( .A1(n724), .A2(r0[6]), .B1(pc_out[6]), .B2(n723), .ZN(
        n699) );
  OAI211D0BWP12T U1416 ( .A1(n1745), .A2(n727), .B(n700), .C(n699), .ZN(n701)
         );
  OA31D0BWP12T U1417 ( .A1(n703), .A2(n702), .A3(n701), .B(n728), .Z(
        regD_out[6]) );
  AOI22D0BWP12T U1418 ( .A1(r8[2]), .A2(n705), .B1(n704), .B2(r4[2]), .ZN(n709) );
  AOI22D0BWP12T U1419 ( .A1(n[2039]), .A2(n707), .B1(n706), .B2(r10[2]), .ZN(
        n708) );
  CKND2D1BWP12T U1420 ( .A1(n709), .A2(n708), .ZN(n731) );
  AOI22D0BWP12T U1421 ( .A1(r7[2]), .A2(n711), .B1(n710), .B2(r5[2]), .ZN(n720) );
  AOI22D0BWP12T U1422 ( .A1(lr[2]), .A2(n713), .B1(n712), .B2(r9[2]), .ZN(n719) );
  AOI22D0BWP12T U1423 ( .A1(r6[2]), .A2(n715), .B1(n714), .B2(r11[2]), .ZN(
        n718) );
  CKND2D0BWP12T U1424 ( .A1(n716), .A2(r12[2]), .ZN(n717) );
  ND4D1BWP12T U1425 ( .A1(n720), .A2(n719), .A3(n718), .A4(n717), .ZN(n730) );
  AOI22D0BWP12T U1426 ( .A1(r3[2]), .A2(n722), .B1(n721), .B2(r2[2]), .ZN(n726) );
  AOI22D0BWP12T U1427 ( .A1(n724), .A2(r0[2]), .B1(pc_out[2]), .B2(n723), .ZN(
        n725) );
  OAI211D0BWP12T U1428 ( .A1(n1969), .A2(n727), .B(n726), .C(n725), .ZN(n729)
         );
  OA31D0BWP12T U1429 ( .A1(n731), .A2(n730), .A3(n729), .B(n728), .Z(
        regD_out[2]) );
  INVD1BWP12T U1430 ( .I(pc_out[6]), .ZN(n1751) );
  OAI22D1BWP12T U1431 ( .A1(n1751), .A2(n1884), .B1(n1883), .B2(n732), .ZN(
        n737) );
  OAI22D1BWP12T U1432 ( .A1(n1746), .A2(n1888), .B1(n1887), .B2(n1736), .ZN(
        n736) );
  AOI22D1BWP12T U1433 ( .A1(n112), .A2(r12[6]), .B1(n1684), .B2(tmp1[6]), .ZN(
        n733) );
  IOA21D1BWP12T U1434 ( .A1(n1891), .A2(r4[6]), .B(n733), .ZN(n735) );
  OAI22D1BWP12T U1435 ( .A1(n1895), .A2(n1738), .B1(n1893), .B2(n1745), .ZN(
        n734) );
  NR4D0BWP12T U1436 ( .A1(n737), .A2(n736), .A3(n735), .A4(n734), .ZN(n745) );
  OAI22D1BWP12T U1437 ( .A1(n1903), .A2(n738), .B1(n1901), .B2(n1750), .ZN(
        n743) );
  INVD1BWP12T U1438 ( .I(n[2035]), .ZN(n1748) );
  OAI22D1BWP12T U1439 ( .A1(n1907), .A2(n1749), .B1(n1905), .B2(n1748), .ZN(
        n742) );
  OAI22D1BWP12T U1440 ( .A1(n1737), .A2(n1910), .B1(n1909), .B2(n1747), .ZN(
        n741) );
  OAI22D1BWP12T U1441 ( .A1(n1915), .A2(n1739), .B1(n1913), .B2(n739), .ZN(
        n740) );
  NR4D0BWP12T U1442 ( .A1(n743), .A2(n742), .A3(n741), .A4(n740), .ZN(n744) );
  AOI22D1BWP12T U1443 ( .A1(r1[21]), .A2(n164), .B1(n1993), .B2(r12[21]), .ZN(
        n749) );
  AOI22D1BWP12T U1444 ( .A1(r3[21]), .A2(n1994), .B1(n168), .B2(lr[21]), .ZN(
        n748) );
  AOI22D1BWP12T U1445 ( .A1(r8[21]), .A2(n171), .B1(n1995), .B2(n[2020]), .ZN(
        n747) );
  AOI22D1BWP12T U1446 ( .A1(pc_out[21]), .A2(n174), .B1(n1996), .B2(r6[21]), 
        .ZN(n746) );
  AN4XD1BWP12T U1447 ( .A1(n749), .A2(n748), .A3(n747), .A4(n746), .Z(n756) );
  AOI22D1BWP12T U1448 ( .A1(tmp1[21]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[21]), .ZN(n752) );
  AOI22D1BWP12T U1449 ( .A1(r9[21]), .A2(n152), .B1(n2002), .B2(r4[21]), .ZN(
        n751) );
  AOI22D1BWP12T U1450 ( .A1(r11[21]), .A2(n1955), .B1(n1954), .B2(r0[21]), 
        .ZN(n750) );
  AN3XD1BWP12T U1451 ( .A1(n752), .A2(n751), .A3(n750), .Z(n755) );
  AOI22D1BWP12T U1452 ( .A1(r5[21]), .A2(n1988), .B1(n158), .B2(r10[21]), .ZN(
        n754) );
  AOI22D1BWP12T U1453 ( .A1(r7[21]), .A2(n1990), .B1(n1989), .B2(r2[21]), .ZN(
        n753) );
  AO222D0BWP12T U1454 ( .A1(n1277), .A2(n1346), .B1(n1276), .B2(r4[28]), .C1(
        write2_in[28]), .C2(n1275), .Z(n2517) );
  AO222D0BWP12T U1455 ( .A1(n1259), .A2(n1346), .B1(n1258), .B2(r8[28]), .C1(
        write2_in[28]), .C2(n1257), .Z(n2389) );
  AO222D0BWP12T U1456 ( .A1(n1271), .A2(n1346), .B1(n1270), .B2(r6[28]), .C1(
        write2_in[28]), .C2(n1269), .Z(n2453) );
  AO222D0BWP12T U1457 ( .A1(n1274), .A2(n1346), .B1(n1273), .B2(r1[28]), .C1(
        write2_in[28]), .C2(n1272), .Z(n2613) );
  AO222D0BWP12T U1458 ( .A1(n1268), .A2(n1346), .B1(n1267), .B2(r5[28]), .C1(
        write2_in[28]), .C2(n1266), .Z(n2485) );
  AO222D0BWP12T U1459 ( .A1(n1283), .A2(n1346), .B1(n1282), .B2(r9[28]), .C1(
        write2_in[28]), .C2(n1281), .Z(n2357) );
  AO222D0BWP12T U1460 ( .A1(n1265), .A2(n1346), .B1(n1264), .B2(r0[28]), .C1(
        write2_in[28]), .C2(n1263), .Z(n2645) );
  AO222D0BWP12T U1461 ( .A1(n1262), .A2(n1346), .B1(n1261), .B2(r7[28]), .C1(
        write2_in[28]), .C2(n1260), .Z(n2421) );
  AO222D0BWP12T U1462 ( .A1(n1292), .A2(n1346), .B1(n1291), .B2(write2_in[28]), 
        .C1(n1290), .C2(r2[28]), .Z(n2581) );
  AO222D0BWP12T U1463 ( .A1(n1298), .A2(n1346), .B1(n1297), .B2(write2_in[28]), 
        .C1(n1296), .C2(r3[28]), .Z(n2549) );
  AO222D0BWP12T U1464 ( .A1(n1289), .A2(n1346), .B1(n1288), .B2(write2_in[28]), 
        .C1(n1287), .C2(r11[28]), .Z(n2293) );
  BUFFD3BWP12T U1465 ( .I(write1_in[16]), .Z(n1247) );
  AO222D0BWP12T U1466 ( .A1(n1262), .A2(n1247), .B1(n1261), .B2(r7[16]), .C1(
        write2_in[16]), .C2(n1260), .Z(n2409) );
  AO222D0BWP12T U1467 ( .A1(n1277), .A2(n1247), .B1(n1276), .B2(r4[16]), .C1(
        write2_in[16]), .C2(n1275), .Z(n2505) );
  AO222D0BWP12T U1468 ( .A1(n1268), .A2(n1247), .B1(n1267), .B2(r5[16]), .C1(
        write2_in[16]), .C2(n1266), .Z(n2473) );
  AO222D0BWP12T U1469 ( .A1(n1280), .A2(n1247), .B1(n1279), .B2(lr[16]), .C1(
        write2_in[16]), .C2(n1278), .Z(n2217) );
  AO222D0BWP12T U1470 ( .A1(n1283), .A2(n1247), .B1(n1282), .B2(r9[16]), .C1(
        write2_in[16]), .C2(n1281), .Z(n2345) );
  AO222D0BWP12T U1471 ( .A1(n1286), .A2(n1247), .B1(n1285), .B2(r12[16]), .C1(
        write2_in[16]), .C2(n1284), .Z(n2249) );
  AO222D0BWP12T U1472 ( .A1(n1259), .A2(n1247), .B1(n1258), .B2(r8[16]), .C1(
        write2_in[16]), .C2(n1257), .Z(n2377) );
  AO222D0BWP12T U1473 ( .A1(n1265), .A2(n1247), .B1(n1264), .B2(r0[16]), .C1(
        write2_in[16]), .C2(n1263), .Z(n2633) );
  AO222D0BWP12T U1474 ( .A1(n1271), .A2(n1247), .B1(n1270), .B2(r6[16]), .C1(
        write2_in[16]), .C2(n1269), .Z(n2441) );
  AO222D0BWP12T U1475 ( .A1(n1274), .A2(n1247), .B1(n1273), .B2(r1[16]), .C1(
        write2_in[16]), .C2(n1272), .Z(n2601) );
  AO222D0BWP12T U1476 ( .A1(n1301), .A2(n1247), .B1(n1300), .B2(n[2025]), .C1(
        write2_in[16]), .C2(n1299), .Z(spin[16]) );
  AO222D0BWP12T U1477 ( .A1(n1303), .A2(n1247), .B1(n757), .B2(write2_in[16]), 
        .C1(n1302), .C2(tmp1[16]), .Z(n2153) );
  AO222D0BWP12T U1478 ( .A1(n1295), .A2(n1247), .B1(n1294), .B2(write2_in[16]), 
        .C1(n1293), .C2(r10[16]), .Z(n2313) );
  AO222D0BWP12T U1479 ( .A1(n1298), .A2(n1247), .B1(n1297), .B2(write2_in[16]), 
        .C1(n1296), .C2(r3[16]), .Z(n2537) );
  AO222D0BWP12T U1480 ( .A1(n1292), .A2(n1247), .B1(n1291), .B2(write2_in[16]), 
        .C1(n1290), .C2(r2[16]), .Z(n2569) );
  AO222D0BWP12T U1481 ( .A1(n1289), .A2(n1247), .B1(n1288), .B2(write2_in[16]), 
        .C1(n1287), .C2(r11[16]), .Z(n2281) );
  AO222D0BWP12T U1482 ( .A1(n1298), .A2(n1352), .B1(n1297), .B2(write2_in[30]), 
        .C1(n1296), .C2(r3[30]), .Z(n2551) );
  AO222D0BWP12T U1483 ( .A1(n1292), .A2(n1352), .B1(n1291), .B2(write2_in[30]), 
        .C1(n1290), .C2(r2[30]), .Z(n2583) );
  AO222D0BWP12T U1484 ( .A1(n1303), .A2(write1_in[2]), .B1(n757), .B2(
        write2_in[2]), .C1(n1302), .C2(tmp1[2]), .Z(n2139) );
  AO222D0BWP12T U1485 ( .A1(write1_in[31]), .A2(n1303), .B1(write2_in[31]), 
        .B2(n757), .C1(n1302), .C2(tmp1[31]), .Z(n2168) );
  AO222D0BWP12T U1486 ( .A1(write1_in[31]), .A2(n1301), .B1(write2_in[31]), 
        .B2(n1299), .C1(n[2010]), .C2(n1300), .Z(spin[31]) );
  AO222D0BWP12T U1487 ( .A1(write1_in[31]), .A2(n1295), .B1(write2_in[31]), 
        .B2(n1294), .C1(n1293), .C2(r10[31]), .Z(n2328) );
  AO222D0BWP12T U1488 ( .A1(write1_in[31]), .A2(n1265), .B1(write2_in[31]), 
        .B2(n1263), .C1(r0[31]), .C2(n1264), .Z(n2648) );
  AO222D0BWP12T U1489 ( .A1(write1_in[31]), .A2(n1277), .B1(write2_in[31]), 
        .B2(n1275), .C1(r4[31]), .C2(n1276), .Z(n2520) );
  AO222D0BWP12T U1490 ( .A1(write1_in[31]), .A2(n1274), .B1(write2_in[31]), 
        .B2(n1272), .C1(r1[31]), .C2(n1273), .Z(n2616) );
  AO222D0BWP12T U1491 ( .A1(write1_in[31]), .A2(n1268), .B1(write2_in[31]), 
        .B2(n1266), .C1(r5[31]), .C2(n1267), .Z(n2488) );
  AO222D0BWP12T U1492 ( .A1(write1_in[31]), .A2(n1271), .B1(write2_in[31]), 
        .B2(n1269), .C1(r6[31]), .C2(n1270), .Z(n2456) );
  AO222D0BWP12T U1493 ( .A1(write1_in[31]), .A2(n1262), .B1(write2_in[31]), 
        .B2(n1260), .C1(r7[31]), .C2(n1261), .Z(n2424) );
  AO222D0BWP12T U1494 ( .A1(write1_in[31]), .A2(n1280), .B1(write2_in[31]), 
        .B2(n1278), .C1(lr[31]), .C2(n1279), .Z(n2232) );
  AO222D0BWP12T U1495 ( .A1(write1_in[31]), .A2(n1259), .B1(write2_in[31]), 
        .B2(n1257), .C1(r8[31]), .C2(n1258), .Z(n2392) );
  AO222D0BWP12T U1496 ( .A1(write1_in[31]), .A2(n1289), .B1(write2_in[31]), 
        .B2(n1288), .C1(n1287), .C2(r11[31]), .Z(n2296) );
  AO222D0BWP12T U1497 ( .A1(write1_in[31]), .A2(n1283), .B1(write2_in[31]), 
        .B2(n1281), .C1(r9[31]), .C2(n1282), .Z(n2360) );
  AO222D0BWP12T U1498 ( .A1(write1_in[31]), .A2(n1286), .B1(write2_in[31]), 
        .B2(n1284), .C1(r12[31]), .C2(n1285), .Z(n2264) );
  AO222D0BWP12T U1499 ( .A1(write1_in[31]), .A2(n1292), .B1(write2_in[31]), 
        .B2(n1291), .C1(n1290), .C2(r2[31]), .Z(n2584) );
  AO222D0BWP12T U1500 ( .A1(write1_in[31]), .A2(n1298), .B1(write2_in[31]), 
        .B2(n1297), .C1(n1296), .C2(r3[31]), .Z(n2552) );
  AOI22D1BWP12T U1501 ( .A1(r1[24]), .A2(n164), .B1(n1993), .B2(r12[24]), .ZN(
        n761) );
  AOI22D1BWP12T U1502 ( .A1(r3[24]), .A2(n1994), .B1(n168), .B2(lr[24]), .ZN(
        n760) );
  AOI22D1BWP12T U1503 ( .A1(r8[24]), .A2(n171), .B1(n1995), .B2(n[2017]), .ZN(
        n759) );
  AOI22D1BWP12T U1504 ( .A1(pc_out[24]), .A2(n174), .B1(n1996), .B2(r6[24]), 
        .ZN(n758) );
  AN4XD1BWP12T U1505 ( .A1(n761), .A2(n760), .A3(n759), .A4(n758), .Z(n768) );
  AOI22D1BWP12T U1506 ( .A1(tmp1[24]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[24]), .ZN(n764) );
  AOI22D1BWP12T U1507 ( .A1(r9[24]), .A2(n152), .B1(n2002), .B2(r4[24]), .ZN(
        n763) );
  AOI22D1BWP12T U1508 ( .A1(r11[24]), .A2(n1571), .B1(n1954), .B2(r0[24]), 
        .ZN(n762) );
  AN3XD1BWP12T U1509 ( .A1(n764), .A2(n763), .A3(n762), .Z(n767) );
  AOI22D1BWP12T U1510 ( .A1(r5[24]), .A2(n1988), .B1(n158), .B2(r10[24]), .ZN(
        n766) );
  AOI22D1BWP12T U1511 ( .A1(r7[24]), .A2(n1990), .B1(n1989), .B2(r2[24]), .ZN(
        n765) );
  AOI22D1BWP12T U1512 ( .A1(r1[25]), .A2(n164), .B1(n1993), .B2(r12[25]), .ZN(
        n772) );
  AOI22D1BWP12T U1513 ( .A1(r3[25]), .A2(n1994), .B1(n168), .B2(lr[25]), .ZN(
        n771) );
  AOI22D1BWP12T U1514 ( .A1(r8[25]), .A2(n171), .B1(n1995), .B2(n[2016]), .ZN(
        n770) );
  AOI22D1BWP12T U1515 ( .A1(pc_out[25]), .A2(n174), .B1(n1996), .B2(r6[25]), 
        .ZN(n769) );
  AN4XD1BWP12T U1516 ( .A1(n772), .A2(n771), .A3(n770), .A4(n769), .Z(n779) );
  AOI22D1BWP12T U1517 ( .A1(tmp1[25]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[25]), .ZN(n775) );
  AOI22D1BWP12T U1518 ( .A1(r9[25]), .A2(n152), .B1(n2002), .B2(r4[25]), .ZN(
        n774) );
  AOI22D1BWP12T U1519 ( .A1(r11[25]), .A2(n1571), .B1(n1954), .B2(r0[25]), 
        .ZN(n773) );
  AN3XD1BWP12T U1520 ( .A1(n775), .A2(n774), .A3(n773), .Z(n778) );
  AOI22D1BWP12T U1521 ( .A1(r5[25]), .A2(n1988), .B1(n158), .B2(r10[25]), .ZN(
        n777) );
  AOI22D1BWP12T U1522 ( .A1(r7[25]), .A2(n1990), .B1(n1989), .B2(r2[25]), .ZN(
        n776) );
  AOI22D1BWP12T U1523 ( .A1(r1[22]), .A2(n164), .B1(n1993), .B2(r12[22]), .ZN(
        n783) );
  AOI22D1BWP12T U1524 ( .A1(r3[22]), .A2(n1994), .B1(n168), .B2(lr[22]), .ZN(
        n782) );
  AOI22D1BWP12T U1525 ( .A1(r8[22]), .A2(n171), .B1(n1995), .B2(n[2019]), .ZN(
        n781) );
  AOI22D1BWP12T U1526 ( .A1(pc_out[22]), .A2(n174), .B1(n1996), .B2(r6[22]), 
        .ZN(n780) );
  AOI22D1BWP12T U1527 ( .A1(tmp1[22]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[22]), .ZN(n786) );
  AOI22D1BWP12T U1528 ( .A1(r9[22]), .A2(n152), .B1(n2002), .B2(r4[22]), .ZN(
        n785) );
  AOI22D1BWP12T U1529 ( .A1(r11[22]), .A2(n1955), .B1(n1954), .B2(r0[22]), 
        .ZN(n784) );
  AOI22D1BWP12T U1530 ( .A1(r1[23]), .A2(n164), .B1(n1993), .B2(r12[23]), .ZN(
        n790) );
  AOI22D1BWP12T U1531 ( .A1(r3[23]), .A2(n1994), .B1(n168), .B2(lr[23]), .ZN(
        n789) );
  AOI22D1BWP12T U1532 ( .A1(r8[23]), .A2(n171), .B1(n1995), .B2(n[2018]), .ZN(
        n788) );
  AOI22D1BWP12T U1533 ( .A1(pc_out[23]), .A2(n174), .B1(n1996), .B2(r6[23]), 
        .ZN(n787) );
  AOI22D1BWP12T U1534 ( .A1(tmp1[23]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[23]), .ZN(n792) );
  AOI22D1BWP12T U1535 ( .A1(r11[23]), .A2(n1955), .B1(n1954), .B2(r0[23]), 
        .ZN(n791) );
  AOI22D1BWP12T U1536 ( .A1(r1[26]), .A2(n164), .B1(n1993), .B2(r12[26]), .ZN(
        n796) );
  AOI22D1BWP12T U1537 ( .A1(r8[26]), .A2(n171), .B1(n1995), .B2(n[2015]), .ZN(
        n794) );
  AN4XD1BWP12T U1538 ( .A1(n796), .A2(n795), .A3(n794), .A4(n793), .Z(n803) );
  AOI22D1BWP12T U1539 ( .A1(tmp1[26]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[26]), .ZN(n799) );
  AOI22D1BWP12T U1540 ( .A1(r9[26]), .A2(n152), .B1(n2002), .B2(r4[26]), .ZN(
        n798) );
  AOI22D1BWP12T U1541 ( .A1(r11[26]), .A2(n1955), .B1(n1954), .B2(r0[26]), 
        .ZN(n797) );
  AOI22D1BWP12T U1542 ( .A1(r5[26]), .A2(n1988), .B1(n158), .B2(r10[26]), .ZN(
        n801) );
  AOI22D1BWP12T U1543 ( .A1(r7[26]), .A2(n1990), .B1(n1989), .B2(r2[26]), .ZN(
        n800) );
  ND4D1BWP12T U1544 ( .A1(n803), .A2(n802), .A3(n801), .A4(n800), .ZN(
        regB_out[26]) );
  OR2XD1BWP12T U1545 ( .A1(readC_sel[0]), .A2(readC_sel[1]), .Z(n818) );
  ND3D1BWP12T U1546 ( .A1(readC_sel[2]), .A2(readC_sel[3]), .A3(n1208), .ZN(
        n815) );
  NR2D1BWP12T U1547 ( .A1(n818), .A2(n815), .ZN(n1199) );
  IND2D1BWP12T U1548 ( .A1(readC_sel[1]), .B1(readC_sel[0]), .ZN(n809) );
  INVD1BWP12T U1549 ( .I(readC_sel[2]), .ZN(n806) );
  ND3D1BWP12T U1550 ( .A1(readC_sel[3]), .A2(n1208), .A3(n806), .ZN(n817) );
  OR2XD1BWP12T U1551 ( .A1(n809), .A2(n817), .Z(n1052) );
  INVD1BWP12T U1552 ( .I(n1052), .ZN(n1194) );
  AOI22D0BWP12T U1553 ( .A1(r12[25]), .A2(n1199), .B1(n1194), .B2(r9[25]), 
        .ZN(n826) );
  IND2D1BWP12T U1554 ( .A1(readC_sel[0]), .B1(readC_sel[1]), .ZN(n807) );
  NR2D1BWP12T U1555 ( .A1(n807), .A2(n815), .ZN(n1197) );
  NR2D1BWP12T U1556 ( .A1(n809), .A2(n815), .ZN(n1196) );
  AOI22D0BWP12T U1557 ( .A1(lr[25]), .A2(n1197), .B1(n1196), .B2(n[2016]), 
        .ZN(n825) );
  OR2XD1BWP12T U1558 ( .A1(n807), .A2(n817), .Z(n1101) );
  INVD1BWP12T U1559 ( .I(n1101), .ZN(n1201) );
  ND2D1BWP12T U1560 ( .A1(readC_sel[1]), .A2(readC_sel[0]), .ZN(n816) );
  OR2XD1BWP12T U1561 ( .A1(n816), .A2(n817), .Z(n1112) );
  INVD1BWP12T U1562 ( .I(n1112), .ZN(n1200) );
  AOI22D0BWP12T U1563 ( .A1(r10[25]), .A2(n1201), .B1(n1200), .B2(r11[25]), 
        .ZN(n824) );
  CKND0BWP12T U1564 ( .I(readC_sel[3]), .ZN(n805) );
  TPND2D0BWP12T U1565 ( .A1(readC_sel[2]), .A2(n805), .ZN(n808) );
  OR2XD1BWP12T U1566 ( .A1(n808), .A2(n816), .Z(n1137) );
  INVD1BWP12T U1567 ( .I(n1137), .ZN(n1183) );
  OR2XD1BWP12T U1568 ( .A1(n808), .A2(n818), .Z(n1136) );
  INVD1BWP12T U1569 ( .I(n1136), .ZN(n1182) );
  AOI22D0BWP12T U1570 ( .A1(r7[25]), .A2(n1183), .B1(n1182), .B2(r4[25]), .ZN(
        n814) );
  CKND2D1BWP12T U1571 ( .A1(n806), .A2(n805), .ZN(n810) );
  OR2XD1BWP12T U1572 ( .A1(n807), .A2(n810), .Z(n1141) );
  INVD1BWP12T U1573 ( .I(n1141), .ZN(n1185) );
  OR2XD1BWP12T U1574 ( .A1(n808), .A2(n807), .Z(n1140) );
  INVD1BWP12T U1575 ( .I(n1140), .ZN(n1184) );
  AOI22D0BWP12T U1576 ( .A1(r2[25]), .A2(n1185), .B1(n1184), .B2(r6[25]), .ZN(
        n813) );
  OR2XD1BWP12T U1577 ( .A1(n809), .A2(n808), .Z(n1139) );
  INVD1BWP12T U1578 ( .I(n1139), .ZN(n1187) );
  OR2XD1BWP12T U1579 ( .A1(n809), .A2(n810), .Z(n1138) );
  INVD1BWP12T U1580 ( .I(n1138), .ZN(n1186) );
  AOI22D0BWP12T U1581 ( .A1(r5[25]), .A2(n1187), .B1(n1186), .B2(r1[25]), .ZN(
        n812) );
  OR2XD1BWP12T U1582 ( .A1(n810), .A2(n818), .Z(n1143) );
  INVD1BWP12T U1583 ( .I(n1143), .ZN(n1189) );
  OR2XD1BWP12T U1584 ( .A1(n810), .A2(n816), .Z(n1142) );
  INVD1BWP12T U1585 ( .I(n1142), .ZN(n1188) );
  AOI22D0BWP12T U1586 ( .A1(r0[25]), .A2(n1189), .B1(n1188), .B2(r3[25]), .ZN(
        n811) );
  ND4D1BWP12T U1587 ( .A1(n814), .A2(n813), .A3(n812), .A4(n811), .ZN(n822) );
  CKND0BWP12T U1588 ( .I(pc_out[25]), .ZN(n820) );
  OR2XD1BWP12T U1589 ( .A1(n816), .A2(n815), .Z(n883) );
  NR2D1BWP12T U1590 ( .A1(n818), .A2(n817), .ZN(n1195) );
  INVD1BWP12T U1591 ( .I(n1195), .ZN(n1116) );
  CKND0BWP12T U1592 ( .I(r8[25]), .ZN(n819) );
  OAI22D0BWP12T U1593 ( .A1(n820), .A2(n883), .B1(n1116), .B2(n819), .ZN(n821)
         );
  AOI21D0BWP12T U1594 ( .A1(n822), .A2(n1208), .B(n821), .ZN(n823) );
  ND4D1BWP12T U1595 ( .A1(n826), .A2(n825), .A3(n824), .A4(n823), .ZN(
        regC_out[25]) );
  OAI22D0BWP12T U1596 ( .A1(n1960), .A2(n1137), .B1(n1136), .B2(n827), .ZN(
        n832) );
  OAI22D0BWP12T U1597 ( .A1(n1950), .A2(n1139), .B1(n1138), .B2(n1969), .ZN(
        n831) );
  OAI22D0BWP12T U1598 ( .A1(n1141), .A2(n1958), .B1(n1140), .B2(n1978), .ZN(
        n830) );
  OAI22D0BWP12T U1599 ( .A1(n828), .A2(n1143), .B1(n1142), .B2(n1973), .ZN(
        n829) );
  NR4D0BWP12T U1600 ( .A1(n832), .A2(n831), .A3(n830), .A4(n829), .ZN(n833) );
  OAI22D0BWP12T U1601 ( .A1(n833), .A2(readC_sel[4]), .B1(n883), .B2(n1980), 
        .ZN(n834) );
  AOI21D0BWP12T U1602 ( .A1(lr[2]), .A2(n1197), .B(n834), .ZN(n838) );
  AOI22D0BWP12T U1603 ( .A1(r9[2]), .A2(n1194), .B1(n1200), .B2(r11[2]), .ZN(
        n837) );
  AOI22D0BWP12T U1604 ( .A1(r8[2]), .A2(n1195), .B1(n1201), .B2(r10[2]), .ZN(
        n836) );
  AOI22D0BWP12T U1605 ( .A1(r12[2]), .A2(n1199), .B1(n1196), .B2(n[2039]), 
        .ZN(n835) );
  ND4D1BWP12T U1606 ( .A1(n838), .A2(n837), .A3(n836), .A4(n835), .ZN(
        regC_out[2]) );
  OAI22D0BWP12T U1607 ( .A1(n1928), .A2(n1137), .B1(n1136), .B2(n839), .ZN(
        n844) );
  OAI22D0BWP12T U1608 ( .A1(n1923), .A2(n1139), .B1(n1138), .B2(n1934), .ZN(
        n843) );
  OAI22D0BWP12T U1609 ( .A1(n1141), .A2(n1927), .B1(n1140), .B2(n1939), .ZN(
        n842) );
  OAI22D0BWP12T U1610 ( .A1(n840), .A2(n1143), .B1(n1142), .B2(n1936), .ZN(
        n841) );
  NR4D0BWP12T U1611 ( .A1(n844), .A2(n843), .A3(n842), .A4(n841), .ZN(n845) );
  OAI22D0BWP12T U1612 ( .A1(n845), .A2(readC_sel[4]), .B1(n883), .B2(n1940), 
        .ZN(n846) );
  AOI21D0BWP12T U1613 ( .A1(lr[3]), .A2(n1197), .B(n846), .ZN(n850) );
  AOI22D0BWP12T U1614 ( .A1(r9[3]), .A2(n1194), .B1(n1200), .B2(r11[3]), .ZN(
        n849) );
  AOI22D0BWP12T U1615 ( .A1(r8[3]), .A2(n1195), .B1(n1201), .B2(r10[3]), .ZN(
        n848) );
  AOI22D0BWP12T U1616 ( .A1(r12[3]), .A2(n1199), .B1(n1196), .B2(n[2038]), 
        .ZN(n847) );
  ND4D1BWP12T U1617 ( .A1(n850), .A2(n849), .A3(n848), .A4(n847), .ZN(
        regC_out[3]) );
  AOI22D0BWP12T U1618 ( .A1(r8[4]), .A2(n1195), .B1(n1201), .B2(r10[4]), .ZN(
        n860) );
  AOI22D0BWP12T U1619 ( .A1(r12[4]), .A2(n1199), .B1(n1196), .B2(n[2037]), 
        .ZN(n859) );
  AOI22D0BWP12T U1620 ( .A1(r9[4]), .A2(n1194), .B1(n1200), .B2(r11[4]), .ZN(
        n858) );
  AOI22D0BWP12T U1621 ( .A1(r7[4]), .A2(n1183), .B1(n1182), .B2(r4[4]), .ZN(
        n854) );
  AOI22D0BWP12T U1622 ( .A1(r2[4]), .A2(n1185), .B1(n1184), .B2(r6[4]), .ZN(
        n853) );
  AOI22D0BWP12T U1623 ( .A1(r5[4]), .A2(n1187), .B1(n1186), .B2(r1[4]), .ZN(
        n852) );
  AOI22D0BWP12T U1624 ( .A1(r0[4]), .A2(n1189), .B1(n1188), .B2(r3[4]), .ZN(
        n851) );
  ND4D1BWP12T U1625 ( .A1(n854), .A2(n853), .A3(n852), .A4(n851), .ZN(n856) );
  INVD1BWP12T U1626 ( .I(n1197), .ZN(n1160) );
  OAI22D0BWP12T U1627 ( .A1(n1885), .A2(n883), .B1(n1160), .B2(n1889), .ZN(
        n855) );
  AOI21D0BWP12T U1628 ( .A1(n856), .A2(n1208), .B(n855), .ZN(n857) );
  ND4D1BWP12T U1629 ( .A1(n860), .A2(n859), .A3(n858), .A4(n857), .ZN(
        regC_out[4]) );
  CKND0BWP12T U1630 ( .I(pc_out[30]), .ZN(n1356) );
  INVD1BWP12T U1631 ( .I(n1199), .ZN(n1172) );
  AOI22D0BWP12T U1632 ( .A1(r8[12]), .A2(n1195), .B1(n1194), .B2(r9[12]), .ZN(
        n870) );
  AOI22D0BWP12T U1633 ( .A1(lr[12]), .A2(n1197), .B1(n1196), .B2(n[2029]), 
        .ZN(n869) );
  AOI22D0BWP12T U1634 ( .A1(r10[12]), .A2(n1201), .B1(n1200), .B2(r11[12]), 
        .ZN(n868) );
  AOI22D0BWP12T U1635 ( .A1(r7[12]), .A2(n1183), .B1(n1182), .B2(r4[12]), .ZN(
        n864) );
  AOI22D0BWP12T U1636 ( .A1(r2[12]), .A2(n1185), .B1(n1184), .B2(r6[12]), .ZN(
        n863) );
  AOI22D0BWP12T U1637 ( .A1(r5[12]), .A2(n1187), .B1(n1186), .B2(r1[12]), .ZN(
        n862) );
  AOI22D0BWP12T U1638 ( .A1(r0[12]), .A2(n1189), .B1(n1188), .B2(r3[12]), .ZN(
        n861) );
  ND4D1BWP12T U1639 ( .A1(n864), .A2(n863), .A3(n862), .A4(n861), .ZN(n866) );
  INVD1BWP12T U1640 ( .I(pc_out[12]), .ZN(n1648) );
  OAI22D0BWP12T U1641 ( .A1(n1648), .A2(n883), .B1(n1172), .B2(n1641), .ZN(
        n865) );
  AOI21D0BWP12T U1642 ( .A1(n866), .A2(n1208), .B(n865), .ZN(n867) );
  ND4D1BWP12T U1643 ( .A1(n870), .A2(n869), .A3(n868), .A4(n867), .ZN(
        regC_out[12]) );
  AOI22D0BWP12T U1644 ( .A1(r8[26]), .A2(n1195), .B1(n1194), .B2(r9[26]), .ZN(
        n882) );
  AOI22D0BWP12T U1645 ( .A1(lr[26]), .A2(n1197), .B1(n1199), .B2(r12[26]), 
        .ZN(n881) );
  AOI22D0BWP12T U1646 ( .A1(r10[26]), .A2(n1201), .B1(n1200), .B2(r11[26]), 
        .ZN(n880) );
  AOI22D0BWP12T U1647 ( .A1(r7[26]), .A2(n1183), .B1(n1182), .B2(r4[26]), .ZN(
        n874) );
  AOI22D0BWP12T U1648 ( .A1(r2[26]), .A2(n1185), .B1(n1184), .B2(r6[26]), .ZN(
        n873) );
  AOI22D0BWP12T U1649 ( .A1(r5[26]), .A2(n1187), .B1(n1186), .B2(r1[26]), .ZN(
        n872) );
  AOI22D0BWP12T U1650 ( .A1(r0[26]), .A2(n1189), .B1(n1188), .B2(r3[26]), .ZN(
        n871) );
  ND4D1BWP12T U1651 ( .A1(n874), .A2(n873), .A3(n872), .A4(n871), .ZN(n878) );
  CKND0BWP12T U1652 ( .I(pc_out[26]), .ZN(n876) );
  CKND0BWP12T U1653 ( .I(n[2015]), .ZN(n875) );
  INVD1BWP12T U1654 ( .I(n1196), .ZN(n1148) );
  OAI22D0BWP12T U1655 ( .A1(n876), .A2(n883), .B1(n875), .B2(n1148), .ZN(n877)
         );
  AOI21D0BWP12T U1656 ( .A1(n878), .A2(n1208), .B(n877), .ZN(n879) );
  ND4D1BWP12T U1657 ( .A1(n882), .A2(n881), .A3(n880), .A4(n879), .ZN(
        regC_out[26]) );
  INVD1BWP12T U1658 ( .I(n883), .ZN(n1198) );
  AOI22D0BWP12T U1659 ( .A1(pc_out[24]), .A2(n1198), .B1(n1195), .B2(r8[24]), 
        .ZN(n897) );
  AOI22D0BWP12T U1660 ( .A1(r9[24]), .A2(n1194), .B1(n1200), .B2(r11[24]), 
        .ZN(n896) );
  AOI22D0BWP12T U1661 ( .A1(r7[24]), .A2(n1183), .B1(n1182), .B2(r4[24]), .ZN(
        n887) );
  AOI22D0BWP12T U1662 ( .A1(r2[24]), .A2(n1185), .B1(n1184), .B2(r6[24]), .ZN(
        n886) );
  AOI22D0BWP12T U1663 ( .A1(r5[24]), .A2(n1187), .B1(n1186), .B2(r1[24]), .ZN(
        n885) );
  AOI22D0BWP12T U1664 ( .A1(r0[24]), .A2(n1189), .B1(n1188), .B2(r3[24]), .ZN(
        n884) );
  ND4D1BWP12T U1665 ( .A1(n887), .A2(n886), .A3(n885), .A4(n884), .ZN(n894) );
  CKND0BWP12T U1666 ( .I(r12[24]), .ZN(n889) );
  CKND0BWP12T U1667 ( .I(r10[24]), .ZN(n888) );
  OAI22D0BWP12T U1668 ( .A1(n1172), .A2(n889), .B1(n888), .B2(n1101), .ZN(n893) );
  CKND0BWP12T U1669 ( .I(n[2017]), .ZN(n891) );
  CKND0BWP12T U1670 ( .I(lr[24]), .ZN(n890) );
  OAI22D0BWP12T U1671 ( .A1(n891), .A2(n1148), .B1(n1160), .B2(n890), .ZN(n892) );
  AOI211D0BWP12T U1672 ( .A1(n894), .A2(n1208), .B(n893), .C(n892), .ZN(n895)
         );
  ND3D1BWP12T U1673 ( .A1(n897), .A2(n896), .A3(n895), .ZN(regC_out[24]) );
  AOI22D0BWP12T U1674 ( .A1(pc_out[27]), .A2(n1198), .B1(n1195), .B2(r8[27]), 
        .ZN(n909) );
  AOI22D0BWP12T U1675 ( .A1(lr[27]), .A2(n1197), .B1(n1199), .B2(r12[27]), 
        .ZN(n908) );
  AOI22D0BWP12T U1676 ( .A1(r9[27]), .A2(n1194), .B1(n1201), .B2(r10[27]), 
        .ZN(n907) );
  AOI22D0BWP12T U1677 ( .A1(r7[27]), .A2(n1183), .B1(n1182), .B2(r4[27]), .ZN(
        n901) );
  AOI22D0BWP12T U1678 ( .A1(r2[27]), .A2(n1185), .B1(n1184), .B2(r6[27]), .ZN(
        n900) );
  AOI22D0BWP12T U1679 ( .A1(r5[27]), .A2(n1187), .B1(n1186), .B2(r1[27]), .ZN(
        n899) );
  AOI22D0BWP12T U1680 ( .A1(r0[27]), .A2(n1189), .B1(n1188), .B2(r3[27]), .ZN(
        n898) );
  ND4D1BWP12T U1681 ( .A1(n901), .A2(n900), .A3(n899), .A4(n898), .ZN(n905) );
  CKND0BWP12T U1682 ( .I(n[2014]), .ZN(n903) );
  CKND0BWP12T U1683 ( .I(r11[27]), .ZN(n902) );
  OAI22D0BWP12T U1684 ( .A1(n903), .A2(n1148), .B1(n1112), .B2(n902), .ZN(n904) );
  AOI21D0BWP12T U1685 ( .A1(n905), .A2(n1208), .B(n904), .ZN(n906) );
  ND4D1BWP12T U1686 ( .A1(n909), .A2(n908), .A3(n907), .A4(n906), .ZN(
        regC_out[27]) );
  AOI22D0BWP12T U1687 ( .A1(pc_out[29]), .A2(n1198), .B1(n1195), .B2(r8[29]), 
        .ZN(n921) );
  AOI22D0BWP12T U1688 ( .A1(lr[29]), .A2(n1197), .B1(n1199), .B2(r12[29]), 
        .ZN(n920) );
  AOI22D0BWP12T U1689 ( .A1(r10[29]), .A2(n1201), .B1(n1200), .B2(r11[29]), 
        .ZN(n919) );
  AOI22D0BWP12T U1690 ( .A1(r7[29]), .A2(n1183), .B1(n1182), .B2(r4[29]), .ZN(
        n913) );
  AOI22D0BWP12T U1691 ( .A1(r2[29]), .A2(n1185), .B1(n1184), .B2(r6[29]), .ZN(
        n912) );
  AOI22D0BWP12T U1692 ( .A1(r5[29]), .A2(n1187), .B1(n1186), .B2(r1[29]), .ZN(
        n911) );
  AOI22D0BWP12T U1693 ( .A1(r0[29]), .A2(n1189), .B1(n1188), .B2(r3[29]), .ZN(
        n910) );
  ND4D1BWP12T U1694 ( .A1(n913), .A2(n912), .A3(n911), .A4(n910), .ZN(n917) );
  CKND0BWP12T U1695 ( .I(n[2012]), .ZN(n915) );
  CKND0BWP12T U1696 ( .I(r9[29]), .ZN(n914) );
  OAI22D0BWP12T U1697 ( .A1(n915), .A2(n1148), .B1(n1052), .B2(n914), .ZN(n916) );
  AOI21D0BWP12T U1698 ( .A1(n917), .A2(n1208), .B(n916), .ZN(n918) );
  ND4D1BWP12T U1699 ( .A1(n921), .A2(n920), .A3(n919), .A4(n918), .ZN(
        regC_out[29]) );
  AOI22D0BWP12T U1700 ( .A1(pc_out[15]), .A2(n1198), .B1(n1201), .B2(r10[15]), 
        .ZN(n932) );
  AOI22D0BWP12T U1701 ( .A1(n[2026]), .A2(n1196), .B1(n1199), .B2(r12[15]), 
        .ZN(n931) );
  AOI22D0BWP12T U1702 ( .A1(r9[15]), .A2(n1194), .B1(n1200), .B2(r11[15]), 
        .ZN(n930) );
  AOI22D0BWP12T U1703 ( .A1(r7[15]), .A2(n1183), .B1(n1182), .B2(r4[15]), .ZN(
        n925) );
  AOI22D0BWP12T U1704 ( .A1(r2[15]), .A2(n1185), .B1(n1184), .B2(r6[15]), .ZN(
        n924) );
  AOI22D0BWP12T U1705 ( .A1(r5[15]), .A2(n1187), .B1(n1186), .B2(r1[15]), .ZN(
        n923) );
  AOI22D0BWP12T U1706 ( .A1(r0[15]), .A2(n1189), .B1(n1188), .B2(r3[15]), .ZN(
        n922) );
  ND4D1BWP12T U1707 ( .A1(n925), .A2(n924), .A3(n923), .A4(n922), .ZN(n928) );
  INVD1BWP12T U1708 ( .I(lr[15]), .ZN(n1557) );
  CKND0BWP12T U1709 ( .I(r8[15]), .ZN(n926) );
  OAI22D0BWP12T U1710 ( .A1(n1160), .A2(n1557), .B1(n926), .B2(n1116), .ZN(
        n927) );
  AOI21D0BWP12T U1711 ( .A1(n928), .A2(n1208), .B(n927), .ZN(n929) );
  ND4D1BWP12T U1712 ( .A1(n932), .A2(n931), .A3(n930), .A4(n929), .ZN(
        regC_out[15]) );
  AOI22D0BWP12T U1713 ( .A1(pc_out[8]), .A2(n1198), .B1(n1194), .B2(r9[8]), 
        .ZN(n943) );
  AOI22D0BWP12T U1714 ( .A1(lr[8]), .A2(n1197), .B1(n1196), .B2(n[2033]), .ZN(
        n942) );
  AOI22D0BWP12T U1715 ( .A1(r10[8]), .A2(n1201), .B1(n1200), .B2(r11[8]), .ZN(
        n941) );
  AOI22D0BWP12T U1716 ( .A1(r7[8]), .A2(n1183), .B1(n1182), .B2(r4[8]), .ZN(
        n936) );
  AOI22D0BWP12T U1717 ( .A1(r2[8]), .A2(n1185), .B1(n1184), .B2(r6[8]), .ZN(
        n935) );
  AOI22D0BWP12T U1718 ( .A1(r5[8]), .A2(n1187), .B1(n1186), .B2(r1[8]), .ZN(
        n934) );
  AOI22D0BWP12T U1719 ( .A1(r0[8]), .A2(n1189), .B1(n1188), .B2(r3[8]), .ZN(
        n933) );
  ND4D1BWP12T U1720 ( .A1(n936), .A2(n935), .A3(n934), .A4(n933), .ZN(n939) );
  OAI22D0BWP12T U1721 ( .A1(n1172), .A2(n937), .B1(n1695), .B2(n1116), .ZN(
        n938) );
  AOI21D0BWP12T U1722 ( .A1(n939), .A2(n1208), .B(n938), .ZN(n940) );
  ND4D1BWP12T U1723 ( .A1(n943), .A2(n942), .A3(n941), .A4(n940), .ZN(
        regC_out[8]) );
  AOI22D0BWP12T U1724 ( .A1(n[2040]), .A2(n1196), .B1(n1201), .B2(r10[1]), 
        .ZN(n954) );
  AOI22D0BWP12T U1725 ( .A1(r9[1]), .A2(n1194), .B1(n1200), .B2(r11[1]), .ZN(
        n953) );
  OAI22D0BWP12T U1726 ( .A1(n1160), .A2(n1859), .B1(n1862), .B2(n1116), .ZN(
        n945) );
  NR2D0BWP12T U1727 ( .A1(n1857), .A2(n1172), .ZN(n944) );
  AOI211D0BWP12T U1728 ( .A1(pc_out[1]), .A2(n1198), .B(n945), .C(n944), .ZN(
        n952) );
  AOI22D0BWP12T U1729 ( .A1(r7[1]), .A2(n1183), .B1(n1182), .B2(r4[1]), .ZN(
        n949) );
  AOI22D0BWP12T U1730 ( .A1(r2[1]), .A2(n1185), .B1(n1184), .B2(r6[1]), .ZN(
        n948) );
  AOI22D0BWP12T U1731 ( .A1(r5[1]), .A2(n1187), .B1(n1186), .B2(r1[1]), .ZN(
        n947) );
  AOI22D0BWP12T U1732 ( .A1(r0[1]), .A2(n1189), .B1(n1188), .B2(r3[1]), .ZN(
        n946) );
  ND4D1BWP12T U1733 ( .A1(n949), .A2(n948), .A3(n947), .A4(n946), .ZN(n950) );
  CKND2D0BWP12T U1734 ( .A1(n950), .A2(n1208), .ZN(n951) );
  ND4D1BWP12T U1735 ( .A1(n954), .A2(n953), .A3(n952), .A4(n951), .ZN(
        regC_out[1]) );
  AOI22D0BWP12T U1736 ( .A1(pc_out[18]), .A2(n1198), .B1(n1194), .B2(r9[18]), 
        .ZN(n966) );
  AOI22D0BWP12T U1737 ( .A1(lr[18]), .A2(n1197), .B1(n1196), .B2(n[2023]), 
        .ZN(n965) );
  AOI22D0BWP12T U1738 ( .A1(r10[18]), .A2(n1201), .B1(n1200), .B2(r11[18]), 
        .ZN(n964) );
  AOI22D0BWP12T U1739 ( .A1(r7[18]), .A2(n1183), .B1(n1182), .B2(r4[18]), .ZN(
        n958) );
  AOI22D0BWP12T U1740 ( .A1(r2[18]), .A2(n1185), .B1(n1184), .B2(r6[18]), .ZN(
        n957) );
  AOI22D0BWP12T U1741 ( .A1(r5[18]), .A2(n1187), .B1(n1186), .B2(r1[18]), .ZN(
        n956) );
  AOI22D0BWP12T U1742 ( .A1(r0[18]), .A2(n1189), .B1(n1188), .B2(r3[18]), .ZN(
        n955) );
  ND4D1BWP12T U1743 ( .A1(n958), .A2(n957), .A3(n956), .A4(n955), .ZN(n962) );
  CKND0BWP12T U1744 ( .I(r12[18]), .ZN(n960) );
  CKND0BWP12T U1745 ( .I(r8[18]), .ZN(n959) );
  TPOAI22D0BWP12T U1746 ( .A1(n1172), .A2(n960), .B1(n959), .B2(n1116), .ZN(
        n961) );
  AOI21D0BWP12T U1747 ( .A1(n962), .A2(n1208), .B(n961), .ZN(n963) );
  ND4D1BWP12T U1748 ( .A1(n966), .A2(n965), .A3(n964), .A4(n963), .ZN(
        regC_out[18]) );
  AOI22D0BWP12T U1749 ( .A1(pc_out[0]), .A2(n1198), .B1(n1195), .B2(r8[0]), 
        .ZN(n978) );
  AOI22D0BWP12T U1750 ( .A1(n[2041]), .A2(n1196), .B1(n1199), .B2(r12[0]), 
        .ZN(n977) );
  AOI22D0BWP12T U1751 ( .A1(r9[0]), .A2(n1194), .B1(n1200), .B2(r11[0]), .ZN(
        n976) );
  AOI22D0BWP12T U1752 ( .A1(r7[0]), .A2(n1183), .B1(n1182), .B2(r4[0]), .ZN(
        n970) );
  AOI22D0BWP12T U1753 ( .A1(r2[0]), .A2(n1185), .B1(n1184), .B2(r6[0]), .ZN(
        n969) );
  AOI22D0BWP12T U1754 ( .A1(r5[0]), .A2(n1187), .B1(n1186), .B2(r1[0]), .ZN(
        n968) );
  AOI22D0BWP12T U1755 ( .A1(r0[0]), .A2(n1189), .B1(n1188), .B2(r3[0]), .ZN(
        n967) );
  ND4D1BWP12T U1756 ( .A1(n970), .A2(n969), .A3(n968), .A4(n967), .ZN(n974) );
  OAI22D0BWP12T U1757 ( .A1(n1160), .A2(n972), .B1(n971), .B2(n1101), .ZN(n973) );
  AOI21D0BWP12T U1758 ( .A1(n974), .A2(n1208), .B(n973), .ZN(n975) );
  ND4D1BWP12T U1759 ( .A1(n978), .A2(n977), .A3(n976), .A4(n975), .ZN(
        regC_out[0]) );
  AOI22D0BWP12T U1760 ( .A1(pc_out[5]), .A2(n1198), .B1(n1195), .B2(r8[5]), 
        .ZN(n989) );
  AOI22D0BWP12T U1761 ( .A1(r12[5]), .A2(n1199), .B1(n1196), .B2(n[2036]), 
        .ZN(n988) );
  AOI22D0BWP12T U1762 ( .A1(r10[5]), .A2(n1201), .B1(n1200), .B2(r11[5]), .ZN(
        n987) );
  AOI22D0BWP12T U1763 ( .A1(r7[5]), .A2(n1183), .B1(n1182), .B2(r4[5]), .ZN(
        n982) );
  AOI22D0BWP12T U1764 ( .A1(r2[5]), .A2(n1185), .B1(n1184), .B2(r6[5]), .ZN(
        n981) );
  AOI22D0BWP12T U1765 ( .A1(r5[5]), .A2(n1187), .B1(n1186), .B2(r1[5]), .ZN(
        n980) );
  AOI22D0BWP12T U1766 ( .A1(r0[5]), .A2(n1189), .B1(n1188), .B2(r3[5]), .ZN(
        n979) );
  ND4D1BWP12T U1767 ( .A1(n982), .A2(n981), .A3(n980), .A4(n979), .ZN(n985) );
  OAI22D0BWP12T U1768 ( .A1(n1160), .A2(n1834), .B1(n983), .B2(n1052), .ZN(
        n984) );
  AOI21D0BWP12T U1769 ( .A1(n985), .A2(n1208), .B(n984), .ZN(n986) );
  ND4D1BWP12T U1770 ( .A1(n989), .A2(n988), .A3(n987), .A4(n986), .ZN(
        regC_out[5]) );
  AOI22D0BWP12T U1771 ( .A1(pc_out[20]), .A2(n1198), .B1(n1195), .B2(r8[20]), 
        .ZN(n1001) );
  AOI22D0BWP12T U1772 ( .A1(lr[20]), .A2(n1197), .B1(n1199), .B2(r12[20]), 
        .ZN(n1000) );
  AOI22D0BWP12T U1773 ( .A1(r9[20]), .A2(n1194), .B1(n1201), .B2(r10[20]), 
        .ZN(n999) );
  AOI22D0BWP12T U1774 ( .A1(r7[20]), .A2(n1183), .B1(n1182), .B2(r4[20]), .ZN(
        n993) );
  AOI22D0BWP12T U1775 ( .A1(r2[20]), .A2(n1185), .B1(n1184), .B2(r6[20]), .ZN(
        n992) );
  AOI22D0BWP12T U1776 ( .A1(r5[20]), .A2(n1187), .B1(n1186), .B2(r1[20]), .ZN(
        n991) );
  AOI22D0BWP12T U1777 ( .A1(r0[20]), .A2(n1189), .B1(n1188), .B2(r3[20]), .ZN(
        n990) );
  ND4D1BWP12T U1778 ( .A1(n993), .A2(n992), .A3(n991), .A4(n990), .ZN(n997) );
  CKND0BWP12T U1779 ( .I(n[2021]), .ZN(n995) );
  OAI22D0BWP12T U1780 ( .A1(n995), .A2(n1148), .B1(n1112), .B2(n994), .ZN(n996) );
  AOI21D0BWP12T U1781 ( .A1(n997), .A2(n1208), .B(n996), .ZN(n998) );
  ND4D1BWP12T U1782 ( .A1(n1001), .A2(n1000), .A3(n999), .A4(n998), .ZN(
        regC_out[20]) );
  AOI22D0BWP12T U1783 ( .A1(pc_out[19]), .A2(n1198), .B1(n1195), .B2(r8[19]), 
        .ZN(n1012) );
  AOI22D0BWP12T U1784 ( .A1(n[2022]), .A2(n1196), .B1(n1199), .B2(r12[19]), 
        .ZN(n1011) );
  AOI22D0BWP12T U1785 ( .A1(r10[19]), .A2(n1201), .B1(n1200), .B2(r11[19]), 
        .ZN(n1010) );
  AOI22D0BWP12T U1786 ( .A1(r7[19]), .A2(n1183), .B1(n1182), .B2(r4[19]), .ZN(
        n1005) );
  AOI22D0BWP12T U1787 ( .A1(r2[19]), .A2(n1185), .B1(n1184), .B2(r6[19]), .ZN(
        n1004) );
  AOI22D0BWP12T U1788 ( .A1(r5[19]), .A2(n1187), .B1(n1186), .B2(r1[19]), .ZN(
        n1003) );
  AOI22D0BWP12T U1789 ( .A1(r0[19]), .A2(n1189), .B1(n1188), .B2(r3[19]), .ZN(
        n1002) );
  ND4D1BWP12T U1790 ( .A1(n1005), .A2(n1004), .A3(n1003), .A4(n1002), .ZN(
        n1008) );
  INVD1BWP12T U1791 ( .I(lr[19]), .ZN(n1462) );
  CKND0BWP12T U1792 ( .I(r9[19]), .ZN(n1006) );
  OAI22D0BWP12T U1793 ( .A1(n1160), .A2(n1462), .B1(n1006), .B2(n1052), .ZN(
        n1007) );
  AOI21D0BWP12T U1794 ( .A1(n1008), .A2(n1208), .B(n1007), .ZN(n1009) );
  ND4D1BWP12T U1795 ( .A1(n1012), .A2(n1011), .A3(n1010), .A4(n1009), .ZN(
        regC_out[19]) );
  CKND0BWP12T U1796 ( .I(r8[23]), .ZN(n1018) );
  AOI22D0BWP12T U1797 ( .A1(r7[23]), .A2(n1183), .B1(n1182), .B2(r4[23]), .ZN(
        n1016) );
  AOI22D0BWP12T U1798 ( .A1(r2[23]), .A2(n1185), .B1(n1184), .B2(r6[23]), .ZN(
        n1015) );
  AOI22D0BWP12T U1799 ( .A1(r5[23]), .A2(n1187), .B1(n1186), .B2(r1[23]), .ZN(
        n1014) );
  AOI22D0BWP12T U1800 ( .A1(r0[23]), .A2(n1189), .B1(n1188), .B2(r3[23]), .ZN(
        n1013) );
  ND4D1BWP12T U1801 ( .A1(n1016), .A2(n1015), .A3(n1014), .A4(n1013), .ZN(
        n1017) );
  MOAI22D0BWP12T U1802 ( .A1(n1116), .A2(n1018), .B1(n1017), .B2(n1208), .ZN(
        n1019) );
  AOI21D0BWP12T U1803 ( .A1(lr[23]), .A2(n1197), .B(n1019), .ZN(n1023) );
  AOI22D0BWP12T U1804 ( .A1(r9[23]), .A2(n1194), .B1(n1200), .B2(r11[23]), 
        .ZN(n1022) );
  AOI22D0BWP12T U1805 ( .A1(pc_out[23]), .A2(n1198), .B1(n1201), .B2(r10[23]), 
        .ZN(n1021) );
  AOI22D0BWP12T U1806 ( .A1(n[2018]), .A2(n1196), .B1(n1199), .B2(r12[23]), 
        .ZN(n1020) );
  ND4D1BWP12T U1807 ( .A1(n1023), .A2(n1022), .A3(n1021), .A4(n1020), .ZN(
        regC_out[23]) );
  AOI22D0BWP12T U1808 ( .A1(r12[31]), .A2(n1199), .B1(n1198), .B2(pc_out[31]), 
        .ZN(n1035) );
  AOI22D0BWP12T U1809 ( .A1(lr[31]), .A2(n1197), .B1(n1196), .B2(n[2010]), 
        .ZN(n1034) );
  AOI22D0BWP12T U1810 ( .A1(r8[31]), .A2(n1195), .B1(n1200), .B2(r11[31]), 
        .ZN(n1033) );
  AOI22D0BWP12T U1811 ( .A1(r7[31]), .A2(n1183), .B1(n1182), .B2(r4[31]), .ZN(
        n1027) );
  AOI22D0BWP12T U1812 ( .A1(r2[31]), .A2(n1185), .B1(n1184), .B2(r6[31]), .ZN(
        n1026) );
  AOI22D0BWP12T U1813 ( .A1(r5[31]), .A2(n1187), .B1(n1186), .B2(r1[31]), .ZN(
        n1025) );
  AOI22D0BWP12T U1814 ( .A1(r0[31]), .A2(n1189), .B1(n1188), .B2(r3[31]), .ZN(
        n1024) );
  ND4D1BWP12T U1815 ( .A1(n1027), .A2(n1026), .A3(n1025), .A4(n1024), .ZN(
        n1031) );
  CKND0BWP12T U1816 ( .I(r9[31]), .ZN(n1029) );
  CKND0BWP12T U1817 ( .I(r10[31]), .ZN(n1028) );
  OAI22D0BWP12T U1818 ( .A1(n1052), .A2(n1029), .B1(n1028), .B2(n1101), .ZN(
        n1030) );
  AOI21D0BWP12T U1819 ( .A1(n1031), .A2(n1208), .B(n1030), .ZN(n1032) );
  ND4D1BWP12T U1820 ( .A1(n1035), .A2(n1034), .A3(n1033), .A4(n1032), .ZN(
        regC_out[31]) );
  AOI22D0BWP12T U1821 ( .A1(r8[28]), .A2(n1195), .B1(n1201), .B2(r10[28]), 
        .ZN(n1047) );
  AOI22D0BWP12T U1822 ( .A1(n[2013]), .A2(n1196), .B1(n1198), .B2(pc_out[28]), 
        .ZN(n1046) );
  AOI22D0BWP12T U1823 ( .A1(r9[28]), .A2(n1194), .B1(n1200), .B2(r11[28]), 
        .ZN(n1045) );
  AOI22D0BWP12T U1824 ( .A1(r7[28]), .A2(n1183), .B1(n1182), .B2(r4[28]), .ZN(
        n1039) );
  AOI22D0BWP12T U1825 ( .A1(r2[28]), .A2(n1185), .B1(n1184), .B2(r6[28]), .ZN(
        n1038) );
  AOI22D0BWP12T U1826 ( .A1(r5[28]), .A2(n1187), .B1(n1186), .B2(r1[28]), .ZN(
        n1037) );
  AOI22D0BWP12T U1827 ( .A1(r0[28]), .A2(n1189), .B1(n1188), .B2(r3[28]), .ZN(
        n1036) );
  ND4D1BWP12T U1828 ( .A1(n1039), .A2(n1038), .A3(n1037), .A4(n1036), .ZN(
        n1043) );
  CKND0BWP12T U1829 ( .I(lr[28]), .ZN(n1041) );
  CKND0BWP12T U1830 ( .I(r12[28]), .ZN(n1040) );
  TPOAI22D0BWP12T U1831 ( .A1(n1160), .A2(n1041), .B1(n1040), .B2(n1172), .ZN(
        n1042) );
  AOI21D0BWP12T U1832 ( .A1(n1043), .A2(n1208), .B(n1042), .ZN(n1044) );
  ND4D1BWP12T U1833 ( .A1(n1047), .A2(n1046), .A3(n1045), .A4(n1044), .ZN(
        regC_out[28]) );
  AOI22D0BWP12T U1834 ( .A1(r12[9]), .A2(n1199), .B1(n1198), .B2(pc_out[9]), 
        .ZN(n1060) );
  AOI22D0BWP12T U1835 ( .A1(lr[9]), .A2(n1197), .B1(n1196), .B2(n[2032]), .ZN(
        n1059) );
  AOI22D0BWP12T U1836 ( .A1(r10[9]), .A2(n1201), .B1(n1200), .B2(r11[9]), .ZN(
        n1058) );
  AOI22D0BWP12T U1837 ( .A1(r7[9]), .A2(n1183), .B1(n1182), .B2(r4[9]), .ZN(
        n1051) );
  AOI22D0BWP12T U1838 ( .A1(r2[9]), .A2(n1185), .B1(n1184), .B2(r6[9]), .ZN(
        n1050) );
  AOI22D0BWP12T U1839 ( .A1(r5[9]), .A2(n1187), .B1(n1186), .B2(r1[9]), .ZN(
        n1049) );
  AOI22D0BWP12T U1840 ( .A1(r0[9]), .A2(n1189), .B1(n1188), .B2(r3[9]), .ZN(
        n1048) );
  ND4D1BWP12T U1841 ( .A1(n1051), .A2(n1050), .A3(n1049), .A4(n1048), .ZN(
        n1056) );
  OAI22D0BWP12T U1842 ( .A1(n1116), .A2(n1054), .B1(n1053), .B2(n1052), .ZN(
        n1055) );
  AOI21D0BWP12T U1843 ( .A1(n1056), .A2(n1208), .B(n1055), .ZN(n1057) );
  ND4D1BWP12T U1844 ( .A1(n1060), .A2(n1059), .A3(n1058), .A4(n1057), .ZN(
        regC_out[9]) );
  AOI22D0BWP12T U1845 ( .A1(r12[14]), .A2(n1199), .B1(n1198), .B2(pc_out[14]), 
        .ZN(n1074) );
  AOI22D0BWP12T U1846 ( .A1(r9[14]), .A2(n1194), .B1(n1200), .B2(r11[14]), 
        .ZN(n1073) );
  AOI22D0BWP12T U1847 ( .A1(r7[14]), .A2(n1183), .B1(n1182), .B2(r4[14]), .ZN(
        n1064) );
  AOI22D0BWP12T U1848 ( .A1(r2[14]), .A2(n1185), .B1(n1184), .B2(r6[14]), .ZN(
        n1063) );
  AOI22D0BWP12T U1849 ( .A1(r5[14]), .A2(n1187), .B1(n1186), .B2(r1[14]), .ZN(
        n1062) );
  AOI22D0BWP12T U1850 ( .A1(r0[14]), .A2(n1189), .B1(n1188), .B2(r3[14]), .ZN(
        n1061) );
  ND4D1BWP12T U1851 ( .A1(n1064), .A2(n1063), .A3(n1062), .A4(n1061), .ZN(
        n1071) );
  CKND0BWP12T U1852 ( .I(r8[14]), .ZN(n1066) );
  OAI22D0BWP12T U1853 ( .A1(n1116), .A2(n1066), .B1(n1065), .B2(n1101), .ZN(
        n1070) );
  CKND0BWP12T U1854 ( .I(n[2027]), .ZN(n1068) );
  OAI22D0BWP12T U1855 ( .A1(n1068), .A2(n1148), .B1(n1160), .B2(n1067), .ZN(
        n1069) );
  AOI211D0BWP12T U1856 ( .A1(n1071), .A2(n1208), .B(n1070), .C(n1069), .ZN(
        n1072) );
  ND3D1BWP12T U1857 ( .A1(n1074), .A2(n1073), .A3(n1072), .ZN(regC_out[14]) );
  AOI22D0BWP12T U1858 ( .A1(r8[6]), .A2(n1195), .B1(n1194), .B2(r9[6]), .ZN(
        n1084) );
  AOI22D0BWP12T U1859 ( .A1(lr[6]), .A2(n1197), .B1(n1198), .B2(pc_out[6]), 
        .ZN(n1083) );
  AOI22D0BWP12T U1860 ( .A1(r10[6]), .A2(n1201), .B1(n1200), .B2(r11[6]), .ZN(
        n1082) );
  AOI22D0BWP12T U1861 ( .A1(r7[6]), .A2(n1183), .B1(n1182), .B2(r4[6]), .ZN(
        n1078) );
  AOI22D0BWP12T U1862 ( .A1(r2[6]), .A2(n1185), .B1(n1184), .B2(r6[6]), .ZN(
        n1077) );
  AOI22D0BWP12T U1863 ( .A1(r5[6]), .A2(n1187), .B1(n1186), .B2(r1[6]), .ZN(
        n1076) );
  AOI22D0BWP12T U1864 ( .A1(r0[6]), .A2(n1189), .B1(n1188), .B2(r3[6]), .ZN(
        n1075) );
  ND4D1BWP12T U1865 ( .A1(n1078), .A2(n1077), .A3(n1076), .A4(n1075), .ZN(
        n1080) );
  OAI22D0BWP12T U1866 ( .A1(n1748), .A2(n1148), .B1(n1172), .B2(n1744), .ZN(
        n1079) );
  AOI21D0BWP12T U1867 ( .A1(n1080), .A2(n1208), .B(n1079), .ZN(n1081) );
  ND4D1BWP12T U1868 ( .A1(n1084), .A2(n1083), .A3(n1082), .A4(n1081), .ZN(
        regC_out[6]) );
  AOI22D0BWP12T U1869 ( .A1(r8[11]), .A2(n1195), .B1(n1194), .B2(r9[11]), .ZN(
        n1096) );
  AOI22D0BWP12T U1870 ( .A1(lr[11]), .A2(n1197), .B1(n1198), .B2(pc_out[11]), 
        .ZN(n1095) );
  AOI22D0BWP12T U1871 ( .A1(r10[11]), .A2(n1201), .B1(n1200), .B2(r11[11]), 
        .ZN(n1094) );
  AOI22D0BWP12T U1872 ( .A1(r7[11]), .A2(n1183), .B1(n1182), .B2(r4[11]), .ZN(
        n1088) );
  AOI22D0BWP12T U1873 ( .A1(r2[11]), .A2(n1185), .B1(n1184), .B2(r6[11]), .ZN(
        n1087) );
  AOI22D0BWP12T U1874 ( .A1(r5[11]), .A2(n1187), .B1(n1186), .B2(r1[11]), .ZN(
        n1086) );
  AOI22D0BWP12T U1875 ( .A1(r0[11]), .A2(n1189), .B1(n1188), .B2(r3[11]), .ZN(
        n1085) );
  ND4D1BWP12T U1876 ( .A1(n1088), .A2(n1087), .A3(n1086), .A4(n1085), .ZN(
        n1092) );
  OAI22D0BWP12T U1877 ( .A1(n1090), .A2(n1148), .B1(n1172), .B2(n1089), .ZN(
        n1091) );
  AOI21D0BWP12T U1878 ( .A1(n1092), .A2(n1208), .B(n1091), .ZN(n1093) );
  ND4D1BWP12T U1879 ( .A1(n1096), .A2(n1095), .A3(n1094), .A4(n1093), .ZN(
        regC_out[11]) );
  AOI22D0BWP12T U1880 ( .A1(n[2034]), .A2(n1196), .B1(n1198), .B2(pc_out[7]), 
        .ZN(n1107) );
  AOI22D0BWP12T U1881 ( .A1(r9[7]), .A2(n1194), .B1(n1200), .B2(r11[7]), .ZN(
        n1106) );
  AOI22D0BWP12T U1882 ( .A1(r7[7]), .A2(n1183), .B1(n1182), .B2(r4[7]), .ZN(
        n1100) );
  AOI22D0BWP12T U1883 ( .A1(r2[7]), .A2(n1185), .B1(n1184), .B2(r6[7]), .ZN(
        n1099) );
  AOI22D0BWP12T U1884 ( .A1(r5[7]), .A2(n1187), .B1(n1186), .B2(r1[7]), .ZN(
        n1098) );
  AOI22D0BWP12T U1885 ( .A1(r0[7]), .A2(n1189), .B1(n1188), .B2(r3[7]), .ZN(
        n1097) );
  ND4D1BWP12T U1886 ( .A1(n1100), .A2(n1099), .A3(n1098), .A4(n1097), .ZN(
        n1104) );
  OAI22D0BWP12T U1887 ( .A1(n1172), .A2(n1717), .B1(n1722), .B2(n1116), .ZN(
        n1103) );
  OAI22D0BWP12T U1888 ( .A1(n1160), .A2(n1719), .B1(n1709), .B2(n1101), .ZN(
        n1102) );
  AOI211D0BWP12T U1889 ( .A1(n1104), .A2(n1208), .B(n1103), .C(n1102), .ZN(
        n1105) );
  ND3D1BWP12T U1890 ( .A1(n1107), .A2(n1106), .A3(n1105), .ZN(regC_out[7]) );
  AOI22D0BWP12T U1891 ( .A1(r12[22]), .A2(n1199), .B1(n1198), .B2(pc_out[22]), 
        .ZN(n1123) );
  AOI22D0BWP12T U1892 ( .A1(r9[22]), .A2(n1194), .B1(n1201), .B2(r10[22]), 
        .ZN(n1122) );
  AOI22D0BWP12T U1893 ( .A1(r7[22]), .A2(n1183), .B1(n1182), .B2(r4[22]), .ZN(
        n1111) );
  AOI22D0BWP12T U1894 ( .A1(r2[22]), .A2(n1185), .B1(n1184), .B2(r6[22]), .ZN(
        n1110) );
  AOI22D0BWP12T U1895 ( .A1(r5[22]), .A2(n1187), .B1(n1186), .B2(r1[22]), .ZN(
        n1109) );
  AOI22D0BWP12T U1896 ( .A1(r0[22]), .A2(n1189), .B1(n1188), .B2(r3[22]), .ZN(
        n1108) );
  ND4D1BWP12T U1897 ( .A1(n1111), .A2(n1110), .A3(n1109), .A4(n1108), .ZN(
        n1120) );
  CKND0BWP12T U1898 ( .I(lr[22]), .ZN(n1114) );
  CKND0BWP12T U1899 ( .I(r11[22]), .ZN(n1113) );
  OAI22D0BWP12T U1900 ( .A1(n1160), .A2(n1114), .B1(n1113), .B2(n1112), .ZN(
        n1119) );
  CKND0BWP12T U1901 ( .I(n[2019]), .ZN(n1117) );
  CKND0BWP12T U1902 ( .I(r8[22]), .ZN(n1115) );
  OAI22D0BWP12T U1903 ( .A1(n1117), .A2(n1148), .B1(n1116), .B2(n1115), .ZN(
        n1118) );
  AOI211D0BWP12T U1904 ( .A1(n1120), .A2(n1208), .B(n1119), .C(n1118), .ZN(
        n1121) );
  ND3D1BWP12T U1905 ( .A1(n1123), .A2(n1122), .A3(n1121), .ZN(regC_out[22]) );
  AOI22D0BWP12T U1906 ( .A1(r8[17]), .A2(n1195), .B1(n1201), .B2(r10[17]), 
        .ZN(n1134) );
  AOI22D0BWP12T U1907 ( .A1(r12[17]), .A2(n1199), .B1(n1198), .B2(pc_out[17]), 
        .ZN(n1133) );
  AOI22D0BWP12T U1908 ( .A1(r9[17]), .A2(n1194), .B1(n1200), .B2(r11[17]), 
        .ZN(n1132) );
  AOI22D0BWP12T U1909 ( .A1(r7[17]), .A2(n1183), .B1(n1182), .B2(r4[17]), .ZN(
        n1127) );
  AOI22D0BWP12T U1910 ( .A1(r2[17]), .A2(n1185), .B1(n1184), .B2(r6[17]), .ZN(
        n1126) );
  AOI22D0BWP12T U1911 ( .A1(r5[17]), .A2(n1187), .B1(n1186), .B2(r1[17]), .ZN(
        n1125) );
  AOI22D0BWP12T U1912 ( .A1(r0[17]), .A2(n1189), .B1(n1188), .B2(r3[17]), .ZN(
        n1124) );
  ND4D1BWP12T U1913 ( .A1(n1127), .A2(n1126), .A3(n1125), .A4(n1124), .ZN(
        n1130) );
  CKND0BWP12T U1914 ( .I(n[2024]), .ZN(n1128) );
  INVD1BWP12T U1915 ( .I(lr[17]), .ZN(n1503) );
  OAI22D0BWP12T U1916 ( .A1(n1128), .A2(n1148), .B1(n1160), .B2(n1503), .ZN(
        n1129) );
  AOI21D0BWP12T U1917 ( .A1(n1130), .A2(n1208), .B(n1129), .ZN(n1131) );
  ND4D1BWP12T U1918 ( .A1(n1134), .A2(n1133), .A3(n1132), .A4(n1131), .ZN(
        regC_out[17]) );
  OAI22D0BWP12T U1919 ( .A1(n1673), .A2(n1137), .B1(n1136), .B2(n1135), .ZN(
        n1147) );
  OAI22D0BWP12T U1920 ( .A1(n1671), .A2(n1139), .B1(n1138), .B2(n1660), .ZN(
        n1146) );
  OAI22D0BWP12T U1921 ( .A1(n1141), .A2(n1661), .B1(n1140), .B2(n1666), .ZN(
        n1145) );
  OAI22D0BWP12T U1922 ( .A1(n1672), .A2(n1143), .B1(n1142), .B2(n1670), .ZN(
        n1144) );
  NR4D0BWP12T U1923 ( .A1(n1147), .A2(n1146), .A3(n1145), .A4(n1144), .ZN(
        n1149) );
  OAI22D0BWP12T U1924 ( .A1(n1149), .A2(readC_sel[4]), .B1(n1148), .B2(n1668), 
        .ZN(n1150) );
  AOI21D0BWP12T U1925 ( .A1(lr[10]), .A2(n1197), .B(n1150), .ZN(n1154) );
  AOI22D0BWP12T U1926 ( .A1(r9[10]), .A2(n1194), .B1(n1200), .B2(r11[10]), 
        .ZN(n1153) );
  AOI22D0BWP12T U1927 ( .A1(r8[10]), .A2(n1195), .B1(n1201), .B2(r10[10]), 
        .ZN(n1152) );
  AOI22D0BWP12T U1928 ( .A1(r12[10]), .A2(n1199), .B1(n1198), .B2(pc_out[10]), 
        .ZN(n1151) );
  ND4D1BWP12T U1929 ( .A1(n1154), .A2(n1153), .A3(n1152), .A4(n1151), .ZN(
        regC_out[10]) );
  INVD1BWP12T U1930 ( .I(lr[13]), .ZN(n1588) );
  AOI22D0BWP12T U1931 ( .A1(r7[13]), .A2(n1183), .B1(n1182), .B2(r4[13]), .ZN(
        n1158) );
  AOI22D0BWP12T U1932 ( .A1(r2[13]), .A2(n1185), .B1(n1184), .B2(r6[13]), .ZN(
        n1157) );
  AOI22D0BWP12T U1933 ( .A1(r5[13]), .A2(n1187), .B1(n1186), .B2(r1[13]), .ZN(
        n1156) );
  AOI22D0BWP12T U1934 ( .A1(r0[13]), .A2(n1189), .B1(n1188), .B2(r3[13]), .ZN(
        n1155) );
  ND4D1BWP12T U1935 ( .A1(n1158), .A2(n1157), .A3(n1156), .A4(n1155), .ZN(
        n1159) );
  MOAI22D0BWP12T U1936 ( .A1(n1160), .A2(n1588), .B1(n1159), .B2(n1208), .ZN(
        n1161) );
  AOI21D0BWP12T U1937 ( .A1(n[2028]), .A2(n1196), .B(n1161), .ZN(n1165) );
  AOI22D0BWP12T U1938 ( .A1(r10[13]), .A2(n1201), .B1(n1200), .B2(r11[13]), 
        .ZN(n1164) );
  AOI22D0BWP12T U1939 ( .A1(r8[13]), .A2(n1195), .B1(n1194), .B2(r9[13]), .ZN(
        n1163) );
  AOI22D0BWP12T U1940 ( .A1(r12[13]), .A2(n1199), .B1(n1198), .B2(pc_out[13]), 
        .ZN(n1162) );
  ND4D1BWP12T U1941 ( .A1(n1165), .A2(n1164), .A3(n1163), .A4(n1162), .ZN(
        regC_out[13]) );
  CKND0BWP12T U1942 ( .I(r12[16]), .ZN(n1171) );
  AOI22D0BWP12T U1943 ( .A1(r7[16]), .A2(n1183), .B1(n1182), .B2(r4[16]), .ZN(
        n1169) );
  AOI22D0BWP12T U1944 ( .A1(r2[16]), .A2(n1185), .B1(n1184), .B2(r6[16]), .ZN(
        n1168) );
  AOI22D0BWP12T U1945 ( .A1(r5[16]), .A2(n1187), .B1(n1186), .B2(r1[16]), .ZN(
        n1167) );
  AOI22D0BWP12T U1946 ( .A1(r0[16]), .A2(n1189), .B1(n1188), .B2(r3[16]), .ZN(
        n1166) );
  ND4D1BWP12T U1947 ( .A1(n1169), .A2(n1168), .A3(n1167), .A4(n1166), .ZN(
        n1170) );
  MOAI22D0BWP12T U1948 ( .A1(n1172), .A2(n1171), .B1(n1170), .B2(n1208), .ZN(
        n1173) );
  AOI21D0BWP12T U1949 ( .A1(lr[16]), .A2(n1197), .B(n1173), .ZN(n1177) );
  AOI22D0BWP12T U1950 ( .A1(r9[16]), .A2(n1194), .B1(n1200), .B2(r11[16]), 
        .ZN(n1176) );
  AOI22D0BWP12T U1951 ( .A1(r8[16]), .A2(n1195), .B1(n1201), .B2(r10[16]), 
        .ZN(n1175) );
  AOI22D0BWP12T U1952 ( .A1(n[2025]), .A2(n1196), .B1(n1198), .B2(pc_out[16]), 
        .ZN(n1174) );
  ND4D1BWP12T U1953 ( .A1(n1177), .A2(n1176), .A3(n1175), .A4(n1174), .ZN(
        regC_out[16]) );
  CKND0BWP12T U1954 ( .I(n1178), .ZN(n1181) );
  TPAOI21D0BWP12T U1955 ( .A1(n1375), .A2(next_pc_in[1]), .B(reset), .ZN(n1180) );
  CKND2D0BWP12T U1956 ( .A1(n1363), .A2(pc_out[1]), .ZN(n1179) );
  OAI211D1BWP12T U1957 ( .A1(n1181), .A2(n1209), .B(n1180), .C(n1179), .ZN(
        n2170) );
  AOI22D0BWP12T U1958 ( .A1(r7[21]), .A2(n1183), .B1(n1182), .B2(r4[21]), .ZN(
        n1193) );
  AOI22D0BWP12T U1959 ( .A1(r2[21]), .A2(n1185), .B1(n1184), .B2(r6[21]), .ZN(
        n1192) );
  AOI22D0BWP12T U1960 ( .A1(r5[21]), .A2(n1187), .B1(n1186), .B2(r1[21]), .ZN(
        n1191) );
  AOI22D0BWP12T U1961 ( .A1(r0[21]), .A2(n1189), .B1(n1188), .B2(r3[21]), .ZN(
        n1190) );
  ND4D1BWP12T U1962 ( .A1(n1193), .A2(n1192), .A3(n1191), .A4(n1190), .ZN(
        n1207) );
  AOI22D0BWP12T U1963 ( .A1(r8[21]), .A2(n1195), .B1(n1194), .B2(r9[21]), .ZN(
        n1205) );
  AOI22D0BWP12T U1964 ( .A1(lr[21]), .A2(n1197), .B1(n1196), .B2(n[2020]), 
        .ZN(n1204) );
  AOI22D0BWP12T U1965 ( .A1(r12[21]), .A2(n1199), .B1(n1198), .B2(pc_out[21]), 
        .ZN(n1203) );
  AOI22D0BWP12T U1966 ( .A1(r10[21]), .A2(n1201), .B1(n1200), .B2(r11[21]), 
        .ZN(n1202) );
  ND4D1BWP12T U1967 ( .A1(n1205), .A2(n1204), .A3(n1203), .A4(n1202), .ZN(
        n1206) );
  AO21D1BWP12T U1968 ( .A1(n1208), .A2(n1207), .B(n1206), .Z(regC_out[21]) );
  AN2XD0BWP12T U1969 ( .A1(write2_in[5]), .A2(n1366), .Z(n1211) );
  AOI21D1BWP12T U1970 ( .A1(write1_in[5]), .A2(n1350), .B(n1211), .ZN(n1217)
         );
  TPND2D1BWP12T U1971 ( .A1(n1213), .A2(n1212), .ZN(n1216) );
  XOR2XD1BWP12T U1972 ( .A1(n1217), .A2(n1216), .Z(n1214) );
  AO222D1BWP12T U1973 ( .A1(n1214), .A2(n1364), .B1(n1375), .B2(next_pc_in[5]), 
        .C1(n1363), .C2(pc_out[5]), .Z(n2174) );
  CKND2D0BWP12T U1974 ( .A1(write2_in[6]), .A2(n1366), .ZN(n1215) );
  IOA21D1BWP12T U1975 ( .A1(write1_in[6]), .A2(n1350), .B(n1215), .ZN(n1221)
         );
  TPNR2D1BWP12T U1976 ( .A1(n1217), .A2(n1216), .ZN(n1220) );
  XOR2XD1BWP12T U1977 ( .A1(n1221), .A2(n1220), .Z(n1218) );
  AO222D1BWP12T U1978 ( .A1(n1218), .A2(n1364), .B1(n1375), .B2(next_pc_in[6]), 
        .C1(n1363), .C2(pc_out[6]), .Z(n2175) );
  AN2XD0BWP12T U1979 ( .A1(write2_in[7]), .A2(n1366), .Z(n1219) );
  AOI21D1BWP12T U1980 ( .A1(write1_in[7]), .A2(n1350), .B(n1219), .ZN(n1223)
         );
  TPND2D1BWP12T U1981 ( .A1(n1221), .A2(n1220), .ZN(n1222) );
  AN2XD0BWP12T U1982 ( .A1(write2_in[9]), .A2(n1366), .Z(n1224) );
  AOI21D1BWP12T U1983 ( .A1(write1_in[9]), .A2(n1350), .B(n1224), .ZN(n1228)
         );
  TPND2D1BWP12T U1984 ( .A1(n1226), .A2(n1225), .ZN(n1227) );
  AO222D1BWP12T U1985 ( .A1(n1301), .A2(write1_in[17]), .B1(n1300), .B2(
        n[2024]), .C1(write2_in[17]), .C2(n1299), .Z(spin[17]) );
  AO222D1BWP12T U1986 ( .A1(n1303), .A2(write1_in[17]), .B1(n757), .B2(
        write2_in[17]), .C1(n1302), .C2(tmp1[17]), .Z(n2154) );
  NR2XD1BWP12T U1987 ( .A1(n1228), .A2(n1227), .ZN(n1231) );
  AO222D1BWP12T U1988 ( .A1(n1301), .A2(n1307), .B1(n1300), .B2(n[2022]), .C1(
        write2_in[19]), .C2(n1299), .Z(spin[19]) );
  AO222D1BWP12T U1989 ( .A1(n1301), .A2(write1_in[21]), .B1(n1300), .B2(
        n[2020]), .C1(write2_in[21]), .C2(n1299), .Z(spin[21]) );
  AO222D1BWP12T U1990 ( .A1(n1274), .A2(n1309), .B1(n1273), .B2(r1[20]), .C1(
        write2_in[20]), .C2(n1272), .Z(n2605) );
  AO222D1BWP12T U1991 ( .A1(n1277), .A2(n1309), .B1(n1276), .B2(r4[20]), .C1(
        write2_in[20]), .C2(n1275), .Z(n2509) );
  AO222D1BWP12T U1992 ( .A1(n1268), .A2(n1309), .B1(n1267), .B2(r5[20]), .C1(
        write2_in[20]), .C2(n1266), .Z(n2477) );
  AO222D1BWP12T U1993 ( .A1(n1286), .A2(n1309), .B1(n1285), .B2(r12[20]), .C1(
        write2_in[20]), .C2(n1284), .Z(n2253) );
  AO222D1BWP12T U1994 ( .A1(n1259), .A2(n1309), .B1(n1258), .B2(r8[20]), .C1(
        write2_in[20]), .C2(n1257), .Z(n2381) );
  AO222D1BWP12T U1995 ( .A1(n1265), .A2(n1309), .B1(n1264), .B2(r0[20]), .C1(
        write2_in[20]), .C2(n1263), .Z(n2637) );
  AO222D1BWP12T U1996 ( .A1(n1283), .A2(n1309), .B1(n1282), .B2(r9[20]), .C1(
        write2_in[20]), .C2(n1281), .Z(n2349) );
  AO222D1BWP12T U1997 ( .A1(n1295), .A2(n1309), .B1(n1294), .B2(write2_in[20]), 
        .C1(n1293), .C2(r10[20]), .Z(n2317) );
  AO222D1BWP12T U1998 ( .A1(n1301), .A2(n1309), .B1(n1300), .B2(n[2021]), .C1(
        write2_in[20]), .C2(n1299), .Z(spin[20]) );
  AO222D1BWP12T U1999 ( .A1(n1303), .A2(n1309), .B1(n757), .B2(write2_in[20]), 
        .C1(n1302), .C2(tmp1[20]), .Z(n2157) );
  AN2XD0BWP12T U2000 ( .A1(write2_in[11]), .A2(n1366), .Z(n1229) );
  AOI21D1BWP12T U2001 ( .A1(write1_in[11]), .A2(n1350), .B(n1229), .ZN(n1235)
         );
  CKND2D2BWP12T U2002 ( .A1(n1231), .A2(n1230), .ZN(n1234) );
  XOR2XD1BWP12T U2003 ( .A1(n1235), .A2(n1234), .Z(n1232) );
  AO222D1BWP12T U2004 ( .A1(n1232), .A2(n1364), .B1(n1375), .B2(next_pc_in[11]), .C1(n1363), .C2(pc_out[11]), .Z(n2180) );
  CKND2D0BWP12T U2005 ( .A1(write2_in[12]), .A2(n1366), .ZN(n1233) );
  IOA21D1BWP12T U2006 ( .A1(write1_in[12]), .A2(n1350), .B(n1233), .ZN(n1238)
         );
  NR2XD1BWP12T U2007 ( .A1(n1235), .A2(n1234), .ZN(n1237) );
  XOR2XD1BWP12T U2008 ( .A1(n1238), .A2(n1237), .Z(n1236) );
  AO222D1BWP12T U2009 ( .A1(n1236), .A2(n1364), .B1(n1375), .B2(next_pc_in[12]), .C1(n1363), .C2(pc_out[12]), .Z(n2181) );
  TPND2D2BWP12T U2010 ( .A1(n1238), .A2(n1237), .ZN(n1241) );
  AN2XD0BWP12T U2011 ( .A1(write2_in[13]), .A2(n1366), .Z(n1239) );
  AOI21D1BWP12T U2012 ( .A1(write1_in[13]), .A2(n1350), .B(n1239), .ZN(n1240)
         );
  BUFFD3BWP12T U2013 ( .I(write1_in[22]), .Z(n1318) );
  AO222D1BWP12T U2014 ( .A1(n1298), .A2(n1318), .B1(n1297), .B2(write2_in[22]), 
        .C1(n1296), .C2(r3[22]), .Z(n2543) );
  AO222D1BWP12T U2015 ( .A1(n1292), .A2(n1318), .B1(n1291), .B2(write2_in[22]), 
        .C1(n1290), .C2(r2[22]), .Z(n2575) );
  AO222D1BWP12T U2016 ( .A1(n1289), .A2(n1318), .B1(n1288), .B2(write2_in[22]), 
        .C1(n1287), .C2(r11[22]), .Z(n2287) );
  AO222D1BWP12T U2017 ( .A1(n1295), .A2(n1318), .B1(n1294), .B2(write2_in[22]), 
        .C1(n1293), .C2(r10[22]), .Z(n2319) );
  AO222D1BWP12T U2018 ( .A1(n1280), .A2(n1318), .B1(n1279), .B2(lr[22]), .C1(
        write2_in[22]), .C2(n1278), .Z(n2223) );
  AO222D1BWP12T U2019 ( .A1(n1283), .A2(n1318), .B1(n1282), .B2(r9[22]), .C1(
        write2_in[22]), .C2(n1281), .Z(n2351) );
  AO222D1BWP12T U2020 ( .A1(n1265), .A2(n1318), .B1(n1264), .B2(r0[22]), .C1(
        write2_in[22]), .C2(n1263), .Z(n2639) );
  AO222D1BWP12T U2021 ( .A1(n1259), .A2(n1318), .B1(n1258), .B2(r8[22]), .C1(
        write2_in[22]), .C2(n1257), .Z(n2383) );
  AO222D1BWP12T U2022 ( .A1(n1268), .A2(n1318), .B1(n1267), .B2(r5[22]), .C1(
        write2_in[22]), .C2(n1266), .Z(n2479) );
  AO222D1BWP12T U2023 ( .A1(n1274), .A2(n1318), .B1(n1273), .B2(r1[22]), .C1(
        write2_in[22]), .C2(n1272), .Z(n2607) );
  AO222D1BWP12T U2024 ( .A1(n1277), .A2(n1318), .B1(n1276), .B2(r4[22]), .C1(
        write2_in[22]), .C2(n1275), .Z(n2511) );
  AO222D1BWP12T U2025 ( .A1(n1286), .A2(n1318), .B1(n1285), .B2(r12[22]), .C1(
        write2_in[22]), .C2(n1284), .Z(n2255) );
  AO222D1BWP12T U2026 ( .A1(n1262), .A2(n1318), .B1(n1261), .B2(r7[22]), .C1(
        write2_in[22]), .C2(n1260), .Z(n2415) );
  AO222D1BWP12T U2027 ( .A1(n1271), .A2(n1318), .B1(n1270), .B2(r6[22]), .C1(
        write2_in[22]), .C2(n1269), .Z(n2447) );
  AO222D1BWP12T U2028 ( .A1(n1301), .A2(n1318), .B1(n1300), .B2(n[2019]), .C1(
        write2_in[22]), .C2(n1299), .Z(spin[22]) );
  AO222D1BWP12T U2029 ( .A1(n1303), .A2(n1318), .B1(n757), .B2(write2_in[22]), 
        .C1(n1302), .C2(tmp1[22]), .Z(n2159) );
  AO222D1BWP12T U2030 ( .A1(n1283), .A2(n1322), .B1(n1282), .B2(r9[23]), .C1(
        write2_in[23]), .C2(n1281), .Z(n2352) );
  AO222D1BWP12T U2031 ( .A1(n1277), .A2(n1322), .B1(n1276), .B2(r4[23]), .C1(
        write2_in[23]), .C2(n1275), .Z(n2512) );
  AO222D1BWP12T U2032 ( .A1(n1268), .A2(n1322), .B1(n1267), .B2(r5[23]), .C1(
        write2_in[23]), .C2(n1266), .Z(n2480) );
  AO222D1BWP12T U2033 ( .A1(n1274), .A2(n1322), .B1(n1273), .B2(r1[23]), .C1(
        write2_in[23]), .C2(n1272), .Z(n2608) );
  AO222D1BWP12T U2034 ( .A1(n1271), .A2(n1322), .B1(n1270), .B2(r6[23]), .C1(
        write2_in[23]), .C2(n1269), .Z(n2448) );
  AO222D1BWP12T U2035 ( .A1(n1265), .A2(n1322), .B1(n1264), .B2(r0[23]), .C1(
        write2_in[23]), .C2(n1263), .Z(n2640) );
  AO222D1BWP12T U2036 ( .A1(n1262), .A2(n1322), .B1(n1261), .B2(r7[23]), .C1(
        write2_in[23]), .C2(n1260), .Z(n2416) );
  AO222D1BWP12T U2037 ( .A1(n1259), .A2(n1322), .B1(n1258), .B2(r8[23]), .C1(
        write2_in[23]), .C2(n1257), .Z(n2384) );
  AO222D1BWP12T U2038 ( .A1(n1286), .A2(n1322), .B1(n1285), .B2(r12[23]), .C1(
        write2_in[23]), .C2(n1284), .Z(n2256) );
  AO222D1BWP12T U2039 ( .A1(n1280), .A2(n1322), .B1(n1279), .B2(lr[23]), .C1(
        write2_in[23]), .C2(n1278), .Z(n2224) );
  AO222D1BWP12T U2040 ( .A1(n1298), .A2(n1322), .B1(n1297), .B2(write2_in[23]), 
        .C1(n1296), .C2(r3[23]), .Z(n2544) );
  AO222D1BWP12T U2041 ( .A1(n1289), .A2(n1322), .B1(n1288), .B2(write2_in[23]), 
        .C1(n1287), .C2(r11[23]), .Z(n2288) );
  AO222D1BWP12T U2042 ( .A1(n1292), .A2(n1322), .B1(n1291), .B2(write2_in[23]), 
        .C1(n1290), .C2(r2[23]), .Z(n2576) );
  NR2D2BWP12T U2043 ( .A1(n1241), .A2(n1240), .ZN(n1242) );
  AO222D1BWP12T U2044 ( .A1(n1301), .A2(n1322), .B1(n1300), .B2(n[2018]), .C1(
        write2_in[23]), .C2(n1299), .Z(spin[23]) );
  AO222D1BWP12T U2045 ( .A1(n1303), .A2(n1322), .B1(n757), .B2(write2_in[23]), 
        .C1(n1302), .C2(tmp1[23]), .Z(n2160) );
  TPND2D1BWP12T U2046 ( .A1(n1243), .A2(n1242), .ZN(n1249) );
  AN2XD0BWP12T U2047 ( .A1(write2_in[15]), .A2(n1366), .Z(n1244) );
  AOI21D1BWP12T U2048 ( .A1(n1245), .A2(n1350), .B(n1244), .ZN(n1248) );
  BUFFXD4BWP12T U2049 ( .I(write1_in[24]), .Z(n1324) );
  AO222D1BWP12T U2050 ( .A1(n1280), .A2(n1324), .B1(n1279), .B2(lr[24]), .C1(
        write2_in[24]), .C2(n1278), .Z(n2225) );
  AO222D1BWP12T U2051 ( .A1(n1286), .A2(n1324), .B1(n1285), .B2(r12[24]), .C1(
        write2_in[24]), .C2(n1284), .Z(n2257) );
  AO222D1BWP12T U2052 ( .A1(n1265), .A2(n1324), .B1(n1264), .B2(r0[24]), .C1(
        write2_in[24]), .C2(n1263), .Z(n2641) );
  AO222D1BWP12T U2053 ( .A1(n1271), .A2(n1324), .B1(n1270), .B2(r6[24]), .C1(
        write2_in[24]), .C2(n1269), .Z(n2449) );
  AO222D1BWP12T U2054 ( .A1(n1268), .A2(n1324), .B1(n1267), .B2(r5[24]), .C1(
        write2_in[24]), .C2(n1266), .Z(n2481) );
  AO222D1BWP12T U2055 ( .A1(n1259), .A2(n1324), .B1(n1258), .B2(r8[24]), .C1(
        write2_in[24]), .C2(n1257), .Z(n2385) );
  AO222D1BWP12T U2056 ( .A1(n1283), .A2(n1324), .B1(n1282), .B2(r9[24]), .C1(
        write2_in[24]), .C2(n1281), .Z(n2353) );
  AO222D1BWP12T U2057 ( .A1(n1277), .A2(n1324), .B1(n1276), .B2(r4[24]), .C1(
        write2_in[24]), .C2(n1275), .Z(n2513) );
  AO222D1BWP12T U2058 ( .A1(n1262), .A2(n1324), .B1(n1261), .B2(r7[24]), .C1(
        write2_in[24]), .C2(n1260), .Z(n2417) );
  AO222D1BWP12T U2059 ( .A1(n1274), .A2(n1324), .B1(n1273), .B2(r1[24]), .C1(
        write2_in[24]), .C2(n1272), .Z(n2609) );
  AO222D1BWP12T U2060 ( .A1(n1295), .A2(n1324), .B1(n1294), .B2(write2_in[24]), 
        .C1(n1293), .C2(r10[24]), .Z(n2321) );
  AO222D1BWP12T U2061 ( .A1(n1298), .A2(n1324), .B1(n1297), .B2(write2_in[24]), 
        .C1(n1296), .C2(r3[24]), .Z(n2545) );
  AO222D1BWP12T U2062 ( .A1(n1292), .A2(n1324), .B1(n1291), .B2(write2_in[24]), 
        .C1(n1290), .C2(r2[24]), .Z(n2577) );
  AO222D1BWP12T U2063 ( .A1(n1289), .A2(n1324), .B1(n1288), .B2(write2_in[24]), 
        .C1(n1287), .C2(r11[24]), .Z(n2289) );
  AO222D1BWP12T U2064 ( .A1(n1301), .A2(n1324), .B1(n1300), .B2(n[2017]), .C1(
        write2_in[24]), .C2(n1299), .Z(spin[24]) );
  AO222D1BWP12T U2065 ( .A1(n1303), .A2(n1324), .B1(n757), .B2(write2_in[24]), 
        .C1(n1302), .C2(tmp1[24]), .Z(n2161) );
  CKND2D0BWP12T U2066 ( .A1(write2_in[16]), .A2(n1366), .ZN(n1246) );
  TPNR2D1BWP12T U2067 ( .A1(n1249), .A2(n1248), .ZN(n1250) );
  AO222D1BWP12T U2068 ( .A1(n1265), .A2(write1_in[25]), .B1(n1264), .B2(r0[25]), .C1(write2_in[25]), .C2(n1263), .Z(n2642) );
  AO222D1BWP12T U2069 ( .A1(n1283), .A2(write1_in[25]), .B1(n1282), .B2(r9[25]), .C1(write2_in[25]), .C2(n1281), .Z(n2354) );
  AO222D1BWP12T U2070 ( .A1(n1277), .A2(write1_in[25]), .B1(n1276), .B2(r4[25]), .C1(write2_in[25]), .C2(n1275), .Z(n2514) );
  AO222D1BWP12T U2071 ( .A1(n1259), .A2(write1_in[25]), .B1(n1258), .B2(r8[25]), .C1(write2_in[25]), .C2(n1257), .Z(n2386) );
  AO222D1BWP12T U2072 ( .A1(n1268), .A2(write1_in[25]), .B1(n1267), .B2(r5[25]), .C1(write2_in[25]), .C2(n1266), .Z(n2482) );
  AO222D1BWP12T U2073 ( .A1(n1280), .A2(write1_in[25]), .B1(n1279), .B2(lr[25]), .C1(write2_in[25]), .C2(n1278), .Z(n2226) );
  AO222D1BWP12T U2074 ( .A1(n1286), .A2(write1_in[25]), .B1(n1285), .B2(
        r12[25]), .C1(write2_in[25]), .C2(n1284), .Z(n2258) );
  AO222D1BWP12T U2075 ( .A1(n1274), .A2(write1_in[25]), .B1(n1273), .B2(r1[25]), .C1(write2_in[25]), .C2(n1272), .Z(n2610) );
  AO222D1BWP12T U2076 ( .A1(n1262), .A2(write1_in[25]), .B1(n1261), .B2(r7[25]), .C1(write2_in[25]), .C2(n1260), .Z(n2418) );
  AO222D1BWP12T U2077 ( .A1(n1271), .A2(write1_in[25]), .B1(n1270), .B2(r6[25]), .C1(write2_in[25]), .C2(n1269), .Z(n2450) );
  AO222D1BWP12T U2078 ( .A1(n1289), .A2(write1_in[25]), .B1(n1288), .B2(
        write2_in[25]), .C1(n1287), .C2(r11[25]), .Z(n2290) );
  AO222D1BWP12T U2079 ( .A1(n1292), .A2(write1_in[25]), .B1(n1291), .B2(
        write2_in[25]), .C1(n1290), .C2(r2[25]), .Z(n2578) );
  AO222D1BWP12T U2080 ( .A1(n1295), .A2(write1_in[25]), .B1(n1294), .B2(
        write2_in[25]), .C1(n1293), .C2(r10[25]), .Z(n2322) );
  AO222D1BWP12T U2081 ( .A1(n1298), .A2(write1_in[25]), .B1(n1297), .B2(
        write2_in[25]), .C1(n1296), .C2(r3[25]), .Z(n2546) );
  AO222D1BWP12T U2082 ( .A1(n1301), .A2(write1_in[25]), .B1(n1300), .B2(
        n[2016]), .C1(write2_in[25]), .C2(n1299), .Z(spin[25]) );
  AO222D1BWP12T U2083 ( .A1(n1303), .A2(write1_in[25]), .B1(n757), .B2(
        write2_in[25]), .C1(n1302), .C2(tmp1[25]), .Z(n2162) );
  BUFFXD3BWP12T U2084 ( .I(write1_in[26]), .Z(n1330) );
  AO222D1BWP12T U2085 ( .A1(n1295), .A2(n1330), .B1(n1294), .B2(write2_in[26]), 
        .C1(n1293), .C2(r10[26]), .Z(n2323) );
  AO222D1BWP12T U2086 ( .A1(n1298), .A2(n1330), .B1(n1297), .B2(write2_in[26]), 
        .C1(n1296), .C2(r3[26]), .Z(n2547) );
  AO222D1BWP12T U2087 ( .A1(n1289), .A2(n1330), .B1(n1288), .B2(write2_in[26]), 
        .C1(n1287), .C2(r11[26]), .Z(n2291) );
  AO222D1BWP12T U2088 ( .A1(n1292), .A2(n1330), .B1(n1291), .B2(write2_in[26]), 
        .C1(n1290), .C2(r2[26]), .Z(n2579) );
  AO222D1BWP12T U2089 ( .A1(n1286), .A2(n1330), .B1(n1285), .B2(r12[26]), .C1(
        write2_in[26]), .C2(n1284), .Z(n2259) );
  AO222D1BWP12T U2090 ( .A1(n1280), .A2(n1330), .B1(n1279), .B2(lr[26]), .C1(
        write2_in[26]), .C2(n1278), .Z(n2227) );
  AO222D1BWP12T U2091 ( .A1(n1283), .A2(n1330), .B1(n1282), .B2(r9[26]), .C1(
        write2_in[26]), .C2(n1281), .Z(n2355) );
  AO222D1BWP12T U2092 ( .A1(n1277), .A2(n1330), .B1(n1276), .B2(r4[26]), .C1(
        write2_in[26]), .C2(n1275), .Z(n2515) );
  AO222D1BWP12T U2093 ( .A1(n1262), .A2(n1330), .B1(n1261), .B2(r7[26]), .C1(
        write2_in[26]), .C2(n1260), .Z(n2419) );
  AO222D1BWP12T U2094 ( .A1(n1259), .A2(n1330), .B1(n1258), .B2(r8[26]), .C1(
        write2_in[26]), .C2(n1257), .Z(n2387) );
  AO222D1BWP12T U2095 ( .A1(n1271), .A2(n1330), .B1(n1270), .B2(r6[26]), .C1(
        write2_in[26]), .C2(n1269), .Z(n2451) );
  AO222D1BWP12T U2096 ( .A1(n1274), .A2(n1330), .B1(n1273), .B2(r1[26]), .C1(
        write2_in[26]), .C2(n1272), .Z(n2611) );
  AO222D1BWP12T U2097 ( .A1(n1265), .A2(n1330), .B1(n1264), .B2(r0[26]), .C1(
        write2_in[26]), .C2(n1263), .Z(n2643) );
  AO222D1BWP12T U2098 ( .A1(n1268), .A2(n1330), .B1(n1267), .B2(r5[26]), .C1(
        write2_in[26]), .C2(n1266), .Z(n2483) );
  AO222D1BWP12T U2099 ( .A1(n1301), .A2(n1330), .B1(n1300), .B2(n[2015]), .C1(
        write2_in[26]), .C2(n1299), .Z(spin[26]) );
  AO222D1BWP12T U2100 ( .A1(n1303), .A2(n1330), .B1(n757), .B2(write2_in[26]), 
        .C1(n1302), .C2(tmp1[26]), .Z(n2163) );
  TPND2D1BWP12T U2101 ( .A1(n1251), .A2(n1250), .ZN(n1254) );
  AN2XD0BWP12T U2102 ( .A1(write2_in[17]), .A2(n1366), .Z(n1252) );
  AOI21D1BWP12T U2103 ( .A1(write1_in[17]), .A2(n1350), .B(n1252), .ZN(n1253)
         );
  AO222D1BWP12T U2104 ( .A1(n1286), .A2(n1337), .B1(n1285), .B2(r12[27]), .C1(
        write2_in[27]), .C2(n1284), .Z(n2260) );
  AO222D1BWP12T U2105 ( .A1(n1268), .A2(n1337), .B1(n1267), .B2(r5[27]), .C1(
        write2_in[27]), .C2(n1266), .Z(n2484) );
  AO222D1BWP12T U2106 ( .A1(n1277), .A2(n1337), .B1(n1276), .B2(r4[27]), .C1(
        write2_in[27]), .C2(n1275), .Z(n2516) );
  AO222D1BWP12T U2107 ( .A1(n1271), .A2(n1337), .B1(n1270), .B2(r6[27]), .C1(
        write2_in[27]), .C2(n1269), .Z(n2452) );
  AO222D1BWP12T U2108 ( .A1(n1259), .A2(n1337), .B1(n1258), .B2(r8[27]), .C1(
        write2_in[27]), .C2(n1257), .Z(n2388) );
  AO222D1BWP12T U2109 ( .A1(n1280), .A2(n1337), .B1(n1279), .B2(lr[27]), .C1(
        write2_in[27]), .C2(n1278), .Z(n2228) );
  AO222D1BWP12T U2110 ( .A1(n1262), .A2(n1337), .B1(n1261), .B2(r7[27]), .C1(
        write2_in[27]), .C2(n1260), .Z(n2420) );
  AO222D1BWP12T U2111 ( .A1(n1265), .A2(n1337), .B1(n1264), .B2(r0[27]), .C1(
        write2_in[27]), .C2(n1263), .Z(n2644) );
  AO222D1BWP12T U2112 ( .A1(n1283), .A2(n1337), .B1(n1282), .B2(r9[27]), .C1(
        write2_in[27]), .C2(n1281), .Z(n2356) );
  AO222D1BWP12T U2113 ( .A1(n1274), .A2(n1337), .B1(n1273), .B2(r1[27]), .C1(
        write2_in[27]), .C2(n1272), .Z(n2612) );
  AO222D1BWP12T U2114 ( .A1(n1292), .A2(n1337), .B1(n1291), .B2(write2_in[27]), 
        .C1(n1290), .C2(r2[27]), .Z(n2580) );
  AO222D1BWP12T U2115 ( .A1(n1289), .A2(n1337), .B1(n1288), .B2(write2_in[27]), 
        .C1(n1287), .C2(r11[27]), .Z(n2292) );
  AO222D1BWP12T U2116 ( .A1(n1295), .A2(n1337), .B1(n1294), .B2(write2_in[27]), 
        .C1(n1293), .C2(r10[27]), .Z(n2324) );
  AO222D1BWP12T U2117 ( .A1(n1298), .A2(n1337), .B1(n1297), .B2(write2_in[27]), 
        .C1(n1296), .C2(r3[27]), .Z(n2548) );
  AO222D1BWP12T U2118 ( .A1(n1301), .A2(n1337), .B1(n1300), .B2(n[2014]), .C1(
        write2_in[27]), .C2(n1299), .Z(spin[27]) );
  NR2D2BWP12T U2119 ( .A1(n1254), .A2(n1253), .ZN(n1305) );
  CKND2D0BWP12T U2120 ( .A1(write2_in[18]), .A2(n1366), .ZN(n1255) );
  IOA21D1BWP12T U2121 ( .A1(n1256), .A2(n1350), .B(n1255), .ZN(n1304) );
  AO222D1BWP12T U2122 ( .A1(n1303), .A2(n1337), .B1(n757), .B2(write2_in[27]), 
        .C1(n1302), .C2(tmp1[27]), .Z(n2164) );
  BUFFD2BWP12T U2123 ( .I(write1_in[29]), .Z(n1351) );
  AO222D1BWP12T U2124 ( .A1(n1259), .A2(n1351), .B1(n1258), .B2(r8[29]), .C1(
        write2_in[29]), .C2(n1257), .Z(n2390) );
  AO222D1BWP12T U2125 ( .A1(n1262), .A2(n1351), .B1(n1261), .B2(r7[29]), .C1(
        write2_in[29]), .C2(n1260), .Z(n2422) );
  AO222D1BWP12T U2126 ( .A1(n1265), .A2(n1351), .B1(n1264), .B2(r0[29]), .C1(
        write2_in[29]), .C2(n1263), .Z(n2646) );
  AO222D1BWP12T U2127 ( .A1(n1268), .A2(n1351), .B1(n1267), .B2(r5[29]), .C1(
        write2_in[29]), .C2(n1266), .Z(n2486) );
  AO222D1BWP12T U2128 ( .A1(n1271), .A2(n1351), .B1(n1270), .B2(r6[29]), .C1(
        write2_in[29]), .C2(n1269), .Z(n2454) );
  AO222D1BWP12T U2129 ( .A1(n1274), .A2(n1351), .B1(n1273), .B2(r1[29]), .C1(
        write2_in[29]), .C2(n1272), .Z(n2614) );
  AO222D1BWP12T U2130 ( .A1(n1277), .A2(n1351), .B1(n1276), .B2(r4[29]), .C1(
        write2_in[29]), .C2(n1275), .Z(n2518) );
  AO222D1BWP12T U2131 ( .A1(n1280), .A2(n1351), .B1(n1279), .B2(lr[29]), .C1(
        write2_in[29]), .C2(n1278), .Z(n2230) );
  AO222D1BWP12T U2132 ( .A1(n1283), .A2(n1351), .B1(n1282), .B2(r9[29]), .C1(
        write2_in[29]), .C2(n1281), .Z(n2358) );
  AO222D1BWP12T U2133 ( .A1(n1286), .A2(n1351), .B1(n1285), .B2(r12[29]), .C1(
        write2_in[29]), .C2(n1284), .Z(n2262) );
  AO222D1BWP12T U2134 ( .A1(n1289), .A2(n1351), .B1(n1288), .B2(write2_in[29]), 
        .C1(n1287), .C2(r11[29]), .Z(n2294) );
  AO222D1BWP12T U2135 ( .A1(n1292), .A2(n1351), .B1(n1291), .B2(write2_in[29]), 
        .C1(n1290), .C2(r2[29]), .Z(n2582) );
  AO222D1BWP12T U2136 ( .A1(n1295), .A2(n1351), .B1(n1294), .B2(write2_in[29]), 
        .C1(n1293), .C2(r10[29]), .Z(n2326) );
  AO222D1BWP12T U2137 ( .A1(n1298), .A2(n1351), .B1(n1297), .B2(write2_in[29]), 
        .C1(n1296), .C2(r3[29]), .Z(n2550) );
  AO222D1BWP12T U2138 ( .A1(n1301), .A2(n1351), .B1(n1300), .B2(n[2012]), .C1(
        write2_in[29]), .C2(n1299), .Z(spin[29]) );
  AO222D1BWP12T U2139 ( .A1(n1303), .A2(n1351), .B1(n757), .B2(write2_in[29]), 
        .C1(n1302), .C2(tmp1[29]), .Z(n2166) );
  CKND2D2BWP12T U2140 ( .A1(n1305), .A2(n1304), .ZN(n1311) );
  AN2XD0BWP12T U2141 ( .A1(write2_in[19]), .A2(n1366), .Z(n1306) );
  AOI21D1BWP12T U2142 ( .A1(n1307), .A2(n1350), .B(n1306), .ZN(n1310) );
  ND2XD0BWP12T U2143 ( .A1(write2_in[20]), .A2(n1366), .ZN(n1308) );
  IOA21D2BWP12T U2144 ( .A1(n1309), .A2(n1350), .B(n1308), .ZN(n1314) );
  TPNR2D2BWP12T U2145 ( .A1(n1311), .A2(n1310), .ZN(n1313) );
  XOR2XD1BWP12T U2146 ( .A1(n1314), .A2(n1313), .Z(n1312) );
  AO222D1BWP12T U2147 ( .A1(n1312), .A2(n1364), .B1(n1375), .B2(next_pc_in[20]), .C1(n1363), .C2(pc_out[20]), .Z(n2189) );
  ND2D3BWP12T U2148 ( .A1(n1314), .A2(n1313), .ZN(n1316) );
  TPNR2D3BWP12T U2149 ( .A1(n1316), .A2(n1315), .ZN(n1320) );
  CKND2D0BWP12T U2150 ( .A1(write2_in[22]), .A2(n1366), .ZN(n1317) );
  IOA21D1BWP12T U2151 ( .A1(n1318), .A2(n1350), .B(n1317), .ZN(n1319) );
  ND2XD3BWP12T U2152 ( .A1(n1320), .A2(n1319), .ZN(n1331) );
  CKAN2D1BWP12T U2153 ( .A1(write2_in[23]), .A2(n1366), .Z(n1321) );
  TPNR2D1BWP12T U2154 ( .A1(n1331), .A2(n1333), .ZN(n1326) );
  CKAN2D0BWP12T U2155 ( .A1(write2_in[24]), .A2(n1366), .Z(n1323) );
  AOI21D1BWP12T U2156 ( .A1(n1324), .A2(n1350), .B(n1323), .ZN(n1332) );
  INVD1BWP12T U2157 ( .I(n1332), .ZN(n1325) );
  ND2D1BWP12T U2158 ( .A1(n1326), .A2(n1325), .ZN(n1339) );
  CKAN2D0BWP12T U2159 ( .A1(write2_in[25]), .A2(n1366), .Z(n1327) );
  AOI21D1BWP12T U2160 ( .A1(write1_in[25]), .A2(n1350), .B(n1327), .ZN(n1338)
         );
  XOR2D1BWP12T U2161 ( .A1(n1339), .A2(n1338), .Z(n1328) );
  AO222D1BWP12T U2162 ( .A1(n1328), .A2(n1364), .B1(n1375), .B2(next_pc_in[25]), .C1(n1363), .C2(pc_out[25]), .Z(n2194) );
  AN2XD0BWP12T U2163 ( .A1(write2_in[26]), .A2(n1366), .Z(n1329) );
  AOI21D1BWP12T U2164 ( .A1(n1330), .A2(n1350), .B(n1329), .ZN(n1340) );
  TPNR2D1BWP12T U2165 ( .A1(n1340), .A2(n1331), .ZN(n1335) );
  NR3D1BWP12T U2166 ( .A1(n1338), .A2(n1333), .A3(n1332), .ZN(n1334) );
  AN2XD0BWP12T U2167 ( .A1(write2_in[27]), .A2(n1366), .Z(n1336) );
  XNR2D1BWP12T U2168 ( .A1(n1341), .A2(n1340), .ZN(n1342) );
  AO222D1BWP12T U2169 ( .A1(n1342), .A2(n1364), .B1(n1375), .B2(next_pc_in[26]), .C1(n1363), .C2(pc_out[26]), .Z(n2195) );
  CKND2D0BWP12T U2170 ( .A1(write2_in[28]), .A2(n1366), .ZN(n1345) );
  IOA21D2BWP12T U2171 ( .A1(n1346), .A2(n1350), .B(n1345), .ZN(n1347) );
  CKAN2D0BWP12T U2172 ( .A1(write2_in[29]), .A2(n1366), .Z(n1349) );
  AOI21D1BWP12T U2173 ( .A1(n1351), .A2(n1350), .B(n1349), .ZN(n1361) );
  NR2D2BWP12T U2174 ( .A1(n1362), .A2(n1361), .ZN(n1368) );
  INVD1BWP12T U2175 ( .I(n1368), .ZN(n1379) );
  TPND2D1BWP12T U2176 ( .A1(n1353), .A2(n1364), .ZN(n1371) );
  INVD1BWP12T U2177 ( .I(n1362), .ZN(n1355) );
  INVD1BWP12T U2178 ( .I(n1353), .ZN(n1354) );
  INVD1BWP12T U2179 ( .I(n1361), .ZN(n1357) );
  TPOAI22D1BWP12T U2180 ( .A1(n1357), .A2(n1377), .B1(n1370), .B2(n1356), .ZN(
        n1358) );
  AOI211XD1BWP12T U2181 ( .A1(n1375), .A2(next_pc_in[30]), .B(n1359), .C(n1358), .ZN(n1360) );
  OAI21D1BWP12T U2182 ( .A1(n1379), .A2(n1371), .B(n1360), .ZN(n2199) );
  XOR2D1BWP12T U2183 ( .A1(n1362), .A2(n1361), .Z(n1365) );
  AO222D1BWP12T U2184 ( .A1(n1365), .A2(n1364), .B1(n1375), .B2(next_pc_in[29]), .C1(pc_out[29]), .C2(n1363), .Z(n2198) );
  MUX2ND4BWP12T U2185 ( .I0(write1_in[31]), .I1(write2_in[31]), .S(n1366), 
        .ZN(n1372) );
  INVD1BWP12T U2186 ( .I(n1372), .ZN(n1378) );
  TPNR3D1BWP12T U2187 ( .A1(n1368), .A2(n1372), .A3(n1367), .ZN(n1374) );
  CKND0BWP12T U2188 ( .I(pc_out[31]), .ZN(n1369) );
  TPOAI22D1BWP12T U2189 ( .A1(n1372), .A2(n1371), .B1(n1370), .B2(n1369), .ZN(
        n1373) );
  AOI211XD1BWP12T U2190 ( .A1(n1375), .A2(next_pc_in[31]), .B(n1374), .C(n1373), .ZN(n1376) );
  OAI31D1BWP12T U2191 ( .A1(n1379), .A2(n1378), .A3(n1377), .B(n1376), .ZN(
        n2200) );
  AOI22D1BWP12T U2192 ( .A1(r1[28]), .A2(n164), .B1(n1993), .B2(r12[28]), .ZN(
        n1383) );
  AOI22D1BWP12T U2193 ( .A1(r3[28]), .A2(n1994), .B1(n168), .B2(lr[28]), .ZN(
        n1382) );
  AOI22D1BWP12T U2194 ( .A1(r8[28]), .A2(n171), .B1(n1995), .B2(n[2013]), .ZN(
        n1381) );
  AOI22D1BWP12T U2195 ( .A1(pc_out[28]), .A2(n174), .B1(n1996), .B2(r6[28]), 
        .ZN(n1380) );
  AN4XD1BWP12T U2196 ( .A1(n1383), .A2(n1382), .A3(n1381), .A4(n1380), .Z(
        n1390) );
  AOI22D1BWP12T U2197 ( .A1(tmp1[28]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[28]), .ZN(n1386) );
  AOI22D1BWP12T U2198 ( .A1(r9[28]), .A2(n152), .B1(n2002), .B2(r4[28]), .ZN(
        n1385) );
  AOI22D1BWP12T U2199 ( .A1(r11[28]), .A2(n1955), .B1(n1954), .B2(r0[28]), 
        .ZN(n1384) );
  AN3XD1BWP12T U2200 ( .A1(n1386), .A2(n1385), .A3(n1384), .Z(n1389) );
  AOI22D1BWP12T U2201 ( .A1(r5[28]), .A2(n1988), .B1(n158), .B2(r10[28]), .ZN(
        n1388) );
  AOI22D1BWP12T U2202 ( .A1(r7[28]), .A2(n1990), .B1(n1989), .B2(r2[28]), .ZN(
        n1387) );
  ND4D1BWP12T U2203 ( .A1(n1390), .A2(n1389), .A3(n1388), .A4(n1387), .ZN(
        regB_out[28]) );
  AOI22D1BWP12T U2204 ( .A1(r1[29]), .A2(n164), .B1(n1993), .B2(r12[29]), .ZN(
        n1394) );
  AOI22D1BWP12T U2205 ( .A1(r3[29]), .A2(n1994), .B1(n168), .B2(lr[29]), .ZN(
        n1393) );
  AOI22D1BWP12T U2206 ( .A1(r8[29]), .A2(n171), .B1(n1995), .B2(n[2012]), .ZN(
        n1392) );
  AOI22D1BWP12T U2207 ( .A1(pc_out[29]), .A2(n174), .B1(n1996), .B2(r6[29]), 
        .ZN(n1391) );
  AN4XD1BWP12T U2208 ( .A1(n1394), .A2(n1393), .A3(n1392), .A4(n1391), .Z(
        n1401) );
  AOI22D1BWP12T U2209 ( .A1(tmp1[29]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[29]), .ZN(n1397) );
  AOI22D1BWP12T U2210 ( .A1(r9[29]), .A2(n152), .B1(n2002), .B2(r4[29]), .ZN(
        n1396) );
  AOI22D1BWP12T U2211 ( .A1(r11[29]), .A2(n1955), .B1(n1954), .B2(r0[29]), 
        .ZN(n1395) );
  AN3XD1BWP12T U2212 ( .A1(n1397), .A2(n1396), .A3(n1395), .Z(n1400) );
  AOI22D1BWP12T U2213 ( .A1(r5[29]), .A2(n1988), .B1(n158), .B2(r10[29]), .ZN(
        n1399) );
  AOI22D1BWP12T U2214 ( .A1(r7[29]), .A2(n1990), .B1(n1989), .B2(r2[29]), .ZN(
        n1398) );
  ND4D1BWP12T U2215 ( .A1(n1401), .A2(n1400), .A3(n1399), .A4(n1398), .ZN(
        regB_out[29]) );
  AOI22D1BWP12T U2216 ( .A1(r1[30]), .A2(n164), .B1(n1993), .B2(r12[30]), .ZN(
        n1405) );
  AOI22D1BWP12T U2217 ( .A1(r3[30]), .A2(n1994), .B1(n168), .B2(lr[30]), .ZN(
        n1404) );
  AOI22D1BWP12T U2218 ( .A1(r8[30]), .A2(n171), .B1(n1995), .B2(n[2011]), .ZN(
        n1403) );
  AOI22D1BWP12T U2219 ( .A1(pc_out[30]), .A2(n174), .B1(n1996), .B2(r6[30]), 
        .ZN(n1402) );
  AN4XD1BWP12T U2220 ( .A1(n1405), .A2(n1404), .A3(n1403), .A4(n1402), .Z(
        n1412) );
  AOI22D1BWP12T U2221 ( .A1(tmp1[30]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[30]), .ZN(n1408) );
  AOI22D1BWP12T U2222 ( .A1(r9[30]), .A2(n152), .B1(n2002), .B2(r4[30]), .ZN(
        n1407) );
  AOI22D1BWP12T U2223 ( .A1(r11[30]), .A2(n1955), .B1(n1954), .B2(r0[30]), 
        .ZN(n1406) );
  AN3XD1BWP12T U2224 ( .A1(n1408), .A2(n1407), .A3(n1406), .Z(n1411) );
  AOI22D1BWP12T U2225 ( .A1(r5[30]), .A2(n1988), .B1(n158), .B2(r10[30]), .ZN(
        n1410) );
  AOI22D1BWP12T U2226 ( .A1(r7[30]), .A2(n1990), .B1(n1989), .B2(r2[30]), .ZN(
        n1409) );
  ND4D1BWP12T U2227 ( .A1(n1412), .A2(n1411), .A3(n1410), .A4(n1409), .ZN(
        regB_out[30]) );
  INVD1BWP12T U2228 ( .I(r4[29]), .ZN(n1415) );
  AOI22D1BWP12T U2229 ( .A1(n112), .A2(r12[29]), .B1(n1801), .B2(tmp1[29]), 
        .ZN(n1414) );
  AOI22D1BWP12T U2230 ( .A1(r2[29]), .A2(n1803), .B1(n1802), .B2(r1[29]), .ZN(
        n1413) );
  OA211D1BWP12T U2231 ( .A1(n1415), .A2(n1806), .B(n1414), .C(n1413), .Z(n1423) );
  AOI22D1BWP12T U2232 ( .A1(r9[29]), .A2(n1808), .B1(n120), .B2(r6[29]), .ZN(
        n1419) );
  AOI22D1BWP12T U2233 ( .A1(r8[29]), .A2(n1810), .B1(n1809), .B2(n[2012]), 
        .ZN(n1418) );
  AOI22D1BWP12T U2234 ( .A1(r5[29]), .A2(n123), .B1(n1811), .B2(r3[29]), .ZN(
        n1417) );
  AOI22D1BWP12T U2235 ( .A1(r7[29]), .A2(n126), .B1(n1812), .B2(r0[29]), .ZN(
        n1416) );
  AN4XD1BWP12T U2236 ( .A1(n1419), .A2(n1418), .A3(n1417), .A4(n1416), .Z(
        n1422) );
  AOI22D1BWP12T U2237 ( .A1(pc_out[29]), .A2(n134), .B1(n1817), .B2(r11[29]), 
        .ZN(n1421) );
  AOI22D1BWP12T U2238 ( .A1(lr[29]), .A2(n1819), .B1(n1818), .B2(r10[29]), 
        .ZN(n1420) );
  ND4D1BWP12T U2239 ( .A1(n1423), .A2(n1422), .A3(n1421), .A4(n1420), .ZN(
        regA_out[29]) );
  INVD1BWP12T U2240 ( .I(r4[27]), .ZN(n1426) );
  AOI22D1BWP12T U2241 ( .A1(n112), .A2(r12[27]), .B1(n1801), .B2(tmp1[27]), 
        .ZN(n1425) );
  AOI22D1BWP12T U2242 ( .A1(r2[27]), .A2(n1803), .B1(n1802), .B2(r1[27]), .ZN(
        n1424) );
  OA211D1BWP12T U2243 ( .A1(n1426), .A2(n1806), .B(n1425), .C(n1424), .Z(n1434) );
  AOI22D1BWP12T U2244 ( .A1(r9[27]), .A2(n1808), .B1(n120), .B2(r6[27]), .ZN(
        n1430) );
  AOI22D1BWP12T U2245 ( .A1(r8[27]), .A2(n1810), .B1(n1809), .B2(n[2014]), 
        .ZN(n1429) );
  AOI22D1BWP12T U2246 ( .A1(r5[27]), .A2(n123), .B1(n1811), .B2(r3[27]), .ZN(
        n1428) );
  AOI22D1BWP12T U2247 ( .A1(r7[27]), .A2(n126), .B1(n1812), .B2(r0[27]), .ZN(
        n1427) );
  AN4XD1BWP12T U2248 ( .A1(n1430), .A2(n1429), .A3(n1428), .A4(n1427), .Z(
        n1433) );
  AOI22D1BWP12T U2249 ( .A1(pc_out[27]), .A2(n134), .B1(n1817), .B2(r11[27]), 
        .ZN(n1432) );
  AOI22D1BWP12T U2250 ( .A1(lr[27]), .A2(n1819), .B1(n1818), .B2(r10[27]), 
        .ZN(n1431) );
  ND4D1BWP12T U2251 ( .A1(n1434), .A2(n1433), .A3(n1432), .A4(n1431), .ZN(
        regA_out[27]) );
  INVD1BWP12T U2252 ( .I(r4[31]), .ZN(n1437) );
  AOI22D1BWP12T U2253 ( .A1(n112), .A2(r12[31]), .B1(n1801), .B2(tmp1[31]), 
        .ZN(n1436) );
  AOI22D0BWP12T U2254 ( .A1(r2[31]), .A2(n1803), .B1(n1802), .B2(r1[31]), .ZN(
        n1435) );
  OA211D1BWP12T U2255 ( .A1(n1437), .A2(n1806), .B(n1436), .C(n1435), .Z(n1445) );
  AOI22D1BWP12T U2256 ( .A1(r9[31]), .A2(n1808), .B1(n120), .B2(r6[31]), .ZN(
        n1441) );
  AOI22D1BWP12T U2257 ( .A1(r8[31]), .A2(n1810), .B1(n1809), .B2(n[2010]), 
        .ZN(n1440) );
  AOI22D1BWP12T U2258 ( .A1(r5[31]), .A2(n123), .B1(n1811), .B2(r3[31]), .ZN(
        n1439) );
  AOI22D1BWP12T U2259 ( .A1(r7[31]), .A2(n126), .B1(n1812), .B2(r0[31]), .ZN(
        n1438) );
  AN4XD1BWP12T U2260 ( .A1(n1441), .A2(n1440), .A3(n1439), .A4(n1438), .Z(
        n1444) );
  AOI22D1BWP12T U2261 ( .A1(pc_out[31]), .A2(n134), .B1(n1817), .B2(r11[31]), 
        .ZN(n1443) );
  AOI22D1BWP12T U2262 ( .A1(lr[31]), .A2(n1819), .B1(n1818), .B2(r10[31]), 
        .ZN(n1442) );
  ND4D1BWP12T U2263 ( .A1(n1445), .A2(n1444), .A3(n1443), .A4(n1442), .ZN(
        regA_out[31]) );
  AOI22D1BWP12T U2264 ( .A1(tmp1[20]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[20]), .ZN(n1452) );
  AOI22D1BWP12T U2265 ( .A1(r5[20]), .A2(n1988), .B1(n158), .B2(r10[20]), .ZN(
        n1447) );
  AOI22D1BWP12T U2266 ( .A1(r7[20]), .A2(n1990), .B1(n1989), .B2(r2[20]), .ZN(
        n1446) );
  ND2D1BWP12T U2267 ( .A1(n1447), .A2(n1446), .ZN(n1451) );
  AOI22D1BWP12T U2268 ( .A1(r9[20]), .A2(n152), .B1(n2002), .B2(r4[20]), .ZN(
        n1449) );
  AOI22D1BWP12T U2269 ( .A1(r11[20]), .A2(n1571), .B1(n1954), .B2(r0[20]), 
        .ZN(n1448) );
  ND2D1BWP12T U2270 ( .A1(n1449), .A2(n1448), .ZN(n1450) );
  INR3D0BWP12T U2271 ( .A1(n1452), .B1(n1451), .B2(n1450), .ZN(n1458) );
  AOI22D1BWP12T U2272 ( .A1(r1[20]), .A2(n164), .B1(n1993), .B2(r12[20]), .ZN(
        n1456) );
  AOI22D1BWP12T U2273 ( .A1(r3[20]), .A2(n1994), .B1(n168), .B2(lr[20]), .ZN(
        n1455) );
  AOI22D1BWP12T U2274 ( .A1(r8[20]), .A2(n171), .B1(n1995), .B2(n[2021]), .ZN(
        n1454) );
  AOI22D1BWP12T U2275 ( .A1(pc_out[20]), .A2(n174), .B1(n1996), .B2(r6[20]), 
        .ZN(n1453) );
  AN4XD1BWP12T U2276 ( .A1(n1456), .A2(n1455), .A3(n1454), .A4(n1453), .Z(
        n1457) );
  ND2D1BWP12T U2277 ( .A1(n1458), .A2(n1457), .ZN(regB_out[20]) );
  INVD1BWP12T U2278 ( .I(pc_out[19]), .ZN(n1460) );
  INVD1BWP12T U2279 ( .I(r11[19]), .ZN(n1459) );
  OAI22D1BWP12T U2280 ( .A1(n1460), .A2(n1884), .B1(n1883), .B2(n1459), .ZN(
        n1469) );
  INVD1BWP12T U2281 ( .I(r10[19]), .ZN(n1461) );
  OAI22D1BWP12T U2282 ( .A1(n1462), .A2(n1888), .B1(n1887), .B2(n1461), .ZN(
        n1468) );
  AOI22D1BWP12T U2283 ( .A1(n112), .A2(r12[19]), .B1(n1801), .B2(tmp1[19]), 
        .ZN(n1463) );
  IOA21D1BWP12T U2284 ( .A1(n1891), .A2(r4[19]), .B(n1463), .ZN(n1467) );
  INVD1BWP12T U2285 ( .I(r2[19]), .ZN(n1465) );
  INVD1BWP12T U2286 ( .I(r1[19]), .ZN(n1464) );
  OAI22D1BWP12T U2287 ( .A1(n1895), .A2(n1465), .B1(n1893), .B2(n1464), .ZN(
        n1466) );
  NR4D0BWP12T U2288 ( .A1(n1469), .A2(n1468), .A3(n1467), .A4(n1466), .ZN(
        n1475) );
  AOI22D1BWP12T U2289 ( .A1(r9[19]), .A2(n1808), .B1(n120), .B2(r6[19]), .ZN(
        n1473) );
  AOI22D1BWP12T U2290 ( .A1(r8[19]), .A2(n1810), .B1(n1809), .B2(n[2022]), 
        .ZN(n1472) );
  AOI22D1BWP12T U2291 ( .A1(r5[19]), .A2(n123), .B1(n1811), .B2(r3[19]), .ZN(
        n1471) );
  AOI22D1BWP12T U2292 ( .A1(r7[19]), .A2(n126), .B1(n1812), .B2(r0[19]), .ZN(
        n1470) );
  AN4XD1BWP12T U2293 ( .A1(n1473), .A2(n1472), .A3(n1471), .A4(n1470), .Z(
        n1474) );
  ND2D1BWP12T U2294 ( .A1(n1475), .A2(n1474), .ZN(regA_out[19]) );
  AOI22D1BWP12T U2295 ( .A1(r9[18]), .A2(n1808), .B1(n120), .B2(r6[18]), .ZN(
        n1479) );
  AOI22D1BWP12T U2296 ( .A1(r8[18]), .A2(n1810), .B1(n1809), .B2(n[2023]), 
        .ZN(n1478) );
  AOI22D1BWP12T U2297 ( .A1(r5[18]), .A2(n123), .B1(n1811), .B2(r3[18]), .ZN(
        n1477) );
  AOI22D1BWP12T U2298 ( .A1(r7[18]), .A2(n126), .B1(n1812), .B2(r0[18]), .ZN(
        n1476) );
  AN4XD1BWP12T U2299 ( .A1(n1479), .A2(n1478), .A3(n1477), .A4(n1476), .Z(
        n1486) );
  AOI22D1BWP12T U2300 ( .A1(n112), .A2(r12[18]), .B1(n1684), .B2(tmp1[18]), 
        .ZN(n1482) );
  AOI22D0BWP12T U2301 ( .A1(r2[18]), .A2(n1803), .B1(n1802), .B2(r1[18]), .ZN(
        n1481) );
  CKND2D1BWP12T U2302 ( .A1(n1891), .A2(r4[18]), .ZN(n1480) );
  AN3XD1BWP12T U2303 ( .A1(n1482), .A2(n1481), .A3(n1480), .Z(n1485) );
  AOI22D1BWP12T U2304 ( .A1(pc_out[18]), .A2(n134), .B1(n1817), .B2(r11[18]), 
        .ZN(n1484) );
  AOI22D1BWP12T U2305 ( .A1(lr[18]), .A2(n1819), .B1(n1818), .B2(r10[18]), 
        .ZN(n1483) );
  ND4D1BWP12T U2306 ( .A1(n1486), .A2(n1485), .A3(n1484), .A4(n1483), .ZN(
        regA_out[18]) );
  AOI22D1BWP12T U2307 ( .A1(tmp1[18]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[18]), .ZN(n1489) );
  AOI22D1BWP12T U2308 ( .A1(r9[18]), .A2(n152), .B1(n1732), .B2(r4[18]), .ZN(
        n1488) );
  AOI22D1BWP12T U2309 ( .A1(r11[18]), .A2(n1571), .B1(n1733), .B2(r0[18]), 
        .ZN(n1487) );
  ND3D1BWP12T U2310 ( .A1(n1489), .A2(n1488), .A3(n1487), .ZN(n1493) );
  AOI22D1BWP12T U2311 ( .A1(r5[18]), .A2(n1988), .B1(n158), .B2(r10[18]), .ZN(
        n1491) );
  AOI22D1BWP12T U2312 ( .A1(r7[18]), .A2(n1990), .B1(n1989), .B2(r2[18]), .ZN(
        n1490) );
  ND2D1BWP12T U2313 ( .A1(n1491), .A2(n1490), .ZN(n1492) );
  NR2D1BWP12T U2314 ( .A1(n1493), .A2(n1492), .ZN(n1499) );
  AOI22D1BWP12T U2315 ( .A1(r1[18]), .A2(n164), .B1(n1993), .B2(r12[18]), .ZN(
        n1497) );
  AOI22D1BWP12T U2316 ( .A1(r3[18]), .A2(n1994), .B1(n168), .B2(lr[18]), .ZN(
        n1496) );
  AOI22D1BWP12T U2317 ( .A1(r8[18]), .A2(n171), .B1(n1995), .B2(n[2023]), .ZN(
        n1495) );
  AOI22D1BWP12T U2318 ( .A1(pc_out[18]), .A2(n174), .B1(n1996), .B2(r6[18]), 
        .ZN(n1494) );
  AN4XD1BWP12T U2319 ( .A1(n1497), .A2(n1496), .A3(n1495), .A4(n1494), .Z(
        n1498) );
  ND2D1BWP12T U2320 ( .A1(n1499), .A2(n1498), .ZN(regB_out[18]) );
  INVD1BWP12T U2321 ( .I(pc_out[17]), .ZN(n1501) );
  INVD1BWP12T U2322 ( .I(r11[17]), .ZN(n1500) );
  OAI22D1BWP12T U2323 ( .A1(n1501), .A2(n1884), .B1(n1883), .B2(n1500), .ZN(
        n1510) );
  INVD1BWP12T U2324 ( .I(r10[17]), .ZN(n1502) );
  OAI22D1BWP12T U2325 ( .A1(n1503), .A2(n1888), .B1(n1887), .B2(n1502), .ZN(
        n1509) );
  AOI22D1BWP12T U2326 ( .A1(n112), .A2(r12[17]), .B1(n1684), .B2(tmp1[17]), 
        .ZN(n1504) );
  IOA21D1BWP12T U2327 ( .A1(n1891), .A2(r4[17]), .B(n1504), .ZN(n1508) );
  INVD1BWP12T U2328 ( .I(r2[17]), .ZN(n1506) );
  INVD1BWP12T U2329 ( .I(r1[17]), .ZN(n1505) );
  OAI22D1BWP12T U2330 ( .A1(n1895), .A2(n1506), .B1(n1893), .B2(n1505), .ZN(
        n1507) );
  NR4D0BWP12T U2331 ( .A1(n1510), .A2(n1509), .A3(n1508), .A4(n1507), .ZN(
        n1516) );
  AOI22D1BWP12T U2332 ( .A1(r9[17]), .A2(n1808), .B1(n120), .B2(r6[17]), .ZN(
        n1514) );
  AOI22D1BWP12T U2333 ( .A1(r8[17]), .A2(n1810), .B1(n1809), .B2(n[2024]), 
        .ZN(n1513) );
  AOI22D1BWP12T U2334 ( .A1(r5[17]), .A2(n123), .B1(n1811), .B2(r3[17]), .ZN(
        n1512) );
  AOI22D1BWP12T U2335 ( .A1(r7[17]), .A2(n126), .B1(n1812), .B2(r0[17]), .ZN(
        n1511) );
  AN4XD1BWP12T U2336 ( .A1(n1514), .A2(n1513), .A3(n1512), .A4(n1511), .Z(
        n1515) );
  ND2D1BWP12T U2337 ( .A1(n1516), .A2(n1515), .ZN(regA_out[17]) );
  AOI22D1BWP12T U2338 ( .A1(tmp1[17]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[17]), .ZN(n1519) );
  AOI22D1BWP12T U2339 ( .A1(r9[17]), .A2(n152), .B1(n1732), .B2(r4[17]), .ZN(
        n1518) );
  AOI22D1BWP12T U2340 ( .A1(r11[17]), .A2(n1571), .B1(n1733), .B2(r0[17]), 
        .ZN(n1517) );
  ND3D1BWP12T U2341 ( .A1(n1519), .A2(n1518), .A3(n1517), .ZN(n1523) );
  AOI22D1BWP12T U2342 ( .A1(r5[17]), .A2(n1988), .B1(n158), .B2(r10[17]), .ZN(
        n1521) );
  AOI22D1BWP12T U2343 ( .A1(r7[17]), .A2(n1990), .B1(n1989), .B2(r2[17]), .ZN(
        n1520) );
  ND2D1BWP12T U2344 ( .A1(n1521), .A2(n1520), .ZN(n1522) );
  NR2D1BWP12T U2345 ( .A1(n1523), .A2(n1522), .ZN(n1529) );
  AOI22D1BWP12T U2346 ( .A1(r1[17]), .A2(n164), .B1(n1993), .B2(r12[17]), .ZN(
        n1527) );
  AOI22D1BWP12T U2347 ( .A1(r3[17]), .A2(n1994), .B1(n168), .B2(lr[17]), .ZN(
        n1526) );
  AOI22D1BWP12T U2348 ( .A1(r8[17]), .A2(n171), .B1(n1995), .B2(n[2024]), .ZN(
        n1525) );
  AOI22D1BWP12T U2349 ( .A1(pc_out[17]), .A2(n174), .B1(n1996), .B2(r6[17]), 
        .ZN(n1524) );
  AN4XD1BWP12T U2350 ( .A1(n1527), .A2(n1526), .A3(n1525), .A4(n1524), .Z(
        n1528) );
  ND2D1BWP12T U2351 ( .A1(n1529), .A2(n1528), .ZN(regB_out[17]) );
  AOI22D1BWP12T U2352 ( .A1(r9[16]), .A2(n1808), .B1(n120), .B2(r6[16]), .ZN(
        n1533) );
  AOI22D1BWP12T U2353 ( .A1(r8[16]), .A2(n1810), .B1(n1809), .B2(n[2025]), 
        .ZN(n1532) );
  AOI22D1BWP12T U2354 ( .A1(r5[16]), .A2(n123), .B1(n1811), .B2(r3[16]), .ZN(
        n1531) );
  AOI22D1BWP12T U2355 ( .A1(r7[16]), .A2(n126), .B1(n1812), .B2(r0[16]), .ZN(
        n1530) );
  AN4XD1BWP12T U2356 ( .A1(n1533), .A2(n1532), .A3(n1531), .A4(n1530), .Z(
        n1540) );
  AOI22D1BWP12T U2357 ( .A1(n112), .A2(r12[16]), .B1(n1684), .B2(tmp1[16]), 
        .ZN(n1536) );
  AOI22D1BWP12T U2358 ( .A1(r2[16]), .A2(n1803), .B1(n1802), .B2(r1[16]), .ZN(
        n1535) );
  CKND2D1BWP12T U2359 ( .A1(n1891), .A2(r4[16]), .ZN(n1534) );
  AN3XD1BWP12T U2360 ( .A1(n1536), .A2(n1535), .A3(n1534), .Z(n1539) );
  AOI22D1BWP12T U2361 ( .A1(pc_out[16]), .A2(n134), .B1(n1817), .B2(r11[16]), 
        .ZN(n1538) );
  AOI22D1BWP12T U2362 ( .A1(lr[16]), .A2(n1819), .B1(n1818), .B2(r10[16]), 
        .ZN(n1537) );
  ND4D1BWP12T U2363 ( .A1(n1540), .A2(n1539), .A3(n1538), .A4(n1537), .ZN(
        regA_out[16]) );
  AOI22D1BWP12T U2364 ( .A1(tmp1[16]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[16]), .ZN(n1543) );
  AOI22D1BWP12T U2365 ( .A1(r9[16]), .A2(n152), .B1(n1732), .B2(r4[16]), .ZN(
        n1542) );
  AOI22D1BWP12T U2366 ( .A1(r11[16]), .A2(n1571), .B1(n1733), .B2(r0[16]), 
        .ZN(n1541) );
  ND3D1BWP12T U2367 ( .A1(n1543), .A2(n1542), .A3(n1541), .ZN(n1547) );
  AOI22D1BWP12T U2368 ( .A1(r5[16]), .A2(n1988), .B1(n158), .B2(r10[16]), .ZN(
        n1545) );
  AOI22D1BWP12T U2369 ( .A1(r7[16]), .A2(n1990), .B1(n1989), .B2(r2[16]), .ZN(
        n1544) );
  ND2D1BWP12T U2370 ( .A1(n1545), .A2(n1544), .ZN(n1546) );
  NR2D1BWP12T U2371 ( .A1(n1547), .A2(n1546), .ZN(n1553) );
  AOI22D1BWP12T U2372 ( .A1(r1[16]), .A2(n164), .B1(n1993), .B2(r12[16]), .ZN(
        n1551) );
  AOI22D1BWP12T U2373 ( .A1(r3[16]), .A2(n1994), .B1(n168), .B2(lr[16]), .ZN(
        n1550) );
  AOI22D1BWP12T U2374 ( .A1(r8[16]), .A2(n171), .B1(n1995), .B2(n[2025]), .ZN(
        n1549) );
  AOI22D1BWP12T U2375 ( .A1(pc_out[16]), .A2(n174), .B1(n1996), .B2(r6[16]), 
        .ZN(n1548) );
  AN4XD1BWP12T U2376 ( .A1(n1551), .A2(n1550), .A3(n1549), .A4(n1548), .Z(
        n1552) );
  ND2D1BWP12T U2377 ( .A1(n1553), .A2(n1552), .ZN(regB_out[16]) );
  INVD0BWP12T U2378 ( .I(pc_out[15]), .ZN(n1555) );
  INVD1BWP12T U2379 ( .I(r11[15]), .ZN(n1554) );
  OAI22D1BWP12T U2380 ( .A1(n1555), .A2(n1884), .B1(n1883), .B2(n1554), .ZN(
        n1564) );
  INVD1BWP12T U2381 ( .I(r10[15]), .ZN(n1556) );
  OAI22D1BWP12T U2382 ( .A1(n1557), .A2(n1888), .B1(n1887), .B2(n1556), .ZN(
        n1563) );
  AOI22D1BWP12T U2383 ( .A1(n112), .A2(r12[15]), .B1(n1684), .B2(tmp1[15]), 
        .ZN(n1558) );
  IOA21D1BWP12T U2384 ( .A1(n1891), .A2(r4[15]), .B(n1558), .ZN(n1562) );
  INVD1BWP12T U2385 ( .I(r2[15]), .ZN(n1560) );
  INVD1BWP12T U2386 ( .I(r1[15]), .ZN(n1559) );
  OAI22D1BWP12T U2387 ( .A1(n1895), .A2(n1560), .B1(n1893), .B2(n1559), .ZN(
        n1561) );
  NR4D0BWP12T U2388 ( .A1(n1564), .A2(n1563), .A3(n1562), .A4(n1561), .ZN(
        n1570) );
  AOI22D1BWP12T U2389 ( .A1(r9[15]), .A2(n1808), .B1(n120), .B2(r6[15]), .ZN(
        n1568) );
  AOI22D1BWP12T U2390 ( .A1(r8[15]), .A2(n1810), .B1(n1809), .B2(n[2026]), 
        .ZN(n1567) );
  AOI22D1BWP12T U2391 ( .A1(r5[15]), .A2(n123), .B1(n1811), .B2(r3[15]), .ZN(
        n1566) );
  AOI22D1BWP12T U2392 ( .A1(r7[15]), .A2(n126), .B1(n1812), .B2(r0[15]), .ZN(
        n1565) );
  AN4XD1BWP12T U2393 ( .A1(n1568), .A2(n1567), .A3(n1566), .A4(n1565), .Z(
        n1569) );
  ND2D1BWP12T U2394 ( .A1(n1570), .A2(n1569), .ZN(regA_out[15]) );
  AOI22D1BWP12T U2395 ( .A1(tmp1[15]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[15]), .ZN(n1574) );
  AOI22D1BWP12T U2396 ( .A1(r9[15]), .A2(n152), .B1(n1732), .B2(r4[15]), .ZN(
        n1573) );
  AOI22D1BWP12T U2397 ( .A1(r11[15]), .A2(n1571), .B1(n1733), .B2(r0[15]), 
        .ZN(n1572) );
  ND3D1BWP12T U2398 ( .A1(n1574), .A2(n1573), .A3(n1572), .ZN(n1578) );
  AOI22D1BWP12T U2399 ( .A1(r5[15]), .A2(n1988), .B1(n158), .B2(r10[15]), .ZN(
        n1576) );
  AOI22D1BWP12T U2400 ( .A1(r7[15]), .A2(n1990), .B1(n1989), .B2(r2[15]), .ZN(
        n1575) );
  ND2D1BWP12T U2401 ( .A1(n1576), .A2(n1575), .ZN(n1577) );
  NR2D1BWP12T U2402 ( .A1(n1578), .A2(n1577), .ZN(n1584) );
  AOI22D1BWP12T U2403 ( .A1(r1[15]), .A2(n164), .B1(n1993), .B2(r12[15]), .ZN(
        n1582) );
  AOI22D1BWP12T U2404 ( .A1(r3[15]), .A2(n1994), .B1(n168), .B2(lr[15]), .ZN(
        n1581) );
  AOI22D1BWP12T U2405 ( .A1(r8[15]), .A2(n171), .B1(n1995), .B2(n[2026]), .ZN(
        n1580) );
  AOI22D1BWP12T U2406 ( .A1(pc_out[15]), .A2(n174), .B1(n1996), .B2(r6[15]), 
        .ZN(n1579) );
  AN4XD1BWP12T U2407 ( .A1(n1582), .A2(n1581), .A3(n1580), .A4(n1579), .Z(
        n1583) );
  ND2D1BWP12T U2408 ( .A1(n1584), .A2(n1583), .ZN(regB_out[15]) );
  INVD0BWP12T U2409 ( .I(pc_out[13]), .ZN(n1586) );
  INVD1BWP12T U2410 ( .I(r11[13]), .ZN(n1585) );
  OAI22D1BWP12T U2411 ( .A1(n1586), .A2(n1884), .B1(n1883), .B2(n1585), .ZN(
        n1595) );
  INVD1BWP12T U2412 ( .I(r10[13]), .ZN(n1587) );
  OAI22D1BWP12T U2413 ( .A1(n1588), .A2(n1888), .B1(n1887), .B2(n1587), .ZN(
        n1594) );
  AOI22D1BWP12T U2414 ( .A1(n112), .A2(r12[13]), .B1(n1684), .B2(tmp1[13]), 
        .ZN(n1589) );
  IOA21D1BWP12T U2415 ( .A1(n1891), .A2(r4[13]), .B(n1589), .ZN(n1593) );
  INVD1BWP12T U2416 ( .I(r2[13]), .ZN(n1591) );
  INVD1BWP12T U2417 ( .I(r1[13]), .ZN(n1590) );
  OAI22D1BWP12T U2418 ( .A1(n1895), .A2(n1591), .B1(n1893), .B2(n1590), .ZN(
        n1592) );
  NR4D0BWP12T U2419 ( .A1(n1595), .A2(n1594), .A3(n1593), .A4(n1592), .ZN(
        n1601) );
  AOI22D1BWP12T U2420 ( .A1(r9[13]), .A2(n1808), .B1(n120), .B2(r6[13]), .ZN(
        n1599) );
  AOI22D1BWP12T U2421 ( .A1(r8[13]), .A2(n1810), .B1(n1809), .B2(n[2028]), 
        .ZN(n1598) );
  AOI22D1BWP12T U2422 ( .A1(r5[13]), .A2(n123), .B1(n1811), .B2(r3[13]), .ZN(
        n1597) );
  AOI22D1BWP12T U2423 ( .A1(r7[13]), .A2(n126), .B1(n1812), .B2(r0[13]), .ZN(
        n1596) );
  AN4XD1BWP12T U2424 ( .A1(n1599), .A2(n1598), .A3(n1597), .A4(n1596), .Z(
        n1600) );
  ND2D1BWP12T U2425 ( .A1(n1601), .A2(n1600), .ZN(regA_out[13]) );
  AOI22D1BWP12T U2426 ( .A1(tmp1[13]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[13]), .ZN(n1604) );
  AOI22D1BWP12T U2427 ( .A1(r9[13]), .A2(n152), .B1(n1732), .B2(r4[13]), .ZN(
        n1603) );
  AOI22D1BWP12T U2428 ( .A1(r11[13]), .A2(n2003), .B1(n1733), .B2(r0[13]), 
        .ZN(n1602) );
  ND3D1BWP12T U2429 ( .A1(n1604), .A2(n1603), .A3(n1602), .ZN(n1614) );
  AOI22D1BWP12T U2430 ( .A1(r1[13]), .A2(n164), .B1(n1993), .B2(r12[13]), .ZN(
        n1606) );
  AOI22D1BWP12T U2431 ( .A1(r8[13]), .A2(n171), .B1(n1995), .B2(n[2028]), .ZN(
        n1605) );
  ND2D1BWP12T U2432 ( .A1(n1606), .A2(n1605), .ZN(n1613) );
  AOI22D1BWP12T U2433 ( .A1(r3[13]), .A2(n1994), .B1(n168), .B2(lr[13]), .ZN(
        n1608) );
  AOI22D1BWP12T U2434 ( .A1(pc_out[13]), .A2(n174), .B1(n1996), .B2(r6[13]), 
        .ZN(n1607) );
  ND2D1BWP12T U2435 ( .A1(n1608), .A2(n1607), .ZN(n1612) );
  AOI22D1BWP12T U2436 ( .A1(r5[13]), .A2(n1988), .B1(n158), .B2(r10[13]), .ZN(
        n1610) );
  AOI22D1BWP12T U2437 ( .A1(r7[13]), .A2(n1990), .B1(n1989), .B2(r2[13]), .ZN(
        n1609) );
  ND2D1BWP12T U2438 ( .A1(n1610), .A2(n1609), .ZN(n1611) );
  NR4D0BWP12T U2439 ( .A1(n1614), .A2(n1613), .A3(n1612), .A4(n1611), .ZN(
        n1615) );
  INVD1BWP12T U2440 ( .I(n1615), .ZN(regB_out[13]) );
  OAI22D1BWP12T U2441 ( .A1(n1648), .A2(n1884), .B1(n1883), .B2(n1616), .ZN(
        n1621) );
  OAI22D1BWP12T U2442 ( .A1(n1643), .A2(n1888), .B1(n1887), .B2(n1633), .ZN(
        n1620) );
  AOI22D1BWP12T U2443 ( .A1(n112), .A2(r12[12]), .B1(n1684), .B2(tmp1[12]), 
        .ZN(n1617) );
  IOA21D1BWP12T U2444 ( .A1(n1891), .A2(r4[12]), .B(n1617), .ZN(n1619) );
  OAI22D1BWP12T U2445 ( .A1(n1895), .A2(n1635), .B1(n1893), .B2(n1642), .ZN(
        n1618) );
  NR4D0BWP12T U2446 ( .A1(n1621), .A2(n1620), .A3(n1619), .A4(n1618), .ZN(
        n1629) );
  OAI22D1BWP12T U2447 ( .A1(n1903), .A2(n1622), .B1(n1901), .B2(n1647), .ZN(
        n1627) );
  INVD1BWP12T U2448 ( .I(n[2029]), .ZN(n1645) );
  OAI22D1BWP12T U2449 ( .A1(n1907), .A2(n1646), .B1(n1905), .B2(n1645), .ZN(
        n1626) );
  OAI22D1BWP12T U2450 ( .A1(n1634), .A2(n1910), .B1(n1909), .B2(n1644), .ZN(
        n1625) );
  OAI22D1BWP12T U2451 ( .A1(n1915), .A2(n1636), .B1(n1913), .B2(n1623), .ZN(
        n1624) );
  NR4D0BWP12T U2452 ( .A1(n1627), .A2(n1626), .A3(n1625), .A4(n1624), .ZN(
        n1628) );
  ND2D1BWP12T U2453 ( .A1(n1629), .A2(n1628), .ZN(regA_out[12]) );
  INVD1BWP12T U2454 ( .I(tmp1[12]), .ZN(n1630) );
  MOAI22D0BWP12T U2455 ( .A1(n1630), .A2(n1951), .B1(n150), .B2(
        immediate2_in[12]), .ZN(n1640) );
  AOI22D1BWP12T U2456 ( .A1(r9[12]), .A2(n152), .B1(n1732), .B2(r4[12]), .ZN(
        n1632) );
  AOI22D1BWP12T U2457 ( .A1(r11[12]), .A2(n1955), .B1(n1733), .B2(r0[12]), 
        .ZN(n1631) );
  ND2D1BWP12T U2458 ( .A1(n1632), .A2(n1631), .ZN(n1639) );
  OAI22D1BWP12T U2459 ( .A1(n1634), .A2(n1949), .B1(n1948), .B2(n1633), .ZN(
        n1638) );
  OAI22D1BWP12T U2460 ( .A1(n1961), .A2(n1636), .B1(n1959), .B2(n1635), .ZN(
        n1637) );
  NR4D0BWP12T U2461 ( .A1(n1640), .A2(n1639), .A3(n1638), .A4(n1637), .ZN(
        n1654) );
  OAI22D1BWP12T U2462 ( .A1(n1642), .A2(n1968), .B1(n1967), .B2(n1641), .ZN(
        n1652) );
  OAI22D1BWP12T U2463 ( .A1(n1644), .A2(n1972), .B1(n1971), .B2(n1643), .ZN(
        n1651) );
  OAI22D1BWP12T U2464 ( .A1(n1977), .A2(n1646), .B1(n1975), .B2(n1645), .ZN(
        n1650) );
  OAI22D1BWP12T U2465 ( .A1(n1981), .A2(n1648), .B1(n1979), .B2(n1647), .ZN(
        n1649) );
  NR4D0BWP12T U2466 ( .A1(n1652), .A2(n1651), .A3(n1650), .A4(n1649), .ZN(
        n1653) );
  ND2D1BWP12T U2467 ( .A1(n1654), .A2(n1653), .ZN(regB_out[12]) );
  OAI22D1BWP12T U2468 ( .A1(n1656), .A2(n1884), .B1(n1883), .B2(n1655), .ZN(
        n1665) );
  OAI22D1BWP12T U2469 ( .A1(n1658), .A2(n1888), .B1(n1887), .B2(n1657), .ZN(
        n1664) );
  AOI22D1BWP12T U2470 ( .A1(n112), .A2(r12[10]), .B1(n1684), .B2(tmp1[10]), 
        .ZN(n1659) );
  IOA21D1BWP12T U2471 ( .A1(n1891), .A2(r4[10]), .B(n1659), .ZN(n1663) );
  OAI22D1BWP12T U2472 ( .A1(n1895), .A2(n1661), .B1(n1893), .B2(n1660), .ZN(
        n1662) );
  NR4D0BWP12T U2473 ( .A1(n1665), .A2(n1664), .A3(n1663), .A4(n1662), .ZN(
        n1679) );
  OAI22D1BWP12T U2474 ( .A1(n1903), .A2(n1667), .B1(n1901), .B2(n1666), .ZN(
        n1677) );
  OAI22D1BWP12T U2475 ( .A1(n1907), .A2(n1669), .B1(n1905), .B2(n1668), .ZN(
        n1676) );
  OAI22D1BWP12T U2476 ( .A1(n1671), .A2(n1910), .B1(n1909), .B2(n1670), .ZN(
        n1675) );
  OAI22D1BWP12T U2477 ( .A1(n1915), .A2(n1673), .B1(n1913), .B2(n1672), .ZN(
        n1674) );
  NR4D0BWP12T U2478 ( .A1(n1677), .A2(n1676), .A3(n1675), .A4(n1674), .ZN(
        n1678) );
  ND2D1BWP12T U2479 ( .A1(n1679), .A2(n1678), .ZN(regA_out[10]) );
  OAI22D1BWP12T U2480 ( .A1(n1681), .A2(n1884), .B1(n1883), .B2(n1680), .ZN(
        n1691) );
  OAI22D1BWP12T U2481 ( .A1(n1683), .A2(n1888), .B1(n1887), .B2(n1682), .ZN(
        n1690) );
  AOI22D1BWP12T U2482 ( .A1(n112), .A2(r12[8]), .B1(n1684), .B2(tmp1[8]), .ZN(
        n1685) );
  IOA21D1BWP12T U2483 ( .A1(n1891), .A2(r4[8]), .B(n1685), .ZN(n1689) );
  OAI22D1BWP12T U2484 ( .A1(n1895), .A2(n1687), .B1(n1893), .B2(n1686), .ZN(
        n1688) );
  NR4D0BWP12T U2485 ( .A1(n1691), .A2(n1690), .A3(n1689), .A4(n1688), .ZN(
        n1705) );
  OAI22D1BWP12T U2486 ( .A1(n1903), .A2(n1693), .B1(n1901), .B2(n1692), .ZN(
        n1703) );
  OAI22D1BWP12T U2487 ( .A1(n1907), .A2(n1695), .B1(n1905), .B2(n1694), .ZN(
        n1702) );
  OAI22D1BWP12T U2488 ( .A1(n1697), .A2(n1910), .B1(n1909), .B2(n1696), .ZN(
        n1701) );
  OAI22D1BWP12T U2489 ( .A1(n1915), .A2(n1699), .B1(n1913), .B2(n1698), .ZN(
        n1700) );
  NR4D0BWP12T U2490 ( .A1(n1703), .A2(n1702), .A3(n1701), .A4(n1700), .ZN(
        n1704) );
  ND2D1BWP12T U2491 ( .A1(n1705), .A2(n1704), .ZN(regA_out[8]) );
  INVD0BWP12T U2492 ( .I(tmp1[7]), .ZN(n1706) );
  MOAI22D0BWP12T U2493 ( .A1(n1706), .A2(n1951), .B1(n150), .B2(
        immediate2_in[7]), .ZN(n1716) );
  AOI22D1BWP12T U2494 ( .A1(r9[7]), .A2(n152), .B1(n1732), .B2(r4[7]), .ZN(
        n1708) );
  AOI22D1BWP12T U2495 ( .A1(r11[7]), .A2(n2003), .B1(n1733), .B2(r0[7]), .ZN(
        n1707) );
  ND2D1BWP12T U2496 ( .A1(n1708), .A2(n1707), .ZN(n1715) );
  OAI22D1BWP12T U2497 ( .A1(n1710), .A2(n1949), .B1(n1948), .B2(n1709), .ZN(
        n1714) );
  OAI22D1BWP12T U2498 ( .A1(n1961), .A2(n1712), .B1(n1959), .B2(n1711), .ZN(
        n1713) );
  NR4D0BWP12T U2499 ( .A1(n1716), .A2(n1715), .A3(n1714), .A4(n1713), .ZN(
        n1730) );
  OAI22D1BWP12T U2500 ( .A1(n1718), .A2(n1968), .B1(n1967), .B2(n1717), .ZN(
        n1728) );
  OAI22D1BWP12T U2501 ( .A1(n1720), .A2(n1972), .B1(n1971), .B2(n1719), .ZN(
        n1727) );
  OAI22D1BWP12T U2502 ( .A1(n1977), .A2(n1722), .B1(n1975), .B2(n1721), .ZN(
        n1726) );
  OAI22D1BWP12T U2503 ( .A1(n1981), .A2(n1724), .B1(n1979), .B2(n1723), .ZN(
        n1725) );
  NR4D0BWP12T U2504 ( .A1(n1728), .A2(n1727), .A3(n1726), .A4(n1725), .ZN(
        n1729) );
  ND2D1BWP12T U2505 ( .A1(n1730), .A2(n1729), .ZN(regB_out[7]) );
  INVD1BWP12T U2506 ( .I(tmp1[6]), .ZN(n1731) );
  MOAI22D0BWP12T U2507 ( .A1(n1731), .A2(n1951), .B1(n150), .B2(
        immediate2_in[6]), .ZN(n1743) );
  AOI22D1BWP12T U2508 ( .A1(r9[6]), .A2(n152), .B1(n1732), .B2(r4[6]), .ZN(
        n1735) );
  AOI22D1BWP12T U2509 ( .A1(r11[6]), .A2(n1955), .B1(n1733), .B2(r0[6]), .ZN(
        n1734) );
  ND2D1BWP12T U2510 ( .A1(n1735), .A2(n1734), .ZN(n1742) );
  OAI22D1BWP12T U2511 ( .A1(n1737), .A2(n1949), .B1(n1948), .B2(n1736), .ZN(
        n1741) );
  OAI22D1BWP12T U2512 ( .A1(n1961), .A2(n1739), .B1(n1959), .B2(n1738), .ZN(
        n1740) );
  NR4D0BWP12T U2513 ( .A1(n1743), .A2(n1742), .A3(n1741), .A4(n1740), .ZN(
        n1757) );
  OAI22D1BWP12T U2514 ( .A1(n1745), .A2(n1968), .B1(n1967), .B2(n1744), .ZN(
        n1755) );
  OAI22D1BWP12T U2515 ( .A1(n1747), .A2(n1972), .B1(n1971), .B2(n1746), .ZN(
        n1754) );
  OAI22D1BWP12T U2516 ( .A1(n1977), .A2(n1749), .B1(n1975), .B2(n1748), .ZN(
        n1753) );
  OAI22D1BWP12T U2517 ( .A1(n1981), .A2(n1751), .B1(n1979), .B2(n1750), .ZN(
        n1752) );
  NR4D0BWP12T U2518 ( .A1(n1755), .A2(n1754), .A3(n1753), .A4(n1752), .ZN(
        n1756) );
  ND2D1BWP12T U2519 ( .A1(n1757), .A2(n1756), .ZN(regB_out[6]) );
  INVD1BWP12T U2520 ( .I(lr[21]), .ZN(n1760) );
  AOI22D1BWP12T U2521 ( .A1(pc_out[21]), .A2(n134), .B1(n1817), .B2(r11[21]), 
        .ZN(n1759) );
  CKND2D1BWP12T U2522 ( .A1(n1818), .A2(r10[21]), .ZN(n1758) );
  OA211D1BWP12T U2523 ( .A1(n1888), .A2(n1760), .B(n1759), .C(n1758), .Z(n1770) );
  INVD1BWP12T U2524 ( .I(r4[21]), .ZN(n1763) );
  AOI22D1BWP12T U2525 ( .A1(n112), .A2(r12[21]), .B1(n1801), .B2(tmp1[21]), 
        .ZN(n1762) );
  AOI22D1BWP12T U2526 ( .A1(r2[21]), .A2(n1803), .B1(n1802), .B2(r1[21]), .ZN(
        n1761) );
  OA211D1BWP12T U2527 ( .A1(n1763), .A2(n1806), .B(n1762), .C(n1761), .Z(n1769) );
  AOI22D1BWP12T U2528 ( .A1(r9[21]), .A2(n1808), .B1(n120), .B2(r6[21]), .ZN(
        n1767) );
  AOI22D1BWP12T U2529 ( .A1(r8[21]), .A2(n1810), .B1(n1809), .B2(n[2020]), 
        .ZN(n1766) );
  AOI22D1BWP12T U2530 ( .A1(r5[21]), .A2(n123), .B1(n1811), .B2(r3[21]), .ZN(
        n1765) );
  AOI22D1BWP12T U2531 ( .A1(r7[21]), .A2(n126), .B1(n1812), .B2(r0[21]), .ZN(
        n1764) );
  AN4XD1BWP12T U2532 ( .A1(n1767), .A2(n1766), .A3(n1765), .A4(n1764), .Z(
        n1768) );
  ND3D1BWP12T U2533 ( .A1(n1770), .A2(n1769), .A3(n1768), .ZN(regA_out[21]) );
  INVD1BWP12T U2534 ( .I(r4[22]), .ZN(n1773) );
  AOI22D1BWP12T U2535 ( .A1(n112), .A2(r12[22]), .B1(n1801), .B2(tmp1[22]), 
        .ZN(n1772) );
  AOI22D1BWP12T U2536 ( .A1(r2[22]), .A2(n1803), .B1(n1802), .B2(r1[22]), .ZN(
        n1771) );
  OA211D1BWP12T U2537 ( .A1(n1773), .A2(n1806), .B(n1772), .C(n1771), .Z(n1781) );
  AOI22D1BWP12T U2538 ( .A1(r9[22]), .A2(n1808), .B1(n120), .B2(r6[22]), .ZN(
        n1777) );
  AOI22D1BWP12T U2539 ( .A1(r8[22]), .A2(n1810), .B1(n1809), .B2(n[2019]), 
        .ZN(n1776) );
  AOI22D1BWP12T U2540 ( .A1(r5[22]), .A2(n123), .B1(n1811), .B2(r3[22]), .ZN(
        n1775) );
  AOI22D1BWP12T U2541 ( .A1(r7[22]), .A2(n126), .B1(n1812), .B2(r0[22]), .ZN(
        n1774) );
  AN4XD1BWP12T U2542 ( .A1(n1777), .A2(n1776), .A3(n1775), .A4(n1774), .Z(
        n1780) );
  AOI22D1BWP12T U2543 ( .A1(pc_out[22]), .A2(n134), .B1(n1817), .B2(r11[22]), 
        .ZN(n1779) );
  AOI22D1BWP12T U2544 ( .A1(lr[22]), .A2(n1819), .B1(n1818), .B2(r10[22]), 
        .ZN(n1778) );
  ND4D1BWP12T U2545 ( .A1(n1781), .A2(n1780), .A3(n1779), .A4(n1778), .ZN(
        regA_out[22]) );
  INVD1BWP12T U2546 ( .I(r4[23]), .ZN(n1784) );
  AOI22D1BWP12T U2547 ( .A1(n112), .A2(r12[23]), .B1(n1801), .B2(tmp1[23]), 
        .ZN(n1783) );
  AOI22D1BWP12T U2548 ( .A1(r2[23]), .A2(n1803), .B1(n1802), .B2(r1[23]), .ZN(
        n1782) );
  AOI22D1BWP12T U2549 ( .A1(r9[23]), .A2(n1808), .B1(n120), .B2(r6[23]), .ZN(
        n1788) );
  AOI22D1BWP12T U2550 ( .A1(r8[23]), .A2(n1810), .B1(n1809), .B2(n[2018]), 
        .ZN(n1787) );
  AOI22D1BWP12T U2551 ( .A1(r5[23]), .A2(n123), .B1(n1811), .B2(r3[23]), .ZN(
        n1786) );
  AOI22D1BWP12T U2552 ( .A1(r7[23]), .A2(n126), .B1(n1812), .B2(r0[23]), .ZN(
        n1785) );
  AN4XD1BWP12T U2553 ( .A1(n1788), .A2(n1787), .A3(n1786), .A4(n1785), .Z(
        n1789) );
  INVD1BWP12T U2554 ( .I(r4[24]), .ZN(n1792) );
  AOI22D1BWP12T U2555 ( .A1(n112), .A2(r12[24]), .B1(n1801), .B2(tmp1[24]), 
        .ZN(n1791) );
  AOI22D1BWP12T U2556 ( .A1(r2[24]), .A2(n1803), .B1(n1802), .B2(r1[24]), .ZN(
        n1790) );
  OA211D1BWP12T U2557 ( .A1(n1792), .A2(n1806), .B(n1791), .C(n1790), .Z(n1800) );
  AOI22D1BWP12T U2558 ( .A1(r9[24]), .A2(n1808), .B1(n120), .B2(r6[24]), .ZN(
        n1796) );
  AOI22D1BWP12T U2559 ( .A1(r8[24]), .A2(n1810), .B1(n1809), .B2(n[2017]), 
        .ZN(n1795) );
  AOI22D1BWP12T U2560 ( .A1(r5[24]), .A2(n123), .B1(n1811), .B2(r3[24]), .ZN(
        n1794) );
  AOI22D1BWP12T U2561 ( .A1(r7[24]), .A2(n126), .B1(n1812), .B2(r0[24]), .ZN(
        n1793) );
  AN4XD1BWP12T U2562 ( .A1(n1796), .A2(n1795), .A3(n1794), .A4(n1793), .Z(
        n1799) );
  AOI22D1BWP12T U2563 ( .A1(pc_out[24]), .A2(n134), .B1(n1817), .B2(r11[24]), 
        .ZN(n1798) );
  AOI22D1BWP12T U2564 ( .A1(lr[24]), .A2(n1819), .B1(n1818), .B2(r10[24]), 
        .ZN(n1797) );
  ND4D1BWP12T U2565 ( .A1(n1800), .A2(n1799), .A3(n1798), .A4(n1797), .ZN(
        regA_out[24]) );
  INVD1BWP12T U2566 ( .I(r4[25]), .ZN(n1807) );
  AOI22D1BWP12T U2567 ( .A1(n112), .A2(r12[25]), .B1(n1801), .B2(tmp1[25]), 
        .ZN(n1805) );
  AOI22D1BWP12T U2568 ( .A1(r2[25]), .A2(n1803), .B1(n1802), .B2(r1[25]), .ZN(
        n1804) );
  AOI22D1BWP12T U2569 ( .A1(r9[25]), .A2(n1808), .B1(n120), .B2(r6[25]), .ZN(
        n1816) );
  AOI22D1BWP12T U2570 ( .A1(r8[25]), .A2(n1810), .B1(n1809), .B2(n[2016]), 
        .ZN(n1815) );
  AOI22D1BWP12T U2571 ( .A1(r5[25]), .A2(n123), .B1(n1811), .B2(r3[25]), .ZN(
        n1814) );
  AOI22D1BWP12T U2572 ( .A1(r7[25]), .A2(n126), .B1(n1812), .B2(r0[25]), .ZN(
        n1813) );
  AN4XD1BWP12T U2573 ( .A1(n1816), .A2(n1815), .A3(n1814), .A4(n1813), .Z(
        n1820) );
  INVD0BWP12T U2574 ( .I(tmp1[5]), .ZN(n1821) );
  MOAI22D0BWP12T U2575 ( .A1(n1821), .A2(n1951), .B1(n150), .B2(
        immediate2_in[5]), .ZN(n1831) );
  AOI22D1BWP12T U2576 ( .A1(r9[5]), .A2(n152), .B1(n1953), .B2(r4[5]), .ZN(
        n1823) );
  AOI22D1BWP12T U2577 ( .A1(r11[5]), .A2(n1955), .B1(n1954), .B2(r0[5]), .ZN(
        n1822) );
  ND2D1BWP12T U2578 ( .A1(n1823), .A2(n1822), .ZN(n1830) );
  OAI22D1BWP12T U2579 ( .A1(n1825), .A2(n1949), .B1(n1948), .B2(n1824), .ZN(
        n1829) );
  OAI22D1BWP12T U2580 ( .A1(n1961), .A2(n1827), .B1(n1959), .B2(n1826), .ZN(
        n1828) );
  NR4D0BWP12T U2581 ( .A1(n1831), .A2(n1830), .A3(n1829), .A4(n1828), .ZN(
        n1845) );
  OAI22D1BWP12T U2582 ( .A1(n1833), .A2(n1968), .B1(n1967), .B2(n1832), .ZN(
        n1843) );
  OAI22D1BWP12T U2583 ( .A1(n1835), .A2(n1972), .B1(n1971), .B2(n1834), .ZN(
        n1842) );
  OAI22D1BWP12T U2584 ( .A1(n1977), .A2(n1837), .B1(n1975), .B2(n1836), .ZN(
        n1841) );
  OAI22D1BWP12T U2585 ( .A1(n1981), .A2(n1839), .B1(n1979), .B2(n1838), .ZN(
        n1840) );
  NR4D0BWP12T U2586 ( .A1(n1843), .A2(n1842), .A3(n1841), .A4(n1840), .ZN(
        n1844) );
  ND2D1BWP12T U2587 ( .A1(n1845), .A2(n1844), .ZN(regB_out[5]) );
  OAI22D1BWP12T U2588 ( .A1(n1847), .A2(n1949), .B1(n1948), .B2(n1846), .ZN(
        n1856) );
  INVD1BWP12T U2589 ( .I(tmp1[1]), .ZN(n1848) );
  MOAI22D0BWP12T U2590 ( .A1(n1848), .A2(n1951), .B1(n150), .B2(
        immediate2_in[1]), .ZN(n1855) );
  AOI22D1BWP12T U2591 ( .A1(r9[1]), .A2(n152), .B1(n1953), .B2(r4[1]), .ZN(
        n1850) );
  AOI22D1BWP12T U2592 ( .A1(r11[1]), .A2(n1955), .B1(n1954), .B2(r0[1]), .ZN(
        n1849) );
  ND2D1BWP12T U2593 ( .A1(n1850), .A2(n1849), .ZN(n1854) );
  OAI22D1BWP12T U2594 ( .A1(n1961), .A2(n1852), .B1(n1959), .B2(n1851), .ZN(
        n1853) );
  NR4D0BWP12T U2595 ( .A1(n1856), .A2(n1855), .A3(n1854), .A4(n1853), .ZN(
        n1870) );
  OAI22D1BWP12T U2596 ( .A1(n1858), .A2(n1968), .B1(n1967), .B2(n1857), .ZN(
        n1868) );
  OAI22D1BWP12T U2597 ( .A1(n1860), .A2(n1972), .B1(n1971), .B2(n1859), .ZN(
        n1867) );
  OAI22D1BWP12T U2598 ( .A1(n1977), .A2(n1862), .B1(n1975), .B2(n1861), .ZN(
        n1866) );
  OAI22D1BWP12T U2599 ( .A1(n1981), .A2(n1864), .B1(n1979), .B2(n1863), .ZN(
        n1865) );
  NR4D0BWP12T U2600 ( .A1(n1868), .A2(n1867), .A3(n1866), .A4(n1865), .ZN(
        n1869) );
  ND2D1BWP12T U2601 ( .A1(n1870), .A2(n1869), .ZN(regB_out[1]) );
  AOI22D1BWP12T U2602 ( .A1(tmp1[0]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[0]), .ZN(n1875) );
  AOI22D1BWP12T U2603 ( .A1(r5[0]), .A2(n1988), .B1(n158), .B2(r10[0]), .ZN(
        n1872) );
  AOI22D1BWP12T U2604 ( .A1(r7[0]), .A2(n1990), .B1(n1989), .B2(r2[0]), .ZN(
        n1871) );
  ND2D1BWP12T U2605 ( .A1(n1872), .A2(n1871), .ZN(n1874) );
  INR3XD0BWP12T U2606 ( .A1(n1875), .B1(n1874), .B2(n1873), .ZN(n1881) );
  AOI22D1BWP12T U2607 ( .A1(r1[0]), .A2(n164), .B1(n1993), .B2(r12[0]), .ZN(
        n1879) );
  AOI22D1BWP12T U2608 ( .A1(r3[0]), .A2(n1994), .B1(n168), .B2(lr[0]), .ZN(
        n1878) );
  AOI22D1BWP12T U2609 ( .A1(r8[0]), .A2(n171), .B1(n1995), .B2(n[2041]), .ZN(
        n1877) );
  AOI22D1BWP12T U2610 ( .A1(pc_out[0]), .A2(n174), .B1(n1996), .B2(r6[0]), 
        .ZN(n1876) );
  AN4XD1BWP12T U2611 ( .A1(n1879), .A2(n1878), .A3(n1877), .A4(n1876), .Z(
        n1880) );
  ND2D1BWP12T U2612 ( .A1(n1881), .A2(n1880), .ZN(regB_out[0]) );
  OAI22D1BWP12T U2613 ( .A1(n1885), .A2(n1884), .B1(n1883), .B2(n1882), .ZN(
        n1899) );
  OAI22D1BWP12T U2614 ( .A1(n1889), .A2(n1888), .B1(n1887), .B2(n1886), .ZN(
        n1898) );
  AOI22D1BWP12T U2615 ( .A1(n112), .A2(r12[4]), .B1(n273), .B2(tmp1[4]), .ZN(
        n1890) );
  IOA21D1BWP12T U2616 ( .A1(n1891), .A2(r4[4]), .B(n1890), .ZN(n1897) );
  OAI22D1BWP12T U2617 ( .A1(n1895), .A2(n1894), .B1(n1893), .B2(n1892), .ZN(
        n1896) );
  NR4D0BWP12T U2618 ( .A1(n1899), .A2(n1898), .A3(n1897), .A4(n1896), .ZN(
        n1921) );
  OAI22D1BWP12T U2619 ( .A1(n1903), .A2(n1902), .B1(n1901), .B2(n1900), .ZN(
        n1919) );
  OAI22D1BWP12T U2620 ( .A1(n1907), .A2(n1906), .B1(n1905), .B2(n1904), .ZN(
        n1918) );
  OAI22D1BWP12T U2621 ( .A1(n1911), .A2(n1910), .B1(n1909), .B2(n1908), .ZN(
        n1917) );
  OAI22D1BWP12T U2622 ( .A1(n1915), .A2(n1914), .B1(n1913), .B2(n1912), .ZN(
        n1916) );
  NR4D0BWP12T U2623 ( .A1(n1919), .A2(n1918), .A3(n1917), .A4(n1916), .ZN(
        n1920) );
  ND2D1BWP12T U2624 ( .A1(n1921), .A2(n1920), .ZN(regA_out[4]) );
  OAI22D1BWP12T U2625 ( .A1(n1923), .A2(n1949), .B1(n1948), .B2(n1922), .ZN(
        n1932) );
  INVD1BWP12T U2626 ( .I(tmp1[3]), .ZN(n1924) );
  MOAI22D0BWP12T U2627 ( .A1(n1924), .A2(n1951), .B1(n150), .B2(
        immediate2_in[3]), .ZN(n1931) );
  AOI22D1BWP12T U2628 ( .A1(r9[3]), .A2(n152), .B1(n1953), .B2(r4[3]), .ZN(
        n1926) );
  AOI22D1BWP12T U2629 ( .A1(r11[3]), .A2(n1955), .B1(n1954), .B2(r0[3]), .ZN(
        n1925) );
  ND2D1BWP12T U2630 ( .A1(n1926), .A2(n1925), .ZN(n1930) );
  OAI22D1BWP12T U2631 ( .A1(n1961), .A2(n1928), .B1(n1959), .B2(n1927), .ZN(
        n1929) );
  NR4D0BWP12T U2632 ( .A1(n1932), .A2(n1931), .A3(n1930), .A4(n1929), .ZN(
        n1946) );
  OAI22D1BWP12T U2633 ( .A1(n1934), .A2(n1968), .B1(n1967), .B2(n1933), .ZN(
        n1944) );
  OAI22D1BWP12T U2634 ( .A1(n1936), .A2(n1972), .B1(n1971), .B2(n1935), .ZN(
        n1943) );
  OAI22D1BWP12T U2635 ( .A1(n1977), .A2(n1938), .B1(n1975), .B2(n1937), .ZN(
        n1942) );
  OAI22D1BWP12T U2636 ( .A1(n1981), .A2(n1940), .B1(n1979), .B2(n1939), .ZN(
        n1941) );
  NR4D0BWP12T U2637 ( .A1(n1944), .A2(n1943), .A3(n1942), .A4(n1941), .ZN(
        n1945) );
  ND2D1BWP12T U2638 ( .A1(n1946), .A2(n1945), .ZN(regB_out[3]) );
  OAI22D1BWP12T U2639 ( .A1(n1950), .A2(n1949), .B1(n1948), .B2(n1947), .ZN(
        n1965) );
  INVD1BWP12T U2640 ( .I(tmp1[2]), .ZN(n1952) );
  MOAI22D0BWP12T U2641 ( .A1(n1952), .A2(n1951), .B1(n150), .B2(
        immediate2_in[2]), .ZN(n1964) );
  AOI22D1BWP12T U2642 ( .A1(r9[2]), .A2(n152), .B1(n1953), .B2(r4[2]), .ZN(
        n1957) );
  AOI22D1BWP12T U2643 ( .A1(r11[2]), .A2(n1955), .B1(n1954), .B2(r0[2]), .ZN(
        n1956) );
  TPND2D0BWP12T U2644 ( .A1(n1957), .A2(n1956), .ZN(n1963) );
  OAI22D1BWP12T U2645 ( .A1(n1961), .A2(n1960), .B1(n1959), .B2(n1958), .ZN(
        n1962) );
  NR4D0BWP12T U2646 ( .A1(n1965), .A2(n1964), .A3(n1963), .A4(n1962), .ZN(
        n1987) );
  OAI22D1BWP12T U2647 ( .A1(n1969), .A2(n1968), .B1(n1967), .B2(n1966), .ZN(
        n1985) );
  OAI22D1BWP12T U2648 ( .A1(n1973), .A2(n1972), .B1(n1971), .B2(n1970), .ZN(
        n1984) );
  OAI22D1BWP12T U2649 ( .A1(n1977), .A2(n1976), .B1(n1975), .B2(n1974), .ZN(
        n1983) );
  OAI22D1BWP12T U2650 ( .A1(n1981), .A2(n1980), .B1(n1979), .B2(n1978), .ZN(
        n1982) );
  NR4D0BWP12T U2651 ( .A1(n1985), .A2(n1984), .A3(n1983), .A4(n1982), .ZN(
        n1986) );
  ND2D1BWP12T U2652 ( .A1(n1987), .A2(n1986), .ZN(regB_out[2]) );
  INR2D1BWP12T U2653 ( .A1(next_cpsr_in[1]), .B1(reset), .ZN(cpsrin[1]) );
  AOI22D1BWP12T U2654 ( .A1(r5[19]), .A2(n1988), .B1(n158), .B2(r10[19]), .ZN(
        n1992) );
  AOI22D1BWP12T U2655 ( .A1(r7[19]), .A2(n1990), .B1(n1989), .B2(r2[19]), .ZN(
        n1991) );
  ND2D1BWP12T U2656 ( .A1(n1992), .A2(n1991), .ZN(n2009) );
  AOI22D1BWP12T U2657 ( .A1(r1[19]), .A2(n164), .B1(n1993), .B2(r12[19]), .ZN(
        n2000) );
  AOI22D1BWP12T U2658 ( .A1(r3[19]), .A2(n1994), .B1(n168), .B2(lr[19]), .ZN(
        n1999) );
  AOI22D1BWP12T U2659 ( .A1(r8[19]), .A2(n171), .B1(n1995), .B2(n[2022]), .ZN(
        n1998) );
  AOI22D1BWP12T U2660 ( .A1(pc_out[19]), .A2(n174), .B1(n1996), .B2(r6[19]), 
        .ZN(n1997) );
  AN4XD1BWP12T U2661 ( .A1(n2000), .A2(n1999), .A3(n1998), .A4(n1997), .Z(
        n2008) );
  AOI22D1BWP12T U2662 ( .A1(tmp1[19]), .A2(n2001), .B1(n150), .B2(
        immediate2_in[19]), .ZN(n2006) );
  AOI22D1BWP12T U2663 ( .A1(r9[19]), .A2(n152), .B1(n2002), .B2(r4[19]), .ZN(
        n2005) );
  AOI22D1BWP12T U2664 ( .A1(r11[19]), .A2(n2003), .B1(n1954), .B2(r0[19]), 
        .ZN(n2004) );
  AN3XD1BWP12T U2665 ( .A1(n2006), .A2(n2005), .A3(n2004), .Z(n2007) );
  IND3D1BWP12T U2666 ( .A1(n2009), .B1(n2008), .B2(n2007), .ZN(regB_out[19])
         );
endmodule


module ALU_VARIABLE ( a, b, op, c_in, result, c_out, z, n, v );
  input [31:0] a;
  input [31:0] b;
  input [3:0] op;
  output [31:0] result;
  input c_in;
  output c_out, z, n, v;
  wire   mult_x_18_n1029, mult_x_18_n1025, mult_x_18_n1021, mult_x_18_n1017,
         mult_x_18_n1013, mult_x_18_n1009, mult_x_18_n1005, mult_x_18_n998,
         mult_x_18_n997, mult_x_18_n994, mult_x_18_n993, mult_x_18_n990,
         mult_x_18_n989, mult_x_18_n986, mult_x_18_n985, mult_x_18_n982,
         mult_x_18_n981, mult_x_18_n978, mult_x_18_n977, mult_x_18_n974,
         mult_x_18_n973, mult_x_18_n969, mult_x_18_n967, mult_x_18_n965,
         mult_x_18_n964, mult_x_18_n963, mult_x_18_n961, mult_x_18_n960,
         mult_x_18_n959, mult_x_18_n958, mult_x_18_n957, mult_x_18_n956,
         mult_x_18_n955, mult_x_18_n954, mult_x_18_n953, mult_x_18_n952,
         mult_x_18_n951, mult_x_18_n950, mult_x_18_n949, mult_x_18_n948,
         mult_x_18_n947, mult_x_18_n946, mult_x_18_n945, mult_x_18_n944,
         mult_x_18_n942, mult_x_18_n941, mult_x_18_n940, mult_x_18_n939,
         mult_x_18_n938, mult_x_18_n937, mult_x_18_n936, mult_x_18_n935,
         mult_x_18_n934, mult_x_18_n933, mult_x_18_n932, mult_x_18_n931,
         mult_x_18_n930, mult_x_18_n929, mult_x_18_n928, mult_x_18_n927,
         mult_x_18_n926, mult_x_18_n925, mult_x_18_n924, mult_x_18_n923,
         mult_x_18_n922, mult_x_18_n921, mult_x_18_n920, mult_x_18_n919,
         mult_x_18_n918, mult_x_18_n917, mult_x_18_n913, mult_x_18_n912,
         mult_x_18_n911, mult_x_18_n910, mult_x_18_n909, mult_x_18_n908,
         mult_x_18_n907, mult_x_18_n906, mult_x_18_n905, mult_x_18_n904,
         mult_x_18_n903, mult_x_18_n902, mult_x_18_n901, mult_x_18_n900,
         mult_x_18_n899, mult_x_18_n898, mult_x_18_n897, mult_x_18_n896,
         mult_x_18_n895, mult_x_18_n894, mult_x_18_n893, mult_x_18_n892,
         mult_x_18_n890, mult_x_18_n889, mult_x_18_n888, mult_x_18_n886,
         mult_x_18_n884, mult_x_18_n882, mult_x_18_n881, mult_x_18_n880,
         mult_x_18_n878, mult_x_18_n877, mult_x_18_n876, mult_x_18_n874,
         mult_x_18_n873, mult_x_18_n872, mult_x_18_n871, mult_x_18_n870,
         mult_x_18_n869, mult_x_18_n866, mult_x_18_n865, mult_x_18_n864,
         mult_x_18_n863, mult_x_18_n862, mult_x_18_n861, mult_x_18_n860,
         mult_x_18_n859, mult_x_18_n858, mult_x_18_n857, mult_x_18_n856,
         mult_x_18_n855, mult_x_18_n854, mult_x_18_n853, mult_x_18_n852,
         mult_x_18_n851, mult_x_18_n850, mult_x_18_n849, mult_x_18_n848,
         mult_x_18_n846, mult_x_18_n845, mult_x_18_n844, mult_x_18_n843,
         mult_x_18_n842, mult_x_18_n841, mult_x_18_n840, mult_x_18_n839,
         mult_x_18_n838, mult_x_18_n837, mult_x_18_n836, mult_x_18_n835,
         mult_x_18_n834, mult_x_18_n833, mult_x_18_n832, mult_x_18_n831,
         mult_x_18_n830, mult_x_18_n829, mult_x_18_n825, mult_x_18_n823,
         mult_x_18_n821, mult_x_18_n819, mult_x_18_n817, mult_x_18_n815,
         mult_x_18_n814, mult_x_18_n813, mult_x_18_n812, mult_x_18_n810,
         mult_x_18_n809, mult_x_18_n808, mult_x_18_n807, mult_x_18_n806,
         mult_x_18_n805, mult_x_18_n804, mult_x_18_n803, mult_x_18_n802,
         mult_x_18_n801, mult_x_18_n800, mult_x_18_n799, mult_x_18_n798,
         mult_x_18_n797, mult_x_18_n794, mult_x_18_n793, mult_x_18_n792,
         mult_x_18_n791, mult_x_18_n790, mult_x_18_n789, mult_x_18_n788,
         mult_x_18_n787, mult_x_18_n786, mult_x_18_n785, mult_x_18_n784,
         mult_x_18_n782, mult_x_18_n781, mult_x_18_n780, mult_x_18_n778,
         mult_x_18_n777, mult_x_18_n776, mult_x_18_n774, mult_x_18_n773,
         mult_x_18_n770, mult_x_18_n769, mult_x_18_n768, mult_x_18_n767,
         mult_x_18_n766, mult_x_18_n765, mult_x_18_n764, mult_x_18_n762,
         mult_x_18_n761, mult_x_18_n760, mult_x_18_n759, mult_x_18_n758,
         mult_x_18_n757, mult_x_18_n753, mult_x_18_n752, mult_x_18_n750,
         mult_x_18_n749, mult_x_18_n744, mult_x_18_n740, mult_x_18_n738,
         mult_x_18_n736, mult_x_18_n735, mult_x_18_n734, mult_x_18_n726,
         mult_x_18_n723, mult_x_18_n722, mult_x_18_n721, mult_x_18_n720,
         mult_x_18_n719, mult_x_18_n718, mult_x_18_n717, mult_x_18_n716,
         mult_x_18_n715, mult_x_18_n714, mult_x_18_n713, mult_x_18_n712,
         mult_x_18_n711, mult_x_18_n710, mult_x_18_n709, mult_x_18_n708,
         mult_x_18_n707, mult_x_18_n706, mult_x_18_n705, mult_x_18_n704,
         mult_x_18_n703, mult_x_18_n702, mult_x_18_n701, mult_x_18_n700,
         mult_x_18_n699, mult_x_18_n698, mult_x_18_n697, mult_x_18_n696,
         mult_x_18_n695, mult_x_18_n694, mult_x_18_n693, mult_x_18_n692,
         mult_x_18_n691, mult_x_18_n690, mult_x_18_n689, mult_x_18_n688,
         mult_x_18_n687, mult_x_18_n686, mult_x_18_n685, mult_x_18_n684,
         mult_x_18_n683, mult_x_18_n682, mult_x_18_n681, mult_x_18_n680,
         mult_x_18_n679, mult_x_18_n678, mult_x_18_n677, mult_x_18_n676,
         mult_x_18_n675, mult_x_18_n674, mult_x_18_n673, mult_x_18_n672,
         mult_x_18_n671, mult_x_18_n670, mult_x_18_n669, mult_x_18_n668,
         mult_x_18_n667, mult_x_18_n666, mult_x_18_n665, mult_x_18_n664,
         mult_x_18_n663, mult_x_18_n662, mult_x_18_n661, mult_x_18_n660,
         mult_x_18_n659, mult_x_18_n658, mult_x_18_n657, mult_x_18_n656,
         mult_x_18_n655, mult_x_18_n654, mult_x_18_n653, mult_x_18_n652,
         mult_x_18_n651, mult_x_18_n650, mult_x_18_n649, mult_x_18_n648,
         mult_x_18_n647, mult_x_18_n646, mult_x_18_n645, mult_x_18_n644,
         mult_x_18_n643, mult_x_18_n642, mult_x_18_n641, mult_x_18_n640,
         mult_x_18_n639, mult_x_18_n638, mult_x_18_n637, mult_x_18_n636,
         mult_x_18_n635, mult_x_18_n634, mult_x_18_n633, mult_x_18_n632,
         mult_x_18_n631, mult_x_18_n630, mult_x_18_n629, mult_x_18_n628,
         mult_x_18_n627, mult_x_18_n626, mult_x_18_n625, mult_x_18_n624,
         mult_x_18_n623, mult_x_18_n622, mult_x_18_n621, mult_x_18_n620,
         mult_x_18_n619, mult_x_18_n618, mult_x_18_n617, mult_x_18_n616,
         mult_x_18_n615, mult_x_18_n614, mult_x_18_n613, mult_x_18_n612,
         mult_x_18_n611, mult_x_18_n610, mult_x_18_n609, mult_x_18_n608,
         mult_x_18_n607, mult_x_18_n606, mult_x_18_n605, mult_x_18_n604,
         mult_x_18_n603, mult_x_18_n602, mult_x_18_n601, mult_x_18_n600,
         mult_x_18_n599, mult_x_18_n598, mult_x_18_n597, mult_x_18_n596,
         mult_x_18_n595, mult_x_18_n594, mult_x_18_n593, mult_x_18_n592,
         mult_x_18_n591, mult_x_18_n590, mult_x_18_n589, mult_x_18_n588,
         mult_x_18_n587, mult_x_18_n586, mult_x_18_n585, mult_x_18_n584,
         mult_x_18_n583, mult_x_18_n582, mult_x_18_n581, mult_x_18_n580,
         mult_x_18_n579, mult_x_18_n578, mult_x_18_n577, mult_x_18_n576,
         mult_x_18_n575, mult_x_18_n574, mult_x_18_n573, mult_x_18_n572,
         mult_x_18_n571, mult_x_18_n570, mult_x_18_n569, mult_x_18_n568,
         mult_x_18_n567, mult_x_18_n566, mult_x_18_n565, mult_x_18_n564,
         mult_x_18_n563, mult_x_18_n562, mult_x_18_n561, mult_x_18_n560,
         mult_x_18_n559, mult_x_18_n558, mult_x_18_n557, mult_x_18_n556,
         mult_x_18_n555, mult_x_18_n554, mult_x_18_n553, mult_x_18_n552,
         mult_x_18_n551, mult_x_18_n550, mult_x_18_n549, mult_x_18_n548,
         mult_x_18_n547, mult_x_18_n546, mult_x_18_n545, mult_x_18_n544,
         mult_x_18_n543, mult_x_18_n542, mult_x_18_n541, mult_x_18_n540,
         mult_x_18_n539, mult_x_18_n538, mult_x_18_n537, mult_x_18_n536,
         mult_x_18_n535, mult_x_18_n534, mult_x_18_n533, mult_x_18_n532,
         mult_x_18_n531, mult_x_18_n530, mult_x_18_n529, mult_x_18_n528,
         mult_x_18_n527, mult_x_18_n526, mult_x_18_n525, mult_x_18_n524,
         mult_x_18_n523, mult_x_18_n522, mult_x_18_n521, mult_x_18_n520,
         mult_x_18_n519, mult_x_18_n518, mult_x_18_n517, mult_x_18_n516,
         mult_x_18_n515, mult_x_18_n514, mult_x_18_n513, mult_x_18_n512,
         mult_x_18_n511, mult_x_18_n510, mult_x_18_n509, mult_x_18_n508,
         mult_x_18_n507, mult_x_18_n506, mult_x_18_n505, mult_x_18_n504,
         mult_x_18_n503, mult_x_18_n502, mult_x_18_n501, mult_x_18_n500,
         mult_x_18_n499, mult_x_18_n498, mult_x_18_n497, mult_x_18_n496,
         mult_x_18_n495, mult_x_18_n494, mult_x_18_n493, mult_x_18_n492,
         mult_x_18_n491, mult_x_18_n490, mult_x_18_n489, mult_x_18_n488,
         mult_x_18_n487, mult_x_18_n486, mult_x_18_n485, mult_x_18_n484,
         mult_x_18_n483, mult_x_18_n482, mult_x_18_n481, mult_x_18_n480,
         mult_x_18_n479, mult_x_18_n478, mult_x_18_n477, mult_x_18_n476,
         mult_x_18_n475, mult_x_18_n474, mult_x_18_n473, mult_x_18_n472,
         mult_x_18_n471, mult_x_18_n470, mult_x_18_n469, mult_x_18_n468,
         mult_x_18_n467, mult_x_18_n466, mult_x_18_n465, mult_x_18_n464,
         mult_x_18_n463, mult_x_18_n462, mult_x_18_n461, mult_x_18_n460,
         mult_x_18_n459, mult_x_18_n458, mult_x_18_n457, mult_x_18_n456,
         mult_x_18_n455, mult_x_18_n454, mult_x_18_n453, mult_x_18_n452,
         mult_x_18_n451, mult_x_18_n450, mult_x_18_n449, mult_x_18_n448,
         mult_x_18_n447, mult_x_18_n446, mult_x_18_n445, mult_x_18_n444,
         mult_x_18_n443, mult_x_18_n442, mult_x_18_n441, mult_x_18_n440,
         mult_x_18_n439, mult_x_18_n438, mult_x_18_n437, mult_x_18_n436,
         mult_x_18_n435, mult_x_18_n434, mult_x_18_n433, mult_x_18_n432,
         mult_x_18_n431, mult_x_18_n430, mult_x_18_n429, mult_x_18_n428,
         mult_x_18_n427, mult_x_18_n426, mult_x_18_n425, mult_x_18_n424,
         mult_x_18_n423, mult_x_18_n422, mult_x_18_n421, mult_x_18_n420,
         mult_x_18_n419, mult_x_18_n418, mult_x_18_n417, mult_x_18_n416,
         mult_x_18_n415, mult_x_18_n414, mult_x_18_n413, mult_x_18_n412,
         mult_x_18_n411, mult_x_18_n410, mult_x_18_n409, mult_x_18_n408,
         mult_x_18_n407, mult_x_18_n406, mult_x_18_n405, mult_x_18_n404,
         mult_x_18_n403, mult_x_18_n402, mult_x_18_n400, mult_x_18_n399,
         mult_x_18_n398, mult_x_18_n397, mult_x_18_n396, mult_x_18_n395,
         mult_x_18_n394, mult_x_18_n393, mult_x_18_n392, mult_x_18_n391,
         mult_x_18_n390, mult_x_18_n389, mult_x_18_n388, mult_x_18_n387,
         mult_x_18_n386, mult_x_18_n385, mult_x_18_n384, mult_x_18_n383,
         mult_x_18_n382, mult_x_18_n381, mult_x_18_n380, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130;

  CMPE42D2BWP12T mult_x_18_U483 ( .A(mult_x_18_n660), .B(mult_x_18_n670), .C(
        mult_x_18_n657), .CIX(mult_x_18_n663), .D(mult_x_18_n667), .CO(
        mult_x_18_n653), .COX(mult_x_18_n652), .S(mult_x_18_n654) );
  CMPE42D1BWP12T mult_x_18_U507 ( .A(mult_x_18_n744), .B(mult_x_18_n941), .C(
        mult_x_18_n997), .CIX(mult_x_18_n721), .D(mult_x_18_n720), .CO(
        mult_x_18_n717), .COX(mult_x_18_n716), .S(mult_x_18_n718) );
  CMPE42D1BWP12T mult_x_18_U502 ( .A(mult_x_18_n710), .B(mult_x_18_n939), .C(
        mult_x_18_n714), .CIX(mult_x_18_n711), .D(mult_x_18_n708), .CO(
        mult_x_18_n705), .COX(mult_x_18_n704), .S(mult_x_18_n706) );
  CMPE42D1BWP12T mult_x_18_U432 ( .A(mult_x_18_n950), .B(mult_x_18_n790), .C(
        mult_x_18_n538), .CIX(mult_x_18_n535), .D(mult_x_18_n520), .CO(
        mult_x_18_n511), .COX(mult_x_18_n510), .S(mult_x_18_n512) );
  CMPE42D1BWP12T mult_x_18_U465 ( .A(mult_x_18_n623), .B(mult_x_18_n610), .C(
        mult_x_18_n620), .CIX(mult_x_18_n616), .D(mult_x_18_n607), .CO(
        mult_x_18_n603), .COX(mult_x_18_n602), .S(mult_x_18_n604) );
  CMPE42D1BWP12T mult_x_18_U490 ( .A(mult_x_18_n679), .B(mult_x_18_n688), .C(
        mult_x_18_n682), .CIX(mult_x_18_n677), .D(mult_x_18_n686), .CO(
        mult_x_18_n673), .COX(mult_x_18_n672), .S(mult_x_18_n674) );
  FA1D0BWP12T U3 ( .A(n817), .B(n816), .CI(n815), .CO(mult_x_18_n714), .S(
        mult_x_18_n715) );
  FA1D0BWP12T U4 ( .A(n820), .B(n819), .CI(n818), .CO(mult_x_18_n688), .S(
        mult_x_18_n689) );
  CKBD1BWP12T U5 ( .I(n2405), .Z(n342) );
  NR2D1BWP12T U6 ( .A1(b[27]), .A2(b[26]), .ZN(n391) );
  INVD3BWP12T U7 ( .I(n2659), .ZN(n2657) );
  AOI21D1BWP12T U8 ( .A1(n352), .A2(n1891), .B(n351), .ZN(n1900) );
  INVD1BWP12T U9 ( .I(n2750), .ZN(n319) );
  INVD1BWP12T U10 ( .I(n2807), .ZN(n321) );
  NR2D1BWP12T U11 ( .A1(n345), .A2(n2766), .ZN(n1878) );
  INVD1BWP12T U12 ( .I(n2404), .ZN(n1937) );
  OR2XD1BWP12T U13 ( .A1(mult_x_18_n674), .A2(mult_x_18_n683), .Z(n1585) );
  OR2XD1BWP12T U14 ( .A1(mult_x_18_n673), .A2(mult_x_18_n665), .Z(n1625) );
  INVD1BWP12T U15 ( .I(n1437), .ZN(n1626) );
  OAI21D1BWP12T U16 ( .A1(n1555), .A2(n286), .B(n285), .ZN(n1561) );
  ND2D1BWP12T U17 ( .A1(n2473), .A2(n3119), .ZN(n1368) );
  INVD1BWP12T U18 ( .I(n2416), .ZN(n2281) );
  OR2XD1BWP12T U19 ( .A1(mult_x_18_n692), .A2(mult_x_18_n699), .Z(n1589) );
  OR2XD1BWP12T U20 ( .A1(mult_x_18_n706), .A2(mult_x_18_n712), .Z(n1595) );
  INVD1BWP12T U21 ( .I(n2799), .ZN(n2802) );
  INVD1BWP12T U22 ( .I(n2748), .ZN(n2749) );
  NR2D1BWP12T U23 ( .A1(n1870), .A2(n1878), .ZN(n1850) );
  OAI21D1BWP12T U24 ( .A1(n615), .A2(n784), .B(n616), .ZN(n343) );
  AOI21D1BWP12T U25 ( .A1(n438), .A2(n778), .B(n437), .ZN(n609) );
  HA1D0BWP12T U26 ( .A(n968), .B(n967), .CO(mult_x_18_n614), .S(mult_x_18_n615) );
  XOR2D1BWP12T U27 ( .A1(n1700), .A2(n1699), .Z(n2827) );
  OAI21D1BWP12T U28 ( .A1(n1271), .A2(n1270), .B(n1269), .ZN(n1276) );
  NR2D1BWP12T U29 ( .A1(n2478), .A2(n2943), .ZN(n1372) );
  CMPE42D1BWP12T U30 ( .A(mult_x_18_n635), .B(mult_x_18_n624), .C(
        mult_x_18_n632), .CIX(mult_x_18_n628), .D(mult_x_18_n621), .CO(
        mult_x_18_n617), .COX(mult_x_18_n616), .S(mult_x_18_n618) );
  CMPE42D1BWP12T U31 ( .A(mult_x_18_n536), .B(mult_x_18_n518), .C(
        mult_x_18_n509), .CIX(mult_x_18_n523), .D(mult_x_18_n527), .CO(
        mult_x_18_n505), .COX(mult_x_18_n504), .S(mult_x_18_n506) );
  INVD1BWP12T U32 ( .I(a[10]), .ZN(n3069) );
  OR2XD1BWP12T U33 ( .A1(n2452), .A2(n2305), .Z(n2114) );
  OAI21D1BWP12T U34 ( .A1(n290), .A2(n1562), .B(n289), .ZN(n699) );
  INVD1BWP12T U35 ( .I(n411), .ZN(n2065) );
  INVD1BWP12T U36 ( .I(b[6]), .ZN(n2259) );
  INVD1BWP12T U37 ( .I(a[14]), .ZN(n2280) );
  OR2XD1BWP12T U38 ( .A1(mult_x_18_n590), .A2(mult_x_18_n603), .Z(n1572) );
  CMPE42D1BWP12T U39 ( .A(mult_x_18_n1013), .B(mult_x_18_n782), .C(
        mult_x_18_n901), .CIX(mult_x_18_n584), .D(mult_x_18_n586), .CO(
        mult_x_18_n570), .COX(mult_x_18_n569), .S(mult_x_18_n571) );
  XNR2D1BWP12T U40 ( .A1(n2633), .A2(n2807), .ZN(n1062) );
  HA1D0BWP12T U41 ( .A(n986), .B(n985), .CO(mult_x_18_n484), .S(mult_x_18_n485) );
  HA1D0BWP12T U42 ( .A(n940), .B(n939), .CO(mult_x_18_n661), .S(mult_x_18_n662) );
  CMPE42D1BWP12T U43 ( .A(mult_x_18_n659), .B(mult_x_18_n649), .C(
        mult_x_18_n656), .CIX(mult_x_18_n652), .D(mult_x_18_n646), .CO(
        mult_x_18_n642), .COX(mult_x_18_n641), .S(mult_x_18_n643) );
  INVD1BWP12T U44 ( .I(n2829), .ZN(n323) );
  INVD1BWP12T U45 ( .I(n559), .ZN(n1538) );
  INVD1BWP12T U46 ( .I(n2522), .ZN(n2247) );
  INVD2BWP12T U47 ( .I(b[0]), .ZN(n2422) );
  INVD2BWP12T U48 ( .I(n3069), .ZN(n3067) );
  INVD3BWP12T U49 ( .I(n386), .ZN(n2750) );
  CKBD1BWP12T U50 ( .I(a[24]), .Z(n2403) );
  INVD2BWP12T U51 ( .I(n2063), .ZN(n1999) );
  DEL025D1BWP12T U52 ( .I(b[14]), .Z(n2522) );
  INVD2BWP12T U53 ( .I(n2261), .ZN(n2766) );
  INVD2BWP12T U54 ( .I(n2252), .ZN(n2501) );
  XNR2D2BWP12T U55 ( .A1(n2494), .A2(n2416), .ZN(n2539) );
  OR2XD1BWP12T U56 ( .A1(mult_x_18_n559), .A2(mult_x_18_n573), .Z(n1637) );
  INVD2BWP12T U57 ( .I(n2998), .ZN(n2993) );
  ND2D1BWP12T U58 ( .A1(n2221), .A2(n2868), .ZN(n2211) );
  INVD1BWP12T U59 ( .I(a[19]), .ZN(n2659) );
  CKBD1BWP12T U60 ( .I(a[18]), .Z(n2689) );
  CKBD1BWP12T U61 ( .I(a[16]), .Z(n2891) );
  INVD1BWP12T U62 ( .I(a[20]), .ZN(n2928) );
  INVD1BWP12T U63 ( .I(n2980), .ZN(n3115) );
  CKBD1BWP12T U64 ( .I(a[22]), .Z(n2963) );
  INVD1BWP12T U65 ( .I(n2996), .ZN(n3105) );
  CMPE42D1BWP12T U66 ( .A(mult_x_18_n548), .B(mult_x_18_n554), .C(
        mult_x_18_n561), .CIX(mult_x_18_n557), .D(mult_x_18_n545), .CO(
        mult_x_18_n541), .COX(mult_x_18_n540), .S(mult_x_18_n542) );
  INVD1BWP12T U67 ( .I(n2501), .ZN(n328) );
  OAI21D1BWP12T U68 ( .A1(n1538), .A2(n313), .B(n312), .ZN(n1455) );
  OR2XD1BWP12T U69 ( .A1(n2249), .A2(n2416), .Z(n1405) );
  OR2XD1BWP12T U70 ( .A1(n3033), .A2(b[13]), .Z(n1908) );
  ND2D1BWP12T U71 ( .A1(n2000), .A2(n1999), .ZN(n537) );
  OR2XD1BWP12T U72 ( .A1(n2405), .A2(n2407), .Z(n2150) );
  OR2XD1BWP12T U73 ( .A1(n3033), .A2(b[13]), .Z(n1690) );
  MOAI22D0BWP12T U74 ( .A1(n595), .A2(n2305), .B1(n2008), .B2(n2297), .ZN(
        n2026) );
  CMPE42D1BWP12T U75 ( .A(mult_x_18_n432), .B(mult_x_18_n449), .C(
        mult_x_18_n429), .CIX(mult_x_18_n446), .D(mult_x_18_n450), .CO(
        mult_x_18_n425), .COX(mult_x_18_n424), .S(mult_x_18_n426) );
  CMPE42D1BWP12T U76 ( .A(mult_x_18_n857), .B(mult_x_18_n821), .C(
        mult_x_18_n926), .CIX(mult_x_18_n578), .D(mult_x_18_n982), .CO(
        mult_x_18_n567), .COX(mult_x_18_n566), .S(mult_x_18_n568) );
  CMPE42D1BWP12T U77 ( .A(mult_x_18_n907), .B(mult_x_18_n884), .C(
        mult_x_18_n932), .CIX(mult_x_18_n655), .D(mult_x_18_n661), .CO(
        mult_x_18_n648), .COX(mult_x_18_n647), .S(mult_x_18_n649) );
  CMPE42D1BWP12T U78 ( .A(mult_x_18_n671), .B(mult_x_18_n961), .C(
        mult_x_18_n668), .CIX(mult_x_18_n672), .D(mult_x_18_n676), .CO(
        mult_x_18_n664), .COX(mult_x_18_n663), .S(mult_x_18_n665) );
  AOI21D1BWP12T U79 ( .A1(n1747), .A2(n1745), .B(n338), .ZN(n1817) );
  AOI21D1BWP12T U80 ( .A1(n1491), .A2(n1489), .B(n338), .ZN(n1487) );
  OAI21D1BWP12T U81 ( .A1(n1150), .A2(n1145), .B(n1148), .ZN(n1842) );
  OAI21D1BWP12T U82 ( .A1(n1668), .A2(n1666), .B(n1835), .ZN(n1665) );
  OAI21D1BWP12T U83 ( .A1(n1697), .A2(n1693), .B(n1694), .ZN(n1724) );
  OAI21D1BWP12T U84 ( .A1(n1487), .A2(n1483), .B(n1484), .ZN(n1482) );
  NR2D1BWP12T U85 ( .A1(n331), .A2(n1804), .ZN(n333) );
  CMPE42D1BWP12T U86 ( .A(mult_x_18_n911), .B(mult_x_18_n888), .C(
        mult_x_18_n936), .CIX(mult_x_18_n693), .D(mult_x_18_n696), .CO(
        mult_x_18_n686), .COX(mult_x_18_n685), .S(mult_x_18_n687) );
  CMPE42D1BWP12T U87 ( .A(mult_x_18_n474), .B(mult_x_18_n480), .C(
        mult_x_18_n471), .CIX(mult_x_18_n486), .D(mult_x_18_n490), .CO(
        mult_x_18_n467), .COX(mult_x_18_n466), .S(mult_x_18_n468) );
  CMPE42D1BWP12T U88 ( .A(mult_x_18_n906), .B(mult_x_18_n958), .C(
        mult_x_18_n931), .CIX(mult_x_18_n644), .D(mult_x_18_n640), .CO(
        mult_x_18_n635), .COX(mult_x_18_n634), .S(mult_x_18_n636) );
  CMPE42D1BWP12T U89 ( .A(mult_x_18_n853), .B(mult_x_18_n817), .C(
        mult_x_18_n897), .CIX(mult_x_18_n516), .D(mult_x_18_n922), .CO(
        mult_x_18_n499), .COX(mult_x_18_n498), .S(mult_x_18_n500) );
  CMPE42D1BWP12T U90 ( .A(mult_x_18_n803), .B(mult_x_18_n735), .C(
        mult_x_18_n835), .CIX(mult_x_18_n532), .D(mult_x_18_n854), .CO(
        mult_x_18_n514), .COX(mult_x_18_n513), .S(mult_x_18_n515) );
  CMPE42D1BWP12T U91 ( .A(mult_x_18_n837), .B(mult_x_18_n781), .C(
        mult_x_18_n856), .CIX(mult_x_18_n566), .D(mult_x_18_n900), .CO(
        mult_x_18_n550), .COX(mult_x_18_n549), .S(mult_x_18_n551) );
  HA1D0BWP12T U92 ( .A(n1011), .B(n1010), .CO(mult_x_18_n696), .S(
        mult_x_18_n697) );
  CMPE42D1BWP12T U93 ( .A(mult_x_18_n1029), .B(mult_x_18_n942), .C(
        mult_x_18_n969), .CIX(mult_x_18_n726), .D(mult_x_18_n998), .CO(
        mult_x_18_n722), .COX(mult_x_18_n721), .S(mult_x_18_n723) );
  CMPE42D1BWP12T U94 ( .A(mult_x_18_n940), .B(mult_x_18_n967), .C(
        mult_x_18_n719), .CIX(mult_x_18_n716), .D(mult_x_18_n715), .CO(
        mult_x_18_n712), .COX(mult_x_18_n711), .S(mult_x_18_n713) );
  HA1D0BWP12T U95 ( .A(n959), .B(n958), .CO(mult_x_18_n521), .S(mult_x_18_n522) );
  HA1D0BWP12T U96 ( .A(n1022), .B(n1021), .CO(mult_x_18_n555), .S(
        mult_x_18_n556) );
  HA1D0BWP12T U97 ( .A(n1039), .B(n1038), .CO(mult_x_18_n639), .S(
        mult_x_18_n640) );
  CMPE42D1BWP12T U98 ( .A(mult_x_18_n938), .B(mult_x_18_n965), .C(
        mult_x_18_n994), .CIX(mult_x_18_n703), .D(mult_x_18_n704), .CO(
        mult_x_18_n699), .COX(mult_x_18_n698), .S(mult_x_18_n700) );
  HA1D0BWP12T U99 ( .A(n875), .B(n874), .CO(mult_x_18_n709), .S(mult_x_18_n710) );
  HA1D0BWP12T U100 ( .A(n245), .B(n244), .CO(n256), .S(n255) );
  CMPE42D1BWP12T U101 ( .A(mult_x_18_n511), .B(mult_x_18_n497), .C(
        mult_x_18_n491), .CIX(mult_x_18_n504), .D(mult_x_18_n508), .CO(
        mult_x_18_n487), .COX(mult_x_18_n486), .S(mult_x_18_n488) );
  OR2XD1BWP12T U102 ( .A1(n1898), .A2(n355), .Z(n357) );
  OR2XD1BWP12T U103 ( .A1(n1753), .A2(n1754), .Z(n335) );
  INVD1BWP12T U104 ( .I(n1831), .ZN(n1266) );
  CKND2D0BWP12T U105 ( .A1(n784), .A2(n785), .ZN(n1) );
  MAOI22D0BWP12T U106 ( .A1(n786), .A2(n1), .B1(n786), .B2(n1), .ZN(n1869) );
  IND4D0BWP12T U107 ( .A1(n2456), .B1(n2457), .B2(n2696), .B3(n2458), .ZN(n2)
         );
  IND4D0BWP12T U108 ( .A1(n2454), .B1(n2668), .B2(n2453), .B3(n2897), .ZN(n3)
         );
  OAI31D0BWP12T U109 ( .A1(n2460), .A2(n2), .A3(n3), .B(n2459), .ZN(n2461) );
  CKND0BWP12T U110 ( .I(n1538), .ZN(n4) );
  AN3D0BWP12T U111 ( .A1(n4), .A2(n1534), .A3(n1536), .Z(n5) );
  AOI211D0BWP12T U112 ( .A1(n1536), .A2(n1537), .B(n1535), .C(n5), .ZN(n6) );
  CKND2D0BWP12T U113 ( .A1(n1539), .A2(n1540), .ZN(n7) );
  MAOI22D0BWP12T U114 ( .A1(n6), .A2(n7), .B1(n6), .B2(n7), .ZN(n3048) );
  IND2D0BWP12T U115 ( .A1(op[0]), .B1(n358), .ZN(n383) );
  NR4D0BWP12T U116 ( .A1(n2846), .A2(n3054), .A3(n2887), .A4(n1682), .ZN(n8)
         );
  NR4D0BWP12T U117 ( .A1(n1712), .A2(n3097), .A3(n2943), .A4(n1713), .ZN(n9)
         );
  NR4D0BWP12T U118 ( .A1(n2741), .A2(n2795), .A3(n1719), .A4(n2827), .ZN(n10)
         );
  IND3D0BWP12T U119 ( .A1(n1720), .B1(n9), .B2(n10), .ZN(n11) );
  OR4D0BWP12T U120 ( .A1(n2781), .A2(n2714), .A3(n1721), .A4(n11), .Z(n12) );
  NR4D0BWP12T U121 ( .A1(n1722), .A2(n3026), .A3(n2683), .A4(n12), .ZN(n13) );
  NR3D0BWP12T U122 ( .A1(n3016), .A2(n2924), .A3(n2655), .ZN(n14) );
  ND4D0BWP12T U123 ( .A1(n2916), .A2(n8), .A3(n13), .A4(n14), .ZN(n15) );
  OR4D0BWP12T U124 ( .A1(n2629), .A2(n1727), .A3(n2983), .A4(n15), .Z(n16) );
  OR4D0BWP12T U125 ( .A1(n1730), .A2(n1728), .A3(n1729), .A4(n16), .Z(n17) );
  NR4D0BWP12T U126 ( .A1(n1732), .A2(n2602), .A3(n1731), .A4(n17), .ZN(n2479)
         );
  OA32D0BWP12T U127 ( .A1(n2149), .A2(n2613), .A3(n2150), .B1(n2750), .B2(
        n2149), .Z(n3037) );
  INR3D0BWP12T U128 ( .A1(n3091), .B1(n2234), .B2(n2216), .ZN(n18) );
  OR4D0BWP12T U129 ( .A1(n3090), .A2(n2212), .A3(n2214), .A4(n2213), .Z(n19)
         );
  AOI211D0BWP12T U130 ( .A1(n2440), .A2(n2776), .B(n2460), .C(n19), .ZN(n20)
         );
  ND4D0BWP12T U131 ( .A1(n2209), .A2(n2800), .A3(n18), .A4(n20), .ZN(n21) );
  OR4D0BWP12T U132 ( .A1(n2926), .A2(n2976), .A3(n2194), .A4(n2616), .Z(n22)
         );
  ND4D0BWP12T U133 ( .A1(n3065), .A2(n2869), .A3(n2669), .A4(n2631), .ZN(n23)
         );
  ND4D0BWP12T U134 ( .A1(n2223), .A2(n2222), .A3(n3013), .A4(n2224), .ZN(n24)
         );
  NR4D0BWP12T U135 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(n25) );
  ND4D0BWP12T U136 ( .A1(n2236), .A2(n2237), .A3(n2235), .A4(n25), .ZN(n2467)
         );
  CKND2D0BWP12T U137 ( .A1(n1385), .A2(n1386), .ZN(n26) );
  MOAI22D0BWP12T U138 ( .A1(n1387), .A2(n26), .B1(n1387), .B2(n26), .ZN(n1713)
         );
  CKND2D0BWP12T U139 ( .A1(n1193), .A2(n1143), .ZN(n27) );
  MAOI22D0BWP12T U140 ( .A1(n1194), .A2(n27), .B1(n1194), .B2(n27), .ZN(n1819)
         );
  CKND2D0BWP12T U141 ( .A1(n1591), .A2(n1592), .ZN(n28) );
  MOAI22D0BWP12T U142 ( .A1(n1593), .A2(n28), .B1(n1593), .B2(n28), .ZN(n3087)
         );
  NR2D0BWP12T U143 ( .A1(n1971), .A2(n1973), .ZN(n29) );
  MOAI22D0BWP12T U144 ( .A1(n2799), .A2(n29), .B1(n2799), .B2(n29), .ZN(n2793)
         );
  IND2D0BWP12T U145 ( .A1(n426), .B1(n358), .ZN(n1867) );
  NR4D0BWP12T U146 ( .A1(n2867), .A2(n2848), .A3(n3051), .A4(n1503), .ZN(n30)
         );
  NR4D0BWP12T U147 ( .A1(n1519), .A2(n1518), .A3(n2787), .A4(n2815), .ZN(n31)
         );
  NR4D0BWP12T U148 ( .A1(n1526), .A2(n3096), .A3(n1525), .A4(n3059), .ZN(n32)
         );
  NR2D0BWP12T U149 ( .A1(n2739), .A2(n2825), .ZN(n33) );
  NR3D0BWP12T U150 ( .A1(n1541), .A2(n2734), .A3(n3048), .ZN(n34) );
  ND4D0BWP12T U151 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(n35) );
  NR4D0BWP12T U152 ( .A1(n1546), .A2(n2918), .A3(n2707), .A4(n35), .ZN(n36) );
  NR3D0BWP12T U153 ( .A1(n3022), .A2(n2946), .A3(n2677), .ZN(n37) );
  NR3D0BWP12T U154 ( .A1(n1548), .A2(n2650), .A3(n2988), .ZN(n38) );
  ND4D0BWP12T U155 ( .A1(n30), .A2(n36), .A3(n37), .A4(n38), .ZN(n39) );
  OR4D0BWP12T U156 ( .A1(n1551), .A2(n1549), .A3(n1550), .A4(n39), .Z(n1553)
         );
  CKND2D0BWP12T U157 ( .A1(n1459), .A2(n1460), .ZN(n40) );
  MOAI22D0BWP12T U158 ( .A1(n1456), .A2(n40), .B1(n1456), .B2(n40), .ZN(n1911)
         );
  IAO21D0BWP12T U159 ( .A1(n2613), .A2(n2133), .B(n2134), .ZN(n3003) );
  IND2D0BWP12T U160 ( .A1(n1737), .B1(n1738), .ZN(n41) );
  MAOI22D0BWP12T U161 ( .A1(n1739), .A2(n41), .B1(n1739), .B2(n41), .ZN(n2991)
         );
  IND3D0BWP12T U162 ( .A1(n1538), .B1(n1534), .B2(n1810), .ZN(n42) );
  AOI211D0BWP12T U163 ( .A1(n1810), .A2(n1537), .B(n1403), .C(n43), .ZN(n44)
         );
  IND2D0BWP12T U164 ( .A1(n1399), .B1(n1400), .ZN(n45) );
  MAOI22D0BWP12T U165 ( .A1(n44), .A2(n45), .B1(n44), .B2(n45), .ZN(n1503) );
  CKND0BWP12T U166 ( .I(n42), .ZN(n43) );
  OAI21D0BWP12T U167 ( .A1(n1700), .A2(n1679), .B(n1678), .ZN(n46) );
  CKND2D0BWP12T U168 ( .A1(n1680), .A2(n1681), .ZN(n47) );
  MOAI22D0BWP12T U169 ( .A1(n46), .A2(n47), .B1(n46), .B2(n47), .ZN(n2887) );
  INR3D0BWP12T U170 ( .A1(n2802), .B1(n1971), .B2(n1973), .ZN(n48) );
  MOAI22D0BWP12T U171 ( .A1(n306), .A2(n48), .B1(n306), .B2(n48), .ZN(n2843)
         );
  IND2D0BWP12T U172 ( .A1(n1602), .B1(n1603), .ZN(n49) );
  MAOI22D0BWP12T U173 ( .A1(n1604), .A2(n49), .B1(n1604), .B2(n49), .ZN(n2791)
         );
  NR2D0BWP12T U174 ( .A1(n2860), .A2(n2310), .ZN(n50) );
  AOI22D0BWP12T U175 ( .A1(n2213), .A2(n3060), .B1(n3095), .B2(n1525), .ZN(n51) );
  MUX2ND0BWP12T U176 ( .I0(n3104), .I1(n3103), .S(n1383), .ZN(n52) );
  AOI31D0BWP12T U177 ( .A1(n3105), .A2(n2980), .A3(n52), .B(n2486), .ZN(n53)
         );
  OAI22D0BWP12T U178 ( .A1(n2262), .A2(n3109), .B1(n2422), .B2(n3105), .ZN(n54) );
  AOI211D0BWP12T U179 ( .A1(n3107), .A2(n2298), .B(n53), .C(n54), .ZN(n55) );
  CKND0BWP12T U180 ( .I(n2951), .ZN(n56) );
  AOI22D0BWP12T U181 ( .A1(n3119), .A2(n1868), .B1(n1614), .B2(n56), .ZN(n57)
         );
  CKND0BWP12T U182 ( .I(n3012), .ZN(n58) );
  AOI22D0BWP12T U183 ( .A1(n1792), .A2(n314), .B1(n2214), .B2(n58), .ZN(n59)
         );
  ND4D0BWP12T U184 ( .A1(n51), .A2(n55), .A3(n57), .A4(n59), .ZN(n60) );
  AOI211D0BWP12T U185 ( .A1(n1713), .A2(n3098), .B(n50), .C(n60), .ZN(n61) );
  OAI21D0BWP12T U186 ( .A1(n2101), .A2(n2438), .B(n3130), .ZN(n62) );
  OAI211D0BWP12T U187 ( .A1(n2103), .A2(n3089), .B(n61), .C(n62), .ZN(
        result[0]) );
  CKND2D0BWP12T U188 ( .A1(n1148), .A2(n1149), .ZN(n63) );
  MAOI22D0BWP12T U189 ( .A1(n1150), .A2(n63), .B1(n1150), .B2(n63), .ZN(n1847)
         );
  CKND0BWP12T U190 ( .I(n1808), .ZN(n64) );
  AOI21D0BWP12T U191 ( .A1(n1806), .A2(n64), .B(n1807), .ZN(n65) );
  CKND2D0BWP12T U192 ( .A1(n1809), .A2(n1810), .ZN(n66) );
  MAOI22D0BWP12T U193 ( .A1(n65), .A2(n66), .B1(n65), .B2(n66), .ZN(n2866) );
  CKND2D0BWP12T U194 ( .A1(n1672), .A2(n1674), .ZN(n67) );
  CKND2D0BWP12T U195 ( .A1(n1675), .A2(n1674), .ZN(n68) );
  OAI211D0BWP12T U196 ( .A1(n1700), .A2(n67), .B(n1673), .C(n68), .ZN(n69) );
  CKND2D0BWP12T U197 ( .A1(n1677), .A2(n1890), .ZN(n70) );
  MOAI22D0BWP12T U198 ( .A1(n69), .A2(n70), .B1(n69), .B2(n70), .ZN(n3054) );
  AOI21D0BWP12T U199 ( .A1(n1598), .A2(n1597), .B(n1596), .ZN(n71) );
  CKND2D0BWP12T U200 ( .A1(n1594), .A2(n1595), .ZN(n72) );
  MAOI22D0BWP12T U201 ( .A1(n71), .A2(n72), .B1(n71), .B2(n72), .ZN(n2865) );
  OAI21D0BWP12T U202 ( .A1(n2095), .A2(n2058), .B(n2431), .ZN(n73) );
  IAO21D0BWP12T U203 ( .A1(n2150), .A2(n2059), .B(n73), .ZN(n74) );
  OAI21D0BWP12T U204 ( .A1(n2349), .A2(n2081), .B(n74), .ZN(n2823) );
  CKND2D0BWP12T U205 ( .A1(n1516), .A2(n1517), .ZN(n75) );
  AOI21D0BWP12T U206 ( .A1(n1511), .A2(n1529), .B(n1512), .ZN(n76) );
  OAI21D0BWP12T U207 ( .A1(n1514), .A2(n76), .B(n1513), .ZN(n77) );
  MOAI22D0BWP12T U208 ( .A1(n75), .A2(n77), .B1(n75), .B2(n77), .ZN(n2815) );
  NR2D0BWP12T U209 ( .A1(n2748), .A2(n1973), .ZN(n78) );
  MOAI22D0BWP12T U210 ( .A1(n2764), .A2(n78), .B1(n2764), .B2(n78), .ZN(n2762)
         );
  OA222D0BWP12T U211 ( .A1(n2097), .A2(n2110), .B1(n2096), .B2(n2095), .C1(
        n2098), .C2(n2133), .Z(n79) );
  OA211D0BWP12T U212 ( .A1(n2099), .A2(n2150), .B(n2431), .C(n79), .Z(n2149)
         );
  CKND0BWP12T U213 ( .I(n1906), .ZN(n80) );
  AOI21D0BWP12T U214 ( .A1(n1888), .A2(n80), .B(n1891), .ZN(n81) );
  CKND2D0BWP12T U215 ( .A1(n1889), .A2(n1890), .ZN(n82) );
  MAOI22D0BWP12T U216 ( .A1(n81), .A2(n82), .B1(n81), .B2(n82), .ZN(n3062) );
  INR2D0BWP12T U217 ( .A1(n1806), .B1(n1808), .ZN(n83) );
  OAI32D0BWP12T U218 ( .A1(n1403), .A2(n1807), .A3(n83), .B1(n1810), .B2(n1403), .ZN(n84) );
  CKND2D0BWP12T U219 ( .A1(n1404), .A2(n1405), .ZN(n85) );
  MAOI22D0BWP12T U220 ( .A1(n84), .A2(n85), .B1(n84), .B2(n85), .ZN(n1758) );
  CKND0BWP12T U221 ( .I(n1700), .ZN(n86) );
  AOI21D0BWP12T U222 ( .A1(n1672), .A2(n86), .B(n1675), .ZN(n87) );
  CKND2D0BWP12T U223 ( .A1(n1673), .A2(n1674), .ZN(n88) );
  MAOI22D0BWP12T U224 ( .A1(n87), .A2(n88), .B1(n87), .B2(n88), .ZN(n2846) );
  CKND0BWP12T U225 ( .I(n2823), .ZN(n89) );
  CKND0BWP12T U226 ( .I(n2452), .ZN(n90) );
  OAI32D0BWP12T U227 ( .A1(n89), .A2(n2822), .A3(n90), .B1(n2448), .B2(n89), 
        .ZN(n2844) );
  IND2D0BWP12T U228 ( .A1(n1615), .B1(n1616), .ZN(n91) );
  MAOI22D0BWP12T U229 ( .A1(n1617), .A2(n91), .B1(n1617), .B2(n91), .ZN(n2760)
         );
  AO222D0BWP12T U230 ( .A1(n2887), .A2(n3098), .B1(n3095), .B2(n2867), .C1(
        n2866), .C2(n314), .Z(n92) );
  AO211D0BWP12T U231 ( .A1(n2886), .A2(n3115), .B(n2885), .C(n92), .Z(n93) );
  AOI211D0BWP12T U232 ( .A1(n3119), .A2(n2873), .B(n2872), .C(n93), .ZN(n94)
         );
  IOA21D0BWP12T U233 ( .A1(n2888), .A2(n3126), .B(n94), .ZN(result[11]) );
  NR2D0BWP12T U234 ( .A1(n2891), .A2(n1964), .ZN(n95) );
  MOAI22D0BWP12T U235 ( .A1(n2560), .A2(n95), .B1(n2560), .B2(n95), .ZN(n1953)
         );
  OAI21D0BWP12T U236 ( .A1(n1906), .A2(n1898), .B(n1900), .ZN(n96) );
  CKND2D0BWP12T U237 ( .A1(n1423), .A2(n1902), .ZN(n97) );
  MOAI22D0BWP12T U238 ( .A1(n96), .A2(n97), .B1(n96), .B2(n97), .ZN(n1912) );
  AOI222D0BWP12T U239 ( .A1(n2406), .A2(n2073), .B1(n2071), .B2(n3110), .C1(
        n2404), .C2(n2072), .ZN(n98) );
  OAI22D0BWP12T U240 ( .A1(n2014), .A2(n2095), .B1(n2015), .B2(n2110), .ZN(n99) );
  AOI211D0BWP12T U241 ( .A1(n2016), .A2(n2200), .B(n1388), .C(n99), .ZN(n100)
         );
  OAI21D0BWP12T U242 ( .A1(n2407), .A2(n98), .B(n100), .ZN(n2213) );
  OAI21D0BWP12T U243 ( .A1(n1808), .A2(n1803), .B(n1802), .ZN(n101) );
  CKND2D0BWP12T U244 ( .A1(n1805), .A2(n1499), .ZN(n102) );
  MOAI22D0BWP12T U245 ( .A1(n101), .A2(n102), .B1(n101), .B2(n102), .ZN(n3085)
         );
  CKND2D0BWP12T U246 ( .A1(n1599), .A2(n1600), .ZN(n103) );
  MOAI22D0BWP12T U247 ( .A1(n1601), .A2(n103), .B1(n1601), .B2(n103), .ZN(
        n2821) );
  CKND2D0BWP12T U248 ( .A1(n1853), .A2(n1849), .ZN(n104) );
  AOI21D0BWP12T U249 ( .A1(n1714), .A2(n1718), .B(n1715), .ZN(n105) );
  OAI21D0BWP12T U250 ( .A1(n1717), .A2(n105), .B(n1716), .ZN(n106) );
  MOAI22D0BWP12T U251 ( .A1(n104), .A2(n106), .B1(n104), .B2(n106), .ZN(n2795)
         );
  AOI21D0BWP12T U252 ( .A1(n1529), .A2(n1511), .B(n1512), .ZN(n107) );
  CKND2D0BWP12T U253 ( .A1(n1513), .A2(n1510), .ZN(n108) );
  MAOI22D0BWP12T U254 ( .A1(n107), .A2(n108), .B1(n107), .B2(n108), .ZN(n2787)
         );
  AOI22D0BWP12T U255 ( .A1(n3115), .A2(n2845), .B1(n2846), .B2(n3098), .ZN(
        n109) );
  INR2D0BWP12T U256 ( .A1(n2848), .B1(n3059), .ZN(n110) );
  AOI211D0BWP12T U257 ( .A1(n314), .A2(n2863), .B(n2862), .C(n110), .ZN(n111)
         );
  AOI22D1BWP12T U258 ( .A1(n2847), .A2(n3130), .B1(n3126), .B2(n2865), .ZN(
        n112) );
  CKND2D0BWP12T U259 ( .A1(n3091), .A2(n2864), .ZN(n113) );
  ND4D1BWP12T U260 ( .A1(n109), .A2(n111), .A3(n112), .A4(n113), .ZN(result[9]) );
  IND2D0BWP12T U261 ( .A1(n2207), .B1(n2750), .ZN(n114) );
  AOI222D0BWP12T U262 ( .A1(n114), .A2(n556), .B1(n2907), .B2(n2904), .C1(
        n2908), .C2(n2905), .ZN(n2223) );
  CKND2D0BWP12T U263 ( .A1(n1390), .A2(n1386), .ZN(n115) );
  MOAI22D0BWP12T U264 ( .A1(n1391), .A2(n115), .B1(n1391), .B2(n115), .ZN(
        n1525) );
  INR3D0BWP12T U265 ( .A1(n1970), .B1(n1968), .B2(n3067), .ZN(n116) );
  MOAI22D0BWP12T U266 ( .A1(n2874), .A2(n116), .B1(n2874), .B2(n116), .ZN(
        n2886) );
  CKND2D0BWP12T U267 ( .A1(n1772), .A2(n1495), .ZN(n117) );
  IOA21D0BWP12T U268 ( .A1(n1769), .A2(n1770), .B(n1768), .ZN(n118) );
  MOAI22D0BWP12T U269 ( .A1(n117), .A2(n118), .B1(n117), .B2(n118), .ZN(n2863)
         );
  CKND2D0BWP12T U270 ( .A1(n1879), .A2(n1880), .ZN(n119) );
  IOA21D0BWP12T U271 ( .A1(n1876), .A2(n1877), .B(n1875), .ZN(n120) );
  MOAI22D0BWP12T U272 ( .A1(n119), .A2(n120), .B1(n119), .B2(n120), .ZN(n2777)
         );
  CKND2D0BWP12T U273 ( .A1(n1605), .A2(n1606), .ZN(n121) );
  MOAI22D0BWP12T U274 ( .A1(n1607), .A2(n121), .B1(n1607), .B2(n121), .ZN(
        n2759) );
  OAI21D0BWP12T U275 ( .A1(n2822), .A2(n3012), .B(n3100), .ZN(n122) );
  AOI22D0BWP12T U276 ( .A1(n2823), .A2(n122), .B1(n314), .B2(n2824), .ZN(n123)
         );
  MOAI22D0BWP12T U277 ( .A1(n2826), .A2(n3044), .B1(n3095), .B2(n2825), .ZN(
        n124) );
  OAI211D0BWP12T U278 ( .A1(n2842), .A2(n2943), .B(n2841), .C(n2840), .ZN(n125) );
  AOI211D0BWP12T U279 ( .A1(n3115), .A2(n2843), .B(n124), .C(n125), .ZN(n126)
         );
  AOI22D0BWP12T U280 ( .A1(n3126), .A2(n2821), .B1(n3052), .B2(n2844), .ZN(
        n127) );
  ND3D0BWP12T U281 ( .A1(n123), .A2(n126), .A3(n127), .ZN(result[7]) );
  MOAI22D0BWP12T U282 ( .A1(n2221), .A2(n2135), .B1(n2221), .B2(n2167), .ZN(
        n128) );
  OAI21D0BWP12T U283 ( .A1(n2217), .A2(n128), .B(n2446), .ZN(n2152) );
  CKND2D0BWP12T U284 ( .A1(n1881), .A2(n548), .ZN(n129) );
  MAOI22D0BWP12T U285 ( .A1(n1906), .A2(n129), .B1(n1906), .B2(n129), .ZN(
        n1885) );
  IAO21D0BWP12T U286 ( .A1(n2406), .A2(n316), .B(n1530), .ZN(n1511) );
  CKND2D0BWP12T U287 ( .A1(n1588), .A2(n1589), .ZN(n130) );
  MOAI22D0BWP12T U288 ( .A1(n1590), .A2(n130), .B1(n1590), .B2(n130), .ZN(
        n2888) );
  CKND2D0BWP12T U289 ( .A1(n2282), .A2(n1970), .ZN(n131) );
  MAOI22D0BWP12T U290 ( .A1(n2851), .A2(n131), .B1(n2851), .B2(n131), .ZN(
        n2845) );
  OR3D0BWP12T U291 ( .A1(op[2]), .A2(op[3]), .A3(n417), .Z(n3089) );
  IND2D0BWP12T U292 ( .A1(n2851), .B1(n2282), .ZN(n1968) );
  CKND2D0BWP12T U293 ( .A1(n1509), .A2(n1785), .ZN(n132) );
  MAOI22D0BWP12T U294 ( .A1(n1538), .A2(n132), .B1(n1538), .B2(n132), .ZN(
        n2825) );
  AOI21D0BWP12T U295 ( .A1(n1877), .A2(n1850), .B(n1852), .ZN(n133) );
  CKND2D0BWP12T U296 ( .A1(n1853), .A2(n1849), .ZN(n134) );
  MAOI22D0BWP12T U297 ( .A1(n133), .A2(n134), .B1(n133), .B2(n134), .ZN(n2794)
         );
  IND2D0BWP12T U298 ( .A1(n579), .B1(n580), .ZN(n135) );
  MAOI22D0BWP12T U299 ( .A1(n581), .A2(n135), .B1(n581), .B2(n135), .ZN(n1619)
         );
  IND3D0BWP12T U300 ( .A1(n2719), .B1(n2141), .B2(n2871), .ZN(n2433) );
  IND2D0BWP12T U301 ( .A1(n2764), .B1(n2749), .ZN(n1971) );
  CKND2D0BWP12T U302 ( .A1(n1937), .A2(n800), .ZN(n136) );
  MAOI22D0BWP12T U303 ( .A1(n2406), .A2(n136), .B1(n2406), .B2(n136), .ZN(
        n1957) );
  MOAI22D0BWP12T U304 ( .A1(n2764), .A2(b[28]), .B1(n2764), .B2(b[28]), .ZN(
        n137) );
  OAI22D0BWP12T U305 ( .A1(n2514), .A2(n2513), .B1(n2512), .B2(n137), .ZN(n138) );
  MOAI22D0BWP12T U306 ( .A1(mult_x_18_n395), .A2(n138), .B1(mult_x_18_n395), 
        .B2(n138), .ZN(n139) );
  MOAI22D0BWP12T U307 ( .A1(n2720), .A2(b[18]), .B1(n2720), .B2(b[18]), .ZN(
        n140) );
  OAI22D0BWP12T U308 ( .A1(n2517), .A2(n2516), .B1(n2515), .B2(n140), .ZN(n141) );
  MOAI22D0BWP12T U309 ( .A1(n2518), .A2(n2807), .B1(n2518), .B2(n2807), .ZN(
        n142) );
  OAI22D0BWP12T U310 ( .A1(n2521), .A2(n2520), .B1(n2519), .B2(n142), .ZN(n143) );
  MOAI22D0BWP12T U311 ( .A1(n141), .A2(n143), .B1(n141), .B2(n143), .ZN(n144)
         );
  MOAI22D0BWP12T U312 ( .A1(n2657), .A2(n2522), .B1(n2657), .B2(n2522), .ZN(
        n145) );
  OAI22D0BWP12T U313 ( .A1(n2525), .A2(n2524), .B1(n2523), .B2(n145), .ZN(n146) );
  MAOI22D0BWP12T U314 ( .A1(n144), .A2(n146), .B1(n144), .B2(n146), .ZN(n147)
         );
  MAOI22D0BWP12T U315 ( .A1(n139), .A2(n147), .B1(n139), .B2(n147), .ZN(n148)
         );
  MAOI22D0BWP12T U316 ( .A1(mult_x_18_n396), .A2(n148), .B1(mult_x_18_n396), 
        .B2(n148), .ZN(n149) );
  MAOI22D0BWP12T U317 ( .A1(mult_x_18_n393), .A2(n149), .B1(mult_x_18_n393), 
        .B2(n149), .ZN(n2526) );
  CKND2D0BWP12T U318 ( .A1(n1888), .A2(n1890), .ZN(n150) );
  CKND2D0BWP12T U319 ( .A1(n1891), .A2(n1890), .ZN(n151) );
  OAI211D0BWP12T U320 ( .A1(n1906), .A2(n150), .B(n1889), .C(n151), .ZN(n152)
         );
  CKND2D0BWP12T U321 ( .A1(n1893), .A2(n1681), .ZN(n153) );
  MOAI22D0BWP12T U322 ( .A1(n152), .A2(n153), .B1(n152), .B2(n153), .ZN(n2873)
         );
  CKND2D0BWP12T U323 ( .A1(n1768), .A2(n1769), .ZN(n154) );
  MAOI22D0BWP12T U324 ( .A1(n1808), .A2(n154), .B1(n1808), .B2(n154), .ZN(
        n1801) );
  AOI21D0BWP12T U325 ( .A1(n1718), .A2(n1714), .B(n1715), .ZN(n155) );
  CKND2D0BWP12T U326 ( .A1(n1716), .A2(n1880), .ZN(n156) );
  MAOI22D0BWP12T U327 ( .A1(n155), .A2(n156), .B1(n155), .B2(n156), .ZN(n2781)
         );
  OR4D0BWP12T U328 ( .A1(n2682), .A2(n1635), .A3(n3024), .A4(n2923), .Z(n157)
         );
  NR4D0BWP12T U329 ( .A1(n2990), .A2(n2628), .A3(n2654), .A4(n157), .ZN(n158)
         );
  NR3D0BWP12T U330 ( .A1(n1640), .A2(n1641), .A3(n1660), .ZN(n159) );
  NR4D0BWP12T U331 ( .A1(n1656), .A2(n1658), .A3(n2601), .A4(n1657), .ZN(n160)
         );
  ND4D0BWP12T U332 ( .A1(n1659), .A2(n158), .A3(n159), .A4(n160), .ZN(n2481)
         );
  MOAI22D0BWP12T U333 ( .A1(a[30]), .A2(n1323), .B1(a[30]), .B2(n1323), .ZN(
        n1988) );
  INR2D0BWP12T U334 ( .A1(n1323), .B1(a[30]), .ZN(n2595) );
  INVD1BWP12T U335 ( .I(a[23]), .ZN(n2636) );
  OA21D0BWP12T U336 ( .A1(n2198), .A2(n2197), .B(n2196), .Z(n2822) );
  IND2D0BWP12T U337 ( .A1(op[2]), .B1(n1358), .ZN(n2994) );
  MAOI22D0BWP12T U338 ( .A1(n2323), .A2(n2185), .B1(n2175), .B2(n2333), .ZN(
        n1287) );
  NR4D0BWP12T U339 ( .A1(n2747), .A2(n2774), .A3(n2808), .A4(n2838), .ZN(n161)
         );
  AN4D0BWP12T U340 ( .A1(n2314), .A2(n2861), .A3(n2310), .A4(n161), .Z(n162)
         );
  CKND2D0BWP12T U341 ( .A1(n2315), .A2(n162), .ZN(n163) );
  OAI31D0BWP12T U342 ( .A1(n2881), .A2(n3077), .A3(n163), .B(n2459), .ZN(n164)
         );
  IND4D0BWP12T U343 ( .A1(n2728), .B1(n2605), .B2(n2344), .B3(n164), .ZN(n2372) );
  CKND2D0BWP12T U344 ( .A1(n1884), .A2(n1674), .ZN(n165) );
  IOA21D0BWP12T U345 ( .A1(n548), .A2(n1882), .B(n1881), .ZN(n166) );
  MOAI22D0BWP12T U346 ( .A1(n165), .A2(n166), .B1(n165), .B2(n166), .ZN(n2850)
         );
  INR3D0BWP12T U347 ( .A1(n375), .B1(n1968), .B2(n3067), .ZN(n1960) );
  AN4D0BWP12T U348 ( .A1(n2453), .A2(n2812), .A3(n2897), .A4(n2458), .Z(n167)
         );
  ND4D0BWP12T U349 ( .A1(n3101), .A2(n2751), .A3(n2668), .A4(n167), .ZN(n168)
         );
  NR3D0BWP12T U350 ( .A1(n2823), .A2(n2456), .A3(n168), .ZN(n169) );
  NR4D0BWP12T U351 ( .A1(n2864), .A2(n2685), .A3(n2164), .A4(n2163), .ZN(n170)
         );
  IAO21D0BWP12T U352 ( .A1(n2750), .A2(n3082), .B(n2715), .ZN(n171) );
  ND4D0BWP12T U353 ( .A1(n2137), .A2(n2744), .A3(n2138), .A4(n171), .ZN(n172)
         );
  NR4D0BWP12T U354 ( .A1(n3025), .A2(n2152), .A3(n2433), .A4(n172), .ZN(n173)
         );
  OAI211D0BWP12T U355 ( .A1(n2750), .A2(n169), .B(n170), .C(n173), .ZN(n2468)
         );
  MOAI22D0BWP12T U356 ( .A1(n2532), .A2(b[24]), .B1(n2532), .B2(b[24]), .ZN(
        n174) );
  OAI22D0BWP12T U357 ( .A1(n2535), .A2(n2534), .B1(n2533), .B2(n174), .ZN(n175) );
  MOAI22D0BWP12T U358 ( .A1(n2633), .A2(n3074), .B1(n2633), .B2(n3074), .ZN(
        n176) );
  OAI22D0BWP12T U359 ( .A1(n2538), .A2(n2537), .B1(n2536), .B2(n176), .ZN(n177) );
  MAOI22D0BWP12T U360 ( .A1(n175), .A2(n177), .B1(n175), .B2(n177), .ZN(n178)
         );
  MOAI22D0BWP12T U361 ( .A1(n3033), .A2(b[20]), .B1(n3033), .B2(b[20]), .ZN(
        n179) );
  OAI22D0BWP12T U362 ( .A1(n2541), .A2(n2540), .B1(n2539), .B2(n179), .ZN(n180) );
  MAOI22D0BWP12T U363 ( .A1(n178), .A2(n180), .B1(n178), .B2(n180), .ZN(n181)
         );
  MAOI22D0BWP12T U364 ( .A1(n2531), .A2(n181), .B1(n2531), .B2(n181), .ZN(n182) );
  MAOI22D0BWP12T U365 ( .A1(mult_x_18_n392), .A2(n182), .B1(mult_x_18_n392), 
        .B2(n182), .ZN(n183) );
  MAOI22D0BWP12T U366 ( .A1(mult_x_18_n383), .A2(n183), .B1(mult_x_18_n383), 
        .B2(n183), .ZN(n2579) );
  CKND2D0BWP12T U367 ( .A1(n1142), .A2(n1143), .ZN(n184) );
  MAOI22D0BWP12T U368 ( .A1(n1144), .A2(n184), .B1(n1144), .B2(n184), .ZN(
        n1546) );
  CKND2D0BWP12T U369 ( .A1(n1794), .A2(n1795), .ZN(n185) );
  MAOI22D0BWP12T U370 ( .A1(n1796), .A2(n185), .B1(n1796), .B2(n185), .ZN(n233) );
  INVD1BWP12T U371 ( .I(a[25]), .ZN(n2292) );
  INR3D0BWP12T U372 ( .A1(op[0]), .B1(op[1]), .B2(n454), .ZN(n3098) );
  OAI21D0BWP12T U373 ( .A1(n1583), .A2(n1138), .B(n1580), .ZN(n186) );
  CKND2D0BWP12T U374 ( .A1(n1139), .A2(n1140), .ZN(n187) );
  MOAI22D0BWP12T U375 ( .A1(n186), .A2(n187), .B1(n186), .B2(n187), .ZN(n1632)
         );
  OA32D0BWP12T U376 ( .A1(n1419), .A2(n2205), .A3(n2150), .B1(n2750), .B2(
        n1419), .Z(n2446) );
  OAI21D0BWP12T U377 ( .A1(n786), .A2(n783), .B(n784), .ZN(n188) );
  CKND2D0BWP12T U378 ( .A1(n616), .A2(n617), .ZN(n189) );
  MOAI22D0BWP12T U379 ( .A1(n188), .A2(n189), .B1(n188), .B2(n189), .ZN(n1874)
         );
  IND4D1BWP12T U380 ( .A1(n1971), .B1(n1955), .B2(n2802), .B3(n2831), .ZN(
        n1464) );
  AO222D0BWP12T U381 ( .A1(n3027), .A2(n314), .B1(n3026), .B2(n3098), .C1(
        n3025), .C2(n3091), .Z(n3047) );
  CKND2D0BWP12T U382 ( .A1(n1493), .A2(n1495), .ZN(n190) );
  CKND2D0BWP12T U383 ( .A1(n1496), .A2(n1495), .ZN(n191) );
  OAI211D0BWP12T U384 ( .A1(n1538), .A2(n190), .B(n1494), .C(n191), .ZN(n192)
         );
  CKND2D0BWP12T U385 ( .A1(n1498), .A2(n1499), .ZN(n193) );
  MOAI22D0BWP12T U386 ( .A1(n192), .A2(n193), .B1(n192), .B2(n193), .ZN(n3051)
         );
  IND2D0BWP12T U387 ( .A1(n426), .B1(n421), .ZN(n2980) );
  IAO21D0BWP12T U388 ( .A1(n2406), .A2(n2407), .B(n1703), .ZN(n1714) );
  INR2D0BWP12T U389 ( .A1(n3088), .B1(n3089), .ZN(n194) );
  AOI22D0BWP12T U390 ( .A1(n3090), .A2(n3091), .B1(n3092), .B2(n194), .ZN(
        n3124) );
  OA21D0BWP12T U391 ( .A1(n1383), .A2(n2262), .B(n1865), .Z(n1868) );
  OAI21D0BWP12T U392 ( .A1(n1538), .A2(n1501), .B(n1500), .ZN(n195) );
  CKND2D0BWP12T U393 ( .A1(n1502), .A2(n1810), .ZN(n196) );
  MOAI22D0BWP12T U394 ( .A1(n195), .A2(n196), .B1(n195), .B2(n196), .ZN(n2867)
         );
  CKND2D0BWP12T U395 ( .A1(n520), .A2(n1597), .ZN(n197) );
  MOAI22D0BWP12T U396 ( .A1(n1598), .A2(n197), .B1(n1598), .B2(n197), .ZN(
        n1620) );
  OAI22D0BWP12T U397 ( .A1(n2113), .A2(n2133), .B1(n2112), .B2(n2150), .ZN(
        n198) );
  AOI211D0BWP12T U398 ( .A1(n2109), .A2(n2108), .B(n2750), .C(n198), .ZN(n199)
         );
  OA21D0BWP12T U399 ( .A1(n2111), .A2(n2110), .B(n199), .Z(n2812) );
  CKND2D0BWP12T U400 ( .A1(n1767), .A2(n1510), .ZN(n200) );
  IOA21D0BWP12T U401 ( .A1(n1795), .A2(n1796), .B(n1794), .ZN(n201) );
  MOAI22D0BWP12T U402 ( .A1(n200), .A2(n201), .B1(n200), .B2(n201), .ZN(n2763)
         );
  AOI21D0BWP12T U403 ( .A1(n2750), .A2(n3103), .B(n2996), .ZN(n202) );
  OAI21D0BWP12T U404 ( .A1(n2995), .A2(n2750), .B(n202), .ZN(n203) );
  MOAI22D0BWP12T U405 ( .A1(n2749), .A2(n203), .B1(n2749), .B2(n3109), .ZN(
        n204) );
  OAI21D0BWP12T U406 ( .A1(n2748), .A2(n3066), .B(n3105), .ZN(n205) );
  AOI22D0BWP12T U407 ( .A1(n3094), .A2(n2747), .B1(n2750), .B2(n205), .ZN(n206) );
  OAI211D0BWP12T U408 ( .A1(n3100), .A2(n2751), .B(n204), .C(n206), .ZN(n2752)
         );
  INR3D0BWP12T U409 ( .A1(n1960), .B1(n1463), .B2(n1464), .ZN(n1972) );
  MUX2ND0BWP12T U410 ( .I0(n1413), .I1(n1414), .S(n2405), .ZN(n2013) );
  OAI22D0BWP12T U411 ( .A1(n2536), .A2(n1131), .B1(n2538), .B2(n1062), .ZN(
        n207) );
  MOAI22D0BWP12T U412 ( .A1(n2608), .A2(n1382), .B1(n2608), .B2(n1382), .ZN(
        n208) );
  OAI22D0BWP12T U413 ( .A1(n2546), .A2(n208), .B1(n2543), .B2(n975), .ZN(n209)
         );
  MAOI22D0BWP12T U414 ( .A1(n207), .A2(n209), .B1(n207), .B2(n209), .ZN(n210)
         );
  OAI22D0BWP12T U415 ( .A1(n2569), .A2(n1059), .B1(n2571), .B2(n862), .ZN(n211) );
  MAOI22D0BWP12T U416 ( .A1(n210), .A2(n211), .B1(n210), .B2(n211), .ZN(
        mult_x_18_n443) );
  MAOI222D0BWP12T U417 ( .A(n211), .B(n207), .C(n209), .ZN(n212) );
  CKND0BWP12T U418 ( .I(n212), .ZN(mult_x_18_n442) );
  CKND0BWP12T U419 ( .I(n2175), .ZN(n213) );
  AO222D0BWP12T U420 ( .A1(n213), .A2(n2311), .B1(n2185), .B2(n2313), .C1(
        n2187), .C2(n2312), .Z(n2216) );
  MAOI22D0BWP12T U421 ( .A1(n2389), .A2(n2388), .B1(n2431), .B2(n2838), .ZN(
        n214) );
  OAI211D0BWP12T U422 ( .A1(n2349), .A2(n2387), .B(n2390), .C(n214), .ZN(n2634) );
  CKND0BWP12T U423 ( .I(n3119), .ZN(n215) );
  AOI22D0BWP12T U424 ( .A1(n3098), .A2(n2957), .B1(n2959), .B2(n3115), .ZN(
        n216) );
  OAI21D0BWP12T U425 ( .A1(n2954), .A2(n215), .B(n216), .ZN(n217) );
  AO211D0BWP12T U426 ( .A1(n2960), .A2(n3126), .B(n2958), .C(n217), .Z(c_out)
         );
  CKND2D0BWP12T U427 ( .A1(n2956), .A2(a[30]), .ZN(n218) );
  OAI211D0BWP12T U428 ( .A1(n2956), .A2(a[30]), .B(n2548), .C(n218), .ZN(n2551) );
  CKND2D0BWP12T U429 ( .A1(n1875), .A2(n1876), .ZN(n219) );
  MOAI22D0BWP12T U430 ( .A1(n1877), .A2(n219), .B1(n1877), .B2(n219), .ZN(
        n2740) );
  AOI22D0BWP12T U431 ( .A1(n3119), .A2(n1911), .B1(n3095), .B2(n1541), .ZN(
        n220) );
  IND2D0BWP12T U432 ( .A1(n3038), .B1(n2434), .ZN(n221) );
  OAI211D0BWP12T U433 ( .A1(n2138), .A2(n3012), .B(n220), .C(n221), .ZN(n1473)
         );
  CKND0BWP12T U434 ( .I(n1538), .ZN(n222) );
  AOI21D0BWP12T U435 ( .A1(n1493), .A2(n222), .B(n1496), .ZN(n223) );
  CKND2D0BWP12T U436 ( .A1(n1494), .A2(n1495), .ZN(n224) );
  MAOI22D0BWP12T U437 ( .A1(n223), .A2(n224), .B1(n223), .B2(n224), .ZN(n2848)
         );
  OAI21D0BWP12T U438 ( .A1(n799), .A2(n795), .B(n796), .ZN(n225) );
  CKND2D0BWP12T U439 ( .A1(n604), .A2(n605), .ZN(n226) );
  MOAI22D0BWP12T U440 ( .A1(n225), .A2(n226), .B1(n225), .B2(n226), .ZN(n1799)
         );
  CKND2D0BWP12T U441 ( .A1(n765), .A2(n766), .ZN(n227) );
  MOAI22D0BWP12T U442 ( .A1(n1610), .A2(n227), .B1(n1610), .B2(n227), .ZN(
        n1613) );
  CKND0BWP12T U443 ( .I(n3095), .ZN(n228) );
  CKND0BWP12T U444 ( .I(n314), .ZN(n229) );
  OAI22D0BWP12T U445 ( .A1(n2589), .A2(n228), .B1(n2591), .B2(n229), .ZN(n2958) );
  AO222D0BWP12T U446 ( .A1(n595), .A2(n2312), .B1(n2313), .B2(n2331), .C1(
        n2334), .C2(n2311), .Z(n2774) );
  OAI21D0BWP12T U447 ( .A1(n1583), .A2(n1576), .B(n1575), .ZN(n230) );
  CKND2D0BWP12T U448 ( .A1(n1578), .A2(n1579), .ZN(n231) );
  MOAI22D0BWP12T U449 ( .A1(n230), .A2(n231), .B1(n230), .B2(n231), .ZN(n2682)
         );
  CKND2D0BWP12T U450 ( .A1(n2280), .A2(n1972), .ZN(n232) );
  MAOI22D0BWP12T U451 ( .A1(n2720), .A2(n232), .B1(n2720), .B2(n232), .ZN(
        n2716) );
  MAOI22D0BWP12T U452 ( .A1(n2349), .A2(n2013), .B1(n2133), .B2(n2205), .ZN(
        n2936) );
  CMPE42D1BWP12T U453 ( .A(mult_x_18_n767), .B(mult_x_18_n760), .C(
        mult_x_18_n787), .CIX(mult_x_18_n481), .D(mult_x_18_n947), .CO(
        mult_x_18_n456), .COX(mult_x_18_n455), .S(mult_x_18_n457) );
  NR2D2BWP12T U454 ( .A1(b[15]), .A2(n2522), .ZN(n400) );
  CMPE42D1BWP12T U455 ( .A(mult_x_18_n648), .B(mult_x_18_n636), .C(
        mult_x_18_n645), .CIX(mult_x_18_n641), .D(mult_x_18_n633), .CO(
        mult_x_18_n629), .COX(mult_x_18_n628), .S(mult_x_18_n630) );
  FA1D2BWP12T U456 ( .A(b[22]), .B(n2963), .CI(n1663), .CO(n1662), .S(n2983)
         );
  AOI21D1BWP12T U457 ( .A1(n1462), .A2(n1460), .B(n450), .ZN(n1697) );
  TPAOI21D1BWP12T U458 ( .A1(n3095), .A2(n1552), .B(n1267), .ZN(n1268) );
  CKND2D2BWP12T U459 ( .A1(n1732), .A2(n3098), .ZN(n1264) );
  INVD2BWP12T U460 ( .I(n545), .ZN(n1700) );
  OAI21D1BWP12T U461 ( .A1(n609), .A2(n442), .B(n441), .ZN(n545) );
  FA1D2BWP12T U462 ( .A(b[30]), .B(a[30]), .CI(n1324), .CO(n2952), .S(n2475)
         );
  TPOAI21D2BWP12T U463 ( .A1(n1897), .A2(n1894), .B(n1895), .ZN(n1846) );
  INVD9BWP12T U464 ( .I(n3111), .ZN(n3102) );
  FA1D2BWP12T U465 ( .A(n2608), .B(n1734), .CI(n1733), .CO(n1321), .S(n2623)
         );
  FA1D2BWP12T U466 ( .A(n1322), .B(a[30]), .CI(n1374), .CO(n2588), .S(n1552)
         );
  DCCKND4BWP12T U467 ( .I(a[11]), .ZN(n2876) );
  NR2D0BWP12T U468 ( .A1(n2253), .A2(n2874), .ZN(n1398) );
  INVD2BWP12T U469 ( .I(n2258), .ZN(n2857) );
  INVD2BWP12T U470 ( .I(n2251), .ZN(n3074) );
  BUFFD6BWP12T U471 ( .I(b[3]), .Z(n2407) );
  INVD1BWP12T U472 ( .I(n3033), .ZN(n834) );
  INVD2BWP12T U473 ( .I(n2876), .ZN(n2874) );
  INVD3BWP12T U474 ( .I(n2722), .ZN(n2720) );
  NR2D1BWP12T U475 ( .A1(n2405), .A2(n2404), .ZN(n779) );
  OR2XD1BWP12T U476 ( .A1(n2489), .A2(n2416), .Z(n1902) );
  NR2D1BWP12T U477 ( .A1(n2764), .A2(n2766), .ZN(n1717) );
  INVD1BWP12T U478 ( .I(n1383), .ZN(n1391) );
  OR2D2BWP12T U479 ( .A1(mult_x_18_n558), .A2(mult_x_18_n542), .Z(n1565) );
  CKND2D1BWP12T U480 ( .A1(n1565), .A2(n1637), .ZN(n290) );
  OR2D2BWP12T U481 ( .A1(mult_x_18_n642), .A2(mult_x_18_n630), .Z(n1140) );
  NR2D1BWP12T U482 ( .A1(mult_x_18_n643), .A2(mult_x_18_n653), .ZN(n1138) );
  INVD1BWP12T U483 ( .I(n1138), .ZN(n1581) );
  ND2D1BWP12T U484 ( .A1(n1140), .A2(n1581), .ZN(n1576) );
  NR2D1BWP12T U485 ( .A1(mult_x_18_n618), .A2(mult_x_18_n629), .ZN(n1577) );
  NR2D1BWP12T U486 ( .A1(n1576), .A2(n1577), .ZN(n283) );
  OR2D2BWP12T U487 ( .A1(mult_x_18_n654), .A2(mult_x_18_n664), .Z(n1628) );
  CKND2D1BWP12T U488 ( .A1(n1628), .A2(n1625), .ZN(n279) );
  OR2D2BWP12T U489 ( .A1(mult_x_18_n684), .A2(mult_x_18_n691), .Z(n1395) );
  CKND2D1BWP12T U490 ( .A1(n1395), .A2(n1589), .ZN(n275) );
  OR2XD1BWP12T U491 ( .A1(mult_x_18_n717), .A2(mult_x_18_n713), .Z(n1597) );
  CKND2D1BWP12T U492 ( .A1(n1595), .A2(n1597), .ZN(n271) );
  BUFFD2BWP12T U493 ( .I(a[2]), .Z(n2404) );
  INVD3BWP12T U494 ( .I(a[1]), .ZN(n3108) );
  INVD15BWP12T U495 ( .I(n3108), .ZN(n3110) );
  XNR2XD4BWP12T U496 ( .A1(n2404), .A2(n3110), .ZN(n2569) );
  INVD2BWP12T U497 ( .I(a[3]), .ZN(n757) );
  INVD6BWP12T U498 ( .I(n757), .ZN(n2406) );
  INVD3BWP12T U499 ( .I(n2406), .ZN(n378) );
  INVD4BWP12T U500 ( .I(n378), .ZN(n2567) );
  XOR2D2BWP12T U501 ( .A1(n2404), .A2(n2567), .Z(n234) );
  ND2D4BWP12T U502 ( .A1(n2569), .A2(n234), .ZN(n2571) );
  CKND4BWP12T U503 ( .I(b[2]), .ZN(n2297) );
  INVD12BWP12T U504 ( .I(n2297), .ZN(n2405) );
  BUFFD2BWP12T U505 ( .I(n2405), .Z(n2547) );
  XNR2D1BWP12T U506 ( .A1(n2547), .A2(n2567), .ZN(n240) );
  XNR2D1BWP12T U507 ( .A1(n2407), .A2(n2567), .ZN(n979) );
  OAI22D1BWP12T U508 ( .A1(n2571), .A2(n240), .B1(n2569), .B2(n979), .ZN(n261)
         );
  INVD3BWP12T U509 ( .I(a[5]), .ZN(n2768) );
  INVD9BWP12T U510 ( .I(n2768), .ZN(n2764) );
  BUFFD2BWP12T U511 ( .I(a[4]), .Z(n2748) );
  XOR2XD1BWP12T U512 ( .A1(n2764), .A2(n2748), .Z(n235) );
  XOR2XD4BWP12T U513 ( .A1(n2748), .A2(n378), .Z(n2512) );
  ND2D4BWP12T U514 ( .A1(n235), .A2(n2512), .ZN(n2514) );
  INVD9BWP12T U515 ( .I(n2422), .ZN(n1383) );
  BUFFXD4BWP12T U516 ( .I(n1383), .Z(n1382) );
  XNR2D1BWP12T U517 ( .A1(n2764), .A2(n1382), .ZN(n236) );
  INVD3BWP12T U518 ( .I(b[1]), .ZN(n3111) );
  XNR2D1BWP12T U519 ( .A1(n2764), .A2(n3102), .ZN(n880) );
  OAI22D1BWP12T U520 ( .A1(n2514), .A2(n236), .B1(n880), .B2(n2512), .ZN(n260)
         );
  BUFFD2BWP12T U521 ( .I(a[0]), .Z(n2262) );
  INVD8BWP12T U522 ( .I(n2262), .ZN(n2486) );
  CKND2D2BWP12T U523 ( .A1(n3110), .A2(n2486), .ZN(n2487) );
  INVD2BWP12T U524 ( .I(b[4]), .ZN(n386) );
  BUFFD2BWP12T U525 ( .I(n2750), .Z(n2542) );
  XNR2XD1BWP12T U526 ( .A1(n2542), .A2(n3110), .ZN(n239) );
  INVD1P75BWP12T U527 ( .I(b[5]), .ZN(n2261) );
  XNR2XD1BWP12T U528 ( .A1(n2766), .A2(n3110), .ZN(n911) );
  OAI22D1BWP12T U529 ( .A1(n2487), .A2(n239), .B1(n911), .B2(n2486), .ZN(n824)
         );
  CKND0BWP12T U530 ( .I(n2764), .ZN(n238) );
  CKBD1BWP12T U531 ( .I(n1383), .Z(n1064) );
  IND2D0BWP12T U532 ( .A1(n1064), .B1(n2764), .ZN(n237) );
  OAI22D1BWP12T U533 ( .A1(n2514), .A2(n238), .B1(n2512), .B2(n237), .ZN(n823)
         );
  NR2D1BWP12T U534 ( .A1(mult_x_18_n723), .A2(n267), .ZN(n1602) );
  XNR2XD1BWP12T U535 ( .A1(n2407), .A2(n3110), .ZN(n241) );
  OAI22D1BWP12T U536 ( .A1(n2487), .A2(n241), .B1(n239), .B2(n2486), .ZN(n264)
         );
  INR2D1BWP12T U537 ( .A1(n1382), .B1(n2512), .ZN(n263) );
  XNR2D1BWP12T U538 ( .A1(n3102), .A2(n2567), .ZN(n242) );
  OAI22D1BWP12T U539 ( .A1(n2571), .A2(n242), .B1(n2569), .B2(n240), .ZN(n262)
         );
  XNR2D1BWP12T U540 ( .A1(n2547), .A2(n3110), .ZN(n247) );
  OAI22D1BWP12T U541 ( .A1(n2487), .A2(n247), .B1(n241), .B2(n2486), .ZN(n245)
         );
  XNR2D1BWP12T U542 ( .A1(n1382), .A2(n2567), .ZN(n243) );
  OAI22D1BWP12T U543 ( .A1(n2571), .A2(n243), .B1(n2569), .B2(n242), .ZN(n244)
         );
  OR2XD1BWP12T U544 ( .A1(n257), .A2(n256), .Z(n1606) );
  IND2XD0BWP12T U545 ( .A1(n1064), .B1(n2567), .ZN(n246) );
  OAI22D1BWP12T U546 ( .A1(n2571), .A2(n378), .B1(n2569), .B2(n246), .ZN(n254)
         );
  NR2D1BWP12T U547 ( .A1(n255), .A2(n254), .ZN(n579) );
  CKBD1BWP12T U548 ( .I(n3102), .Z(n998) );
  XNR2XD1BWP12T U549 ( .A1(n998), .A2(n3110), .ZN(n249) );
  OAI22D1BWP12T U550 ( .A1(n2487), .A2(n249), .B1(n247), .B2(n2486), .ZN(n252)
         );
  INR2D1BWP12T U551 ( .A1(n1382), .B1(n2569), .ZN(n251) );
  OR2XD1BWP12T U552 ( .A1(n252), .A2(n251), .Z(n766) );
  IND2D0BWP12T U553 ( .A1(n1064), .B1(n3110), .ZN(n248) );
  ND2D1BWP12T U554 ( .A1(n248), .A2(n2487), .ZN(n1608) );
  OAI22D1BWP12T U555 ( .A1(n2487), .A2(n1382), .B1(n249), .B2(n2486), .ZN(
        n1609) );
  INVD1BWP12T U556 ( .I(n1609), .ZN(n250) );
  INR2D1BWP12T U557 ( .A1(n1608), .B1(n250), .ZN(n1610) );
  ND2D1BWP12T U558 ( .A1(n252), .A2(n251), .ZN(n765) );
  INVD1BWP12T U559 ( .I(n765), .ZN(n253) );
  AOI21D1BWP12T U560 ( .A1(n766), .A2(n1610), .B(n253), .ZN(n581) );
  ND2D1BWP12T U561 ( .A1(n255), .A2(n254), .ZN(n580) );
  OAI21D1BWP12T U562 ( .A1(n579), .A2(n581), .B(n580), .ZN(n1607) );
  ND2D1BWP12T U563 ( .A1(n257), .A2(n256), .ZN(n1605) );
  INVD1BWP12T U564 ( .I(n1605), .ZN(n258) );
  AOI21D1BWP12T U565 ( .A1(n1606), .A2(n1607), .B(n258), .ZN(n1617) );
  FA1D0BWP12T U566 ( .A(n261), .B(n260), .CI(n259), .CO(n267), .S(n266) );
  FA1D0BWP12T U567 ( .A(n264), .B(n263), .CI(n262), .CO(n265), .S(n257) );
  NR2D1BWP12T U568 ( .A1(n266), .A2(n265), .ZN(n1615) );
  ND2D1BWP12T U569 ( .A1(n266), .A2(n265), .ZN(n1616) );
  OA21D1BWP12T U570 ( .A1(n1617), .A2(n1615), .B(n1616), .Z(n1604) );
  ND2D1BWP12T U571 ( .A1(mult_x_18_n723), .A2(n267), .ZN(n1603) );
  OAI21D1BWP12T U572 ( .A1(n1602), .A2(n1604), .B(n1603), .ZN(n1601) );
  OR2D1BWP12T U573 ( .A1(mult_x_18_n718), .A2(mult_x_18_n722), .Z(n1600) );
  ND2D1BWP12T U574 ( .A1(mult_x_18_n718), .A2(mult_x_18_n722), .ZN(n1599) );
  INVD1BWP12T U575 ( .I(n1599), .ZN(n268) );
  AOI21D1BWP12T U576 ( .A1(n1601), .A2(n1600), .B(n268), .ZN(n519) );
  ND2D1BWP12T U577 ( .A1(mult_x_18_n717), .A2(mult_x_18_n713), .ZN(n520) );
  INVD1BWP12T U578 ( .I(n520), .ZN(n1596) );
  ND2D1BWP12T U579 ( .A1(mult_x_18_n706), .A2(mult_x_18_n712), .ZN(n1594) );
  INVD1BWP12T U580 ( .I(n1594), .ZN(n269) );
  AOI21D1BWP12T U581 ( .A1(n1595), .A2(n1596), .B(n269), .ZN(n270) );
  OAI21D1BWP12T U582 ( .A1(n271), .A2(n519), .B(n270), .ZN(n1593) );
  OR2D1BWP12T U583 ( .A1(mult_x_18_n700), .A2(mult_x_18_n705), .Z(n1592) );
  ND2D1BWP12T U584 ( .A1(mult_x_18_n700), .A2(mult_x_18_n705), .ZN(n1591) );
  INVD1BWP12T U585 ( .I(n1591), .ZN(n272) );
  AOI21D1BWP12T U586 ( .A1(n1593), .A2(n1592), .B(n272), .ZN(n1392) );
  ND2D1BWP12T U587 ( .A1(mult_x_18_n692), .A2(mult_x_18_n699), .ZN(n1588) );
  INVD1BWP12T U588 ( .I(n1588), .ZN(n1393) );
  ND2D1BWP12T U589 ( .A1(mult_x_18_n684), .A2(mult_x_18_n691), .ZN(n1394) );
  INVD1BWP12T U590 ( .I(n1394), .ZN(n273) );
  AOI21D1BWP12T U591 ( .A1(n1395), .A2(n1393), .B(n273), .ZN(n274) );
  OAI21D1BWP12T U592 ( .A1(n275), .A2(n1392), .B(n274), .ZN(n1586) );
  ND2D1BWP12T U593 ( .A1(mult_x_18_n674), .A2(mult_x_18_n683), .ZN(n1584) );
  INVD1BWP12T U594 ( .I(n1584), .ZN(n276) );
  TPAOI21D1BWP12T U595 ( .A1(n1586), .A2(n1585), .B(n276), .ZN(n1437) );
  ND2D1BWP12T U596 ( .A1(mult_x_18_n673), .A2(mult_x_18_n665), .ZN(n1438) );
  INVD1BWP12T U597 ( .I(n1438), .ZN(n1624) );
  ND2D1BWP12T U598 ( .A1(mult_x_18_n654), .A2(mult_x_18_n664), .ZN(n1627) );
  INVD1BWP12T U599 ( .I(n1627), .ZN(n277) );
  AOI21D1BWP12T U600 ( .A1(n1628), .A2(n1624), .B(n277), .ZN(n278) );
  OAI21D1BWP12T U601 ( .A1(n279), .A2(n1437), .B(n278), .ZN(n1137) );
  ND2D1BWP12T U602 ( .A1(mult_x_18_n643), .A2(mult_x_18_n653), .ZN(n1580) );
  CKND1BWP12T U603 ( .I(n1580), .ZN(n281) );
  ND2D1BWP12T U604 ( .A1(mult_x_18_n642), .A2(mult_x_18_n630), .ZN(n1139) );
  INVD1BWP12T U605 ( .I(n1139), .ZN(n280) );
  AOI21D1BWP12T U606 ( .A1(n1140), .A2(n281), .B(n280), .ZN(n1575) );
  ND2D1BWP12T U607 ( .A1(mult_x_18_n618), .A2(mult_x_18_n629), .ZN(n1578) );
  OAI21D1BWP12T U608 ( .A1(n1575), .A2(n1577), .B(n1578), .ZN(n282) );
  AOI21D1BWP12T U609 ( .A1(n283), .A2(n1137), .B(n282), .ZN(n1555) );
  OR2XD1BWP12T U610 ( .A1(mult_x_18_n604), .A2(mult_x_18_n617), .Z(n1569) );
  CKND2D1BWP12T U611 ( .A1(n1572), .A2(n1569), .ZN(n286) );
  ND2D1BWP12T U612 ( .A1(mult_x_18_n604), .A2(mult_x_18_n617), .ZN(n1556) );
  INVD1BWP12T U613 ( .I(n1556), .ZN(n1568) );
  ND2D1BWP12T U614 ( .A1(mult_x_18_n590), .A2(mult_x_18_n603), .ZN(n1571) );
  INVD1BWP12T U615 ( .I(n1571), .ZN(n284) );
  AOI21D1BWP12T U616 ( .A1(n1572), .A2(n1568), .B(n284), .ZN(n285) );
  OR2D1BWP12T U617 ( .A1(mult_x_18_n574), .A2(mult_x_18_n589), .Z(n1559) );
  ND2D1BWP12T U618 ( .A1(mult_x_18_n574), .A2(mult_x_18_n589), .ZN(n1558) );
  INVD1BWP12T U619 ( .I(n1558), .ZN(n287) );
  AOI21D1BWP12T U620 ( .A1(n1561), .A2(n1559), .B(n287), .ZN(n1562) );
  ND2D1BWP12T U621 ( .A1(mult_x_18_n559), .A2(mult_x_18_n573), .ZN(n1636) );
  INVD1BWP12T U622 ( .I(n1636), .ZN(n1563) );
  ND2D1BWP12T U623 ( .A1(mult_x_18_n558), .A2(mult_x_18_n542), .ZN(n1564) );
  INVD1BWP12T U624 ( .I(n1564), .ZN(n288) );
  TPAOI21D1BWP12T U625 ( .A1(n1565), .A2(n1563), .B(n288), .ZN(n289) );
  TPNR2D1BWP12T U626 ( .A1(mult_x_18_n506), .A2(mult_x_18_n524), .ZN(n1272) );
  NR2D1BWP12T U627 ( .A1(mult_x_18_n525), .A2(mult_x_18_n541), .ZN(n1270) );
  NR2D1BWP12T U628 ( .A1(n1272), .A2(n1270), .ZN(n292) );
  ND2D1BWP12T U629 ( .A1(mult_x_18_n525), .A2(mult_x_18_n541), .ZN(n1269) );
  ND2D1BWP12T U630 ( .A1(mult_x_18_n506), .A2(mult_x_18_n524), .ZN(n1273) );
  OAI21D1BWP12T U631 ( .A1(n1272), .A2(n1269), .B(n1273), .ZN(n291) );
  TPAOI21D1BWP12T U632 ( .A1(n699), .A2(n292), .B(n291), .ZN(n1202) );
  INVD1P75BWP12T U633 ( .I(n1202), .ZN(n1650) );
  NR2D1BWP12T U634 ( .A1(mult_x_18_n505), .A2(mult_x_18_n488), .ZN(n643) );
  INVD1BWP12T U635 ( .I(n643), .ZN(n467) );
  ND2D1BWP12T U636 ( .A1(mult_x_18_n505), .A2(mult_x_18_n488), .ZN(n645) );
  INVD1BWP12T U637 ( .I(n645), .ZN(n293) );
  AOI21D1BWP12T U638 ( .A1(n1650), .A2(n467), .B(n293), .ZN(n296) );
  TPNR2D1BWP12T U639 ( .A1(mult_x_18_n487), .A2(mult_x_18_n468), .ZN(n646) );
  INVD1BWP12T U640 ( .I(n646), .ZN(n294) );
  ND2D1BWP12T U641 ( .A1(mult_x_18_n487), .A2(mult_x_18_n468), .ZN(n644) );
  ND2D1BWP12T U642 ( .A1(n294), .A2(n644), .ZN(n295) );
  XOR2XD1BWP12T U643 ( .A1(n296), .A2(n295), .Z(n1658) );
  ND2D1BWP12T U644 ( .A1(op[3]), .A2(op[0]), .ZN(n426) );
  INR3D2BWP12T U645 ( .A1(op[2]), .B1(op[1]), .B2(n426), .ZN(n3126) );
  IND2XD1BWP12T U646 ( .A1(op[3]), .B1(op[2]), .ZN(n454) );
  IND2D1BWP12T U647 ( .A1(op[0]), .B1(op[1]), .ZN(n423) );
  NR2D2BWP12T U648 ( .A1(n454), .A2(n423), .ZN(n3095) );
  INVD1BWP12T U649 ( .I(a[27]), .ZN(n2291) );
  INVD2BWP12T U650 ( .I(n2291), .ZN(n2518) );
  INVD4BWP12T U651 ( .I(n2292), .ZN(n2502) );
  INVD3BWP12T U652 ( .I(n2636), .ZN(n2633) );
  INVD2BWP12T U653 ( .I(a[21]), .ZN(n2998) );
  INVD1P75BWP12T U654 ( .I(n2405), .ZN(n315) );
  NR2D1BWP12T U655 ( .A1(n315), .A2(n2404), .ZN(n774) );
  CKND1BWP12T U656 ( .I(n3102), .ZN(n298) );
  CKBD1BWP12T U657 ( .I(n3110), .Z(n297) );
  NR2D1BWP12T U658 ( .A1(n298), .A2(n297), .ZN(n1520) );
  TPNR2D0BWP12T U659 ( .A1(n774), .A2(n1520), .ZN(n300) );
  NR2D1BWP12T U660 ( .A1(n2262), .A2(c_in), .ZN(n1389) );
  CKND2D1BWP12T U661 ( .A1(n2262), .A2(c_in), .ZN(n1390) );
  TPOAI21D0BWP12T U662 ( .A1(n1383), .A2(n1389), .B(n1390), .ZN(n773) );
  ND2D1BWP12T U663 ( .A1(n298), .A2(n297), .ZN(n1521) );
  CKND2D1BWP12T U664 ( .A1(n315), .A2(n2404), .ZN(n775) );
  OAI21D1BWP12T U665 ( .A1(n774), .A2(n1521), .B(n775), .ZN(n299) );
  AOI21D1BWP12T U666 ( .A1(n300), .A2(n773), .B(n299), .ZN(n606) );
  INVD1P75BWP12T U667 ( .I(n2407), .ZN(n316) );
  NR2D1BWP12T U668 ( .A1(n319), .A2(n2748), .ZN(n1530) );
  INVD1P75BWP12T U669 ( .I(n2766), .ZN(n320) );
  CKBD1BWP12T U670 ( .I(n2764), .Z(n301) );
  NR2D1BWP12T U671 ( .A1(n320), .A2(n301), .ZN(n1514) );
  INVD4BWP12T U672 ( .I(n2259), .ZN(n2807) );
  BUFFD2BWP12T U673 ( .I(a[6]), .Z(n2799) );
  NR2D1BWP12T U674 ( .A1(n321), .A2(n2799), .ZN(n1515) );
  NR2D1BWP12T U675 ( .A1(n1514), .A2(n1515), .ZN(n303) );
  CKND2D1BWP12T U676 ( .A1(n1511), .A2(n303), .ZN(n305) );
  CKND2D1BWP12T U677 ( .A1(n316), .A2(n2406), .ZN(n1527) );
  CKND2D1BWP12T U678 ( .A1(n319), .A2(n2748), .ZN(n1531) );
  OAI21D1BWP12T U679 ( .A1(n1530), .A2(n1527), .B(n1531), .ZN(n1512) );
  ND2D1BWP12T U680 ( .A1(n320), .A2(n301), .ZN(n1513) );
  CKND2D1BWP12T U681 ( .A1(n321), .A2(n2799), .ZN(n1516) );
  OAI21D1BWP12T U682 ( .A1(n1515), .A2(n1513), .B(n1516), .ZN(n302) );
  AOI21D1BWP12T U683 ( .A1(n1512), .A2(n303), .B(n302), .ZN(n304) );
  OAI21D1BWP12T U684 ( .A1(n606), .A2(n305), .B(n304), .ZN(n559) );
  INVD1P75BWP12T U685 ( .I(b[7]), .ZN(n2260) );
  INVD4BWP12T U686 ( .I(n2260), .ZN(n2829) );
  CKBD1BWP12T U687 ( .I(a[7]), .Z(n306) );
  NR2D1BWP12T U688 ( .A1(n323), .A2(n306), .ZN(n557) );
  INVD1BWP12T U689 ( .I(b[8]), .ZN(n2252) );
  BUFFD2BWP12T U690 ( .I(a[8]), .Z(n2398) );
  NR2D1BWP12T U691 ( .A1(n328), .A2(n2398), .ZN(n560) );
  NR2D1BWP12T U692 ( .A1(n557), .A2(n560), .ZN(n1493) );
  INVD1BWP12T U693 ( .I(b[9]), .ZN(n2258) );
  INVD3BWP12T U694 ( .I(a[9]), .ZN(n2853) );
  INVD8BWP12T U695 ( .I(n2853), .ZN(n2851) );
  NR2D1BWP12T U696 ( .A1(n2258), .A2(n2851), .ZN(n1492) );
  INVD1BWP12T U697 ( .I(b[10]), .ZN(n2251) );
  NR2D1BWP12T U698 ( .A1(n2251), .A2(n3067), .ZN(n1497) );
  NR2D1BWP12T U699 ( .A1(n1492), .A2(n1497), .ZN(n308) );
  ND2D1BWP12T U700 ( .A1(n1493), .A2(n308), .ZN(n1501) );
  BUFFD6BWP12T U701 ( .I(b[11]), .Z(n2880) );
  INVD3BWP12T U702 ( .I(n2880), .ZN(n2253) );
  BUFFD3BWP12T U703 ( .I(b[12]), .Z(n2489) );
  INVD1P75BWP12T U704 ( .I(n2489), .ZN(n2249) );
  BUFFD2BWP12T U705 ( .I(a[12]), .Z(n2416) );
  NR2D1BWP12T U706 ( .A1(n2249), .A2(n2416), .ZN(n1399) );
  NR2D1BWP12T U707 ( .A1(n1398), .A2(n1399), .ZN(n1536) );
  INVD1P75BWP12T U708 ( .I(b[13]), .ZN(n2250) );
  INVD2BWP12T U709 ( .I(a[13]), .ZN(n3031) );
  INVD3BWP12T U710 ( .I(n3031), .ZN(n3033) );
  OR2XD1BWP12T U711 ( .A1(n2250), .A2(n3033), .Z(n1540) );
  CKND2D1BWP12T U712 ( .A1(n1536), .A2(n1540), .ZN(n311) );
  OR2XD1BWP12T U713 ( .A1(n1501), .A2(n311), .Z(n313) );
  ND2D1BWP12T U714 ( .A1(n323), .A2(n306), .ZN(n1509) );
  CKND2D1BWP12T U715 ( .A1(n328), .A2(n2398), .ZN(n561) );
  OAI21D1BWP12T U716 ( .A1(n560), .A2(n1509), .B(n561), .ZN(n1496) );
  CKND2D1BWP12T U717 ( .A1(n2258), .A2(n2851), .ZN(n1494) );
  CKND2D1BWP12T U718 ( .A1(n2251), .A2(n3067), .ZN(n1498) );
  OAI21D1BWP12T U719 ( .A1(n1497), .A2(n1494), .B(n1498), .ZN(n307) );
  AOI21D1BWP12T U720 ( .A1(n308), .A2(n1496), .B(n307), .ZN(n1500) );
  ND2D1BWP12T U721 ( .A1(n2253), .A2(n2874), .ZN(n1502) );
  CKND2D1BWP12T U722 ( .A1(n2249), .A2(n2416), .ZN(n1400) );
  OAI21D1BWP12T U723 ( .A1(n1399), .A2(n1502), .B(n1400), .ZN(n1535) );
  CKND2D1BWP12T U724 ( .A1(n2250), .A2(n3033), .ZN(n1539) );
  INVD1BWP12T U725 ( .I(n1539), .ZN(n309) );
  AOI21D1BWP12T U726 ( .A1(n1535), .A2(n1540), .B(n309), .ZN(n310) );
  OA21D1BWP12T U727 ( .A1(n1500), .A2(n311), .B(n310), .Z(n312) );
  OR2XD1BWP12T U728 ( .A1(n2247), .A2(a[14]), .Z(n1453) );
  CKND2D1BWP12T U729 ( .A1(n2247), .A2(a[14]), .ZN(n1452) );
  AOI21D1BWP12T U730 ( .A1(n1455), .A2(n1453), .B(n336), .ZN(n1508) );
  INVD1BWP12T U731 ( .I(b[15]), .ZN(n2248) );
  INVD2BWP12T U732 ( .I(a[15]), .ZN(n2722) );
  TPNR2D0BWP12T U733 ( .A1(n2248), .A2(n2720), .ZN(n1504) );
  CKND2D1BWP12T U734 ( .A1(n2248), .A2(n2720), .ZN(n1505) );
  OAI21D1BWP12T U735 ( .A1(n1508), .A2(n1504), .B(n1505), .ZN(n1545) );
  INVD1BWP12T U736 ( .I(b[16]), .ZN(n2241) );
  OR2XD1BWP12T U737 ( .A1(n2241), .A2(n2891), .Z(n1543) );
  CKND2D1BWP12T U738 ( .A1(n2241), .A2(n2891), .ZN(n1542) );
  AOI21D1BWP12T U739 ( .A1(n1545), .A2(n1543), .B(n337), .ZN(n1144) );
  INVD1BWP12T U740 ( .I(b[17]), .ZN(n2246) );
  INVD2BWP12T U741 ( .I(a[17]), .ZN(n2275) );
  INVD6BWP12T U742 ( .I(n2275), .ZN(n2560) );
  NR2XD0BWP12T U743 ( .A1(n2246), .A2(n2560), .ZN(n1141) );
  CKND2D1BWP12T U744 ( .A1(n2246), .A2(n2560), .ZN(n1142) );
  OAI21D1BWP12T U745 ( .A1(n1144), .A2(n1141), .B(n1142), .ZN(n1491) );
  INVD1BWP12T U746 ( .I(b[18]), .ZN(n2239) );
  OR2XD1BWP12T U747 ( .A1(n2239), .A2(n2689), .Z(n1489) );
  CKND2D1BWP12T U748 ( .A1(n2239), .A2(n2689), .ZN(n1488) );
  BUFFD2BWP12T U749 ( .I(b[19]), .Z(n2663) );
  INVD1BWP12T U750 ( .I(n2663), .ZN(n2240) );
  NR2D1BWP12T U751 ( .A1(n2240), .A2(n2657), .ZN(n1483) );
  ND2D1BWP12T U752 ( .A1(n2240), .A2(n2657), .ZN(n1484) );
  INVD1BWP12T U753 ( .I(b[20]), .ZN(n2238) );
  OR2XD1BWP12T U754 ( .A1(n2238), .A2(a[20]), .Z(n1480) );
  ND2D1BWP12T U755 ( .A1(n2238), .A2(a[20]), .ZN(n1479) );
  AO21D1BWP12T U756 ( .A1(n1482), .A2(n1480), .B(n339), .Z(n1547) );
  INR2D1BWP12T U757 ( .A1(op[1]), .B1(op[2]), .ZN(n358) );
  INR2D1BWP12T U758 ( .A1(op[3]), .B1(n383), .ZN(n314) );
  INVD1BWP12T U759 ( .I(n314), .ZN(n3020) );
  INVD1BWP12T U760 ( .I(b[27]), .ZN(n651) );
  CKND0BWP12T U761 ( .I(b[26]), .ZN(n471) );
  INVD1BWP12T U762 ( .I(b[25]), .ZN(n1279) );
  INVD1BWP12T U763 ( .I(b[24]), .ZN(n703) );
  INVD1BWP12T U764 ( .I(b[23]), .ZN(n1736) );
  INVD1BWP12T U765 ( .I(b[22]), .ZN(n1821) );
  NR2D1BWP12T U766 ( .A1(n1391), .A2(n2262), .ZN(n1790) );
  NR2D1BWP12T U767 ( .A1(n298), .A2(n3110), .ZN(n1788) );
  CKND2D1BWP12T U768 ( .A1(n298), .A2(n3110), .ZN(n1789) );
  OAI21D1BWP12T U769 ( .A1(n1790), .A2(n1788), .B(n1789), .ZN(n602) );
  NR2D1BWP12T U770 ( .A1(n316), .A2(n2406), .ZN(n603) );
  NR2D1BWP12T U771 ( .A1(n315), .A2(n2404), .ZN(n795) );
  NR2D1BWP12T U772 ( .A1(n603), .A2(n795), .ZN(n318) );
  CKND2D1BWP12T U773 ( .A1(n315), .A2(n2404), .ZN(n796) );
  CKND2D1BWP12T U774 ( .A1(n316), .A2(n2406), .ZN(n604) );
  OAI21D1BWP12T U775 ( .A1(n603), .A2(n796), .B(n604), .ZN(n317) );
  AOI21D1BWP12T U776 ( .A1(n602), .A2(n318), .B(n317), .ZN(n1764) );
  NR2D1BWP12T U777 ( .A1(n319), .A2(n2748), .ZN(n1765) );
  NR2D1BWP12T U778 ( .A1(n320), .A2(n2764), .ZN(n1766) );
  NR2D1BWP12T U779 ( .A1(n1765), .A2(n1766), .ZN(n1775) );
  CKBD1BWP12T U780 ( .I(a[7]), .Z(n322) );
  NR2D1BWP12T U781 ( .A1(n323), .A2(n322), .ZN(n1783) );
  NR2D1BWP12T U782 ( .A1(n321), .A2(n2799), .ZN(n1779) );
  NR2D1BWP12T U783 ( .A1(n1783), .A2(n1779), .ZN(n325) );
  CKND2D1BWP12T U784 ( .A1(n1775), .A2(n325), .ZN(n327) );
  CKND2D1BWP12T U785 ( .A1(n319), .A2(n2748), .ZN(n1794) );
  CKND2D1BWP12T U786 ( .A1(n320), .A2(n2764), .ZN(n1767) );
  OAI21D1BWP12T U787 ( .A1(n1794), .A2(n1766), .B(n1767), .ZN(n1777) );
  CKND2D1BWP12T U788 ( .A1(n321), .A2(n2799), .ZN(n1778) );
  ND2D1BWP12T U789 ( .A1(n323), .A2(n322), .ZN(n1784) );
  OAI21D1BWP12T U790 ( .A1(n1783), .A2(n1778), .B(n1784), .ZN(n324) );
  AOI21D1BWP12T U791 ( .A1(n1777), .A2(n325), .B(n324), .ZN(n326) );
  OAI21D1BWP12T U792 ( .A1(n1764), .A2(n327), .B(n326), .ZN(n1770) );
  INVD1P75BWP12T U793 ( .I(n1770), .ZN(n1808) );
  OR2D2BWP12T U794 ( .A1(n2253), .A2(n2874), .Z(n1810) );
  ND2D1BWP12T U795 ( .A1(n1810), .A2(n1405), .ZN(n331) );
  NR2D1BWP12T U796 ( .A1(n2251), .A2(n3067), .ZN(n1804) );
  NR2D1BWP12T U797 ( .A1(n2258), .A2(n2851), .ZN(n1771) );
  NR2D1BWP12T U798 ( .A1(n328), .A2(n2398), .ZN(n553) );
  NR2D1BWP12T U799 ( .A1(n1771), .A2(n553), .ZN(n1401) );
  ND2D1BWP12T U800 ( .A1(n333), .A2(n1401), .ZN(n1753) );
  NR2D1BWP12T U801 ( .A1(n2250), .A2(n3033), .ZN(n1754) );
  CKND2D1BWP12T U802 ( .A1(n328), .A2(n2398), .ZN(n1768) );
  CKND2D1BWP12T U803 ( .A1(n2258), .A2(n2851), .ZN(n1772) );
  OAI21D1BWP12T U804 ( .A1(n1771), .A2(n1768), .B(n1772), .ZN(n1402) );
  ND2D1BWP12T U805 ( .A1(n2251), .A2(n3067), .ZN(n1805) );
  ND2D1BWP12T U806 ( .A1(n2253), .A2(n2874), .ZN(n1809) );
  INVD1BWP12T U807 ( .I(n1809), .ZN(n1403) );
  ND2D1BWP12T U808 ( .A1(n2249), .A2(n2416), .ZN(n1404) );
  INVD1BWP12T U809 ( .I(n1404), .ZN(n329) );
  AOI21D1BWP12T U810 ( .A1(n1405), .A2(n1403), .B(n329), .ZN(n330) );
  OAI21D1BWP12T U811 ( .A1(n331), .A2(n1805), .B(n330), .ZN(n332) );
  TPAOI21D1BWP12T U812 ( .A1(n333), .A2(n1402), .B(n332), .ZN(n1752) );
  ND2D1BWP12T U813 ( .A1(n2250), .A2(n3033), .ZN(n1755) );
  OA21D1BWP12T U814 ( .A1(n1752), .A2(n1754), .B(n1755), .Z(n334) );
  TPOAI21D1BWP12T U815 ( .A1(n1808), .A2(n335), .B(n334), .ZN(n1443) );
  OR2XD1BWP12T U816 ( .A1(n2247), .A2(a[14]), .Z(n1441) );
  ND2D1BWP12T U817 ( .A1(n2247), .A2(a[14]), .ZN(n1440) );
  INVD1BWP12T U818 ( .I(n1440), .ZN(n336) );
  TPAOI21D1BWP12T U819 ( .A1(n1443), .A2(n1441), .B(n336), .ZN(n1763) );
  NR2D1BWP12T U820 ( .A1(n2248), .A2(n2720), .ZN(n1760) );
  ND2D1BWP12T U821 ( .A1(n2248), .A2(n2720), .ZN(n1761) );
  TPOAI21D1BWP12T U822 ( .A1(n1763), .A2(n1760), .B(n1761), .ZN(n1751) );
  OR2XD1BWP12T U823 ( .A1(n2241), .A2(n2891), .Z(n1749) );
  ND2D1BWP12T U824 ( .A1(n2241), .A2(n2891), .ZN(n1748) );
  INVD1BWP12T U825 ( .I(n1748), .ZN(n337) );
  TPAOI21D1BWP12T U826 ( .A1(n1751), .A2(n1749), .B(n337), .ZN(n1194) );
  NR2D1BWP12T U827 ( .A1(n2246), .A2(n2560), .ZN(n1192) );
  ND2D1BWP12T U828 ( .A1(n2246), .A2(n2560), .ZN(n1193) );
  TPOAI21D1BWP12T U829 ( .A1(n1194), .A2(n1192), .B(n1193), .ZN(n1747) );
  OR2XD1BWP12T U830 ( .A1(n2239), .A2(n2689), .Z(n1745) );
  ND2D1BWP12T U831 ( .A1(n2239), .A2(n2689), .ZN(n1744) );
  INVD1BWP12T U832 ( .I(n1744), .ZN(n338) );
  NR2D1BWP12T U833 ( .A1(n2240), .A2(n2657), .ZN(n1814) );
  ND2D1BWP12T U834 ( .A1(n2240), .A2(n2657), .ZN(n1815) );
  TPOAI21D1BWP12T U835 ( .A1(n1817), .A2(n1814), .B(n1815), .ZN(n1743) );
  OR2XD1BWP12T U836 ( .A1(n2238), .A2(a[20]), .Z(n1741) );
  CKND2D1BWP12T U837 ( .A1(n2238), .A2(a[20]), .ZN(n1740) );
  INVD1BWP12T U838 ( .I(n1740), .ZN(n339) );
  TPAOI21D1BWP12T U839 ( .A1(n1743), .A2(n1741), .B(n339), .ZN(n1739) );
  INVD1BWP12T U840 ( .I(b[21]), .ZN(n340) );
  NR2XD0BWP12T U841 ( .A1(n340), .A2(n2993), .ZN(n1737) );
  ND2D1BWP12T U842 ( .A1(n340), .A2(n2993), .ZN(n1738) );
  OAI21D1BWP12T U843 ( .A1(n1739), .A2(n1737), .B(n1738), .ZN(n1820) );
  INVD1BWP12T U844 ( .I(n1829), .ZN(n457) );
  CKND2D1BWP12T U845 ( .A1(n1383), .A2(n2262), .ZN(n1865) );
  CKBD1BWP12T U846 ( .I(n3110), .Z(n341) );
  NR2D1BWP12T U847 ( .A1(n998), .A2(n341), .ZN(n1863) );
  ND2D1BWP12T U848 ( .A1(n998), .A2(n341), .ZN(n1864) );
  OAI21D1BWP12T U849 ( .A1(n1865), .A2(n1863), .B(n1864), .ZN(n614) );
  NR2D1BWP12T U850 ( .A1(n2407), .A2(n2406), .ZN(n615) );
  NR2D1BWP12T U851 ( .A1(n342), .A2(n2404), .ZN(n783) );
  NR2D1BWP12T U852 ( .A1(n615), .A2(n783), .ZN(n344) );
  ND2D1BWP12T U853 ( .A1(n342), .A2(n2404), .ZN(n784) );
  CKND2D1BWP12T U854 ( .A1(n2407), .A2(n2406), .ZN(n616) );
  AOI21D1BWP12T U855 ( .A1(n614), .A2(n344), .B(n343), .ZN(n1848) );
  NR2D1BWP12T U856 ( .A1(n2750), .A2(n2748), .ZN(n1870) );
  CKBD1BWP12T U857 ( .I(n2764), .Z(n345) );
  CKBD1BWP12T U858 ( .I(a[7]), .Z(n346) );
  NR2D1BWP12T U859 ( .A1(n346), .A2(n2829), .ZN(n1858) );
  TPNR2D1BWP12T U860 ( .A1(n2807), .A2(n2799), .ZN(n1854) );
  NR2D1BWP12T U861 ( .A1(n1858), .A2(n1854), .ZN(n348) );
  CKND2D1BWP12T U862 ( .A1(n1850), .A2(n348), .ZN(n350) );
  ND2D1BWP12T U863 ( .A1(n2750), .A2(n2748), .ZN(n1875) );
  CKND2D1BWP12T U864 ( .A1(n345), .A2(n2766), .ZN(n1879) );
  OAI21D1BWP12T U865 ( .A1(n1878), .A2(n1875), .B(n1879), .ZN(n1852) );
  ND2D1BWP12T U866 ( .A1(n2807), .A2(n2799), .ZN(n1853) );
  CKND2D1BWP12T U867 ( .A1(n346), .A2(n2829), .ZN(n1859) );
  OAI21D1BWP12T U868 ( .A1(n1858), .A2(n1853), .B(n1859), .ZN(n347) );
  AOI21D1BWP12T U869 ( .A1(n1852), .A2(n348), .B(n347), .ZN(n349) );
  TPOAI21D1BWP12T U870 ( .A1(n1848), .A2(n350), .B(n349), .ZN(n1882) );
  INVD3BWP12T U871 ( .I(n1882), .ZN(n1906) );
  NR2D1BWP12T U872 ( .A1(n2851), .A2(n2857), .ZN(n1883) );
  NR2D1BWP12T U873 ( .A1(n2501), .A2(n2398), .ZN(n542) );
  NR2D1BWP12T U874 ( .A1(n1883), .A2(n542), .ZN(n1888) );
  NR2D1BWP12T U875 ( .A1(n2874), .A2(n2880), .ZN(n1892) );
  NR2D1BWP12T U876 ( .A1(n3074), .A2(n3067), .ZN(n1887) );
  NR2D1BWP12T U877 ( .A1(n1892), .A2(n1887), .ZN(n352) );
  ND2D1BWP12T U878 ( .A1(n1888), .A2(n352), .ZN(n1898) );
  ND2D1BWP12T U879 ( .A1(n1908), .A2(n1902), .ZN(n355) );
  CKND2D1BWP12T U880 ( .A1(n2501), .A2(n2398), .ZN(n1881) );
  CKND2D1BWP12T U881 ( .A1(n2851), .A2(n2857), .ZN(n1884) );
  OAI21D1BWP12T U882 ( .A1(n1883), .A2(n1881), .B(n1884), .ZN(n1891) );
  CKND2D1BWP12T U883 ( .A1(n3074), .A2(n3067), .ZN(n1889) );
  CKND2D1BWP12T U884 ( .A1(n2874), .A2(n2880), .ZN(n1893) );
  OAI21D1BWP12T U885 ( .A1(n1892), .A2(n1889), .B(n1893), .ZN(n351) );
  ND2D1BWP12T U886 ( .A1(n2489), .A2(n2416), .ZN(n1423) );
  CKND1BWP12T U887 ( .I(n1423), .ZN(n1901) );
  CKND2D1BWP12T U888 ( .A1(n3033), .A2(b[13]), .ZN(n1907) );
  INVD1BWP12T U889 ( .I(n1907), .ZN(n353) );
  AOI21D1BWP12T U890 ( .A1(n1908), .A2(n1901), .B(n353), .ZN(n354) );
  OA21D1BWP12T U891 ( .A1(n1900), .A2(n355), .B(n354), .Z(n356) );
  RCOAI21D2BWP12T U892 ( .A1(n1906), .A2(n357), .B(n356), .ZN(n1456) );
  OR2XD1BWP12T U893 ( .A1(n2522), .A2(a[14]), .Z(n1460) );
  ND2D1BWP12T U894 ( .A1(n2522), .A2(a[14]), .ZN(n1459) );
  INVD1BWP12T U895 ( .I(n1459), .ZN(n450) );
  TPAOI21D2BWP12T U896 ( .A1(n1456), .A2(n1460), .B(n450), .ZN(n1897) );
  NR2D1BWP12T U897 ( .A1(n2720), .A2(b[15]), .ZN(n1894) );
  ND2D1BWP12T U898 ( .A1(n2720), .A2(b[15]), .ZN(n1895) );
  OR2XD1BWP12T U899 ( .A1(b[16]), .A2(n2891), .Z(n1844) );
  ND2D1BWP12T U900 ( .A1(b[16]), .A2(n2891), .ZN(n1843) );
  INVD1BWP12T U901 ( .I(n1843), .ZN(n451) );
  TPAOI21D1BWP12T U902 ( .A1(n1846), .A2(n1844), .B(n451), .ZN(n1150) );
  NR2D1BWP12T U903 ( .A1(n2560), .A2(b[17]), .ZN(n1145) );
  ND2D1BWP12T U904 ( .A1(n2560), .A2(b[17]), .ZN(n1148) );
  OR2XD1BWP12T U905 ( .A1(b[18]), .A2(n2689), .Z(n1840) );
  ND2D1BWP12T U906 ( .A1(b[18]), .A2(n2689), .ZN(n1839) );
  INVD1BWP12T U907 ( .I(n1839), .ZN(n452) );
  TPAOI21D1BWP12T U908 ( .A1(n1842), .A2(n1840), .B(n452), .ZN(n1838) );
  NR2D1BWP12T U909 ( .A1(n2657), .A2(n2663), .ZN(n1666) );
  ND2D1BWP12T U910 ( .A1(n2657), .A2(n2663), .ZN(n1835) );
  TPOAI21D1BWP12T U911 ( .A1(n1838), .A2(n1666), .B(n1835), .ZN(n1920) );
  OR2XD1BWP12T U912 ( .A1(b[20]), .A2(a[20]), .Z(n1918) );
  ND2D1BWP12T U913 ( .A1(b[20]), .A2(a[20]), .ZN(n1917) );
  INVD1BWP12T U914 ( .I(n1917), .ZN(n453) );
  AO21D1BWP12T U915 ( .A1(n1920), .A2(n1918), .B(n453), .Z(n1834) );
  INVD2BWP12T U916 ( .I(n1867), .ZN(n3119) );
  MUX2XD0BWP12T U917 ( .I0(n2720), .I1(a[14]), .S(n1383), .Z(n2323) );
  NR2D4BWP12T U918 ( .A1(n3102), .A2(n1383), .ZN(n2064) );
  INVD6BWP12T U919 ( .I(n2064), .ZN(n2000) );
  INR2XD2BWP12T U920 ( .A1(n2297), .B1(n2000), .ZN(n2070) );
  ND2D1BWP12T U921 ( .A1(n2000), .A2(n2405), .ZN(n415) );
  INVD1BWP12T U922 ( .I(n415), .ZN(n359) );
  TPNR2D1BWP12T U923 ( .A1(n2070), .A2(n359), .ZN(n1207) );
  AN2XD2BWP12T U924 ( .A1(n3102), .A2(n1383), .Z(n2063) );
  ND2D1BWP12T U925 ( .A1(n1207), .A2(n537), .ZN(n2175) );
  NR2D1BWP12T U926 ( .A1(n415), .A2(n537), .ZN(n2185) );
  MUX2ND0BWP12T U927 ( .I0(n2560), .I1(n2891), .S(n1383), .ZN(n2319) );
  NR2D1BWP12T U928 ( .A1(n537), .A2(n359), .ZN(n2183) );
  MUX2ND0BWP12T U929 ( .I0(n3033), .I1(n2416), .S(n1383), .ZN(n2333) );
  AOI22D0BWP12T U930 ( .A1(n2185), .A2(n2319), .B1(n2183), .B2(n2333), .ZN(
        n362) );
  INVD1BWP12T U931 ( .I(n537), .ZN(n360) );
  OR2XD2BWP12T U932 ( .A1(n1207), .A2(n360), .Z(n1282) );
  INVD4BWP12T U933 ( .I(n1282), .ZN(n2187) );
  MUX2XD0BWP12T U934 ( .I0(n2657), .I1(n2689), .S(n1383), .Z(n1347) );
  INVD1BWP12T U935 ( .I(n1347), .ZN(n2318) );
  TPND2D0BWP12T U936 ( .A1(n2187), .A2(n2318), .ZN(n361) );
  OAI211D0BWP12T U937 ( .A1(n2323), .A2(n2175), .B(n362), .C(n361), .ZN(n2226)
         );
  INVD0BWP12T U938 ( .I(n2226), .ZN(n374) );
  INVD1BWP12T U939 ( .I(n2070), .ZN(n2198) );
  XNR2D2BWP12T U940 ( .A1(n2198), .A2(n2407), .ZN(n2221) );
  INVD1BWP12T U941 ( .I(n2221), .ZN(n2229) );
  ND2D1BWP12T U942 ( .A1(n2198), .A2(n2750), .ZN(n363) );
  ND2D1BWP12T U943 ( .A1(n2407), .A2(n2750), .ZN(n2343) );
  ND2D2BWP12T U944 ( .A1(n363), .A2(n2343), .ZN(n2868) );
  ND2D1BWP12T U945 ( .A1(n2229), .A2(n2868), .ZN(n2170) );
  NR2D1BWP12T U946 ( .A1(n1207), .A2(n537), .ZN(n1153) );
  TPNR2D0BWP12T U947 ( .A1(n2422), .A2(n2262), .ZN(n2298) );
  TPNR2D0BWP12T U948 ( .A1(n1383), .A2(n3110), .ZN(n364) );
  NR2D1BWP12T U949 ( .A1(n2298), .A2(n364), .ZN(n2311) );
  TPND2D0BWP12T U950 ( .A1(n1153), .A2(n2311), .ZN(n366) );
  MUX2ND0BWP12T U951 ( .I0(n2406), .I1(n2404), .S(n1383), .ZN(n1344) );
  INVD1BWP12T U952 ( .I(n1344), .ZN(n2313) );
  ND2D1BWP12T U953 ( .A1(n2187), .A2(n2313), .ZN(n365) );
  ND2D1BWP12T U954 ( .A1(n366), .A2(n365), .ZN(n2228) );
  INVD1BWP12T U955 ( .I(n2228), .ZN(n2209) );
  INVD1BWP12T U956 ( .I(n2175), .ZN(n2181) );
  CKMUX2D1BWP12T U957 ( .I0(a[7]), .I1(n2799), .S(n1383), .Z(n2143) );
  INVD1BWP12T U958 ( .I(n2143), .ZN(n2337) );
  MUX2ND0BWP12T U959 ( .I0(n2851), .I1(n2398), .S(n1383), .ZN(n2335) );
  AOI22D0BWP12T U960 ( .A1(n2181), .A2(n2337), .B1(n1153), .B2(n2335), .ZN(
        n368) );
  MUX2ND0BWP12T U961 ( .I0(n2874), .I1(n3067), .S(n1383), .ZN(n2332) );
  MUX2XD1BWP12T U962 ( .I0(n2764), .I1(n2748), .S(n1383), .Z(n2312) );
  INVD1BWP12T U963 ( .I(n2312), .ZN(n1152) );
  AOI22D0BWP12T U964 ( .A1(n2187), .A2(n2332), .B1(n2183), .B2(n1152), .ZN(
        n367) );
  CKND2D1BWP12T U965 ( .A1(n368), .A2(n367), .ZN(n2225) );
  MUX2D1BWP12T U966 ( .I0(n2209), .I1(n2225), .S(n2221), .Z(n2869) );
  INVD1BWP12T U967 ( .I(n2868), .ZN(n2217) );
  ND2XD0BWP12T U968 ( .A1(n2869), .A2(n2217), .ZN(n373) );
  MUX2NXD0BWP12T U969 ( .I0(n2518), .I1(a[26]), .S(n1383), .ZN(n2324) );
  INVD0BWP12T U970 ( .I(n2324), .ZN(n2184) );
  MUX2NXD0BWP12T U971 ( .I0(n2633), .I1(n2963), .S(n1383), .ZN(n2327) );
  CKND2D0BWP12T U972 ( .A1(n2181), .A2(n2327), .ZN(n370) );
  MUX2NXD0BWP12T U973 ( .I0(n2502), .I1(n2403), .S(n1383), .ZN(n2326) );
  MUX2NXD0BWP12T U974 ( .I0(n2993), .I1(a[20]), .S(n1383), .ZN(n2317) );
  AOI22D0BWP12T U975 ( .A1(n2185), .A2(n2326), .B1(n2183), .B2(n2317), .ZN(
        n369) );
  OAI211D0BWP12T U976 ( .A1(n2184), .A2(n1282), .B(n370), .C(n369), .ZN(n371)
         );
  INVD1BWP12T U977 ( .I(n2211), .ZN(n2908) );
  OR2XD1BWP12T U978 ( .A1(n2407), .A2(n2750), .Z(n2375) );
  NR2D1BWP12T U979 ( .A1(n2198), .A2(n2375), .ZN(n2157) );
  AOI21D0BWP12T U980 ( .A1(n371), .A2(n2908), .B(n2157), .ZN(n372) );
  OAI211D1BWP12T U981 ( .A1(n374), .A2(n2170), .B(n373), .C(n372), .ZN(n2235)
         );
  TPND2D0BWP12T U982 ( .A1(op[0]), .A2(op[1]), .ZN(n417) );
  NR2D1BWP12T U983 ( .A1(n454), .A2(n417), .ZN(n3091) );
  INVD2BWP12T U984 ( .I(n3091), .ZN(n3012) );
  INVD1BWP12T U985 ( .I(n2502), .ZN(n1293) );
  INVD1BWP12T U986 ( .I(n2403), .ZN(n2293) );
  INVD1BWP12T U987 ( .I(n2633), .ZN(n1944) );
  INVD1BWP12T U988 ( .I(n2963), .ZN(n2965) );
  INVD1BWP12T U989 ( .I(n2993), .ZN(n1952) );
  CKND2BWP12T U990 ( .I(n2398), .ZN(n2282) );
  CKND1BWP12T U991 ( .I(n2874), .ZN(n375) );
  TPND2D0BWP12T U992 ( .A1(n834), .A2(n2281), .ZN(n1463) );
  CKND2D1BWP12T U993 ( .A1(n1024), .A2(n2280), .ZN(n376) );
  NR2XD0BWP12T U994 ( .A1(n1463), .A2(n376), .ZN(n377) );
  CKND2D1BWP12T U995 ( .A1(n1960), .A2(n377), .ZN(n381) );
  ND2D1BWP12T U996 ( .A1(n378), .A2(n1937), .ZN(n380) );
  INVD1BWP12T U997 ( .I(n3110), .ZN(n379) );
  ND2D1BWP12T U998 ( .A1(n379), .A2(n2486), .ZN(n608) );
  NR2D1BWP12T U999 ( .A1(n380), .A2(n608), .ZN(n1955) );
  NR2D1BWP12T U1000 ( .A1(n381), .A2(n1464), .ZN(n1151) );
  NR2XD0BWP12T U1001 ( .A1(n2560), .A2(n2891), .ZN(n1946) );
  INVD1BWP12T U1002 ( .I(n2689), .ZN(n2687) );
  CKND2D1BWP12T U1003 ( .A1(n1946), .A2(n2687), .ZN(n1949) );
  NR2XD0BWP12T U1004 ( .A1(n1949), .A2(n2657), .ZN(n382) );
  CKND2D1BWP12T U1005 ( .A1(n1151), .A2(n382), .ZN(n1954) );
  TPNR2D0BWP12T U1006 ( .A1(op[1]), .A2(op[2]), .ZN(n421) );
  ND2D1BWP12T U1007 ( .A1(n1986), .A2(n3115), .ZN(n434) );
  CKND0BWP12T U1008 ( .I(op[3]), .ZN(n420) );
  INR2D1BWP12T U1009 ( .A1(n420), .B1(n383), .ZN(n3040) );
  IND2D1BWP12T U1010 ( .A1(n3102), .B1(n2405), .ZN(n1335) );
  ND2D1BWP12T U1011 ( .A1(n3102), .A2(n2405), .ZN(n2322) );
  OA22XD1BWP12T U1012 ( .A1(n2143), .A2(n1335), .B1(n2312), .B2(n2322), .Z(
        n385) );
  OR2D2BWP12T U1013 ( .A1(n2405), .A2(n3102), .Z(n1329) );
  INVD1BWP12T U1014 ( .I(n1329), .ZN(n595) );
  IND2D1BWP12T U1015 ( .A1(n2405), .B1(n3102), .ZN(n1333) );
  INVD1BWP12T U1016 ( .I(n1333), .ZN(n2331) );
  AOI22D0BWP12T U1017 ( .A1(n595), .A2(n2332), .B1(n2335), .B2(n2331), .ZN(
        n384) );
  ND2D1BWP12T U1018 ( .A1(n385), .A2(n384), .ZN(n2366) );
  AOI22D1BWP12T U1019 ( .A1(n2313), .A2(n595), .B1(n2331), .B2(n2311), .ZN(
        n2315) );
  MUX2NXD0BWP12T U1020 ( .I0(n2366), .I1(n2315), .S(n2407), .ZN(n2881) );
  BUFFD2BWP12T U1021 ( .I(n386), .Z(n2431) );
  AOI22D0BWP12T U1022 ( .A1(n2318), .A2(n595), .B1(n2331), .B2(n2319), .ZN(
        n388) );
  INVD1BWP12T U1023 ( .I(n2322), .ZN(n2336) );
  TPND2D0BWP12T U1024 ( .A1(n2333), .A2(n2336), .ZN(n387) );
  OAI211D1BWP12T U1025 ( .A1(n2323), .A2(n1335), .B(n388), .C(n387), .ZN(n2365) );
  INVD1BWP12T U1026 ( .I(n2407), .ZN(n2349) );
  NR2D1BWP12T U1027 ( .A1(n2349), .A2(n2750), .ZN(n2381) );
  AOI22D0BWP12T U1028 ( .A1(n595), .A2(n2324), .B1(n2326), .B2(n2331), .ZN(
        n390) );
  INVD1BWP12T U1029 ( .I(n1335), .ZN(n2334) );
  AOI22D0BWP12T U1030 ( .A1(n2336), .A2(n2317), .B1(n2327), .B2(n2334), .ZN(
        n389) );
  AOI21D0BWP12T U1031 ( .A1(n390), .A2(n389), .B(n2375), .ZN(n409) );
  NR2XD0BWP12T U1032 ( .A1(b[31]), .A2(b[30]), .ZN(n393) );
  NR2XD0BWP12T U1033 ( .A1(b[29]), .A2(b[28]), .ZN(n392) );
  ND4D1BWP12T U1034 ( .A1(n393), .A2(n392), .A3(n391), .A4(n2261), .ZN(n407)
         );
  TPNR2D0BWP12T U1035 ( .A1(b[25]), .A2(b[24]), .ZN(n397) );
  TPNR2D1BWP12T U1036 ( .A1(b[23]), .A2(b[22]), .ZN(n396) );
  NR2XD0BWP12T U1037 ( .A1(b[21]), .A2(b[20]), .ZN(n395) );
  NR2D1BWP12T U1038 ( .A1(n2663), .A2(b[18]), .ZN(n394) );
  ND4D1BWP12T U1039 ( .A1(n397), .A2(n396), .A3(n395), .A4(n394), .ZN(n406) );
  TPNR2D0BWP12T U1040 ( .A1(b[17]), .A2(b[16]), .ZN(n401) );
  NR2D1BWP12T U1041 ( .A1(b[13]), .A2(n2489), .ZN(n399) );
  NR2D1BWP12T U1042 ( .A1(n2880), .A2(n3074), .ZN(n398) );
  ND4D1BWP12T U1043 ( .A1(n401), .A2(n400), .A3(n399), .A4(n398), .ZN(n405) );
  NR2D1BWP12T U1044 ( .A1(n2857), .A2(n2501), .ZN(n403) );
  NR2D1BWP12T U1045 ( .A1(n2829), .A2(n2807), .ZN(n402) );
  ND2D1BWP12T U1046 ( .A1(n403), .A2(n402), .ZN(n404) );
  NR4D1BWP12T U1047 ( .A1(n407), .A2(n406), .A3(n405), .A4(n404), .ZN(n408) );
  CKND1BWP12T U1048 ( .I(n408), .ZN(n2437) );
  AOI211D0BWP12T U1049 ( .A1(n2365), .A2(n2381), .B(n409), .C(n2437), .ZN(n410) );
  OA21XD0BWP12T U1050 ( .A1(n2881), .A2(n2431), .B(n410), .Z(n2394) );
  INVD1BWP12T U1051 ( .I(a[31]), .ZN(n2305) );
  CKND2BWP12T U1052 ( .I(a[30]), .ZN(n2289) );
  OAI22D0BWP12T U1053 ( .A1(n2000), .A2(n2291), .B1(n1999), .B2(n2289), .ZN(
        n413) );
  IND2D2BWP12T U1054 ( .A1(n1383), .B1(n3102), .ZN(n2002) );
  INVD1BWP12T U1055 ( .I(a[29]), .ZN(n2607) );
  IND2XD1BWP12T U1056 ( .A1(n3102), .B1(n1383), .ZN(n411) );
  INVD4BWP12T U1057 ( .I(n2065), .ZN(n2001) );
  CKND1BWP12T U1058 ( .I(a[28]), .ZN(n2287) );
  OAI22D0BWP12T U1059 ( .A1(n2002), .A2(n2607), .B1(n2001), .B2(n2287), .ZN(
        n412) );
  NR2D1BWP12T U1060 ( .A1(n413), .A2(n412), .ZN(n2011) );
  MUX2XD0BWP12T U1061 ( .I0(n2305), .I1(n2011), .S(n2297), .Z(n414) );
  INR2D1BWP12T U1062 ( .A1(n415), .B1(n414), .ZN(n588) );
  INVD1BWP12T U1063 ( .I(n588), .ZN(n416) );
  NR2D1BWP12T U1064 ( .A1(n416), .A2(n2407), .ZN(n2140) );
  INVD1BWP12T U1065 ( .I(n2140), .ZN(n2458) );
  INVD3BWP12T U1066 ( .I(n408), .ZN(n2090) );
  INVD9BWP12T U1067 ( .I(n2090), .ZN(n2452) );
  ND2XD16BWP12T U1068 ( .A1(n2452), .A2(n2431), .ZN(n2448) );
  NR2D1BWP12T U1069 ( .A1(n2448), .A2(n3089), .ZN(n1306) );
  NR2D1BWP12T U1070 ( .A1(n2750), .A2(n3012), .ZN(n3060) );
  NR2D1BWP12T U1071 ( .A1(n1306), .A2(n3060), .ZN(n3004) );
  NR2XD0BWP12T U1072 ( .A1(n2458), .A2(n3004), .ZN(n432) );
  INVD1BWP12T U1073 ( .I(n2305), .ZN(n2956) );
  IND2D0BWP12T U1074 ( .A1(n2956), .B1(n2750), .ZN(n418) );
  ND2D1BWP12T U1075 ( .A1(n2452), .A2(n418), .ZN(n2040) );
  INVD1BWP12T U1076 ( .I(n2040), .ZN(n2054) );
  IND2D1BWP12T U1077 ( .A1(n2407), .B1(n2405), .ZN(n2095) );
  INVD1BWP12T U1078 ( .I(n2095), .ZN(n2108) );
  ND2D1BWP12T U1079 ( .A1(n2407), .A2(n2956), .ZN(n2197) );
  INVD1BWP12T U1080 ( .I(n2197), .ZN(n2093) );
  AOI21D0BWP12T U1081 ( .A1(n2108), .A2(n2956), .B(n2093), .ZN(n419) );
  OAI21D0BWP12T U1082 ( .A1(n2011), .A2(n2150), .B(n419), .ZN(n2048) );
  TPND2D0BWP12T U1083 ( .A1(n2054), .A2(n2048), .ZN(n2051) );
  NR2D1BWP12T U1084 ( .A1(op[0]), .A2(op[1]), .ZN(n1358) );
  INR2D1BWP12T U1085 ( .A1(n1358), .B1(n454), .ZN(n3130) );
  INVD1BWP12T U1086 ( .I(n3130), .ZN(n3044) );
  ND2D1BWP12T U1087 ( .A1(n2448), .A2(n2956), .ZN(n2039) );
  INVD1BWP12T U1088 ( .I(n2039), .ZN(n2084) );
  ND2D1BWP12T U1089 ( .A1(n2084), .A2(n3130), .ZN(n2970) );
  AN3D1BWP12T U1090 ( .A1(n421), .A2(op[0]), .A3(n420), .Z(n3107) );
  INVD1BWP12T U1091 ( .I(n3107), .ZN(n3066) );
  CKND2D0BWP12T U1092 ( .A1(op[3]), .A2(op[2]), .ZN(n422) );
  INR2D1BWP12T U1093 ( .A1(n1358), .B1(n422), .ZN(n2996) );
  OAI21D0BWP12T U1094 ( .A1(n2518), .A2(n3066), .B(n3105), .ZN(n429) );
  NR2D0BWP12T U1095 ( .A1(n423), .A2(n422), .ZN(n2304) );
  NR2D1BWP12T U1096 ( .A1(n3107), .A2(n2304), .ZN(n2995) );
  MUX2ND0BWP12T U1097 ( .I0(n2995), .I1(n2994), .S(b[27]), .ZN(n424) );
  NR2D0BWP12T U1098 ( .A1(n424), .A2(n2996), .ZN(n427) );
  CKND2D0BWP12T U1099 ( .A1(op[2]), .A2(op[1]), .ZN(n425) );
  NR2D1BWP12T U1100 ( .A1(n426), .A2(n425), .ZN(n3070) );
  INVD1BWP12T U1101 ( .I(n3070), .ZN(n3109) );
  MUX2ND0BWP12T U1102 ( .I0(n427), .I1(n3109), .S(n2291), .ZN(n428) );
  AOI21D0BWP12T U1103 ( .A1(b[27]), .A2(n429), .B(n428), .ZN(n430) );
  OAI211D0BWP12T U1104 ( .A1(n2051), .A2(n3044), .B(n2970), .C(n430), .ZN(n431) );
  RCAOI211D0BWP12T U1105 ( .A1(n3040), .A2(n2394), .B(n432), .C(n431), .ZN(
        n433) );
  OAI211D1BWP12T U1106 ( .A1(n2235), .A2(n3012), .B(n434), .C(n433), .ZN(n435)
         );
  AOI21D1BWP12T U1107 ( .A1(n1930), .A2(n3119), .B(n435), .ZN(n456) );
  CKBD1BWP12T U1108 ( .I(n3102), .Z(n436) );
  NR2D1BWP12T U1109 ( .A1(n436), .A2(n3110), .ZN(n1707) );
  NR2D1BWP12T U1110 ( .A1(n779), .A2(n1707), .ZN(n438) );
  CKBD1BWP12T U1111 ( .I(n1383), .Z(n1387) );
  NR2D1BWP12T U1112 ( .A1(n2262), .A2(c_in), .ZN(n1384) );
  CKND2D1BWP12T U1113 ( .A1(n2262), .A2(c_in), .ZN(n1385) );
  OAI21D1BWP12T U1114 ( .A1(n1391), .A2(n1384), .B(n1385), .ZN(n778) );
  ND2D1BWP12T U1115 ( .A1(n436), .A2(n3110), .ZN(n1708) );
  CKND2D1BWP12T U1116 ( .A1(n2405), .A2(n2404), .ZN(n780) );
  OAI21D1BWP12T U1117 ( .A1(n779), .A2(n1708), .B(n780), .ZN(n437) );
  NR2D1BWP12T U1118 ( .A1(n2750), .A2(n2748), .ZN(n1703) );
  NR2D1BWP12T U1119 ( .A1(n1717), .A2(n1854), .ZN(n440) );
  ND2D1BWP12T U1120 ( .A1(n1714), .A2(n440), .ZN(n442) );
  ND2D1BWP12T U1121 ( .A1(n2407), .A2(n2406), .ZN(n1701) );
  CKND2D1BWP12T U1122 ( .A1(n2750), .A2(n2748), .ZN(n1704) );
  OAI21D1BWP12T U1123 ( .A1(n1703), .A2(n1701), .B(n1704), .ZN(n1715) );
  ND2D1BWP12T U1124 ( .A1(n2764), .A2(n2766), .ZN(n1716) );
  OAI21D1BWP12T U1125 ( .A1(n1854), .A2(n1716), .B(n1853), .ZN(n439) );
  AOI21D1BWP12T U1126 ( .A1(n1715), .A2(n440), .B(n439), .ZN(n441) );
  CKBD1BWP12T U1127 ( .I(a[7]), .Z(n443) );
  NR2D1BWP12T U1128 ( .A1(n443), .A2(n2829), .ZN(n543) );
  NR2D1BWP12T U1129 ( .A1(n2501), .A2(n2398), .ZN(n546) );
  NR2D1BWP12T U1130 ( .A1(n543), .A2(n546), .ZN(n1672) );
  NR2D1BWP12T U1131 ( .A1(n2851), .A2(n2857), .ZN(n1671) );
  NR2D1BWP12T U1132 ( .A1(n3074), .A2(n3067), .ZN(n1676) );
  NR2D1BWP12T U1133 ( .A1(n1671), .A2(n1676), .ZN(n445) );
  ND2D1BWP12T U1134 ( .A1(n1672), .A2(n445), .ZN(n1679) );
  NR2D1BWP12T U1135 ( .A1(n2874), .A2(n2880), .ZN(n1406) );
  NR2D1BWP12T U1136 ( .A1(n2489), .A2(n2416), .ZN(n1410) );
  NR2D1BWP12T U1137 ( .A1(n1406), .A2(n1410), .ZN(n1685) );
  CKND2D1BWP12T U1138 ( .A1(n1685), .A2(n1690), .ZN(n447) );
  OR2XD1BWP12T U1139 ( .A1(n1679), .A2(n447), .Z(n449) );
  ND2D1BWP12T U1140 ( .A1(n443), .A2(n2829), .ZN(n1698) );
  CKND2D1BWP12T U1141 ( .A1(n2501), .A2(n2398), .ZN(n547) );
  OAI21D1BWP12T U1142 ( .A1(n546), .A2(n1698), .B(n547), .ZN(n1675) );
  CKND2D1BWP12T U1143 ( .A1(n2851), .A2(n2857), .ZN(n1673) );
  CKND2D1BWP12T U1144 ( .A1(n3074), .A2(n3067), .ZN(n1677) );
  OAI21D1BWP12T U1145 ( .A1(n1676), .A2(n1673), .B(n1677), .ZN(n444) );
  AOI21D1BWP12T U1146 ( .A1(n445), .A2(n1675), .B(n444), .ZN(n1678) );
  ND2D1BWP12T U1147 ( .A1(n2874), .A2(n2880), .ZN(n1680) );
  OAI21D1BWP12T U1148 ( .A1(n1410), .A2(n1680), .B(n1423), .ZN(n1684) );
  CKND2D1BWP12T U1149 ( .A1(n3033), .A2(b[13]), .ZN(n1689) );
  AOI21D1BWP12T U1150 ( .A1(n1684), .A2(n1690), .B(n353), .ZN(n446) );
  OA21D1BWP12T U1151 ( .A1(n1678), .A2(n447), .B(n446), .Z(n448) );
  RCOAI21D1BWP12T U1152 ( .A1(n1700), .A2(n449), .B(n448), .ZN(n1462) );
  NR2XD0BWP12T U1153 ( .A1(n2720), .A2(b[15]), .ZN(n1693) );
  CKND2D1BWP12T U1154 ( .A1(n2720), .A2(b[15]), .ZN(n1694) );
  TPAOI21D1BWP12T U1155 ( .A1(n1724), .A2(n1844), .B(n451), .ZN(n1147) );
  TPOAI21D1BWP12T U1156 ( .A1(n1147), .A2(n1145), .B(n1148), .ZN(n1670) );
  TPAOI21D1BWP12T U1157 ( .A1(n1670), .A2(n1840), .B(n452), .ZN(n1668) );
  AO21D1BWP12T U1158 ( .A1(n1665), .A2(n1918), .B(n453), .Z(n1726) );
  CKND2D1BWP12T U1159 ( .A1(n1728), .A2(n3098), .ZN(n455) );
  OAI211D1BWP12T U1160 ( .A1(n3020), .A2(n457), .B(n456), .C(n455), .ZN(n458)
         );
  AOI21D1BWP12T U1161 ( .A1(n3095), .A2(n1549), .B(n458), .ZN(n459) );
  IOA21D1BWP12T U1162 ( .A1(n1658), .A2(n3126), .B(n459), .ZN(result[27]) );
  INVD2BWP12T U1163 ( .I(a[7]), .ZN(n896) );
  INVD8BWP12T U1164 ( .I(n896), .ZN(n2555) );
  XNR2XD8BWP12T U1165 ( .A1(n2398), .A2(n2555), .ZN(n2533) );
  INVD2BWP12T U1166 ( .I(n2851), .ZN(n844) );
  INVD6BWP12T U1167 ( .I(n844), .ZN(n2532) );
  XOR2XD1BWP12T U1168 ( .A1(n2398), .A2(n2532), .Z(n460) );
  TPND2D3BWP12T U1169 ( .A1(n2533), .A2(n460), .ZN(n2535) );
  XNR2D0BWP12T U1170 ( .A1(n2532), .A2(b[21]), .ZN(n944) );
  XNR2D0BWP12T U1171 ( .A1(n2532), .A2(b[22]), .ZN(n1104) );
  OAI22D0BWP12T U1172 ( .A1(n2535), .A2(n944), .B1(n2533), .B2(n1104), .ZN(
        mult_x_18_n893) );
  XNR2XD4BWP12T U1173 ( .A1(a[20]), .A2(n2657), .ZN(n2491) );
  XOR2XD1BWP12T U1174 ( .A1(a[20]), .A2(n2993), .Z(n461) );
  TPND2D2BWP12T U1175 ( .A1(n2491), .A2(n461), .ZN(n2493) );
  XNR2XD1BWP12T U1176 ( .A1(n2993), .A2(n3074), .ZN(n827) );
  XNR2XD0BWP12T U1177 ( .A1(n2993), .A2(n2880), .ZN(n2492) );
  OAI22D0BWP12T U1178 ( .A1(n2493), .A2(n827), .B1(n2491), .B2(n2492), .ZN(
        mult_x_18_n784) );
  XNR2XD1BWP12T U1179 ( .A1(n3110), .A2(b[28]), .ZN(n861) );
  XNR2XD1BWP12T U1180 ( .A1(n3110), .A2(b[29]), .ZN(n1088) );
  OAI22D1BWP12T U1181 ( .A1(n2487), .A2(n861), .B1(n1088), .B2(n2486), .ZN(
        n465) );
  INVD1BWP12T U1182 ( .I(n2607), .ZN(n2608) );
  XOR2D0BWP12T U1183 ( .A1(n2608), .A2(a[28]), .Z(n462) );
  XNR2XD1BWP12T U1184 ( .A1(a[28]), .A2(n2518), .ZN(n2543) );
  ND2D1BWP12T U1185 ( .A1(n462), .A2(n2543), .ZN(n2546) );
  IND2D1BWP12T U1186 ( .A1(n1382), .B1(n2608), .ZN(n463) );
  OAI22D1BWP12T U1187 ( .A1(n2546), .A2(n2607), .B1(n2543), .B2(n463), .ZN(
        n464) );
  HA1D0BWP12T U1188 ( .A(n465), .B(n464), .CO(mult_x_18_n444), .S(
        mult_x_18_n445) );
  XNR2D2BWP12T U1189 ( .A1(n2764), .A2(n2799), .ZN(n2557) );
  XOR2D2BWP12T U1190 ( .A1(n2555), .A2(n2799), .Z(n466) );
  CKND2D8BWP12T U1191 ( .A1(n2557), .A2(n466), .ZN(n2559) );
  XNR2XD1BWP12T U1192 ( .A1(n2555), .A2(b[23]), .ZN(n1004) );
  XNR2XD0BWP12T U1193 ( .A1(n2555), .A2(b[24]), .ZN(n642) );
  TPOAI22D0BWP12T U1194 ( .A1(n2559), .A2(n1004), .B1(n2557), .B2(n642), .ZN(
        mult_x_18_n918) );
  CKND2D1BWP12T U1195 ( .A1(n467), .A2(n645), .ZN(n468) );
  XNR2D1BWP12T U1196 ( .A1(n1650), .A2(n468), .ZN(n1660) );
  INVD1BWP12T U1197 ( .I(n1660), .ZN(n518) );
  INVD2BWP12T U1198 ( .I(n3126), .ZN(n2951) );
  FA1D1BWP12T U1199 ( .A(n471), .B(a[26]), .CI(n469), .CO(n695), .S(n1551) );
  FA1D0BWP12T U1200 ( .A(n471), .B(a[26]), .CI(n470), .CO(n650), .S(n1828) );
  INVD1BWP12T U1201 ( .I(n1828), .ZN(n515) );
  FA1D2BWP12T U1202 ( .A(b[26]), .B(a[26]), .CI(n472), .CO(n653), .S(n1924) );
  OAI22D1BWP12T U1203 ( .A1(n2000), .A2(n2289), .B1(n2001), .B2(n2305), .ZN(
        n2201) );
  MUX2D1BWP12T U1204 ( .I0(a[26]), .I1(n2518), .S(n1383), .Z(n522) );
  NR2D1BWP12T U1205 ( .A1(n2002), .A2(a[28]), .ZN(n474) );
  NR2D1BWP12T U1206 ( .A1(n1999), .A2(n2608), .ZN(n473) );
  NR2D1BWP12T U1207 ( .A1(n474), .A2(n473), .ZN(n475) );
  OAI21D1BWP12T U1208 ( .A1(n3102), .A2(n522), .B(n475), .ZN(n2029) );
  INVD1BWP12T U1209 ( .I(n2029), .ZN(n747) );
  MUX2D1BWP12T U1210 ( .I0(n2201), .I1(n747), .S(n2297), .Z(n2212) );
  INVD1BWP12T U1211 ( .I(n2212), .ZN(n807) );
  INR2D1BWP12T U1212 ( .A1(n2262), .B1(n2002), .ZN(n1226) );
  CKND1BWP12T U1213 ( .I(n1226), .ZN(n1209) );
  TPNR2D0BWP12T U1214 ( .A1(n1207), .A2(n1209), .ZN(n477) );
  MUX2ND0BWP12T U1215 ( .I0(n2404), .I1(n3110), .S(n1383), .ZN(n1211) );
  INVD1BWP12T U1216 ( .I(n1211), .ZN(n674) );
  NR2D1BWP12T U1217 ( .A1(n674), .A2(n1226), .ZN(n1231) );
  INVD1BWP12T U1218 ( .I(n1231), .ZN(n476) );
  OAI21D1BWP12T U1219 ( .A1(n2187), .A2(n477), .B(n476), .ZN(n804) );
  MUX2ND0BWP12T U1220 ( .I0(n2799), .I1(n2764), .S(n1383), .ZN(n682) );
  MUX2ND0BWP12T U1221 ( .I0(n2748), .I1(n2406), .S(n1383), .ZN(n1208) );
  AOI22D0BWP12T U1222 ( .A1(n2181), .A2(n682), .B1(n2183), .B2(n1208), .ZN(
        n479) );
  MUX2ND0BWP12T U1223 ( .I0(n3067), .I1(n2851), .S(n1383), .ZN(n1244) );
  MUX2ND0BWP12T U1224 ( .I0(n2398), .I1(a[7]), .S(n1383), .ZN(n1247) );
  AOI22D0BWP12T U1225 ( .A1(n2187), .A2(n1244), .B1(n1153), .B2(n1247), .ZN(
        n478) );
  ND2D1BWP12T U1226 ( .A1(n479), .A2(n478), .ZN(n2155) );
  MUX2D1BWP12T U1227 ( .I0(n804), .I1(n2155), .S(n2221), .Z(n3065) );
  CKND0BWP12T U1228 ( .I(n3065), .ZN(n488) );
  MUX2ND0BWP12T U1229 ( .I0(a[14]), .I1(n3033), .S(n1383), .ZN(n1245) );
  CKND2D0BWP12T U1230 ( .A1(n2181), .A2(n1245), .ZN(n482) );
  MUX2NXD0BWP12T U1231 ( .I0(n2891), .I1(n2720), .S(n1383), .ZN(n1240) );
  MUX2NXD0BWP12T U1232 ( .I0(n2416), .I1(n2874), .S(n1383), .ZN(n1246) );
  AOI22D0BWP12T U1233 ( .A1(n2185), .A2(n1240), .B1(n2183), .B2(n1246), .ZN(
        n481) );
  MUX2NXD0BWP12T U1234 ( .I0(n2689), .I1(n2560), .S(n1383), .ZN(n1238) );
  CKND2D0BWP12T U1235 ( .A1(n2187), .A2(n1238), .ZN(n480) );
  ND3D1BWP12T U1236 ( .A1(n482), .A2(n481), .A3(n480), .ZN(n2156) );
  INVD1BWP12T U1237 ( .I(n2170), .ZN(n2904) );
  MUX2NXD0BWP12T U1238 ( .I0(n2963), .I1(n2993), .S(n1383), .ZN(n1241) );
  CKND2D0BWP12T U1239 ( .A1(n2181), .A2(n1241), .ZN(n485) );
  MUX2NXD0BWP12T U1240 ( .I0(n2403), .I1(n2633), .S(n1383), .ZN(n1233) );
  MUX2NXD0BWP12T U1241 ( .I0(a[20]), .I1(n2657), .S(n1383), .ZN(n1239) );
  AOI22D0BWP12T U1242 ( .A1(n2185), .A2(n1233), .B1(n2183), .B2(n1239), .ZN(
        n484) );
  MUX2NXD0BWP12T U1243 ( .I0(a[26]), .I1(n2502), .S(n1383), .ZN(n1232) );
  CKND2D0BWP12T U1244 ( .A1(n2187), .A2(n1232), .ZN(n483) );
  AOI31D0BWP12T U1245 ( .A1(n485), .A2(n484), .A3(n483), .B(n2211), .ZN(n486)
         );
  AOI211D0BWP12T U1246 ( .A1(n2156), .A2(n2904), .B(n2157), .C(n486), .ZN(n487) );
  TPOAI21D0BWP12T U1247 ( .A1(n488), .A2(n2868), .B(n487), .ZN(n2236) );
  OA21D1BWP12T U1248 ( .A1(n807), .A2(n2375), .B(n2236), .Z(n510) );
  HA1D1BWP12T U1249 ( .A(n2290), .B(n489), .CO(n689), .S(n1985) );
  ND2D1BWP12T U1250 ( .A1(n1985), .A2(n3115), .ZN(n509) );
  AOI22D0BWP12T U1251 ( .A1(n2336), .A2(n1208), .B1(n682), .B2(n2334), .ZN(
        n491) );
  AOI22D0BWP12T U1252 ( .A1(n595), .A2(n1244), .B1(n1247), .B2(n2331), .ZN(
        n490) );
  ND2D1BWP12T U1253 ( .A1(n491), .A2(n490), .ZN(n2380) );
  AOI21D0BWP12T U1254 ( .A1(n1226), .A2(n2297), .B(n595), .ZN(n492) );
  NR2D1BWP12T U1255 ( .A1(n1231), .A2(n492), .ZN(n2350) );
  INVD1BWP12T U1256 ( .I(n2350), .ZN(n792) );
  MUX2NXD0BWP12T U1257 ( .I0(n2380), .I1(n792), .S(n2407), .ZN(n3077) );
  NR2D0BWP12T U1258 ( .A1(n3077), .A2(n2431), .ZN(n497) );
  OAI22D0BWP12T U1259 ( .A1(n1329), .A2(n1238), .B1(n1240), .B2(n1333), .ZN(
        n2377) );
  OAI22D0BWP12T U1260 ( .A1(n2322), .A2(n1246), .B1(n1245), .B2(n1335), .ZN(
        n2376) );
  INVD1BWP12T U1261 ( .I(n2381), .ZN(n2082) );
  TPNR3D0BWP12T U1262 ( .A1(n2377), .A2(n2376), .A3(n2082), .ZN(n496) );
  AOI22D0BWP12T U1263 ( .A1(n2336), .A2(n1239), .B1(n1241), .B2(n2334), .ZN(
        n494) );
  AOI22D0BWP12T U1264 ( .A1(n595), .A2(n1232), .B1(n1233), .B2(n2331), .ZN(
        n493) );
  AOI21D0BWP12T U1265 ( .A1(n494), .A2(n493), .B(n2375), .ZN(n495) );
  NR4D0BWP12T U1266 ( .A1(n497), .A2(n496), .A3(n495), .A4(n2090), .ZN(n2395)
         );
  ND2XD0BWP12T U1267 ( .A1(n2000), .A2(n2956), .ZN(n498) );
  INR2XD0BWP12T U1268 ( .A1(n498), .B1(n2201), .ZN(n1225) );
  CKND0BWP12T U1269 ( .I(n1225), .ZN(n499) );
  MUX2ND0BWP12T U1270 ( .I0(n499), .I1(n747), .S(n2297), .ZN(n500) );
  OA21XD1BWP12T U1271 ( .A1(n500), .A2(n2407), .B(n2197), .Z(n2033) );
  INVD1BWP12T U1272 ( .I(n2114), .ZN(n2101) );
  NR2D1BWP12T U1273 ( .A1(n2054), .A2(n2101), .ZN(n2009) );
  INVD1BWP12T U1274 ( .I(n2009), .ZN(n2022) );
  CKND2D0BWP12T U1275 ( .A1(n2022), .A2(n3130), .ZN(n1309) );
  AOI21D0BWP12T U1276 ( .A1(n2033), .A2(n2039), .B(n1309), .ZN(n507) );
  CKND0BWP12T U1277 ( .I(n1306), .ZN(n2697) );
  INR2D1BWP12T U1278 ( .A1(n2349), .B1(n807), .ZN(n3061) );
  INVD1BWP12T U1279 ( .I(n3061), .ZN(n2457) );
  INVD1BWP12T U1280 ( .I(n2995), .ZN(n3104) );
  INVD1BWP12T U1281 ( .I(n2994), .ZN(n3103) );
  MUX2ND0BWP12T U1282 ( .I0(n3104), .I1(n3103), .S(b[26]), .ZN(n501) );
  CKND2D0BWP12T U1283 ( .A1(n501), .A2(n3105), .ZN(n502) );
  CKND1BWP12T U1284 ( .I(a[26]), .ZN(n2290) );
  MUX2NXD0BWP12T U1285 ( .I0(n502), .I1(n3070), .S(n2290), .ZN(n505) );
  OAI21D0BWP12T U1286 ( .A1(a[26]), .A2(n3066), .B(n3105), .ZN(n503) );
  CKND2D0BWP12T U1287 ( .A1(n503), .A2(b[26]), .ZN(n504) );
  OAI211D1BWP12T U1288 ( .A1(n2697), .A2(n2457), .B(n505), .C(n504), .ZN(n506)
         );
  AOI211XD0BWP12T U1289 ( .A1(n3040), .A2(n2395), .B(n507), .C(n506), .ZN(n508) );
  OAI211D1BWP12T U1290 ( .A1(n510), .A2(n3012), .B(n509), .C(n508), .ZN(n511)
         );
  AOI21D1BWP12T U1291 ( .A1(n1924), .A2(n3119), .B(n511), .ZN(n514) );
  FA1D0BWP12T U1292 ( .A(b[26]), .B(a[26]), .CI(n512), .CO(n652), .S(n1730) );
  CKND2D1BWP12T U1293 ( .A1(n1730), .A2(n3098), .ZN(n513) );
  OAI211D1BWP12T U1294 ( .A1(n3020), .A2(n515), .B(n514), .C(n513), .ZN(n516)
         );
  AOI21D1BWP12T U1295 ( .A1(n3095), .A2(n1551), .B(n516), .ZN(n517) );
  OAI21D1BWP12T U1296 ( .A1(n518), .A2(n2951), .B(n517), .ZN(result[26]) );
  INVD1BWP12T U1297 ( .I(n519), .ZN(n1598) );
  INVD1BWP12T U1298 ( .I(n1620), .ZN(n578) );
  INVD1BWP12T U1299 ( .I(n1464), .ZN(n1970) );
  XNR2XD1BWP12T U1300 ( .A1(n1970), .A2(n2398), .ZN(n1958) );
  OAI22D1BWP12T U1301 ( .A1(n2000), .A2(n2293), .B1(n2001), .B2(n2292), .ZN(
        n521) );
  AOI21D1BWP12T U1302 ( .A1(n3102), .A2(n522), .B(n521), .ZN(n1414) );
  OAI22D0BWP12T U1303 ( .A1(n2000), .A2(n2287), .B1(n2305), .B2(n1999), .ZN(
        n524) );
  OAI22D1BWP12T U1304 ( .A1(n2002), .A2(n2289), .B1(n2001), .B2(n2607), .ZN(
        n523) );
  NR2D1BWP12T U1305 ( .A1(n524), .A2(n523), .ZN(n2205) );
  OAI22D1BWP12T U1306 ( .A1(n1414), .A2(n2150), .B1(n2205), .B2(n2095), .ZN(
        n2207) );
  OAI22D1BWP12T U1307 ( .A1(n2000), .A2(n2398), .B1(n2874), .B2(n1999), .ZN(
        n526) );
  OAI22D0BWP12T U1308 ( .A1(n3067), .A2(n2002), .B1(n2001), .B2(n2851), .ZN(
        n525) );
  NR2D1BWP12T U1309 ( .A1(n526), .A2(n525), .ZN(n2016) );
  INVD0BWP12T U1310 ( .I(n2016), .ZN(n529) );
  OAI22D1BWP12T U1311 ( .A1(n2000), .A2(n2928), .B1(n2002), .B2(n2965), .ZN(
        n528) );
  OAI22D0BWP12T U1312 ( .A1(n2001), .A2(n2998), .B1(n1999), .B2(n2636), .ZN(
        n527) );
  NR2D1BWP12T U1313 ( .A1(n528), .A2(n527), .ZN(n1413) );
  ND2D1BWP12T U1314 ( .A1(n2407), .A2(n2405), .ZN(n2110) );
  OAI22D0BWP12T U1315 ( .A1(n529), .A2(n2150), .B1(n1413), .B2(n2110), .ZN(
        n536) );
  OAI22D0BWP12T U1316 ( .A1(n2000), .A2(n2281), .B1(n1999), .B2(n2722), .ZN(
        n531) );
  OAI22D1BWP12T U1317 ( .A1(n2002), .A2(n2280), .B1(n2001), .B2(n3031), .ZN(
        n530) );
  NR2D1BWP12T U1318 ( .A1(n531), .A2(n530), .ZN(n2015) );
  OAI21D0BWP12T U1319 ( .A1(n2015), .A2(n2095), .B(n2431), .ZN(n535) );
  CKND1BWP12T U1320 ( .I(n2891), .ZN(n2893) );
  OAI22D0BWP12T U1321 ( .A1(n2000), .A2(n2893), .B1(n2001), .B2(n2275), .ZN(
        n533) );
  OAI22D0BWP12T U1322 ( .A1(n2002), .A2(n2687), .B1(n1999), .B2(n2659), .ZN(
        n532) );
  NR2D1BWP12T U1323 ( .A1(n533), .A2(n532), .ZN(n2019) );
  NR2D1BWP12T U1324 ( .A1(n2349), .A2(n2405), .ZN(n2200) );
  INVD1BWP12T U1325 ( .I(n2200), .ZN(n2133) );
  TPNR2D0BWP12T U1326 ( .A1(n2019), .A2(n2133), .ZN(n534) );
  NR3D1BWP12T U1327 ( .A1(n536), .A2(n535), .A3(n534), .ZN(n554) );
  INVD1BWP12T U1328 ( .I(n554), .ZN(n556) );
  INR2D1BWP12T U1329 ( .A1(n2262), .B1(n2000), .ZN(n1379) );
  INR2D1BWP12T U1330 ( .A1(n1379), .B1(n2405), .ZN(n2907) );
  INVD1BWP12T U1331 ( .I(n1208), .ZN(n1228) );
  INVD1BWP12T U1332 ( .I(n682), .ZN(n1227) );
  AOI22D1BWP12T U1333 ( .A1(n2181), .A2(n1228), .B1(n1227), .B2(n1153), .ZN(
        n541) );
  INVD0BWP12T U1334 ( .I(n1247), .ZN(n539) );
  NR2D0BWP12T U1335 ( .A1(n537), .A2(n1211), .ZN(n538) );
  AOI22D0BWP12T U1336 ( .A1(n2187), .A2(n539), .B1(n1207), .B2(n538), .ZN(n540) );
  ND2D1BWP12T U1337 ( .A1(n541), .A2(n540), .ZN(n2905) );
  INVD1BWP12T U1338 ( .I(n1698), .ZN(n544) );
  AOI21D1BWP12T U1339 ( .A1(n545), .A2(n1860), .B(n544), .ZN(n550) );
  INVD0BWP12T U1340 ( .I(n546), .ZN(n548) );
  CKND2D1BWP12T U1341 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2XD1BWP12T U1342 ( .A1(n550), .A2(n549), .Z(n1719) );
  AOI22D0BWP12T U1343 ( .A1(n3119), .A2(n1885), .B1(n1719), .B2(n3098), .ZN(
        n551) );
  OAI21D1BWP12T U1344 ( .A1(n2223), .A2(n3012), .B(n551), .ZN(n552) );
  AOI21D1BWP12T U1345 ( .A1(n3115), .A2(n1958), .B(n552), .ZN(n577) );
  INVD1BWP12T U1346 ( .I(n553), .ZN(n1769) );
  ND2D1BWP12T U1347 ( .A1(n2207), .A2(n2452), .ZN(n555) );
  AOI21D1BWP12T U1348 ( .A1(n2448), .A2(n555), .B(n554), .ZN(n564) );
  AOI211XD0BWP12T U1349 ( .A1(n2093), .A2(n556), .B(n564), .C(n2101), .ZN(
        n2061) );
  INVD1BWP12T U1350 ( .I(n1509), .ZN(n558) );
  TPAOI21D0BWP12T U1351 ( .A1(n559), .A2(n1785), .B(n558), .ZN(n563) );
  CKND2D1BWP12T U1352 ( .A1(n1769), .A2(n561), .ZN(n562) );
  XOR2XD1BWP12T U1353 ( .A1(n563), .A2(n562), .Z(n1518) );
  MOAI22D0BWP12T U1354 ( .A1(n2061), .A2(n3044), .B1(n1518), .B2(n3095), .ZN(
        n575) );
  INVD1BWP12T U1355 ( .I(n564), .ZN(n2442) );
  AOI22D0BWP12T U1356 ( .A1(n2336), .A2(n1211), .B1(n1208), .B2(n2334), .ZN(
        n566) );
  AOI22D0BWP12T U1357 ( .A1(n595), .A2(n1247), .B1(n682), .B2(n2331), .ZN(n565) );
  ND2D1BWP12T U1358 ( .A1(n566), .A2(n565), .ZN(n2351) );
  INVD1BWP12T U1359 ( .I(n2351), .ZN(n725) );
  MUX2NXD0BWP12T U1360 ( .I0(n725), .I1(n2907), .S(n2407), .ZN(n567) );
  NR2D1BWP12T U1361 ( .A1(n567), .A2(n2448), .ZN(n2386) );
  TPND2D0BWP12T U1362 ( .A1(n2386), .A2(n3040), .ZN(n573) );
  OAI21D0BWP12T U1363 ( .A1(n2398), .A2(n3066), .B(n3105), .ZN(n571) );
  MUX2ND0BWP12T U1364 ( .I0(n2995), .I1(n2994), .S(n2501), .ZN(n568) );
  NR2D0BWP12T U1365 ( .A1(n568), .A2(n2996), .ZN(n569) );
  MUX2ND0BWP12T U1366 ( .I0(n569), .I1(n3109), .S(n2282), .ZN(n570) );
  RCAOI21D0BWP12T U1367 ( .A1(n2501), .A2(n571), .B(n570), .ZN(n572) );
  OAI211D1BWP12T U1368 ( .A1(n3089), .A2(n2442), .B(n573), .C(n572), .ZN(n574)
         );
  AOI211XD0BWP12T U1369 ( .A1(n314), .A2(n1801), .B(n575), .C(n574), .ZN(n576)
         );
  OAI211D1BWP12T U1370 ( .A1(n2951), .A2(n578), .B(n577), .C(n576), .ZN(
        result[8]) );
  INVD1BWP12T U1371 ( .I(n3089), .ZN(n3052) );
  ND2D1BWP12T U1372 ( .A1(n2452), .A2(n3052), .ZN(n3038) );
  CKND2D1BWP12T U1373 ( .A1(n3038), .A2(n3012), .ZN(n2717) );
  INVD1BWP12T U1374 ( .I(n2717), .ZN(n2870) );
  TPOAI22D0BWP12T U1375 ( .A1(n2000), .A2(n2659), .B1(n1999), .B2(n2965), .ZN(
        n583) );
  OAI22D1BWP12T U1376 ( .A1(n2998), .A2(n2002), .B1(n2001), .B2(n2928), .ZN(
        n582) );
  NR2D1BWP12T U1377 ( .A1(n583), .A2(n582), .ZN(n2056) );
  OAI22D1BWP12T U1378 ( .A1(n2000), .A2(n2636), .B1(n1999), .B2(n2290), .ZN(
        n585) );
  OAI22D1BWP12T U1379 ( .A1(n2002), .A2(n2292), .B1(n2001), .B2(n2293), .ZN(
        n584) );
  NR2D1BWP12T U1380 ( .A1(n585), .A2(n584), .ZN(n2044) );
  MUX2NXD0BWP12T U1381 ( .I0(n2056), .I1(n2044), .S(n2405), .ZN(n586) );
  NR2D1BWP12T U1382 ( .A1(n586), .A2(n2407), .ZN(n627) );
  INVD1BWP12T U1383 ( .I(n627), .ZN(n587) );
  OAI21D1BWP12T U1384 ( .A1(n588), .A2(n2349), .B(n587), .ZN(n2668) );
  OAI22D1BWP12T U1385 ( .A1(n2000), .A2(n2876), .B1(n1999), .B2(n2280), .ZN(
        n590) );
  OAI22D0BWP12T U1386 ( .A1(n2002), .A2(n3031), .B1(n2001), .B2(n2281), .ZN(
        n589) );
  NR2D1BWP12T U1387 ( .A1(n590), .A2(n589), .ZN(n2058) );
  OAI22D0BWP12T U1388 ( .A1(n2000), .A2(n2722), .B1(n1999), .B2(n2687), .ZN(
        n592) );
  OAI22D0BWP12T U1389 ( .A1(n2002), .A2(n2275), .B1(n2001), .B2(n2893), .ZN(
        n591) );
  NR2D1BWP12T U1390 ( .A1(n592), .A2(n591), .ZN(n2057) );
  OAI22D0BWP12T U1391 ( .A1(n2058), .A2(n2133), .B1(n2057), .B2(n2110), .ZN(
        n601) );
  CKND1BWP12T U1392 ( .I(a[7]), .ZN(n2831) );
  OAI22D0BWP12T U1393 ( .A1(n2000), .A2(n2831), .B1(n1999), .B2(n3069), .ZN(
        n594) );
  OAI22D0BWP12T U1394 ( .A1(n2002), .A2(n2853), .B1(n2001), .B2(n2282), .ZN(
        n593) );
  NR2D1BWP12T U1395 ( .A1(n594), .A2(n593), .ZN(n2059) );
  OAI21D0BWP12T U1396 ( .A1(n2059), .A2(n2095), .B(n2431), .ZN(n600) );
  NR2D1BWP12T U1397 ( .A1(n1333), .A2(n1383), .ZN(n2072) );
  INR2D1BWP12T U1398 ( .A1(n1383), .B1(n1333), .ZN(n2073) );
  AOI22D0BWP12T U1399 ( .A1(n2764), .A2(n2072), .B1(n2073), .B2(n2799), .ZN(
        n598) );
  CKND2D1BWP12T U1400 ( .A1(n595), .A2(n1383), .ZN(n1334) );
  INVD1BWP12T U1401 ( .I(n1334), .ZN(n2071) );
  CKND2D0BWP12T U1402 ( .A1(n2071), .A2(n2748), .ZN(n597) );
  CKND2D0BWP12T U1403 ( .A1(n2070), .A2(n2406), .ZN(n596) );
  TPAOI31D0BWP12T U1404 ( .A1(n598), .A2(n597), .A3(n596), .B(n2407), .ZN(n599) );
  NR3D1BWP12T U1405 ( .A1(n601), .A2(n600), .A3(n599), .ZN(n629) );
  AO21D1BWP12T U1406 ( .A1(n2668), .A2(n2750), .B(n629), .Z(n2141) );
  INVD1BWP12T U1407 ( .I(n602), .ZN(n799) );
  CKND0BWP12T U1408 ( .I(n603), .ZN(n605) );
  CKND1BWP12T U1409 ( .I(n3095), .ZN(n3059) );
  INVD1BWP12T U1410 ( .I(n606), .ZN(n1529) );
  CKND2D0BWP12T U1411 ( .A1(n605), .A2(n1527), .ZN(n607) );
  XNR2D1BWP12T U1412 ( .A1(n1529), .A2(n607), .ZN(n1519) );
  INVD1BWP12T U1413 ( .I(n1519), .ZN(n613) );
  CKND0BWP12T U1414 ( .I(n608), .ZN(n800) );
  INVD1BWP12T U1415 ( .I(n3040), .ZN(n2903) );
  NR2XD2BWP12T U1416 ( .A1(n2448), .A2(n2903), .ZN(n3078) );
  INVD1P75BWP12T U1417 ( .I(n3078), .ZN(n2860) );
  TPNR2D1BWP12T U1418 ( .A1(n2860), .A2(n2407), .ZN(n3094) );
  INVD1BWP12T U1419 ( .I(n2315), .ZN(n2364) );
  AOI22D1BWP12T U1420 ( .A1(n3115), .A2(n1957), .B1(n3094), .B2(n2364), .ZN(
        n612) );
  INVD1BWP12T U1421 ( .I(n609), .ZN(n1718) );
  CKND2D1BWP12T U1422 ( .A1(n617), .A2(n1701), .ZN(n610) );
  XNR2D1BWP12T U1423 ( .A1(n1718), .A2(n610), .ZN(n1720) );
  CKND2D0BWP12T U1424 ( .A1(n1720), .A2(n3098), .ZN(n611) );
  OAI211D1BWP12T U1425 ( .A1(n3059), .A2(n613), .B(n612), .C(n611), .ZN(n625)
         );
  CKND2D1BWP12T U1426 ( .A1(n2908), .A2(n3091), .ZN(n2836) );
  INVD1BWP12T U1427 ( .I(n614), .ZN(n786) );
  INVD0BWP12T U1428 ( .I(n615), .ZN(n617) );
  CKND2D0BWP12T U1429 ( .A1(n1874), .A2(n3119), .ZN(n623) );
  OAI21D0BWP12T U1430 ( .A1(n2406), .A2(n3066), .B(n3105), .ZN(n621) );
  MUX2ND0BWP12T U1431 ( .I0(n2995), .I1(n2994), .S(n2407), .ZN(n618) );
  NR2D0BWP12T U1432 ( .A1(n618), .A2(n2996), .ZN(n619) );
  MUX2ND0BWP12T U1433 ( .I0(n619), .I1(n3109), .S(n757), .ZN(n620) );
  RCAOI21D0BWP12T U1434 ( .A1(n2407), .A2(n621), .B(n620), .ZN(n622) );
  OAI211D1BWP12T U1435 ( .A1(n2209), .A2(n2836), .B(n623), .C(n622), .ZN(n624)
         );
  AOI211D1BWP12T U1436 ( .A1(n314), .A2(n1799), .B(n625), .C(n624), .ZN(n632)
         );
  NR2D0BWP12T U1437 ( .A1(n2110), .A2(n2956), .ZN(n626) );
  AO211D1BWP12T U1438 ( .A1(n2200), .A2(n2011), .B(n627), .C(n626), .Z(n2667)
         );
  INVD1BWP12T U1439 ( .I(n2667), .ZN(n628) );
  INVD1BWP12T U1440 ( .I(n2448), .ZN(n2459) );
  AOI21D1BWP12T U1441 ( .A1(n628), .A2(n2452), .B(n2459), .ZN(n630) );
  OAI21D1BWP12T U1442 ( .A1(n630), .A2(n629), .B(n2114), .ZN(n2106) );
  ND2XD0BWP12T U1443 ( .A1(n2106), .A2(n3130), .ZN(n631) );
  OAI211D1BWP12T U1444 ( .A1(n2870), .A2(n2141), .B(n632), .C(n631), .ZN(n633)
         );
  AO21D1BWP12T U1445 ( .A1(n1619), .A2(n3126), .B(n633), .Z(result[3]) );
  XNR2XD1BWP12T U1446 ( .A1(n2532), .A2(n2829), .ZN(n1095) );
  XNR2XD1BWP12T U1447 ( .A1(n2532), .A2(n2501), .ZN(n950) );
  OAI22D1BWP12T U1448 ( .A1(n2535), .A2(n1095), .B1(n2533), .B2(n950), .ZN(
        mult_x_18_n907) );
  XNR2XD0BWP12T U1449 ( .A1(n2567), .A2(b[28]), .ZN(n1058) );
  XNR2XD1BWP12T U1450 ( .A1(n2567), .A2(b[29]), .ZN(n2570) );
  OAI22D0BWP12T U1451 ( .A1(n2571), .A2(n1058), .B1(n2569), .B2(n2570), .ZN(
        mult_x_18_n973) );
  XNR2D1BWP12T U1452 ( .A1(n2407), .A2(n2532), .ZN(n1040) );
  XNR2XD1BWP12T U1453 ( .A1(n2542), .A2(n2532), .ZN(n972) );
  OAI22D1BWP12T U1454 ( .A1(n2535), .A2(n1040), .B1(n2533), .B2(n972), .ZN(
        mult_x_18_n911) );
  XNR2D1BWP12T U1455 ( .A1(n2807), .A2(n3110), .ZN(n910) );
  XNR2D1BWP12T U1456 ( .A1(n2829), .A2(n3110), .ZN(n814) );
  OAI22D1BWP12T U1457 ( .A1(n2487), .A2(n910), .B1(n814), .B2(n2486), .ZN(n635) );
  CKBD1BWP12T U1458 ( .I(n2405), .Z(n965) );
  XNR2D1BWP12T U1459 ( .A1(n2764), .A2(n965), .ZN(n879) );
  XNR2D1BWP12T U1460 ( .A1(n2764), .A2(n2407), .ZN(n901) );
  OAI22D1BWP12T U1461 ( .A1(n2514), .A2(n879), .B1(n901), .B2(n2512), .ZN(n634) );
  HA1D0BWP12T U1462 ( .A(n635), .B(n634), .CO(mult_x_18_n719), .S(
        mult_x_18_n720) );
  XNR2XD1BWP12T U1463 ( .A1(n2567), .A2(n2880), .ZN(n835) );
  XNR2XD1BWP12T U1464 ( .A1(n2567), .A2(n2489), .ZN(n905) );
  OAI22D1BWP12T U1465 ( .A1(n2571), .A2(n835), .B1(n2569), .B2(n905), .ZN(
        mult_x_18_n990) );
  XNR2D2BWP12T U1466 ( .A1(n2560), .A2(n2689), .ZN(n2523) );
  XOR2XD1BWP12T U1467 ( .A1(n2689), .A2(n2657), .Z(n636) );
  CKND2D2BWP12T U1468 ( .A1(n2523), .A2(n636), .ZN(n2525) );
  XNR2D0BWP12T U1469 ( .A1(n2657), .A2(n2489), .ZN(n637) );
  XNR2XD1BWP12T U1470 ( .A1(n2657), .A2(b[13]), .ZN(n2524) );
  OAI22D0BWP12T U1471 ( .A1(n2525), .A2(n637), .B1(n2523), .B2(n2524), .ZN(
        mult_x_18_n797) );
  XNR2XD1BWP12T U1472 ( .A1(n2657), .A2(n2880), .ZN(n1071) );
  OAI22D0BWP12T U1473 ( .A1(n2525), .A2(n1071), .B1(n2523), .B2(n637), .ZN(
        mult_x_18_n798) );
  XNR2D2BWP12T U1474 ( .A1(n2633), .A2(n2403), .ZN(n2504) );
  XOR2XD1BWP12T U1475 ( .A1(n2502), .A2(n2403), .Z(n638) );
  CKND2D2BWP12T U1476 ( .A1(n2504), .A2(n638), .ZN(n2506) );
  IND2D0BWP12T U1477 ( .A1(n1064), .B1(n2502), .ZN(n639) );
  OAI22D1BWP12T U1478 ( .A1(n2506), .A2(n1293), .B1(n2504), .B2(n639), .ZN(
        mult_x_18_n735) );
  XNR2XD1BWP12T U1479 ( .A1(n2555), .A2(n2501), .ZN(n1073) );
  XNR2XD1BWP12T U1480 ( .A1(n2555), .A2(n2857), .ZN(n1025) );
  OAI22D1BWP12T U1481 ( .A1(n2559), .A2(n1073), .B1(n2557), .B2(n1025), .ZN(
        mult_x_18_n933) );
  XNR2D1BWP12T U1482 ( .A1(n2502), .A2(n2807), .ZN(n828) );
  XNR2XD1BWP12T U1483 ( .A1(n2502), .A2(n2829), .ZN(n2505) );
  OAI22D0BWP12T U1484 ( .A1(n2506), .A2(n828), .B1(n2504), .B2(n2505), .ZN(
        mult_x_18_n764) );
  XNR2D2BWP12T U1485 ( .A1(n2963), .A2(n2993), .ZN(n2536) );
  XOR2XD1BWP12T U1486 ( .A1(n2633), .A2(n2963), .Z(n640) );
  ND2D3BWP12T U1487 ( .A1(n2536), .A2(n640), .ZN(n2538) );
  XNR2XD1BWP12T U1488 ( .A1(n2633), .A2(n2501), .ZN(n1130) );
  XNR2XD0BWP12T U1489 ( .A1(n2633), .A2(n2857), .ZN(n2537) );
  OAI22D0BWP12T U1490 ( .A1(n2538), .A2(n1130), .B1(n2537), .B2(n2536), .ZN(
        mult_x_18_n773) );
  XNR2XD1BWP12T U1491 ( .A1(a[26]), .A2(n2502), .ZN(n2519) );
  XOR2XD1BWP12T U1492 ( .A1(a[26]), .A2(n2518), .Z(n641) );
  TPND2D1BWP12T U1493 ( .A1(n2519), .A2(n641), .ZN(n2521) );
  XNR2XD0BWP12T U1494 ( .A1(n2542), .A2(n2518), .ZN(n1133) );
  XNR2XD0BWP12T U1495 ( .A1(n2518), .A2(n2766), .ZN(n2520) );
  OAI22D0BWP12T U1496 ( .A1(n2521), .A2(n1133), .B1(n2519), .B2(n2520), .ZN(
        mult_x_18_n757) );
  XNR2XD0BWP12T U1497 ( .A1(n2555), .A2(b[25]), .ZN(n2558) );
  OAI22D0BWP12T U1498 ( .A1(n2559), .A2(n642), .B1(n2557), .B2(n2558), .ZN(
        mult_x_18_n917) );
  NR2D1BWP12T U1499 ( .A1(n643), .A2(n646), .ZN(n1642) );
  OAI21D1BWP12T U1500 ( .A1(n646), .A2(n645), .B(n644), .ZN(n1644) );
  AOI21D1BWP12T U1501 ( .A1(n1650), .A2(n1642), .B(n1644), .ZN(n649) );
  NR2D1BWP12T U1502 ( .A1(mult_x_18_n467), .A2(mult_x_18_n448), .ZN(n1646) );
  INVD1BWP12T U1503 ( .I(n1646), .ZN(n647) );
  ND2D1BWP12T U1504 ( .A1(mult_x_18_n467), .A2(mult_x_18_n448), .ZN(n1645) );
  ND2D1BWP12T U1505 ( .A1(n647), .A2(n1645), .ZN(n648) );
  XOR2XD1BWP12T U1506 ( .A1(n649), .A2(n648), .Z(n1656) );
  INVD1BWP12T U1507 ( .I(n1656), .ZN(n698) );
  CKND0BWP12T U1508 ( .I(b[28]), .ZN(n1205) );
  FA1D0BWP12T U1509 ( .A(n651), .B(n2518), .CI(n650), .CO(n1204), .S(n1829) );
  FA1D2BWP12T U1510 ( .A(n2518), .B(b[27]), .CI(n652), .CO(n1263), .S(n1728)
         );
  CKND2D1BWP12T U1511 ( .A1(n1731), .A2(n3098), .ZN(n693) );
  FA1D2BWP12T U1512 ( .A(n2518), .B(b[27]), .CI(n653), .CO(n1206), .S(n1930)
         );
  ND2D1BWP12T U1513 ( .A1(n1931), .A2(n3119), .ZN(n692) );
  NR2D1BWP12T U1514 ( .A1(n2221), .A2(n2868), .ZN(n2178) );
  AOI222D1BWP12T U1515 ( .A1(n2198), .A2(n1379), .B1(n2187), .B2(n1228), .C1(
        n674), .C2(n2185), .ZN(n2166) );
  INVD1BWP12T U1516 ( .I(n2166), .ZN(n2135) );
  CKND0BWP12T U1517 ( .I(n1246), .ZN(n656) );
  INVD1BWP12T U1518 ( .I(n2183), .ZN(n1351) );
  INVD1BWP12T U1519 ( .I(n2185), .ZN(n1350) );
  OAI22D0BWP12T U1520 ( .A1(n1351), .A2(n682), .B1(n1350), .B2(n1244), .ZN(
        n655) );
  NR2D0BWP12T U1521 ( .A1(n2175), .A2(n1247), .ZN(n654) );
  AOI211D1BWP12T U1522 ( .A1(n656), .A2(n2187), .B(n655), .C(n654), .ZN(n2167)
         );
  NR2D0BWP12T U1523 ( .A1(n2868), .A2(n2157), .ZN(n657) );
  ND2D1BWP12T U1524 ( .A1(n657), .A2(n2221), .ZN(n2179) );
  CKND0BWP12T U1525 ( .I(n1239), .ZN(n660) );
  OAI22D0BWP12T U1526 ( .A1(n1350), .A2(n1238), .B1(n1351), .B2(n1245), .ZN(
        n659) );
  NR2D0BWP12T U1527 ( .A1(n2175), .A2(n1240), .ZN(n658) );
  AOI211XD0BWP12T U1528 ( .A1(n660), .A2(n2187), .B(n659), .C(n658), .ZN(n2165) );
  OAI22D0BWP12T U1529 ( .A1(n2167), .A2(n2179), .B1(n2165), .B2(n2170), .ZN(
        n666) );
  CKND0BWP12T U1530 ( .I(n1233), .ZN(n663) );
  OAI22D0BWP12T U1531 ( .A1(n1350), .A2(n1232), .B1(n1351), .B2(n1241), .ZN(
        n662) );
  MUX2NXD0BWP12T U1532 ( .I0(a[28]), .I1(n2518), .S(n1383), .ZN(n1234) );
  NR2D0BWP12T U1533 ( .A1(n1282), .A2(n1234), .ZN(n661) );
  AOI211D0BWP12T U1534 ( .A1(n663), .A2(n2181), .B(n662), .C(n661), .ZN(n664)
         );
  NR2D0BWP12T U1535 ( .A1(n664), .A2(n2211), .ZN(n665) );
  AO211D1BWP12T U1536 ( .A1(n2178), .A2(n2135), .B(n666), .C(n665), .Z(n2164)
         );
  AOI21D0BWP12T U1537 ( .A1(n2287), .A2(n3107), .B(n2996), .ZN(n672) );
  CKND0BWP12T U1538 ( .I(n2205), .ZN(n667) );
  INVD1BWP12T U1539 ( .I(n2150), .ZN(n2089) );
  MUX2NXD0BWP12T U1540 ( .I0(n2956), .I1(n667), .S(n2089), .ZN(n1420) );
  AOI21D0BWP12T U1541 ( .A1(n2039), .A2(n1420), .B(n2009), .ZN(n2053) );
  CKND2D0BWP12T U1542 ( .A1(n2053), .A2(n3130), .ZN(n671) );
  MUX2ND0BWP12T U1543 ( .I0(n3104), .I1(n3103), .S(b[28]), .ZN(n668) );
  CKND2D0BWP12T U1544 ( .A1(n668), .A2(n3105), .ZN(n669) );
  MUX2NXD0BWP12T U1545 ( .I0(n669), .I1(n3070), .S(n2287), .ZN(n670) );
  OAI211D1BWP12T U1546 ( .A1(n672), .A2(n1205), .B(n671), .C(n670), .ZN(n688)
         );
  INVD0BWP12T U1547 ( .I(n3004), .ZN(n673) );
  ND2D1BWP12T U1548 ( .A1(n673), .A2(n2089), .ZN(n2612) );
  OAI22D0BWP12T U1549 ( .A1(n674), .A2(n1333), .B1(n1379), .B2(n2297), .ZN(
        n676) );
  NR2XD0BWP12T U1550 ( .A1(n1228), .A2(n1329), .ZN(n675) );
  NR2D1BWP12T U1551 ( .A1(n676), .A2(n675), .ZN(n2747) );
  AOI22D0BWP12T U1552 ( .A1(n595), .A2(n1239), .B1(n1238), .B2(n2331), .ZN(
        n678) );
  AOI22D0BWP12T U1553 ( .A1(n2336), .A2(n1245), .B1(n1240), .B2(n2334), .ZN(
        n677) );
  ND2D1BWP12T U1554 ( .A1(n678), .A2(n677), .ZN(n2362) );
  AOI22D0BWP12T U1555 ( .A1(n595), .A2(n1234), .B1(n1241), .B2(n2336), .ZN(
        n680) );
  AOI22D0BWP12T U1556 ( .A1(n2331), .A2(n1232), .B1(n1233), .B2(n2334), .ZN(
        n679) );
  AOI21D0BWP12T U1557 ( .A1(n680), .A2(n679), .B(n2375), .ZN(n681) );
  AOI211D0BWP12T U1558 ( .A1(n2381), .A2(n2362), .B(n681), .C(n2437), .ZN(n686) );
  AOI22D0BWP12T U1559 ( .A1(n595), .A2(n1246), .B1(n682), .B2(n2336), .ZN(n684) );
  AOI22D0BWP12T U1560 ( .A1(n2331), .A2(n1244), .B1(n1247), .B2(n2334), .ZN(
        n683) );
  ND2D1BWP12T U1561 ( .A1(n684), .A2(n683), .ZN(n2361) );
  IND2D1BWP12T U1562 ( .A1(n2407), .B1(n2750), .ZN(n1332) );
  INVD1BWP12T U1563 ( .I(n1332), .ZN(n2340) );
  TPND2D0BWP12T U1564 ( .A1(n2361), .A2(n2340), .ZN(n685) );
  OAI211D0BWP12T U1565 ( .A1(n2747), .A2(n2343), .B(n686), .C(n685), .ZN(n2344) );
  OAI22D1BWP12T U1566 ( .A1(n2612), .A2(n2205), .B1(n2344), .B2(n2903), .ZN(
        n687) );
  RCAOI211D0BWP12T U1567 ( .A1(n2164), .A2(n3091), .B(n688), .C(n687), .ZN(
        n691) );
  HA1D1BWP12T U1568 ( .A(n2291), .B(n689), .CO(n1224), .S(n1986) );
  ND2D1BWP12T U1569 ( .A1(n1983), .A2(n3115), .ZN(n690) );
  ND4D1BWP12T U1570 ( .A1(n693), .A2(n692), .A3(n691), .A4(n690), .ZN(n694) );
  AOI21D1BWP12T U1571 ( .A1(n314), .A2(n1826), .B(n694), .ZN(n697) );
  FA1D1BWP12T U1572 ( .A(n651), .B(n2518), .CI(n695), .CO(n1203), .S(n1549) );
  ND2D1BWP12T U1573 ( .A1(n1554), .A2(n3095), .ZN(n696) );
  OAI211D1BWP12T U1574 ( .A1(n2951), .A2(n698), .B(n697), .C(n696), .ZN(
        result[28]) );
  INVD1P75BWP12T U1575 ( .I(n699), .ZN(n1271) );
  INVD1BWP12T U1576 ( .I(n1270), .ZN(n700) );
  CKND2D1BWP12T U1577 ( .A1(n700), .A2(n1269), .ZN(n701) );
  XOR2XD1BWP12T U1578 ( .A1(n1271), .A2(n701), .Z(n1640) );
  INVD1BWP12T U1579 ( .I(n1640), .ZN(n742) );
  FA1D0BWP12T U1580 ( .A(n703), .B(n2403), .CI(n702), .CO(n1278), .S(n1825) );
  FA1D0BWP12T U1581 ( .A(b[24]), .B(n2403), .CI(n704), .CO(n1314), .S(n1727)
         );
  INVD1BWP12T U1582 ( .I(n1727), .ZN(n737) );
  INVD1BWP12T U1583 ( .I(n3098), .ZN(n2943) );
  FA1D0BWP12T U1584 ( .A(b[24]), .B(n2403), .CI(n705), .CO(n1280), .S(n1926)
         );
  CKND2D1BWP12T U1585 ( .A1(n1926), .A2(n3119), .ZN(n736) );
  HA1D0BWP12T U1586 ( .A(n2293), .B(n706), .CO(n1292), .S(n1982) );
  INVD1BWP12T U1587 ( .I(n1245), .ZN(n1219) );
  CKND0BWP12T U1588 ( .I(n1244), .ZN(n707) );
  AOI22D0BWP12T U1589 ( .A1(n2185), .A2(n1219), .B1(n2183), .B2(n707), .ZN(
        n710) );
  INVD0BWP12T U1590 ( .I(n1240), .ZN(n708) );
  ND2D1BWP12T U1591 ( .A1(n2187), .A2(n708), .ZN(n709) );
  OAI211D1BWP12T U1592 ( .A1(n2175), .A2(n1246), .B(n710), .C(n709), .ZN(n2909) );
  OR3D0BWP12T U1593 ( .A1(n2868), .A2(n2229), .A3(n2905), .Z(n716) );
  CKND0BWP12T U1594 ( .I(n2907), .ZN(n720) );
  CKND2D0BWP12T U1595 ( .A1(n2181), .A2(n1239), .ZN(n713) );
  AOI22D0BWP12T U1596 ( .A1(n2185), .A2(n1241), .B1(n2183), .B2(n1238), .ZN(
        n712) );
  CKND2D0BWP12T U1597 ( .A1(n2187), .A2(n1233), .ZN(n711) );
  TPAOI31D0BWP12T U1598 ( .A1(n713), .A2(n712), .A3(n711), .B(n2211), .ZN(n714) );
  AOI211XD0BWP12T U1599 ( .A1(n2178), .A2(n720), .B(n714), .C(n2157), .ZN(n715) );
  OAI211D1BWP12T U1600 ( .A1(n2170), .A2(n2909), .B(n716), .C(n715), .ZN(n2224) );
  NR2D1BWP12T U1601 ( .A1(n2224), .A2(n3012), .ZN(n734) );
  CKND0BWP12T U1602 ( .I(n2343), .ZN(n808) );
  AOI22D0BWP12T U1603 ( .A1(n2336), .A2(n1238), .B1(n1239), .B2(n2334), .ZN(
        n718) );
  AOI22D0BWP12T U1604 ( .A1(n595), .A2(n1233), .B1(n1241), .B2(n2331), .ZN(
        n717) );
  AOI21D0BWP12T U1605 ( .A1(n718), .A2(n717), .B(n2375), .ZN(n719) );
  AOI211D0BWP12T U1606 ( .A1(n808), .A2(n720), .B(n719), .C(n2437), .ZN(n724)
         );
  AOI22D0BWP12T U1607 ( .A1(n2336), .A2(n1244), .B1(n1246), .B2(n2334), .ZN(
        n722) );
  AOI22D0BWP12T U1608 ( .A1(n595), .A2(n1240), .B1(n1245), .B2(n2331), .ZN(
        n721) );
  ND2D1BWP12T U1609 ( .A1(n722), .A2(n721), .ZN(n2352) );
  ND2XD0BWP12T U1610 ( .A1(n2352), .A2(n2381), .ZN(n723) );
  OAI211D1BWP12T U1611 ( .A1(n725), .A2(n1332), .B(n724), .C(n723), .ZN(n2391)
         );
  OAI21D0BWP12T U1612 ( .A1(n2403), .A2(n3066), .B(n3105), .ZN(n730) );
  CKND2D1BWP12T U1613 ( .A1(n2039), .A2(n2197), .ZN(n1301) );
  INVD1BWP12T U1614 ( .I(n1301), .ZN(n2021) );
  NR2D0BWP12T U1615 ( .A1(n2021), .A2(n3044), .ZN(n729) );
  MUX2ND0BWP12T U1616 ( .I0(n2995), .I1(n2994), .S(b[24]), .ZN(n726) );
  NR2D0BWP12T U1617 ( .A1(n726), .A2(n2996), .ZN(n727) );
  MUX2ND0BWP12T U1618 ( .I0(n727), .I1(n3109), .S(n2293), .ZN(n728) );
  RCAOI211D0BWP12T U1619 ( .A1(b[24]), .A2(n730), .B(n729), .C(n728), .ZN(n732) );
  NR2D1BWP12T U1620 ( .A1(n2040), .A2(n3044), .ZN(n1258) );
  INVD1BWP12T U1621 ( .I(n1258), .ZN(n3005) );
  CKND2D1BWP12T U1622 ( .A1(n3004), .A2(n3005), .ZN(n2899) );
  CKND2D1BWP12T U1623 ( .A1(n2899), .A2(n2207), .ZN(n731) );
  OAI211D1BWP12T U1624 ( .A1(n2903), .A2(n2391), .B(n732), .C(n731), .ZN(n733)
         );
  AOI211D1BWP12T U1625 ( .A1(n1982), .A2(n3115), .B(n734), .C(n733), .ZN(n735)
         );
  OAI211D1BWP12T U1626 ( .A1(n737), .A2(n2943), .B(n736), .C(n735), .ZN(n738)
         );
  AOI21D1BWP12T U1627 ( .A1(n314), .A2(n1825), .B(n738), .ZN(n741) );
  FA1D0BWP12T U1628 ( .A(n703), .B(n2403), .CI(n739), .CO(n1277), .S(n1548) );
  CKND2D1BWP12T U1629 ( .A1(n1548), .A2(n3095), .ZN(n740) );
  OAI211D1BWP12T U1630 ( .A1(n2951), .A2(n742), .B(n741), .C(n740), .ZN(
        result[24]) );
  TPOAI22D0BWP12T U1631 ( .A1(n2000), .A2(n2687), .B1(n1999), .B2(n2998), .ZN(
        n744) );
  OAI22D1BWP12T U1632 ( .A1(n2002), .A2(n2928), .B1(n2001), .B2(n2659), .ZN(
        n743) );
  NR2D1BWP12T U1633 ( .A1(n744), .A2(n743), .ZN(n2111) );
  OAI22D1BWP12T U1634 ( .A1(n2000), .A2(n2965), .B1(n1999), .B2(n2292), .ZN(
        n746) );
  OAI22D1BWP12T U1635 ( .A1(n2002), .A2(n2293), .B1(n2001), .B2(n2636), .ZN(
        n745) );
  NR2D1BWP12T U1636 ( .A1(n746), .A2(n745), .ZN(n2028) );
  MUX2NXD0BWP12T U1637 ( .I0(n2111), .I1(n2028), .S(n2405), .ZN(n2037) );
  NR2D1BWP12T U1638 ( .A1(n2037), .A2(n2407), .ZN(n2162) );
  NR2XD0BWP12T U1639 ( .A1(n747), .A2(n2133), .ZN(n748) );
  NR2D1BWP12T U1640 ( .A1(n2162), .A2(n748), .ZN(n768) );
  INVD0BWP12T U1641 ( .I(n2110), .ZN(n767) );
  CKND2D1BWP12T U1642 ( .A1(n1225), .A2(n767), .ZN(n749) );
  ND2D1BWP12T U1643 ( .A1(n768), .A2(n749), .ZN(n2041) );
  TPOAI21D0BWP12T U1644 ( .A1(n2041), .A2(n2437), .B(n2448), .ZN(n764) );
  OAI22D1BWP12T U1645 ( .A1(n2000), .A2(n3067), .B1(n3033), .B2(n1999), .ZN(
        n751) );
  OAI22D1BWP12T U1646 ( .A1(n2416), .A2(n2002), .B1(n2001), .B2(n2874), .ZN(
        n750) );
  NR2D1BWP12T U1647 ( .A1(n751), .A2(n750), .ZN(n2109) );
  OAI22D1BWP12T U1648 ( .A1(n2000), .A2(n2280), .B1(n1999), .B2(n2275), .ZN(
        n753) );
  OAI22D1BWP12T U1649 ( .A1(n2002), .A2(n2893), .B1(n2001), .B2(n2722), .ZN(
        n752) );
  NR2D1BWP12T U1650 ( .A1(n753), .A2(n752), .ZN(n2113) );
  TPNR2D0BWP12T U1651 ( .A1(n2113), .A2(n2110), .ZN(n754) );
  AOI211D1BWP12T U1652 ( .A1(n2109), .A2(n2200), .B(n754), .C(n2750), .ZN(n763) );
  OAI22D1BWP12T U1653 ( .A1(n2000), .A2(n2802), .B1(n1999), .B2(n2853), .ZN(
        n756) );
  OAI22D1BWP12T U1654 ( .A1(n2002), .A2(n2282), .B1(n2001), .B2(n2831), .ZN(
        n755) );
  NR2D1BWP12T U1655 ( .A1(n756), .A2(n755), .ZN(n2112) );
  CKND2D0BWP12T U1656 ( .A1(n2112), .A2(n2405), .ZN(n761) );
  AOI21D1BWP12T U1657 ( .A1(n2070), .A2(n1937), .B(n2407), .ZN(n760) );
  AOI22D1BWP12T U1658 ( .A1(n2071), .A2(n757), .B1(n2073), .B2(n2768), .ZN(
        n759) );
  ND2XD0BWP12T U1659 ( .A1(n2072), .A2(n2749), .ZN(n758) );
  ND4D1BWP12T U1660 ( .A1(n761), .A2(n760), .A3(n759), .A4(n758), .ZN(n762) );
  CKND2D1BWP12T U1661 ( .A1(n763), .A2(n762), .ZN(n771) );
  AOI21D1BWP12T U1662 ( .A1(n764), .A2(n771), .B(n2101), .ZN(n2118) );
  CKND2D1BWP12T U1663 ( .A1(n1613), .A2(n3126), .ZN(n813) );
  INVD1BWP12T U1664 ( .I(n2201), .ZN(n2204) );
  TPND2D0BWP12T U1665 ( .A1(n2204), .A2(n767), .ZN(n770) );
  INVD1BWP12T U1666 ( .I(n768), .ZN(n769) );
  INR2D1BWP12T U1667 ( .A1(n770), .B1(n769), .ZN(n2455) );
  ND2D1BWP12T U1668 ( .A1(n2455), .A2(n2452), .ZN(n772) );
  INVD1BWP12T U1669 ( .I(n771), .ZN(n805) );
  AOI21D1BWP12T U1670 ( .A1(n772), .A2(n2448), .B(n805), .ZN(n2450) );
  INVD1BWP12T U1671 ( .I(n773), .ZN(n1524) );
  OAI21D1BWP12T U1672 ( .A1(n1524), .A2(n1520), .B(n1521), .ZN(n777) );
  CKND2D1BWP12T U1673 ( .A1(n797), .A2(n775), .ZN(n776) );
  XNR2D1BWP12T U1674 ( .A1(n777), .A2(n776), .ZN(n1526) );
  INVD1BWP12T U1675 ( .I(n1526), .ZN(n803) );
  INVD1BWP12T U1676 ( .I(n778), .ZN(n1711) );
  OAI21D1BWP12T U1677 ( .A1(n1711), .A2(n1707), .B(n1708), .ZN(n782) );
  ND2XD0BWP12T U1678 ( .A1(n785), .A2(n780), .ZN(n781) );
  XNR2D1BWP12T U1679 ( .A1(n782), .A2(n781), .ZN(n1712) );
  INVD1BWP12T U1680 ( .I(n3094), .ZN(n793) );
  CKND0BWP12T U1681 ( .I(n783), .ZN(n785) );
  MUX2ND0BWP12T U1682 ( .I0(n3104), .I1(n3103), .S(n2405), .ZN(n787) );
  AOI21D0BWP12T U1683 ( .A1(n3105), .A2(n787), .B(n1937), .ZN(n790) );
  AOI21D0BWP12T U1684 ( .A1(n3107), .A2(n1937), .B(n2996), .ZN(n788) );
  OAI22D0BWP12T U1685 ( .A1(n788), .A2(n2297), .B1(n2404), .B2(n3109), .ZN(
        n789) );
  RCAOI211D0BWP12T U1686 ( .A1(n1869), .A2(n3119), .B(n790), .C(n789), .ZN(
        n791) );
  OAI21D1BWP12T U1687 ( .A1(n793), .A2(n792), .B(n791), .ZN(n794) );
  AOI21D1BWP12T U1688 ( .A1(n3098), .A2(n1712), .B(n794), .ZN(n802) );
  INVD0BWP12T U1689 ( .I(n795), .ZN(n797) );
  CKND2D1BWP12T U1690 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2XD1BWP12T U1691 ( .A1(n799), .A2(n798), .Z(n1793) );
  XNR2D0BWP12T U1692 ( .A1(n800), .A2(n2404), .ZN(n1956) );
  AOI22D0BWP12T U1693 ( .A1(n1793), .A2(n314), .B1(n3115), .B2(n1956), .ZN(
        n801) );
  OAI211D1BWP12T U1694 ( .A1(n3059), .A2(n803), .B(n802), .C(n801), .ZN(n811)
         );
  INVD1BWP12T U1695 ( .I(n804), .ZN(n2159) );
  TPNR2D0BWP12T U1696 ( .A1(n2037), .A2(n1332), .ZN(n806) );
  AOI211D1BWP12T U1697 ( .A1(n808), .A2(n807), .B(n806), .C(n805), .ZN(n809)
         );
  AOI21D1BWP12T U1698 ( .A1(n2159), .A2(n2908), .B(n809), .ZN(n2137) );
  NR2D1BWP12T U1699 ( .A1(n2137), .A2(n3012), .ZN(n810) );
  AOI211D1BWP12T U1700 ( .A1(n2450), .A2(n3052), .B(n811), .C(n810), .ZN(n812)
         );
  OAI211D2BWP12T U1701 ( .A1(n2118), .A2(n3044), .B(n813), .C(n812), .ZN(
        result[2]) );
  XNR2D1BWP12T U1702 ( .A1(n3110), .A2(n2501), .ZN(n873) );
  OAI22D1BWP12T U1703 ( .A1(n2487), .A2(n814), .B1(n873), .B2(n2486), .ZN(n817) );
  INR2D1BWP12T U1704 ( .A1(n1382), .B1(n2533), .ZN(n816) );
  XNR2XD1BWP12T U1705 ( .A1(n2567), .A2(n2766), .ZN(n872) );
  XNR2D1BWP12T U1706 ( .A1(n2567), .A2(n2807), .ZN(n846) );
  OAI22D1BWP12T U1707 ( .A1(n2571), .A2(n872), .B1(n2569), .B2(n846), .ZN(n815) );
  XNR2XD1BWP12T U1708 ( .A1(n3110), .A2(n2880), .ZN(n1007) );
  XNR2D1BWP12T U1709 ( .A1(n3110), .A2(n2489), .ZN(n913) );
  OAI22D1BWP12T U1710 ( .A1(n2487), .A2(n1007), .B1(n913), .B2(n2486), .ZN(
        n820) );
  INVD12BWP12T U1711 ( .I(n2876), .ZN(n2494) );
  INR2D1BWP12T U1712 ( .A1(n1382), .B1(n2539), .ZN(n819) );
  XNR2XD1BWP12T U1713 ( .A1(n2567), .A2(n2857), .ZN(n930) );
  XNR2XD1BWP12T U1714 ( .A1(n2567), .A2(n3074), .ZN(n836) );
  OAI22D1BWP12T U1715 ( .A1(n2571), .A2(n930), .B1(n2569), .B2(n836), .ZN(n818) );
  XOR2XD1BWP12T U1716 ( .A1(n2494), .A2(n3067), .Z(n821) );
  XNR2XD4BWP12T U1717 ( .A1(n2532), .A2(n3067), .ZN(n2495) );
  CKND2D8BWP12T U1718 ( .A1(n821), .A2(n2495), .ZN(n2498) );
  XNR2D0BWP12T U1719 ( .A1(n2494), .A2(b[20]), .ZN(n1116) );
  XNR2D0BWP12T U1720 ( .A1(n2494), .A2(b[21]), .ZN(n2497) );
  OAI22D0BWP12T U1721 ( .A1(n2498), .A2(n1116), .B1(n2497), .B2(n2495), .ZN(
        mult_x_18_n869) );
  XOR2D1BWP12T U1722 ( .A1(n3033), .A2(n2416), .Z(n822) );
  CKND2D2BWP12T U1723 ( .A1(n2539), .A2(n822), .ZN(n2541) );
  XNR2D0BWP12T U1724 ( .A1(n3033), .A2(b[18]), .ZN(n1097) );
  XNR2XD0BWP12T U1725 ( .A1(n3033), .A2(n2663), .ZN(n2540) );
  OAI22D0BWP12T U1726 ( .A1(n2541), .A2(n1097), .B1(n2539), .B2(n2540), .ZN(
        mult_x_18_n848) );
  HA1D0BWP12T U1727 ( .A(n824), .B(n823), .CO(mult_x_18_n726), .S(n259) );
  XNR2XD1BWP12T U1728 ( .A1(n3110), .A2(b[30]), .ZN(n1087) );
  XNR2XD1BWP12T U1729 ( .A1(n3110), .A2(b[31]), .ZN(n2485) );
  OAI22D1BWP12T U1730 ( .A1(n2487), .A2(n1087), .B1(n2485), .B2(n2486), .ZN(
        n2530) );
  XNR2XD1BWP12T U1731 ( .A1(n2608), .A2(a[30]), .ZN(n2548) );
  IND2D0BWP12T U1732 ( .A1(n1382), .B1(n2956), .ZN(n825) );
  OAI22D1BWP12T U1733 ( .A1(n2551), .A2(n2305), .B1(n2548), .B2(n825), .ZN(
        n2529) );
  XNR2XD4BWP12T U1734 ( .A1(a[14]), .A2(n3033), .ZN(n2515) );
  XOR2XD1BWP12T U1735 ( .A1(a[14]), .A2(n2720), .Z(n826) );
  ND2D3BWP12T U1736 ( .A1(n2515), .A2(n826), .ZN(n2517) );
  XNR2D0BWP12T U1737 ( .A1(n2720), .A2(b[15]), .ZN(n1089) );
  XNR2XD0BWP12T U1738 ( .A1(n2720), .A2(b[16]), .ZN(n1129) );
  TPOAI22D0BWP12T U1739 ( .A1(n2517), .A2(n1089), .B1(n2515), .B2(n1129), .ZN(
        mult_x_18_n830) );
  XNR2XD1BWP12T U1740 ( .A1(n2993), .A2(n2857), .ZN(n995) );
  TPOAI22D0BWP12T U1741 ( .A1(n2493), .A2(n995), .B1(n2491), .B2(n827), .ZN(
        mult_x_18_n785) );
  XNR2XD1BWP12T U1742 ( .A1(n2764), .A2(b[26]), .ZN(n1098) );
  XNR2XD1BWP12T U1743 ( .A1(n2764), .A2(b[27]), .ZN(n2513) );
  OAI22D0BWP12T U1744 ( .A1(n2514), .A2(n1098), .B1(n2513), .B2(n2512), .ZN(
        mult_x_18_n944) );
  XNR2XD1BWP12T U1745 ( .A1(n2502), .A2(n2766), .ZN(n988) );
  TPOAI22D0BWP12T U1746 ( .A1(n2506), .A2(n988), .B1(n2504), .B2(n828), .ZN(
        mult_x_18_n765) );
  IND2D0BWP12T U1747 ( .A1(n1064), .B1(n2993), .ZN(n829) );
  OAI22D1BWP12T U1748 ( .A1(n2493), .A2(n1952), .B1(n2491), .B2(n829), .ZN(
        n832) );
  XNR2D1BWP12T U1749 ( .A1(n2494), .A2(n3074), .ZN(n954) );
  XNR2XD1BWP12T U1750 ( .A1(n2494), .A2(n2880), .ZN(n907) );
  OAI22D1BWP12T U1751 ( .A1(n2498), .A2(n954), .B1(n907), .B2(n2495), .ZN(n831) );
  XNR2XD1BWP12T U1752 ( .A1(n2567), .A2(b[18]), .ZN(n854) );
  XNR2XD1BWP12T U1753 ( .A1(n2567), .A2(n2663), .ZN(n908) );
  OAI22D1BWP12T U1754 ( .A1(n2571), .A2(n854), .B1(n2569), .B2(n908), .ZN(n830) );
  FA1D0BWP12T U1755 ( .A(n832), .B(n831), .CI(n830), .CO(mult_x_18_n584), .S(
        mult_x_18_n585) );
  IND2D0BWP12T U1756 ( .A1(n1064), .B1(n3033), .ZN(n833) );
  OAI22D1BWP12T U1757 ( .A1(n2541), .A2(n834), .B1(n2539), .B2(n833), .ZN(n839) );
  XNR2D1BWP12T U1758 ( .A1(n2764), .A2(n2501), .ZN(n1050) );
  XNR2D1BWP12T U1759 ( .A1(n2764), .A2(n2857), .ZN(n1125) );
  OAI22D1BWP12T U1760 ( .A1(n2514), .A2(n1050), .B1(n1125), .B2(n2512), .ZN(
        n838) );
  OAI22D1BWP12T U1761 ( .A1(n2571), .A2(n836), .B1(n2569), .B2(n835), .ZN(n837) );
  FA1D0BWP12T U1762 ( .A(n839), .B(n838), .CI(n837), .CO(mult_x_18_n678), .S(
        mult_x_18_n679) );
  INR2D1BWP12T U1763 ( .A1(n1382), .B1(n2536), .ZN(mult_x_18_n782) );
  XNR2XD1BWP12T U1764 ( .A1(n3110), .A2(b[23]), .ZN(n1017) );
  XNR2XD1BWP12T U1765 ( .A1(n3110), .A2(b[24]), .ZN(n956) );
  OAI22D1BWP12T U1766 ( .A1(n2487), .A2(n1017), .B1(n956), .B2(n2486), .ZN(
        n842) );
  INR2D1BWP12T U1767 ( .A1(n1382), .B1(n2504), .ZN(n841) );
  XNR2D0BWP12T U1768 ( .A1(n2567), .A2(b[21]), .ZN(n1067) );
  XNR2D0BWP12T U1769 ( .A1(n2567), .A2(b[22]), .ZN(n850) );
  OAI22D1BWP12T U1770 ( .A1(n2571), .A2(n1067), .B1(n2569), .B2(n850), .ZN(
        n840) );
  FA1D0BWP12T U1771 ( .A(n842), .B(n841), .CI(n840), .CO(mult_x_18_n538), .S(
        mult_x_18_n539) );
  IND2D0BWP12T U1772 ( .A1(n1064), .B1(n2532), .ZN(n843) );
  OAI22D1BWP12T U1773 ( .A1(n2535), .A2(n844), .B1(n2533), .B2(n843), .ZN(n849) );
  XNR2XD1BWP12T U1774 ( .A1(n1382), .A2(n2532), .ZN(n845) );
  XNR2D1BWP12T U1775 ( .A1(n3102), .A2(n2532), .ZN(n886) );
  OAI22D1BWP12T U1776 ( .A1(n2535), .A2(n845), .B1(n2533), .B2(n886), .ZN(n848) );
  XNR2XD1BWP12T U1777 ( .A1(n2567), .A2(n2829), .ZN(n1044) );
  OAI22D1BWP12T U1778 ( .A1(n2571), .A2(n846), .B1(n2569), .B2(n1044), .ZN(
        n847) );
  FA1D0BWP12T U1779 ( .A(n849), .B(n848), .CI(n847), .CO(mult_x_18_n707), .S(
        mult_x_18_n708) );
  INR2D1BWP12T U1780 ( .A1(n1382), .B1(n2495), .ZN(mult_x_18_n890) );
  XNR2XD1BWP12T U1781 ( .A1(n2633), .A2(n2829), .ZN(n1131) );
  XNR2XD1BWP12T U1782 ( .A1(n2608), .A2(n998), .ZN(n975) );
  XNR2XD1BWP12T U1783 ( .A1(n2567), .A2(b[26]), .ZN(n862) );
  XNR2D0BWP12T U1784 ( .A1(n2567), .A2(b[27]), .ZN(n1059) );
  XNR2XD1BWP12T U1785 ( .A1(n2494), .A2(n2522), .ZN(n927) );
  XNR2XD1BWP12T U1786 ( .A1(n2494), .A2(b[15]), .ZN(n934) );
  OAI22D1BWP12T U1787 ( .A1(n2498), .A2(n927), .B1(n934), .B2(n2495), .ZN(n853) );
  XNR2XD1BWP12T U1788 ( .A1(n2633), .A2(n965), .ZN(n883) );
  XNR2XD1BWP12T U1789 ( .A1(n2407), .A2(n2633), .ZN(n947) );
  OAI22D1BWP12T U1790 ( .A1(n2538), .A2(n883), .B1(n947), .B2(n2536), .ZN(n852) );
  XNR2D0BWP12T U1791 ( .A1(n2567), .A2(b[23]), .ZN(n877) );
  OAI22D1BWP12T U1792 ( .A1(n2571), .A2(n850), .B1(n2569), .B2(n877), .ZN(n851) );
  FA1D0BWP12T U1793 ( .A(n853), .B(n852), .CI(n851), .CO(mult_x_18_n519), .S(
        mult_x_18_n520) );
  XNR2XD1BWP12T U1794 ( .A1(n3110), .A2(n2663), .ZN(n963) );
  XNR2XD1BWP12T U1795 ( .A1(n3110), .A2(b[20]), .ZN(n892) );
  OAI22D1BWP12T U1796 ( .A1(n2487), .A2(n963), .B1(n892), .B2(n2486), .ZN(n857) );
  INR2D1BWP12T U1797 ( .A1(n1382), .B1(n2491), .ZN(n856) );
  XNR2XD1BWP12T U1798 ( .A1(n2567), .A2(b[17]), .ZN(n1029) );
  OAI22D1BWP12T U1799 ( .A1(n2571), .A2(n1029), .B1(n2569), .B2(n854), .ZN(
        n855) );
  FA1D0BWP12T U1800 ( .A(n857), .B(n856), .CI(n855), .CO(mult_x_18_n600), .S(
        mult_x_18_n601) );
  XNR2D1BWP12T U1801 ( .A1(n3110), .A2(b[15]), .ZN(n935) );
  XNR2D1BWP12T U1802 ( .A1(n3110), .A2(b[16]), .ZN(n1035) );
  OAI22D1BWP12T U1803 ( .A1(n2487), .A2(n935), .B1(n1035), .B2(n2486), .ZN(
        n860) );
  XNR2XD4BWP12T U1804 ( .A1(n2720), .A2(n2891), .ZN(n2561) );
  INR2D1BWP12T U1805 ( .A1(n1382), .B1(n2561), .ZN(n859) );
  XNR2XD1BWP12T U1806 ( .A1(n2567), .A2(b[13]), .ZN(n904) );
  XNR2XD1BWP12T U1807 ( .A1(n2567), .A2(n2522), .ZN(n868) );
  OAI22D1BWP12T U1808 ( .A1(n2571), .A2(n904), .B1(n2569), .B2(n868), .ZN(n858) );
  FA1D0BWP12T U1809 ( .A(n860), .B(n859), .CI(n858), .CO(mult_x_18_n650), .S(
        mult_x_18_n651) );
  XNR2XD1BWP12T U1810 ( .A1(n3110), .A2(b[27]), .ZN(n981) );
  OAI22D1BWP12T U1811 ( .A1(n2487), .A2(n981), .B1(n861), .B2(n2486), .ZN(n865) );
  INR2D1BWP12T U1812 ( .A1(n1382), .B1(n2543), .ZN(n864) );
  XNR2D0BWP12T U1813 ( .A1(n2567), .A2(b[25]), .ZN(n888) );
  OAI22D1BWP12T U1814 ( .A1(n2571), .A2(n888), .B1(n2569), .B2(n862), .ZN(n863) );
  FA1D0BWP12T U1815 ( .A(n865), .B(n864), .CI(n863), .CO(mult_x_18_n464), .S(
        mult_x_18_n465) );
  INR2D1BWP12T U1816 ( .A1(n1382), .B1(n2515), .ZN(mult_x_18_n846) );
  INR2D1BWP12T U1817 ( .A1(n1382), .B1(n2548), .ZN(mult_x_18_n750) );
  INR2D1BWP12T U1818 ( .A1(n1382), .B1(n2557), .ZN(mult_x_18_n942) );
  INR2D1BWP12T U1819 ( .A1(n1382), .B1(n2523), .ZN(mult_x_18_n810) );
  XNR2D1BWP12T U1820 ( .A1(n2494), .A2(n2807), .ZN(n931) );
  XNR2XD1BWP12T U1821 ( .A1(n2494), .A2(n2829), .ZN(n1048) );
  OAI22D1BWP12T U1822 ( .A1(n2498), .A2(n931), .B1(n1048), .B2(n2495), .ZN(
        n871) );
  XOR2XD1BWP12T U1823 ( .A1(n2560), .A2(n2891), .Z(n866) );
  CKND2D2BWP12T U1824 ( .A1(n2561), .A2(n866), .ZN(n2564) );
  XNR2D1BWP12T U1825 ( .A1(n2560), .A2(n1382), .ZN(n867) );
  XNR2D1BWP12T U1826 ( .A1(n2560), .A2(n3102), .ZN(n974) );
  OAI22D1BWP12T U1827 ( .A1(n2564), .A2(n867), .B1(n974), .B2(n2561), .ZN(n870) );
  XNR2XD1BWP12T U1828 ( .A1(n2567), .A2(b[15]), .ZN(n887) );
  OAI22D1BWP12T U1829 ( .A1(n2571), .A2(n868), .B1(n2569), .B2(n887), .ZN(n869) );
  FA1D0BWP12T U1830 ( .A(n871), .B(n870), .CI(n869), .CO(mult_x_18_n637), .S(
        mult_x_18_n638) );
  INR2D1BWP12T U1831 ( .A1(n1382), .B1(n2519), .ZN(mult_x_18_n762) );
  XNR2XD1BWP12T U1832 ( .A1(n2764), .A2(b[16]), .ZN(n1077) );
  XNR2XD1BWP12T U1833 ( .A1(n2764), .A2(b[17]), .ZN(n882) );
  OAI22D1BWP12T U1834 ( .A1(n2514), .A2(n1077), .B1(n882), .B2(n2512), .ZN(
        mult_x_18_n954) );
  XNR2XD1BWP12T U1835 ( .A1(n3110), .A2(b[21]), .ZN(n891) );
  XNR2XD1BWP12T U1836 ( .A1(n3110), .A2(b[22]), .ZN(n1018) );
  OAI22D1BWP12T U1837 ( .A1(n2487), .A2(n891), .B1(n1018), .B2(n2486), .ZN(
        mult_x_18_n1013) );
  XNR2XD1BWP12T U1838 ( .A1(n2532), .A2(b[13]), .ZN(n922) );
  XNR2XD1BWP12T U1839 ( .A1(n2532), .A2(n2522), .ZN(n1003) );
  OAI22D1BWP12T U1840 ( .A1(n2535), .A2(n922), .B1(n2533), .B2(n1003), .ZN(
        mult_x_18_n901) );
  XNR2XD1BWP12T U1841 ( .A1(n2542), .A2(n2567), .ZN(n978) );
  OAI22D1BWP12T U1842 ( .A1(n2571), .A2(n978), .B1(n2569), .B2(n872), .ZN(
        mult_x_18_n997) );
  XNR2D1BWP12T U1843 ( .A1(n2764), .A2(n3074), .ZN(n1124) );
  XNR2XD1BWP12T U1844 ( .A1(n2764), .A2(n2880), .ZN(n903) );
  OAI22D1BWP12T U1845 ( .A1(n2514), .A2(n1124), .B1(n903), .B2(n2512), .ZN(
        mult_x_18_n960) );
  XNR2D1BWP12T U1846 ( .A1(n3110), .A2(n2857), .ZN(n878) );
  OAI22D1BWP12T U1847 ( .A1(n2487), .A2(n873), .B1(n878), .B2(n2486), .ZN(n875) );
  XNR2D1BWP12T U1848 ( .A1(n2764), .A2(n2542), .ZN(n900) );
  XNR2D1BWP12T U1849 ( .A1(n2764), .A2(n2766), .ZN(n899) );
  OAI22D1BWP12T U1850 ( .A1(n2514), .A2(n900), .B1(n899), .B2(n2512), .ZN(n874) );
  XNR2XD1BWP12T U1851 ( .A1(n1382), .A2(n2657), .ZN(n876) );
  XNR2XD1BWP12T U1852 ( .A1(n998), .A2(n2657), .ZN(n881) );
  OAI22D1BWP12T U1853 ( .A1(n2525), .A2(n876), .B1(n2523), .B2(n881), .ZN(
        mult_x_18_n809) );
  XNR2D0BWP12T U1854 ( .A1(n2567), .A2(b[24]), .ZN(n889) );
  OAI22D1BWP12T U1855 ( .A1(n2571), .A2(n877), .B1(n2569), .B2(n889), .ZN(
        mult_x_18_n978) );
  XNR2D1BWP12T U1856 ( .A1(n3110), .A2(n3074), .ZN(n1008) );
  OAI22D1BWP12T U1857 ( .A1(n2487), .A2(n878), .B1(n1008), .B2(n2486), .ZN(
        mult_x_18_n1025) );
  OAI22D1BWP12T U1858 ( .A1(n2514), .A2(n880), .B1(n879), .B2(n2512), .ZN(
        mult_x_18_n969) );
  XNR2XD1BWP12T U1859 ( .A1(n3033), .A2(n2857), .ZN(n1122) );
  XNR2XD1BWP12T U1860 ( .A1(n3033), .A2(n3074), .ZN(n921) );
  OAI22D1BWP12T U1861 ( .A1(n2541), .A2(n1122), .B1(n2539), .B2(n921), .ZN(
        mult_x_18_n857) );
  XNR2D1BWP12T U1862 ( .A1(n2547), .A2(n2657), .ZN(n898) );
  OAI22D1BWP12T U1863 ( .A1(n2525), .A2(n881), .B1(n2523), .B2(n898), .ZN(
        mult_x_18_n808) );
  XNR2XD1BWP12T U1864 ( .A1(n2764), .A2(b[22]), .ZN(n897) );
  XNR2XD1BWP12T U1865 ( .A1(n2764), .A2(b[23]), .ZN(n953) );
  OAI22D1BWP12T U1866 ( .A1(n2514), .A2(n897), .B1(n953), .B2(n2512), .ZN(
        mult_x_18_n948) );
  XNR2XD1BWP12T U1867 ( .A1(n2764), .A2(n2522), .ZN(n1000) );
  XNR2XD1BWP12T U1868 ( .A1(n2764), .A2(b[15]), .ZN(n1078) );
  OAI22D1BWP12T U1869 ( .A1(n2514), .A2(n1000), .B1(n1078), .B2(n2512), .ZN(
        mult_x_18_n956) );
  XNR2D1BWP12T U1870 ( .A1(n2764), .A2(n2489), .ZN(n902) );
  XNR2D1BWP12T U1871 ( .A1(n2764), .A2(b[13]), .ZN(n1001) );
  OAI22D1BWP12T U1872 ( .A1(n2514), .A2(n902), .B1(n1001), .B2(n2512), .ZN(
        mult_x_18_n958) );
  XNR2XD1BWP12T U1873 ( .A1(n3102), .A2(n2518), .ZN(n1053) );
  XNR2D1BWP12T U1874 ( .A1(n2547), .A2(n2518), .ZN(n1033) );
  OAI22D1BWP12T U1875 ( .A1(n2521), .A2(n1053), .B1(n1033), .B2(n2519), .ZN(
        mult_x_18_n760) );
  XNR2XD1BWP12T U1876 ( .A1(n2764), .A2(b[18]), .ZN(n993) );
  OAI22D1BWP12T U1877 ( .A1(n2514), .A2(n882), .B1(n993), .B2(n2512), .ZN(
        mult_x_18_n953) );
  XNR2XD1BWP12T U1878 ( .A1(n2633), .A2(n3102), .ZN(n884) );
  OAI22D1BWP12T U1879 ( .A1(n2538), .A2(n884), .B1(n883), .B2(n2536), .ZN(
        mult_x_18_n780) );
  XNR2XD1BWP12T U1880 ( .A1(n1382), .A2(n2633), .ZN(n885) );
  OAI22D1BWP12T U1881 ( .A1(n2538), .A2(n885), .B1(n884), .B2(n2536), .ZN(
        mult_x_18_n781) );
  XNR2D1BWP12T U1882 ( .A1(n2547), .A2(n2532), .ZN(n1041) );
  OAI22D1BWP12T U1883 ( .A1(n2535), .A2(n886), .B1(n2533), .B2(n1041), .ZN(
        mult_x_18_n913) );
  XNR2XD1BWP12T U1884 ( .A1(n2567), .A2(b[16]), .ZN(n1030) );
  OAI22D1BWP12T U1885 ( .A1(n2571), .A2(n887), .B1(n2569), .B2(n1030), .ZN(
        mult_x_18_n986) );
  OAI22D1BWP12T U1886 ( .A1(n2571), .A2(n889), .B1(n2569), .B2(n888), .ZN(
        mult_x_18_n977) );
  XNR2XD1BWP12T U1887 ( .A1(n1382), .A2(n2555), .ZN(n890) );
  XNR2D1BWP12T U1888 ( .A1(n3102), .A2(n2555), .ZN(n951) );
  OAI22D1BWP12T U1889 ( .A1(n2559), .A2(n890), .B1(n2557), .B2(n951), .ZN(
        mult_x_18_n941) );
  OAI22D1BWP12T U1890 ( .A1(n2487), .A2(n892), .B1(n891), .B2(n2486), .ZN(n894) );
  XNR2D1BWP12T U1891 ( .A1(n2560), .A2(n2542), .ZN(n928) );
  XNR2D1BWP12T U1892 ( .A1(n2560), .A2(n2766), .ZN(n906) );
  OAI22D1BWP12T U1893 ( .A1(n2564), .A2(n928), .B1(n906), .B2(n2561), .ZN(n893) );
  HA1D1BWP12T U1894 ( .A(n894), .B(n893), .CO(mult_x_18_n586), .S(
        mult_x_18_n587) );
  XNR2XD1BWP12T U1895 ( .A1(n2532), .A2(n2663), .ZN(n1119) );
  XNR2XD1BWP12T U1896 ( .A1(n2532), .A2(b[20]), .ZN(n945) );
  OAI22D1BWP12T U1897 ( .A1(n2535), .A2(n1119), .B1(n2533), .B2(n945), .ZN(
        mult_x_18_n895) );
  XNR2XD1BWP12T U1898 ( .A1(n2555), .A2(b[20]), .ZN(n1031) );
  XNR2XD1BWP12T U1899 ( .A1(n2555), .A2(b[21]), .ZN(n948) );
  OAI22D1BWP12T U1900 ( .A1(n2559), .A2(n1031), .B1(n2557), .B2(n948), .ZN(
        mult_x_18_n921) );
  IND2D0BWP12T U1901 ( .A1(n1064), .B1(n2555), .ZN(n895) );
  OAI22D1BWP12T U1902 ( .A1(n2559), .A2(n896), .B1(n2557), .B2(n895), .ZN(
        mult_x_18_n744) );
  XNR2XD1BWP12T U1903 ( .A1(n2764), .A2(b[21]), .ZN(n918) );
  OAI22D1BWP12T U1904 ( .A1(n2514), .A2(n918), .B1(n897), .B2(n2512), .ZN(
        mult_x_18_n949) );
  XNR2XD1BWP12T U1905 ( .A1(n2555), .A2(b[15]), .ZN(n980) );
  XNR2XD1BWP12T U1906 ( .A1(n2555), .A2(b[16]), .ZN(n1056) );
  OAI22D1BWP12T U1907 ( .A1(n2559), .A2(n980), .B1(n2557), .B2(n1056), .ZN(
        mult_x_18_n926) );
  XNR2XD1BWP12T U1908 ( .A1(n3033), .A2(b[13]), .ZN(n1057) );
  XNR2XD1BWP12T U1909 ( .A1(n3033), .A2(n2522), .ZN(n1086) );
  OAI22D1BWP12T U1910 ( .A1(n2541), .A2(n1057), .B1(n2539), .B2(n1086), .ZN(
        mult_x_18_n853) );
  XNR2XD1BWP12T U1911 ( .A1(n2407), .A2(n2657), .ZN(n1028) );
  OAI22D1BWP12T U1912 ( .A1(n2525), .A2(n898), .B1(n2523), .B2(n1028), .ZN(
        mult_x_18_n807) );
  XNR2D1BWP12T U1913 ( .A1(n2993), .A2(n2807), .ZN(n1079) );
  XNR2XD1BWP12T U1914 ( .A1(n2993), .A2(n2829), .ZN(n949) );
  OAI22D1BWP12T U1915 ( .A1(n2493), .A2(n1079), .B1(n2491), .B2(n949), .ZN(
        mult_x_18_n788) );
  XNR2D1BWP12T U1916 ( .A1(n2764), .A2(n2807), .ZN(n917) );
  OAI22D1BWP12T U1917 ( .A1(n2514), .A2(n899), .B1(n917), .B2(n2512), .ZN(
        mult_x_18_n965) );
  XNR2D1BWP12T U1918 ( .A1(n3110), .A2(b[17]), .ZN(n1034) );
  XNR2D1BWP12T U1919 ( .A1(n3110), .A2(b[18]), .ZN(n964) );
  OAI22D1BWP12T U1920 ( .A1(n2487), .A2(n1034), .B1(n964), .B2(n2486), .ZN(
        mult_x_18_n1017) );
  XNR2XD1BWP12T U1921 ( .A1(n2633), .A2(n2542), .ZN(n946) );
  XNR2XD1BWP12T U1922 ( .A1(n2633), .A2(n2766), .ZN(n1063) );
  OAI22D1BWP12T U1923 ( .A1(n2538), .A2(n946), .B1(n1063), .B2(n2536), .ZN(
        mult_x_18_n777) );
  OAI22D1BWP12T U1924 ( .A1(n2514), .A2(n901), .B1(n900), .B2(n2512), .ZN(
        mult_x_18_n967) );
  OAI22D1BWP12T U1925 ( .A1(n2514), .A2(n903), .B1(n902), .B2(n2512), .ZN(
        mult_x_18_n959) );
  OAI22D1BWP12T U1926 ( .A1(n2571), .A2(n905), .B1(n2569), .B2(n904), .ZN(
        mult_x_18_n989) );
  XNR2D1BWP12T U1927 ( .A1(n2720), .A2(n2501), .ZN(n1091) );
  XNR2D1BWP12T U1928 ( .A1(n2720), .A2(n2857), .ZN(n962) );
  OAI22D1BWP12T U1929 ( .A1(n2517), .A2(n1091), .B1(n2515), .B2(n962), .ZN(
        mult_x_18_n837) );
  XNR2XD1BWP12T U1930 ( .A1(n3110), .A2(b[25]), .ZN(n955) );
  XNR2XD1BWP12T U1931 ( .A1(n3110), .A2(b[26]), .ZN(n982) );
  OAI22D1BWP12T U1932 ( .A1(n2487), .A2(n955), .B1(n982), .B2(n2486), .ZN(
        mult_x_18_n1009) );
  XNR2D1BWP12T U1933 ( .A1(n2560), .A2(n2807), .ZN(n1020) );
  OAI22D1BWP12T U1934 ( .A1(n2564), .A2(n906), .B1(n1020), .B2(n2561), .ZN(
        mult_x_18_n821) );
  XNR2D1BWP12T U1935 ( .A1(n2494), .A2(n2489), .ZN(n933) );
  OAI22D1BWP12T U1936 ( .A1(n2498), .A2(n907), .B1(n933), .B2(n2495), .ZN(
        mult_x_18_n878) );
  XNR2XD1BWP12T U1937 ( .A1(n2567), .A2(b[20]), .ZN(n1068) );
  OAI22D1BWP12T U1938 ( .A1(n2571), .A2(n908), .B1(n2569), .B2(n1068), .ZN(
        mult_x_18_n982) );
  XNR2D0BWP12T U1939 ( .A1(n1382), .A2(n2993), .ZN(n909) );
  XNR2XD1BWP12T U1940 ( .A1(n3102), .A2(n2993), .ZN(n1106) );
  OAI22D1BWP12T U1941 ( .A1(n2493), .A2(n909), .B1(n2491), .B2(n1106), .ZN(
        mult_x_18_n794) );
  XNR2D1BWP12T U1942 ( .A1(n3110), .A2(b[13]), .ZN(n912) );
  XNR2D1BWP12T U1943 ( .A1(n3110), .A2(n2522), .ZN(n936) );
  OAI22D1BWP12T U1944 ( .A1(n2487), .A2(n912), .B1(n936), .B2(n2486), .ZN(
        mult_x_18_n1021) );
  XNR2XD1BWP12T U1945 ( .A1(n2494), .A2(b[18]), .ZN(n1100) );
  XNR2XD1BWP12T U1946 ( .A1(n2494), .A2(n2663), .ZN(n1117) );
  OAI22D1BWP12T U1947 ( .A1(n2498), .A2(n1100), .B1(n1117), .B2(n2495), .ZN(
        mult_x_18_n871) );
  XNR2XD1BWP12T U1948 ( .A1(n2494), .A2(n2407), .ZN(n914) );
  XNR2D1BWP12T U1949 ( .A1(n2494), .A2(n2542), .ZN(n938) );
  OAI22D1BWP12T U1950 ( .A1(n2498), .A2(n914), .B1(n938), .B2(n2495), .ZN(
        mult_x_18_n886) );
  OAI22D1BWP12T U1951 ( .A1(n2487), .A2(n911), .B1(n910), .B2(n2486), .ZN(
        mult_x_18_n1029) );
  XNR2XD1BWP12T U1952 ( .A1(n2532), .A2(b[15]), .ZN(n1002) );
  XNR2XD1BWP12T U1953 ( .A1(n2532), .A2(b[16]), .ZN(n920) );
  OAI22D1BWP12T U1954 ( .A1(n2535), .A2(n1002), .B1(n2533), .B2(n920), .ZN(
        mult_x_18_n899) );
  XNR2D1BWP12T U1955 ( .A1(n3102), .A2(n3033), .ZN(n942) );
  XNR2D1BWP12T U1956 ( .A1(n2547), .A2(n3033), .ZN(n1049) );
  OAI22D1BWP12T U1957 ( .A1(n2541), .A2(n942), .B1(n2539), .B2(n1049), .ZN(
        mult_x_18_n865) );
  OAI22D1BWP12T U1958 ( .A1(n2487), .A2(n913), .B1(n912), .B2(n2486), .ZN(n916) );
  XNR2D1BWP12T U1959 ( .A1(n2494), .A2(n965), .ZN(n1135) );
  OAI22D1BWP12T U1960 ( .A1(n2498), .A2(n1135), .B1(n914), .B2(n2495), .ZN(
        n915) );
  HA1D1BWP12T U1961 ( .A(n916), .B(n915), .CO(mult_x_18_n680), .S(
        mult_x_18_n681) );
  XNR2D1BWP12T U1962 ( .A1(n2764), .A2(n2829), .ZN(n1051) );
  OAI22D1BWP12T U1963 ( .A1(n2514), .A2(n917), .B1(n1051), .B2(n2512), .ZN(
        mult_x_18_n964) );
  XNR2D0BWP12T U1964 ( .A1(n2764), .A2(b[20]), .ZN(n941) );
  OAI22D1BWP12T U1965 ( .A1(n2514), .A2(n941), .B1(n918), .B2(n2512), .ZN(
        mult_x_18_n950) );
  XNR2XD1BWP12T U1966 ( .A1(n2407), .A2(n2502), .ZN(n1014) );
  XNR2XD1BWP12T U1967 ( .A1(n2542), .A2(n2502), .ZN(n989) );
  OAI22D1BWP12T U1968 ( .A1(n2506), .A2(n1014), .B1(n2504), .B2(n989), .ZN(
        mult_x_18_n767) );
  XNR2XD1BWP12T U1969 ( .A1(n2532), .A2(n2880), .ZN(n1107) );
  XNR2XD1BWP12T U1970 ( .A1(n2532), .A2(n2489), .ZN(n923) );
  OAI22D1BWP12T U1971 ( .A1(n2535), .A2(n1107), .B1(n2533), .B2(n923), .ZN(
        mult_x_18_n903) );
  XNR2XD1BWP12T U1972 ( .A1(n2532), .A2(b[17]), .ZN(n919) );
  XNR2D0BWP12T U1973 ( .A1(n2532), .A2(b[18]), .ZN(n1120) );
  OAI22D1BWP12T U1974 ( .A1(n2535), .A2(n919), .B1(n2533), .B2(n1120), .ZN(
        mult_x_18_n897) );
  OAI22D1BWP12T U1975 ( .A1(n2535), .A2(n920), .B1(n2533), .B2(n919), .ZN(
        mult_x_18_n898) );
  XNR2XD1BWP12T U1976 ( .A1(n3033), .A2(n2880), .ZN(n1085) );
  OAI22D1BWP12T U1977 ( .A1(n2541), .A2(n921), .B1(n2539), .B2(n1085), .ZN(
        mult_x_18_n856) );
  XNR2D1BWP12T U1978 ( .A1(n2657), .A2(n2807), .ZN(n926) );
  XNR2D0BWP12T U1979 ( .A1(n2657), .A2(n2829), .ZN(n1052) );
  OAI22D1BWP12T U1980 ( .A1(n2525), .A2(n926), .B1(n2523), .B2(n1052), .ZN(
        mult_x_18_n803) );
  XNR2D1BWP12T U1981 ( .A1(n2560), .A2(n2857), .ZN(n957) );
  XNR2D1BWP12T U1982 ( .A1(n2560), .A2(n3074), .ZN(n984) );
  OAI22D1BWP12T U1983 ( .A1(n2564), .A2(n957), .B1(n984), .B2(n2561), .ZN(
        mult_x_18_n817) );
  OAI22D1BWP12T U1984 ( .A1(n2535), .A2(n923), .B1(n2533), .B2(n922), .ZN(
        mult_x_18_n902) );
  XNR2D0BWP12T U1985 ( .A1(n1382), .A2(n2502), .ZN(n924) );
  XNR2XD1BWP12T U1986 ( .A1(n3102), .A2(n2502), .ZN(n960) );
  OAI22D1BWP12T U1987 ( .A1(n2506), .A2(n924), .B1(n2504), .B2(n960), .ZN(
        mult_x_18_n770) );
  IND2D0BWP12T U1988 ( .A1(n1382), .B1(n2518), .ZN(n925) );
  OAI22D1BWP12T U1989 ( .A1(n2521), .A2(n2291), .B1(n2519), .B2(n925), .ZN(
        mult_x_18_n734) );
  XNR2XD1BWP12T U1990 ( .A1(n2657), .A2(n2766), .ZN(n1126) );
  OAI22D1BWP12T U1991 ( .A1(n2525), .A2(n1126), .B1(n2523), .B2(n926), .ZN(
        mult_x_18_n804) );
  XNR2XD1BWP12T U1992 ( .A1(n2494), .A2(b[13]), .ZN(n932) );
  OAI22D1BWP12T U1993 ( .A1(n2498), .A2(n932), .B1(n927), .B2(n2495), .ZN(
        mult_x_18_n876) );
  XNR2XD1BWP12T U1994 ( .A1(n2560), .A2(n2880), .ZN(n983) );
  XNR2D1BWP12T U1995 ( .A1(n2560), .A2(n2489), .ZN(n1016) );
  OAI22D1BWP12T U1996 ( .A1(n2564), .A2(n983), .B1(n1016), .B2(n2561), .ZN(
        mult_x_18_n815) );
  XNR2D1BWP12T U1997 ( .A1(n2560), .A2(n2407), .ZN(n966) );
  OAI22D1BWP12T U1998 ( .A1(n2564), .A2(n966), .B1(n928), .B2(n2561), .ZN(
        mult_x_18_n823) );
  XNR2D1BWP12T U1999 ( .A1(n2494), .A2(n1382), .ZN(n929) );
  XNR2XD1BWP12T U2000 ( .A1(n2494), .A2(n3102), .ZN(n1136) );
  OAI22D1BWP12T U2001 ( .A1(n2498), .A2(n929), .B1(n1136), .B2(n2495), .ZN(
        mult_x_18_n889) );
  XNR2XD1BWP12T U2002 ( .A1(n2567), .A2(n2501), .ZN(n1043) );
  OAI22D1BWP12T U2003 ( .A1(n2571), .A2(n1043), .B1(n2569), .B2(n930), .ZN(
        mult_x_18_n993) );
  XNR2D1BWP12T U2004 ( .A1(n2494), .A2(n2766), .ZN(n937) );
  OAI22D1BWP12T U2005 ( .A1(n2498), .A2(n937), .B1(n931), .B2(n2495), .ZN(
        mult_x_18_n884) );
  OAI22D1BWP12T U2006 ( .A1(n2498), .A2(n933), .B1(n932), .B2(n2495), .ZN(
        mult_x_18_n877) );
  XNR2XD1BWP12T U2007 ( .A1(n2494), .A2(b[16]), .ZN(n952) );
  OAI22D1BWP12T U2008 ( .A1(n2498), .A2(n934), .B1(n952), .B2(n2495), .ZN(
        mult_x_18_n874) );
  OAI22D1BWP12T U2009 ( .A1(n2487), .A2(n936), .B1(n935), .B2(n2486), .ZN(n940) );
  OAI22D1BWP12T U2010 ( .A1(n2498), .A2(n938), .B1(n937), .B2(n2495), .ZN(n939) );
  XNR2XD1BWP12T U2011 ( .A1(n2764), .A2(n2663), .ZN(n992) );
  OAI22D1BWP12T U2012 ( .A1(n2514), .A2(n992), .B1(n941), .B2(n2512), .ZN(
        mult_x_18_n951) );
  XNR2XD1BWP12T U2013 ( .A1(n1382), .A2(n3033), .ZN(n943) );
  OAI22D1BWP12T U2014 ( .A1(n2541), .A2(n943), .B1(n2539), .B2(n942), .ZN(
        mult_x_18_n866) );
  OAI22D1BWP12T U2015 ( .A1(n2535), .A2(n945), .B1(n2533), .B2(n944), .ZN(
        mult_x_18_n894) );
  OAI22D1BWP12T U2016 ( .A1(n2538), .A2(n947), .B1(n946), .B2(n2536), .ZN(
        mult_x_18_n778) );
  XNR2XD1BWP12T U2017 ( .A1(n2555), .A2(b[22]), .ZN(n1005) );
  OAI22D1BWP12T U2018 ( .A1(n2559), .A2(n948), .B1(n2557), .B2(n1005), .ZN(
        mult_x_18_n920) );
  XNR2XD1BWP12T U2019 ( .A1(n2993), .A2(n2501), .ZN(n996) );
  OAI22D1BWP12T U2020 ( .A1(n2493), .A2(n949), .B1(n2491), .B2(n996), .ZN(
        mult_x_18_n787) );
  XNR2XD1BWP12T U2021 ( .A1(n2542), .A2(n2555), .ZN(n1012) );
  XNR2XD1BWP12T U2022 ( .A1(n2555), .A2(n2766), .ZN(n991) );
  OAI22D1BWP12T U2023 ( .A1(n2559), .A2(n1012), .B1(n2557), .B2(n991), .ZN(
        mult_x_18_n937) );
  XNR2XD1BWP12T U2024 ( .A1(n2532), .A2(n2857), .ZN(n1069) );
  OAI22D1BWP12T U2025 ( .A1(n2535), .A2(n950), .B1(n2533), .B2(n1069), .ZN(
        mult_x_18_n906) );
  XNR2D1BWP12T U2026 ( .A1(n2720), .A2(n3074), .ZN(n961) );
  XNR2XD1BWP12T U2027 ( .A1(n2720), .A2(n2880), .ZN(n1110) );
  OAI22D1BWP12T U2028 ( .A1(n2517), .A2(n961), .B1(n2515), .B2(n1110), .ZN(
        mult_x_18_n835) );
  XNR2D1BWP12T U2029 ( .A1(n2547), .A2(n2555), .ZN(n969) );
  OAI22D1BWP12T U2030 ( .A1(n2559), .A2(n951), .B1(n2557), .B2(n969), .ZN(
        mult_x_18_n940) );
  XNR2D1BWP12T U2031 ( .A1(n2547), .A2(n2993), .ZN(n1105) );
  XNR2XD1BWP12T U2032 ( .A1(n2407), .A2(n2993), .ZN(n971) );
  OAI22D1BWP12T U2033 ( .A1(n2493), .A2(n1105), .B1(n2491), .B2(n971), .ZN(
        mult_x_18_n792) );
  XNR2XD1BWP12T U2034 ( .A1(n2494), .A2(b[17]), .ZN(n1101) );
  OAI22D1BWP12T U2035 ( .A1(n2498), .A2(n952), .B1(n1101), .B2(n2495), .ZN(
        mult_x_18_n873) );
  XNR2XD1BWP12T U2036 ( .A1(n2555), .A2(b[17]), .ZN(n1055) );
  XNR2XD1BWP12T U2037 ( .A1(n2555), .A2(b[18]), .ZN(n997) );
  OAI22D1BWP12T U2038 ( .A1(n2559), .A2(n1055), .B1(n2557), .B2(n997), .ZN(
        mult_x_18_n924) );
  XNR2XD1BWP12T U2039 ( .A1(n2764), .A2(b[24]), .ZN(n1027) );
  OAI22D1BWP12T U2040 ( .A1(n2514), .A2(n953), .B1(n1027), .B2(n2512), .ZN(
        mult_x_18_n947) );
  XNR2D1BWP12T U2041 ( .A1(n2494), .A2(n2857), .ZN(n1006) );
  OAI22D1BWP12T U2042 ( .A1(n2498), .A2(n1006), .B1(n954), .B2(n2495), .ZN(
        mult_x_18_n880) );
  OAI22D1BWP12T U2043 ( .A1(n2487), .A2(n956), .B1(n955), .B2(n2486), .ZN(n959) );
  XNR2D1BWP12T U2044 ( .A1(n2560), .A2(n2501), .ZN(n970) );
  OAI22D1BWP12T U2045 ( .A1(n2564), .A2(n970), .B1(n957), .B2(n2561), .ZN(n958) );
  XNR2XD1BWP12T U2046 ( .A1(n2547), .A2(n2502), .ZN(n1015) );
  OAI22D1BWP12T U2047 ( .A1(n2506), .A2(n960), .B1(n2504), .B2(n1015), .ZN(
        mult_x_18_n769) );
  OAI22D1BWP12T U2048 ( .A1(n2517), .A2(n962), .B1(n2515), .B2(n961), .ZN(
        mult_x_18_n836) );
  OAI22D1BWP12T U2049 ( .A1(n2487), .A2(n964), .B1(n963), .B2(n2486), .ZN(n968) );
  XNR2D1BWP12T U2050 ( .A1(n2560), .A2(n965), .ZN(n973) );
  OAI22D1BWP12T U2051 ( .A1(n2564), .A2(n973), .B1(n966), .B2(n2561), .ZN(n967) );
  XNR2D1BWP12T U2052 ( .A1(n2407), .A2(n2555), .ZN(n1013) );
  OAI22D1BWP12T U2053 ( .A1(n2559), .A2(n969), .B1(n2557), .B2(n1013), .ZN(
        mult_x_18_n939) );
  XNR2D1BWP12T U2054 ( .A1(n2560), .A2(n2829), .ZN(n1019) );
  OAI22D1BWP12T U2055 ( .A1(n2564), .A2(n1019), .B1(n970), .B2(n2561), .ZN(
        mult_x_18_n819) );
  XNR2XD1BWP12T U2056 ( .A1(n2542), .A2(n2993), .ZN(n977) );
  OAI22D1BWP12T U2057 ( .A1(n2493), .A2(n971), .B1(n2491), .B2(n977), .ZN(
        mult_x_18_n791) );
  XNR2XD1BWP12T U2058 ( .A1(n2532), .A2(n2766), .ZN(n990) );
  OAI22D1BWP12T U2059 ( .A1(n2535), .A2(n972), .B1(n2533), .B2(n990), .ZN(
        mult_x_18_n910) );
  OAI22D1BWP12T U2060 ( .A1(n2564), .A2(n974), .B1(n973), .B2(n2561), .ZN(
        mult_x_18_n825) );
  XNR2XD1BWP12T U2061 ( .A1(n2547), .A2(n2608), .ZN(n1121) );
  OAI22D1BWP12T U2062 ( .A1(n2546), .A2(n975), .B1(n1121), .B2(n2543), .ZN(
        mult_x_18_n753) );
  XNR2XD1BWP12T U2063 ( .A1(n1382), .A2(n2720), .ZN(n976) );
  XNR2XD1BWP12T U2064 ( .A1(n3102), .A2(n2720), .ZN(n994) );
  OAI22D1BWP12T U2065 ( .A1(n2517), .A2(n976), .B1(n2515), .B2(n994), .ZN(
        mult_x_18_n845) );
  XNR2XD1BWP12T U2066 ( .A1(n2993), .A2(n2766), .ZN(n1080) );
  OAI22D1BWP12T U2067 ( .A1(n2493), .A2(n977), .B1(n2491), .B2(n1080), .ZN(
        mult_x_18_n790) );
  OAI22D1BWP12T U2068 ( .A1(n2571), .A2(n979), .B1(n2569), .B2(n978), .ZN(
        mult_x_18_n998) );
  XNR2XD1BWP12T U2069 ( .A1(n2555), .A2(n2522), .ZN(n987) );
  OAI22D1BWP12T U2070 ( .A1(n2559), .A2(n987), .B1(n2557), .B2(n980), .ZN(
        mult_x_18_n927) );
  OAI22D1BWP12T U2071 ( .A1(n2487), .A2(n982), .B1(n981), .B2(n2486), .ZN(n986) );
  OAI22D1BWP12T U2072 ( .A1(n2564), .A2(n984), .B1(n983), .B2(n2561), .ZN(n985) );
  XNR2XD1BWP12T U2073 ( .A1(n2555), .A2(b[13]), .ZN(n1042) );
  OAI22D1BWP12T U2074 ( .A1(n2559), .A2(n1042), .B1(n2557), .B2(n987), .ZN(
        mult_x_18_n928) );
  OAI22D1BWP12T U2075 ( .A1(n2506), .A2(n989), .B1(n2504), .B2(n988), .ZN(
        mult_x_18_n766) );
  XNR2D1BWP12T U2076 ( .A1(n2532), .A2(n2807), .ZN(n1096) );
  OAI22D1BWP12T U2077 ( .A1(n2535), .A2(n990), .B1(n2533), .B2(n1096), .ZN(
        mult_x_18_n909) );
  XNR2XD1BWP12T U2078 ( .A1(n2542), .A2(n2720), .ZN(n1112) );
  XNR2XD1BWP12T U2079 ( .A1(n2720), .A2(n2766), .ZN(n1094) );
  OAI22D1BWP12T U2080 ( .A1(n2517), .A2(n1112), .B1(n2515), .B2(n1094), .ZN(
        mult_x_18_n841) );
  XNR2D1BWP12T U2081 ( .A1(n2555), .A2(n2807), .ZN(n1061) );
  OAI22D1BWP12T U2082 ( .A1(n2559), .A2(n991), .B1(n2557), .B2(n1061), .ZN(
        mult_x_18_n936) );
  OAI22D1BWP12T U2083 ( .A1(n2514), .A2(n993), .B1(n992), .B2(n2512), .ZN(
        mult_x_18_n952) );
  XNR2D1BWP12T U2084 ( .A1(n2547), .A2(n2720), .ZN(n1060) );
  OAI22D1BWP12T U2085 ( .A1(n2517), .A2(n994), .B1(n2515), .B2(n1060), .ZN(
        mult_x_18_n844) );
  OAI22D1BWP12T U2086 ( .A1(n2493), .A2(n996), .B1(n2491), .B2(n995), .ZN(
        mult_x_18_n786) );
  XNR2D0BWP12T U2087 ( .A1(n2555), .A2(n2663), .ZN(n1032) );
  OAI22D1BWP12T U2088 ( .A1(n2559), .A2(n997), .B1(n2557), .B2(n1032), .ZN(
        mult_x_18_n923) );
  XNR2XD1BWP12T U2089 ( .A1(n1382), .A2(n2956), .ZN(n999) );
  XNR2XD1BWP12T U2090 ( .A1(n2956), .A2(n998), .ZN(n2550) );
  OAI22D1BWP12T U2091 ( .A1(n2551), .A2(n999), .B1(n2550), .B2(n2548), .ZN(
        mult_x_18_n749) );
  OAI22D1BWP12T U2092 ( .A1(n2514), .A2(n1001), .B1(n1000), .B2(n2512), .ZN(
        mult_x_18_n957) );
  OAI22D1BWP12T U2093 ( .A1(n2535), .A2(n1003), .B1(n2533), .B2(n1002), .ZN(
        mult_x_18_n900) );
  OAI22D1BWP12T U2094 ( .A1(n2559), .A2(n1005), .B1(n2557), .B2(n1004), .ZN(
        mult_x_18_n919) );
  XNR2D1BWP12T U2095 ( .A1(n2494), .A2(n2501), .ZN(n1047) );
  OAI22D1BWP12T U2096 ( .A1(n2498), .A2(n1047), .B1(n1006), .B2(n2495), .ZN(
        mult_x_18_n881) );
  OAI22D1BWP12T U2097 ( .A1(n2487), .A2(n1008), .B1(n1007), .B2(n2486), .ZN(
        n1011) );
  IND2D0BWP12T U2098 ( .A1(n1064), .B1(n2494), .ZN(n1009) );
  OAI22D1BWP12T U2099 ( .A1(n2498), .A2(n375), .B1(n2495), .B2(n1009), .ZN(
        n1010) );
  OAI22D1BWP12T U2100 ( .A1(n2559), .A2(n1013), .B1(n2557), .B2(n1012), .ZN(
        mult_x_18_n938) );
  OAI22D1BWP12T U2101 ( .A1(n2506), .A2(n1015), .B1(n1014), .B2(n2504), .ZN(
        mult_x_18_n768) );
  XNR2D1BWP12T U2102 ( .A1(n2560), .A2(b[13]), .ZN(n1128) );
  OAI22D1BWP12T U2103 ( .A1(n2564), .A2(n1016), .B1(n1128), .B2(n2561), .ZN(
        mult_x_18_n814) );
  OAI22D1BWP12T U2104 ( .A1(n2487), .A2(n1018), .B1(n1017), .B2(n2486), .ZN(
        n1022) );
  OAI22D1BWP12T U2105 ( .A1(n2564), .A2(n1020), .B1(n1019), .B2(n2561), .ZN(
        n1021) );
  CKND0BWP12T U2106 ( .I(n2720), .ZN(n1024) );
  IND2D0BWP12T U2107 ( .A1(n1064), .B1(n2720), .ZN(n1023) );
  OAI22D1BWP12T U2108 ( .A1(n2517), .A2(n1024), .B1(n2515), .B2(n1023), .ZN(
        mult_x_18_n740) );
  XNR2XD1BWP12T U2109 ( .A1(n2555), .A2(n3074), .ZN(n1026) );
  OAI22D1BWP12T U2110 ( .A1(n2559), .A2(n1025), .B1(n2557), .B2(n1026), .ZN(
        mult_x_18_n932) );
  XNR2XD1BWP12T U2111 ( .A1(n2555), .A2(n2880), .ZN(n1103) );
  OAI22D1BWP12T U2112 ( .A1(n2559), .A2(n1026), .B1(n2557), .B2(n1103), .ZN(
        mult_x_18_n931) );
  XNR2XD1BWP12T U2113 ( .A1(n2764), .A2(b[25]), .ZN(n1099) );
  OAI22D1BWP12T U2114 ( .A1(n2514), .A2(n1027), .B1(n1099), .B2(n2512), .ZN(
        mult_x_18_n946) );
  XNR2XD1BWP12T U2115 ( .A1(n2542), .A2(n2657), .ZN(n1127) );
  OAI22D1BWP12T U2116 ( .A1(n2525), .A2(n1028), .B1(n2523), .B2(n1127), .ZN(
        mult_x_18_n806) );
  XNR2D1BWP12T U2117 ( .A1(n2720), .A2(n2807), .ZN(n1093) );
  XNR2XD1BWP12T U2118 ( .A1(n2720), .A2(n2829), .ZN(n1092) );
  OAI22D1BWP12T U2119 ( .A1(n2517), .A2(n1093), .B1(n2515), .B2(n1092), .ZN(
        mult_x_18_n839) );
  OAI22D1BWP12T U2120 ( .A1(n2571), .A2(n1030), .B1(n2569), .B2(n1029), .ZN(
        mult_x_18_n985) );
  OAI22D1BWP12T U2121 ( .A1(n2559), .A2(n1032), .B1(n2557), .B2(n1031), .ZN(
        mult_x_18_n922) );
  XNR2XD1BWP12T U2122 ( .A1(n2407), .A2(n2518), .ZN(n1134) );
  OAI22D1BWP12T U2123 ( .A1(n2521), .A2(n1033), .B1(n1134), .B2(n2519), .ZN(
        mult_x_18_n759) );
  OAI22D1BWP12T U2124 ( .A1(n2487), .A2(n1035), .B1(n1034), .B2(n2486), .ZN(
        n1039) );
  CKND0BWP12T U2125 ( .I(n2560), .ZN(n1037) );
  IND2D0BWP12T U2126 ( .A1(n1064), .B1(n2560), .ZN(n1036) );
  OAI22D1BWP12T U2127 ( .A1(n2564), .A2(n1037), .B1(n2561), .B2(n1036), .ZN(
        n1038) );
  OAI22D1BWP12T U2128 ( .A1(n2535), .A2(n1041), .B1(n2533), .B2(n1040), .ZN(
        mult_x_18_n912) );
  XNR2XD1BWP12T U2129 ( .A1(n2555), .A2(n2489), .ZN(n1102) );
  OAI22D1BWP12T U2130 ( .A1(n2559), .A2(n1102), .B1(n2557), .B2(n1042), .ZN(
        mult_x_18_n929) );
  XNR2XD1BWP12T U2131 ( .A1(n3033), .A2(n2766), .ZN(n1082) );
  XNR2D1BWP12T U2132 ( .A1(n3033), .A2(n2807), .ZN(n1066) );
  OAI22D1BWP12T U2133 ( .A1(n2541), .A2(n1082), .B1(n2539), .B2(n1066), .ZN(
        mult_x_18_n861) );
  OAI22D1BWP12T U2134 ( .A1(n2571), .A2(n1044), .B1(n2569), .B2(n1043), .ZN(
        mult_x_18_n994) );
  CKND0BWP12T U2135 ( .I(n2657), .ZN(n1046) );
  IND2D0BWP12T U2136 ( .A1(n1064), .B1(n2657), .ZN(n1045) );
  OAI22D1BWP12T U2137 ( .A1(n2525), .A2(n1046), .B1(n2523), .B2(n1045), .ZN(
        mult_x_18_n738) );
  OAI22D1BWP12T U2138 ( .A1(n2498), .A2(n1048), .B1(n1047), .B2(n2495), .ZN(
        mult_x_18_n882) );
  XNR2D1BWP12T U2139 ( .A1(n2407), .A2(n3033), .ZN(n1070) );
  OAI22D1BWP12T U2140 ( .A1(n2541), .A2(n1049), .B1(n2539), .B2(n1070), .ZN(
        mult_x_18_n864) );
  OAI22D1BWP12T U2141 ( .A1(n2514), .A2(n1051), .B1(n1050), .B2(n2512), .ZN(
        mult_x_18_n963) );
  XNR2XD1BWP12T U2142 ( .A1(n2657), .A2(n2501), .ZN(n1076) );
  OAI22D1BWP12T U2143 ( .A1(n2525), .A2(n1052), .B1(n2523), .B2(n1076), .ZN(
        mult_x_18_n802) );
  XNR2XD1BWP12T U2144 ( .A1(n1382), .A2(n2518), .ZN(n1054) );
  OAI22D1BWP12T U2145 ( .A1(n2521), .A2(n1054), .B1(n2519), .B2(n1053), .ZN(
        mult_x_18_n761) );
  OAI22D1BWP12T U2146 ( .A1(n2559), .A2(n1056), .B1(n2557), .B2(n1055), .ZN(
        mult_x_18_n925) );
  XNR2XD1BWP12T U2147 ( .A1(n3033), .A2(n2489), .ZN(n1084) );
  OAI22D1BWP12T U2148 ( .A1(n2541), .A2(n1084), .B1(n2539), .B2(n1057), .ZN(
        mult_x_18_n854) );
  XNR2XD1BWP12T U2149 ( .A1(n2657), .A2(n2857), .ZN(n1075) );
  XNR2XD1BWP12T U2150 ( .A1(n2657), .A2(n3074), .ZN(n1072) );
  OAI22D1BWP12T U2151 ( .A1(n2525), .A2(n1075), .B1(n2523), .B2(n1072), .ZN(
        mult_x_18_n800) );
  OAI22D1BWP12T U2152 ( .A1(n2571), .A2(n1059), .B1(n2569), .B2(n1058), .ZN(
        mult_x_18_n974) );
  XNR2XD1BWP12T U2153 ( .A1(n2407), .A2(n2720), .ZN(n1113) );
  OAI22D1BWP12T U2154 ( .A1(n2517), .A2(n1060), .B1(n2515), .B2(n1113), .ZN(
        mult_x_18_n843) );
  XNR2XD1BWP12T U2155 ( .A1(n2555), .A2(n2829), .ZN(n1074) );
  OAI22D1BWP12T U2156 ( .A1(n2559), .A2(n1061), .B1(n2557), .B2(n1074), .ZN(
        mult_x_18_n935) );
  OAI22D1BWP12T U2157 ( .A1(n2538), .A2(n1063), .B1(n1062), .B2(n2536), .ZN(
        mult_x_18_n776) );
  IND2D0BWP12T U2158 ( .A1(n1064), .B1(n2633), .ZN(n1065) );
  OAI22D1BWP12T U2159 ( .A1(n2538), .A2(n1944), .B1(n2536), .B2(n1065), .ZN(
        mult_x_18_n736) );
  XNR2XD1BWP12T U2160 ( .A1(n3033), .A2(n2829), .ZN(n1118) );
  OAI22D1BWP12T U2161 ( .A1(n2541), .A2(n1066), .B1(n2539), .B2(n1118), .ZN(
        mult_x_18_n860) );
  OAI22D1BWP12T U2162 ( .A1(n2571), .A2(n1068), .B1(n2569), .B2(n1067), .ZN(
        mult_x_18_n981) );
  XNR2XD1BWP12T U2163 ( .A1(n2720), .A2(n2489), .ZN(n1109) );
  XNR2XD1BWP12T U2164 ( .A1(n2720), .A2(b[13]), .ZN(n1081) );
  OAI22D1BWP12T U2165 ( .A1(n2517), .A2(n1109), .B1(n2515), .B2(n1081), .ZN(
        mult_x_18_n833) );
  XNR2XD1BWP12T U2166 ( .A1(n2532), .A2(n3074), .ZN(n1108) );
  OAI22D1BWP12T U2167 ( .A1(n2535), .A2(n1069), .B1(n2533), .B2(n1108), .ZN(
        mult_x_18_n905) );
  XNR2XD1BWP12T U2168 ( .A1(n2542), .A2(n3033), .ZN(n1083) );
  OAI22D1BWP12T U2169 ( .A1(n2541), .A2(n1070), .B1(n2539), .B2(n1083), .ZN(
        mult_x_18_n863) );
  OAI22D1BWP12T U2170 ( .A1(n2525), .A2(n1072), .B1(n2523), .B2(n1071), .ZN(
        mult_x_18_n799) );
  OAI22D1BWP12T U2171 ( .A1(n2559), .A2(n1074), .B1(n2557), .B2(n1073), .ZN(
        mult_x_18_n934) );
  OAI22D1BWP12T U2172 ( .A1(n2525), .A2(n1076), .B1(n2523), .B2(n1075), .ZN(
        mult_x_18_n801) );
  OAI22D1BWP12T U2173 ( .A1(n2514), .A2(n1078), .B1(n1077), .B2(n2512), .ZN(
        mult_x_18_n955) );
  OAI22D1BWP12T U2174 ( .A1(n2493), .A2(n1080), .B1(n2491), .B2(n1079), .ZN(
        mult_x_18_n789) );
  XNR2XD1BWP12T U2175 ( .A1(n2720), .A2(n2522), .ZN(n1090) );
  OAI22D1BWP12T U2176 ( .A1(n2517), .A2(n1081), .B1(n2515), .B2(n1090), .ZN(
        mult_x_18_n832) );
  OAI22D1BWP12T U2177 ( .A1(n2541), .A2(n1083), .B1(n2539), .B2(n1082), .ZN(
        mult_x_18_n862) );
  OAI22D1BWP12T U2178 ( .A1(n2541), .A2(n1085), .B1(n2539), .B2(n1084), .ZN(
        mult_x_18_n855) );
  XNR2XD0BWP12T U2179 ( .A1(n3033), .A2(b[15]), .ZN(n1111) );
  OAI22D1BWP12T U2180 ( .A1(n2541), .A2(n1086), .B1(n2539), .B2(n1111), .ZN(
        mult_x_18_n852) );
  OAI22D1BWP12T U2181 ( .A1(n2487), .A2(n1088), .B1(n1087), .B2(n2486), .ZN(
        mult_x_18_n1005) );
  OAI22D1BWP12T U2182 ( .A1(n2517), .A2(n1090), .B1(n2515), .B2(n1089), .ZN(
        mult_x_18_n831) );
  OAI22D1BWP12T U2183 ( .A1(n2517), .A2(n1092), .B1(n2515), .B2(n1091), .ZN(
        mult_x_18_n838) );
  OAI22D1BWP12T U2184 ( .A1(n2517), .A2(n1094), .B1(n2515), .B2(n1093), .ZN(
        mult_x_18_n840) );
  OAI22D1BWP12T U2185 ( .A1(n2535), .A2(n1096), .B1(n2533), .B2(n1095), .ZN(
        mult_x_18_n908) );
  XNR2XD0BWP12T U2186 ( .A1(n3033), .A2(b[17]), .ZN(n1114) );
  OAI22D1BWP12T U2187 ( .A1(n2541), .A2(n1114), .B1(n2539), .B2(n1097), .ZN(
        mult_x_18_n849) );
  OAI22D1BWP12T U2188 ( .A1(n2514), .A2(n1099), .B1(n1098), .B2(n2512), .ZN(
        mult_x_18_n945) );
  OAI22D1BWP12T U2189 ( .A1(n2498), .A2(n1101), .B1(n1100), .B2(n2495), .ZN(
        mult_x_18_n872) );
  OAI22D1BWP12T U2190 ( .A1(n2559), .A2(n1103), .B1(n2557), .B2(n1102), .ZN(
        mult_x_18_n930) );
  XNR2D0BWP12T U2191 ( .A1(n2532), .A2(b[23]), .ZN(n2534) );
  OAI22D1BWP12T U2192 ( .A1(n2535), .A2(n1104), .B1(n2533), .B2(n2534), .ZN(
        mult_x_18_n892) );
  OAI22D1BWP12T U2193 ( .A1(n2493), .A2(n1106), .B1(n2491), .B2(n1105), .ZN(
        mult_x_18_n793) );
  OAI22D1BWP12T U2194 ( .A1(n2535), .A2(n1108), .B1(n2533), .B2(n1107), .ZN(
        mult_x_18_n904) );
  OAI22D1BWP12T U2195 ( .A1(n2517), .A2(n1110), .B1(n2515), .B2(n1109), .ZN(
        mult_x_18_n834) );
  XNR2XD0BWP12T U2196 ( .A1(n3033), .A2(b[16]), .ZN(n1115) );
  OAI22D1BWP12T U2197 ( .A1(n2541), .A2(n1111), .B1(n2539), .B2(n1115), .ZN(
        mult_x_18_n851) );
  OAI22D1BWP12T U2198 ( .A1(n2517), .A2(n1113), .B1(n2515), .B2(n1112), .ZN(
        mult_x_18_n842) );
  OAI22D1BWP12T U2199 ( .A1(n2541), .A2(n1115), .B1(n2539), .B2(n1114), .ZN(
        mult_x_18_n850) );
  OAI22D1BWP12T U2200 ( .A1(n2498), .A2(n1117), .B1(n1116), .B2(n2495), .ZN(
        mult_x_18_n870) );
  XNR2XD1BWP12T U2201 ( .A1(n3033), .A2(n2501), .ZN(n1123) );
  OAI22D1BWP12T U2202 ( .A1(n2541), .A2(n1118), .B1(n2539), .B2(n1123), .ZN(
        mult_x_18_n859) );
  OAI22D1BWP12T U2203 ( .A1(n2535), .A2(n1120), .B1(n2533), .B2(n1119), .ZN(
        mult_x_18_n896) );
  XNR2XD1BWP12T U2204 ( .A1(n2407), .A2(n2608), .ZN(n2545) );
  OAI22D1BWP12T U2205 ( .A1(n2546), .A2(n1121), .B1(n2545), .B2(n2543), .ZN(
        mult_x_18_n752) );
  OAI22D1BWP12T U2206 ( .A1(n2541), .A2(n1123), .B1(n2539), .B2(n1122), .ZN(
        mult_x_18_n858) );
  OAI22D1BWP12T U2207 ( .A1(n2514), .A2(n1125), .B1(n1124), .B2(n2512), .ZN(
        mult_x_18_n961) );
  OAI22D1BWP12T U2208 ( .A1(n2525), .A2(n1127), .B1(n2523), .B2(n1126), .ZN(
        mult_x_18_n805) );
  XNR2D0BWP12T U2209 ( .A1(n2560), .A2(n2522), .ZN(n1132) );
  OAI22D1BWP12T U2210 ( .A1(n2564), .A2(n1128), .B1(n1132), .B2(n2561), .ZN(
        mult_x_18_n813) );
  XNR2XD0BWP12T U2211 ( .A1(n2720), .A2(b[17]), .ZN(n2516) );
  OAI22D1BWP12T U2212 ( .A1(n2517), .A2(n1129), .B1(n2515), .B2(n2516), .ZN(
        mult_x_18_n829) );
  OAI22D1BWP12T U2213 ( .A1(n2538), .A2(n1131), .B1(n1130), .B2(n2536), .ZN(
        mult_x_18_n774) );
  XNR2D0BWP12T U2214 ( .A1(n2560), .A2(b[15]), .ZN(n2563) );
  OAI22D1BWP12T U2215 ( .A1(n2564), .A2(n1132), .B1(n2563), .B2(n2561), .ZN(
        mult_x_18_n812) );
  OAI22D1BWP12T U2216 ( .A1(n2521), .A2(n1134), .B1(n1133), .B2(n2519), .ZN(
        mult_x_18_n758) );
  TPOAI22D1BWP12T U2217 ( .A1(n2498), .A2(n1136), .B1(n1135), .B2(n2495), .ZN(
        mult_x_18_n888) );
  INVD1BWP12T U2218 ( .I(n1137), .ZN(n1583) );
  INVD1BWP12T U2219 ( .I(n1632), .ZN(n1197) );
  CKND0BWP12T U2220 ( .I(n1141), .ZN(n1143) );
  INVD1BWP12T U2221 ( .I(n1145), .ZN(n1149) );
  CKND2D0BWP12T U2222 ( .A1(n1149), .A2(n1148), .ZN(n1146) );
  XOR2XD0BWP12T U2223 ( .A1(n1147), .A2(n1146), .Z(n1722) );
  INVD1BWP12T U2224 ( .I(n1722), .ZN(n1190) );
  CKND2D1BWP12T U2225 ( .A1(n1847), .A2(n3119), .ZN(n1189) );
  INVD1BWP12T U2226 ( .I(n1151), .ZN(n1964) );
  AOI22D0BWP12T U2227 ( .A1(n2181), .A2(n1152), .B1(n2183), .B2(n1344), .ZN(
        n1155) );
  AOI22D0BWP12T U2228 ( .A1(n2187), .A2(n2335), .B1(n1153), .B2(n2337), .ZN(
        n1154) );
  ND2D1BWP12T U2229 ( .A1(n1155), .A2(n1154), .ZN(n1281) );
  ND2D1BWP12T U2230 ( .A1(n2187), .A2(n2311), .ZN(n2210) );
  OAI22D0BWP12T U2231 ( .A1(n1281), .A2(n2170), .B1(n2210), .B2(n2179), .ZN(
        n1157) );
  INVD0BWP12T U2232 ( .I(n2319), .ZN(n2174) );
  CKND0BWP12T U2233 ( .I(n2332), .ZN(n2144) );
  AOI22D0BWP12T U2234 ( .A1(n2187), .A2(n2174), .B1(n2183), .B2(n2144), .ZN(
        n1288) );
  AOI21D0BWP12T U2235 ( .A1(n1287), .A2(n1288), .B(n2211), .ZN(n1156) );
  NR2D1BWP12T U2236 ( .A1(n1157), .A2(n1156), .ZN(n2222) );
  ND2D1BWP12T U2237 ( .A1(n2311), .A2(n595), .ZN(n2314) );
  INVD0BWP12T U2238 ( .I(n2335), .ZN(n2142) );
  OAI22D0BWP12T U2239 ( .A1(n2142), .A2(n1329), .B1(n2143), .B2(n1333), .ZN(
        n1159) );
  OAI22D0BWP12T U2240 ( .A1(n2313), .A2(n2322), .B1(n2312), .B2(n1335), .ZN(
        n1158) );
  NR2D1BWP12T U2241 ( .A1(n1159), .A2(n1158), .ZN(n1294) );
  INVD1BWP12T U2242 ( .I(n2375), .ZN(n2388) );
  CKND0BWP12T U2243 ( .I(n2323), .ZN(n2171) );
  AOI22D0BWP12T U2244 ( .A1(n2331), .A2(n2171), .B1(n595), .B2(n2319), .ZN(
        n1161) );
  AOI22D0BWP12T U2245 ( .A1(n2336), .A2(n2332), .B1(n2333), .B2(n2334), .ZN(
        n1160) );
  ND2D1BWP12T U2246 ( .A1(n1161), .A2(n1160), .ZN(n1298) );
  MOAI22D0BWP12T U2247 ( .A1(n1294), .A2(n2082), .B1(n2388), .B2(n1298), .ZN(
        n1162) );
  ND2D1BWP12T U2248 ( .A1(n2452), .A2(n2343), .ZN(n2359) );
  RCAOI211D0BWP12T U2249 ( .A1(n2750), .A2(n2314), .B(n1162), .C(n2359), .ZN(
        n2368) );
  MUX2ND0BWP12T U2250 ( .I0(n2995), .I1(n2994), .S(b[17]), .ZN(n1163) );
  NR2D0BWP12T U2251 ( .A1(n1163), .A2(n2996), .ZN(n1166) );
  OAI21D0BWP12T U2252 ( .A1(n2560), .A2(n3066), .B(n3105), .ZN(n1164) );
  AOI22D0BWP12T U2253 ( .A1(n3070), .A2(n2275), .B1(n1164), .B2(b[17]), .ZN(
        n1165) );
  OAI211D0BWP12T U2254 ( .A1(n1166), .A2(n2275), .B(n2970), .C(n1165), .ZN(
        n1181) );
  OAI22D1BWP12T U2255 ( .A1(n2000), .A2(n2998), .B1(n1999), .B2(n2293), .ZN(
        n1168) );
  OAI22D1BWP12T U2256 ( .A1(n2002), .A2(n2636), .B1(n2001), .B2(n2965), .ZN(
        n1167) );
  NR2D1BWP12T U2257 ( .A1(n1168), .A2(n1167), .ZN(n2098) );
  OAI22D1BWP12T U2258 ( .A1(n2000), .A2(n2275), .B1(n2001), .B2(n2687), .ZN(
        n1170) );
  OAI22D1BWP12T U2259 ( .A1(n2002), .A2(n2659), .B1(n1999), .B2(n2928), .ZN(
        n1169) );
  NR2D1BWP12T U2260 ( .A1(n1170), .A2(n1169), .ZN(n2096) );
  OAI22D1BWP12T U2261 ( .A1(n2098), .A2(n2095), .B1(n2096), .B2(n2150), .ZN(
        n1184) );
  INR2XD0BWP12T U2262 ( .A1(n2502), .B1(n2000), .ZN(n1172) );
  NR2D1BWP12T U2263 ( .A1(n2001), .A2(n2290), .ZN(n1171) );
  NR2D1BWP12T U2264 ( .A1(n1172), .A2(n1171), .ZN(n1176) );
  NR2D1BWP12T U2265 ( .A1(n2002), .A2(n2291), .ZN(n1174) );
  NR2D1BWP12T U2266 ( .A1(n1999), .A2(n2287), .ZN(n1173) );
  NR2D1BWP12T U2267 ( .A1(n1174), .A2(n1173), .ZN(n1175) );
  ND2D1BWP12T U2268 ( .A1(n1176), .A2(n1175), .ZN(n1182) );
  INVD1BWP12T U2269 ( .I(n1182), .ZN(n2097) );
  AOI21D0BWP12T U2270 ( .A1(n2097), .A2(n2297), .B(n2349), .ZN(n1179) );
  OAI22D1BWP12T U2271 ( .A1(n2000), .A2(n2607), .B1(n2001), .B2(n2289), .ZN(
        n2008) );
  NR2D1BWP12T U2272 ( .A1(n2002), .A2(n2305), .ZN(n1177) );
  NR2D2BWP12T U2273 ( .A1(n2008), .A2(n1177), .ZN(n2613) );
  INVD0BWP12T U2274 ( .I(n2613), .ZN(n1178) );
  OAI22D1BWP12T U2275 ( .A1(n1184), .A2(n1179), .B1(n2110), .B2(n1178), .ZN(
        n2453) );
  TPNR2D0BWP12T U2276 ( .A1(n3004), .A2(n2453), .ZN(n1180) );
  AOI211XD0BWP12T U2277 ( .A1(n2368), .A2(n3040), .B(n1181), .C(n1180), .ZN(
        n1186) );
  MUX2NXD0BWP12T U2278 ( .I0(n1182), .I1(n2008), .S(n2405), .ZN(n1183) );
  OAI21D0BWP12T U2279 ( .A1(n2305), .A2(n2322), .B(n1183), .ZN(n1992) );
  AOI21D1BWP12T U2280 ( .A1(n1992), .A2(n2407), .B(n1184), .ZN(n2027) );
  INVD1BWP12T U2281 ( .I(n2027), .ZN(n2078) );
  CKND2D1BWP12T U2282 ( .A1(n2078), .A2(n1258), .ZN(n1185) );
  OAI211D1BWP12T U2283 ( .A1(n2222), .A2(n3012), .B(n1186), .C(n1185), .ZN(
        n1187) );
  AOI21D1BWP12T U2284 ( .A1(n1953), .A2(n3115), .B(n1187), .ZN(n1188) );
  OAI211D1BWP12T U2285 ( .A1(n1190), .A2(n2943), .B(n1189), .C(n1188), .ZN(
        n1191) );
  AOI21D1BWP12T U2286 ( .A1(n3095), .A2(n1546), .B(n1191), .ZN(n1196) );
  ND2D1BWP12T U2287 ( .A1(n1819), .A2(n314), .ZN(n1195) );
  OAI211D2BWP12T U2288 ( .A1(n2951), .A2(n1197), .B(n1196), .C(n1195), .ZN(
        result[17]) );
  TPNR2D1BWP12T U2289 ( .A1(mult_x_18_n447), .A2(mult_x_18_n426), .ZN(n1651)
         );
  NR2D1BWP12T U2290 ( .A1(n1651), .A2(n1646), .ZN(n1199) );
  TPND2D0BWP12T U2291 ( .A1(n1199), .A2(n1642), .ZN(n1201) );
  ND2D1BWP12T U2292 ( .A1(mult_x_18_n447), .A2(mult_x_18_n426), .ZN(n1652) );
  TPOAI21D0BWP12T U2293 ( .A1(n1651), .A2(n1645), .B(n1652), .ZN(n1198) );
  TPAOI21D0BWP12T U2294 ( .A1(n1199), .A2(n1644), .B(n1198), .ZN(n1200) );
  OAI21D1BWP12T U2295 ( .A1(n1202), .A2(n1201), .B(n1200), .ZN(n1320) );
  FA1D1BWP12T U2296 ( .A(n1205), .B(a[28]), .CI(n1203), .CO(n1476), .S(n1554)
         );
  CKND0BWP12T U2297 ( .I(b[30]), .ZN(n1322) );
  CKND1BWP12T U2298 ( .I(b[29]), .ZN(n1734) );
  FA1D0BWP12T U2299 ( .A(n1205), .B(a[28]), .CI(n1204), .CO(n1733), .S(n1826)
         );
  FA1D2BWP12T U2300 ( .A(b[28]), .B(a[28]), .CI(n1206), .CO(n1928), .S(n1931)
         );
  CKND0BWP12T U2301 ( .I(n1207), .ZN(n1210) );
  OAI22D1BWP12T U2302 ( .A1(n1210), .A2(n1209), .B1(n1350), .B2(n1208), .ZN(
        n1213) );
  NR2D1BWP12T U2303 ( .A1(n2175), .A2(n1211), .ZN(n1212) );
  AOI211D1BWP12T U2304 ( .A1(n1227), .A2(n2187), .B(n1213), .C(n1212), .ZN(
        n2800) );
  CKND0BWP12T U2305 ( .I(n2800), .ZN(n1223) );
  INVD0BWP12T U2306 ( .I(n1241), .ZN(n1216) );
  OAI22D0BWP12T U2307 ( .A1(n1350), .A2(n1239), .B1(n1351), .B2(n1240), .ZN(
        n1215) );
  TPNR2D0BWP12T U2308 ( .A1(n2175), .A2(n1238), .ZN(n1214) );
  AOI211D1BWP12T U2309 ( .A1(n1216), .A2(n2187), .B(n1215), .C(n1214), .ZN(
        n2168) );
  OAI22D0BWP12T U2310 ( .A1(n1351), .A2(n1247), .B1(n1350), .B2(n1246), .ZN(
        n1218) );
  NR2D0BWP12T U2311 ( .A1(n2175), .A2(n1244), .ZN(n1217) );
  AOI211D1BWP12T U2312 ( .A1(n1219), .A2(n2187), .B(n1218), .C(n1217), .ZN(
        n2169) );
  OAI22D0BWP12T U2313 ( .A1(n1350), .A2(n1234), .B1(n1351), .B2(n1233), .ZN(
        n1221) );
  NR2D0BWP12T U2314 ( .A1(n2175), .A2(n1232), .ZN(n1220) );
  AOI211D0BWP12T U2315 ( .A1(n2187), .A2(n2608), .B(n1221), .C(n1220), .ZN(
        n1222) );
  OAI222D0BWP12T U2316 ( .A1(n2170), .A2(n2168), .B1(n2179), .B2(n2169), .C1(
        n2211), .C2(n1222), .ZN(n2194) );
  AOI21D1BWP12T U2317 ( .A1(n2178), .A2(n1223), .B(n2194), .ZN(n1261) );
  HA1D1BWP12T U2318 ( .A(n2287), .B(n1224), .CO(n1942), .S(n1983) );
  ND2D1BWP12T U2319 ( .A1(n1988), .A2(n3115), .ZN(n1260) );
  MUX2NXD0BWP12T U2320 ( .I0(n1225), .I1(n2305), .S(n2405), .ZN(n2030) );
  TPAOI21D0BWP12T U2321 ( .A1(n2030), .A2(n2349), .B(n2093), .ZN(n2031) );
  INVD1BWP12T U2322 ( .I(n2031), .ZN(n1447) );
  OAI22D0BWP12T U2323 ( .A1(n1227), .A2(n1329), .B1(n1226), .B2(n2322), .ZN(
        n1230) );
  NR2D0BWP12T U2324 ( .A1(n1228), .A2(n1333), .ZN(n1229) );
  AOI211D1BWP12T U2325 ( .A1(n1231), .A2(n2405), .B(n1230), .C(n1229), .ZN(
        n2808) );
  AOI22D0BWP12T U2326 ( .A1(n2336), .A2(n1233), .B1(n1232), .B2(n2334), .ZN(
        n1236) );
  CKND2D0BWP12T U2327 ( .A1(n1234), .A2(n2331), .ZN(n1235) );
  OAI211D0BWP12T U2328 ( .A1(n2608), .A2(n1334), .B(n1236), .C(n1235), .ZN(
        n1237) );
  CKND0BWP12T U2329 ( .I(n2157), .ZN(n1339) );
  NR2D0BWP12T U2330 ( .A1(n1339), .A2(a[30]), .ZN(n1941) );
  AOI211D0BWP12T U2331 ( .A1(n1237), .A2(n2388), .B(n1941), .C(n2437), .ZN(
        n1251) );
  AOI22D0BWP12T U2332 ( .A1(n2331), .A2(n1239), .B1(n1238), .B2(n2334), .ZN(
        n1243) );
  AOI22D0BWP12T U2333 ( .A1(n595), .A2(n1241), .B1(n1240), .B2(n2336), .ZN(
        n1242) );
  ND2D1BWP12T U2334 ( .A1(n1243), .A2(n1242), .ZN(n2345) );
  AOI22D0BWP12T U2335 ( .A1(n595), .A2(n1245), .B1(n1244), .B2(n2334), .ZN(
        n1249) );
  AOI22D0BWP12T U2336 ( .A1(n2336), .A2(n1247), .B1(n1246), .B2(n2331), .ZN(
        n1248) );
  ND2D1BWP12T U2337 ( .A1(n1249), .A2(n1248), .ZN(n2348) );
  AOI22D0BWP12T U2338 ( .A1(n2381), .A2(n2345), .B1(n2348), .B2(n2340), .ZN(
        n1250) );
  OA211D0BWP12T U2339 ( .A1(n2808), .A2(n2343), .B(n1251), .C(n1250), .Z(n2356) );
  MOAI22D0BWP12T U2340 ( .A1(n2204), .A2(n2612), .B1(n2356), .B2(n3040), .ZN(
        n1257) );
  MUX2ND0BWP12T U2341 ( .I0(n2995), .I1(n2994), .S(b[30]), .ZN(n1252) );
  NR2D0BWP12T U2342 ( .A1(n1252), .A2(n2996), .ZN(n1255) );
  OAI21D0BWP12T U2343 ( .A1(a[30]), .A2(n3066), .B(n3105), .ZN(n1253) );
  AOI22D0BWP12T U2344 ( .A1(n3070), .A2(n2289), .B1(n1253), .B2(b[30]), .ZN(
        n1254) );
  OAI211D1BWP12T U2345 ( .A1(n1255), .A2(n2289), .B(n2970), .C(n1254), .ZN(
        n1256) );
  AOI211XD0BWP12T U2346 ( .A1(n1258), .A2(n1447), .B(n1257), .C(n1256), .ZN(
        n1259) );
  OAI211D1BWP12T U2347 ( .A1(n1261), .A2(n3012), .B(n1260), .C(n1259), .ZN(
        n1262) );
  AOI21D1BWP12T U2348 ( .A1(n2475), .A2(n3119), .B(n1262), .ZN(n1265) );
  FA1D0BWP12T U2349 ( .A(b[28]), .B(a[28]), .CI(n1263), .CO(n1661), .S(n1731)
         );
  OAI211D2BWP12T U2350 ( .A1(n3020), .A2(n1266), .B(n1265), .C(n1264), .ZN(
        n1267) );
  IOA21D2BWP12T U2351 ( .A1(n1657), .A2(n3126), .B(n1268), .ZN(result[30]) );
  INVD1BWP12T U2352 ( .I(n1272), .ZN(n1274) );
  AN2XD1BWP12T U2353 ( .A1(n1274), .A2(n1273), .Z(n1275) );
  CKXOR2D1BWP12T U2354 ( .A1(n1276), .A2(n1275), .Z(n1641) );
  FA1D1BWP12T U2355 ( .A(n1279), .B(n2502), .CI(n1277), .CO(n469), .S(n1550)
         );
  FA1D0BWP12T U2356 ( .A(n1279), .B(n2502), .CI(n1278), .CO(n470), .S(n1823)
         );
  INVD1BWP12T U2357 ( .I(n1823), .ZN(n1317) );
  FA1D2BWP12T U2358 ( .A(n2502), .B(b[25]), .CI(n1280), .CO(n472), .S(n1927)
         );
  MUX2D1BWP12T U2359 ( .I0(n2210), .I1(n1281), .S(n2221), .Z(n2154) );
  CKND2D0BWP12T U2360 ( .A1(n2154), .A2(n2217), .ZN(n1291) );
  CKND0BWP12T U2361 ( .I(n2327), .ZN(n2182) );
  OAI22D0BWP12T U2362 ( .A1(n1350), .A2(n2182), .B1(n1351), .B2(n1347), .ZN(
        n1284) );
  INVD0BWP12T U2363 ( .I(n2326), .ZN(n2180) );
  NR2D0BWP12T U2364 ( .A1(n1282), .A2(n2180), .ZN(n1283) );
  AOI211D0BWP12T U2365 ( .A1(n2181), .A2(n2317), .B(n1284), .C(n1283), .ZN(
        n1285) );
  OAI21D0BWP12T U2366 ( .A1(n1285), .A2(n2211), .B(n1339), .ZN(n1286) );
  AOI31D0BWP12T U2367 ( .A1(n2904), .A2(n1288), .A3(n1287), .B(n1286), .ZN(
        n1290) );
  MUX2ND0BWP12T U2368 ( .I0(n2613), .I1(n2097), .S(n2297), .ZN(n1289) );
  AOI22D1BWP12T U2369 ( .A1(n1291), .A2(n1290), .B1(n2388), .B2(n1289), .ZN(
        n2237) );
  HA1D0BWP12T U2370 ( .A(n1293), .B(n1292), .CO(n489), .S(n1980) );
  CKND2D1BWP12T U2371 ( .A1(n1980), .A2(n3115), .ZN(n1312) );
  INVD1BWP12T U2372 ( .I(n2314), .ZN(n3093) );
  MUX2NXD0BWP12T U2373 ( .I0(n1294), .I1(n3093), .S(n2407), .ZN(n2861) );
  CKND0BWP12T U2374 ( .I(n2861), .ZN(n1300) );
  AOI22D0BWP12T U2375 ( .A1(n595), .A2(n2326), .B1(n2327), .B2(n2331), .ZN(
        n1296) );
  AOI22D0BWP12T U2376 ( .A1(n2318), .A2(n2336), .B1(n2317), .B2(n2334), .ZN(
        n1295) );
  AOI21D0BWP12T U2377 ( .A1(n1296), .A2(n1295), .B(n2375), .ZN(n1297) );
  AOI211XD0BWP12T U2378 ( .A1(n1298), .A2(n2381), .B(n1297), .C(n2437), .ZN(
        n1299) );
  TPOAI21D0BWP12T U2379 ( .A1(n1300), .A2(n2431), .B(n1299), .ZN(n2369) );
  AOI21D0BWP12T U2380 ( .A1(n1992), .A2(n2349), .B(n1301), .ZN(n2010) );
  OAI21D0BWP12T U2381 ( .A1(n2502), .A2(n3066), .B(n3105), .ZN(n1305) );
  MUX2ND0BWP12T U2382 ( .I0(n2995), .I1(n2994), .S(b[25]), .ZN(n1302) );
  NR2D0BWP12T U2383 ( .A1(n1302), .A2(n2996), .ZN(n1303) );
  MUX2ND0BWP12T U2384 ( .I0(n1303), .I1(n3109), .S(n2292), .ZN(n1304) );
  AOI21D0BWP12T U2385 ( .A1(b[25]), .A2(n1305), .B(n1304), .ZN(n1308) );
  OAI22D1BWP12T U2386 ( .A1(n2613), .A2(n2095), .B1(n2097), .B2(n2150), .ZN(
        n2454) );
  TPND2D0BWP12T U2387 ( .A1(n1306), .A2(n2454), .ZN(n1307) );
  OAI211D1BWP12T U2388 ( .A1(n1309), .A2(n2010), .B(n1308), .C(n1307), .ZN(
        n1310) );
  IAO21D1BWP12T U2389 ( .A1(n2369), .A2(n2903), .B(n1310), .ZN(n1311) );
  OAI211D1BWP12T U2390 ( .A1(n2237), .A2(n3012), .B(n1312), .C(n1311), .ZN(
        n1313) );
  AOI21D1BWP12T U2391 ( .A1(n1927), .A2(n3119), .B(n1313), .ZN(n1316) );
  FA1D2BWP12T U2392 ( .A(n2502), .B(b[25]), .CI(n1314), .CO(n512), .S(n1729)
         );
  CKND2D1BWP12T U2393 ( .A1(n1729), .A2(n3098), .ZN(n1315) );
  OAI211D1BWP12T U2394 ( .A1(n3020), .A2(n1317), .B(n1316), .C(n1315), .ZN(
        n1318) );
  AOI21D1BWP12T U2395 ( .A1(n3095), .A2(n1550), .B(n1318), .ZN(n1319) );
  IOA21D2BWP12T U2396 ( .A1(n1641), .A2(n3126), .B(n1319), .ZN(result[25]) );
  FA1D1BWP12T U2397 ( .A(mult_x_18_n425), .B(mult_x_18_n405), .CI(n1320), .CO(
        n2484), .S(n1657) );
  INVD1BWP12T U2398 ( .I(n2587), .ZN(n1659) );
  FA1D2BWP12T U2399 ( .A(n1322), .B(a[30]), .CI(n1321), .CO(n2590), .S(n1831)
         );
  XNR2D1BWP12T U2400 ( .A1(n2595), .A2(n2956), .ZN(n2596) );
  INVD1BWP12T U2401 ( .I(n2596), .ZN(n1369) );
  INVD1BWP12T U2402 ( .I(b[31]), .ZN(n2953) );
  AOI22D0BWP12T U2403 ( .A1(n595), .A2(n2327), .B1(n2317), .B2(n2331), .ZN(
        n1326) );
  AOI22D0BWP12T U2404 ( .A1(n2336), .A2(n2319), .B1(n2318), .B2(n2334), .ZN(
        n1325) );
  ND2D1BWP12T U2405 ( .A1(n1326), .A2(n1325), .ZN(n2389) );
  OAI22D0BWP12T U2406 ( .A1(n2311), .A2(n2322), .B1(n2312), .B2(n1333), .ZN(
        n1328) );
  OAI22D0BWP12T U2407 ( .A1(n2313), .A2(n1335), .B1(n2143), .B2(n1329), .ZN(
        n1327) );
  NR2D1BWP12T U2408 ( .A1(n1328), .A2(n1327), .ZN(n2838) );
  INVD0BWP12T U2409 ( .I(n2333), .ZN(n2145) );
  OAI22D0BWP12T U2410 ( .A1(n2323), .A2(n1329), .B1(n2145), .B2(n1333), .ZN(
        n1331) );
  OAI22D0BWP12T U2411 ( .A1(n2144), .A2(n1335), .B1(n2142), .B2(n2322), .ZN(
        n1330) );
  NR2D1BWP12T U2412 ( .A1(n1331), .A2(n1330), .ZN(n2387) );
  OAI22D0BWP12T U2413 ( .A1(n2838), .A2(n2343), .B1(n2387), .B2(n1332), .ZN(
        n1341) );
  MUX2NXD0BWP12T U2414 ( .I0(n2608), .I1(a[28]), .S(n1383), .ZN(n2325) );
  CKND0BWP12T U2415 ( .I(n2325), .ZN(n2186) );
  OAI22D0BWP12T U2416 ( .A1(n2180), .A2(n2322), .B1(n2186), .B2(n1333), .ZN(
        n1337) );
  OAI22D0BWP12T U2417 ( .A1(n2184), .A2(n1335), .B1(n1334), .B2(a[30]), .ZN(
        n1336) );
  OAI21D0BWP12T U2418 ( .A1(n1337), .A2(n1336), .B(n2388), .ZN(n1338) );
  OAI211D1BWP12T U2419 ( .A1(n2956), .A2(n1339), .B(n1338), .C(n2452), .ZN(
        n1340) );
  AOI211D1BWP12T U2420 ( .A1(n2381), .A2(n2389), .B(n1341), .C(n1340), .ZN(
        n2355) );
  AOI22D0BWP12T U2421 ( .A1(n2312), .A2(n2185), .B1(n2183), .B2(n2311), .ZN(
        n1343) );
  CKND2D1BWP12T U2422 ( .A1(n2187), .A2(n2143), .ZN(n1342) );
  OAI211D1BWP12T U2423 ( .A1(n2175), .A2(n1344), .B(n1343), .C(n1342), .ZN(
        n2234) );
  AOI22D0BWP12T U2424 ( .A1(n2185), .A2(n2317), .B1(n2183), .B2(n2319), .ZN(
        n1346) );
  TPND2D0BWP12T U2425 ( .A1(n2187), .A2(n2327), .ZN(n1345) );
  OAI211D0BWP12T U2426 ( .A1(n1347), .A2(n2175), .B(n1346), .C(n1345), .ZN(
        n2231) );
  NR2D0BWP12T U2427 ( .A1(n2175), .A2(n2332), .ZN(n1349) );
  OAI22D0BWP12T U2428 ( .A1(n1351), .A2(n2335), .B1(n1350), .B2(n2333), .ZN(
        n1348) );
  AOI211D1BWP12T U2429 ( .A1(n2323), .A2(n2187), .B(n1349), .C(n1348), .ZN(
        n2230) );
  NR2D0BWP12T U2430 ( .A1(n2175), .A2(n2324), .ZN(n1353) );
  OAI22D0BWP12T U2431 ( .A1(n1351), .A2(n2326), .B1(n1350), .B2(n2325), .ZN(
        n1352) );
  AOI211D0BWP12T U2432 ( .A1(n2187), .A2(a[30]), .B(n1353), .C(n1352), .ZN(
        n1354) );
  OAI222D1BWP12T U2433 ( .A1(n2170), .A2(n2231), .B1(n2179), .B2(n2230), .C1(
        n2211), .C2(n1354), .ZN(n2163) );
  AOI21D1BWP12T U2434 ( .A1(n2178), .A2(n2234), .B(n2163), .ZN(n1355) );
  NR2D1BWP12T U2435 ( .A1(n1355), .A2(n3012), .ZN(n1366) );
  NR2D0BWP12T U2436 ( .A1(n2305), .A2(n2407), .ZN(n1356) );
  TPND2D0BWP12T U2437 ( .A1(n2070), .A2(n1356), .ZN(n2432) );
  XNR2XD1BWP12T U2438 ( .A1(b[31]), .A2(n2956), .ZN(n2593) );
  INVD1BWP12T U2439 ( .I(n2593), .ZN(n1357) );
  AOI22D0BWP12T U2440 ( .A1(n1357), .A2(n3107), .B1(b[31]), .B2(n2996), .ZN(
        n1364) );
  NR2D0BWP12T U2441 ( .A1(b[31]), .A2(op[2]), .ZN(n1361) );
  CKND0BWP12T U2442 ( .I(n1358), .ZN(n1360) );
  CKND0BWP12T U2443 ( .I(n2304), .ZN(n1359) );
  OAI22D0BWP12T U2444 ( .A1(n1361), .A2(n1360), .B1(b[31]), .B2(n1359), .ZN(
        n1362) );
  MUX2ND0BWP12T U2445 ( .I0(n3070), .I1(n1362), .S(n2956), .ZN(n1363) );
  OAI211D1BWP12T U2446 ( .A1(n2432), .A2(n3004), .B(n1364), .C(n1363), .ZN(
        n1365) );
  RCAOI211D0BWP12T U2447 ( .A1(n3040), .A2(n2355), .B(n1366), .C(n1365), .ZN(
        n1367) );
  OAI211D1BWP12T U2448 ( .A1(n1369), .A2(n2980), .B(n1368), .C(n1367), .ZN(
        n1373) );
  FA1D2BWP12T U2449 ( .A(b[30]), .B(a[30]), .CI(n1370), .CO(n2955), .S(n1732)
         );
  CKND2BWP12T U2450 ( .I(n1371), .ZN(n2478) );
  AOI211XD1BWP12T U2451 ( .A1(n1832), .A2(n314), .B(n1373), .C(n1372), .ZN(
        n1376) );
  CKND2D2BWP12T U2452 ( .A1(n2483), .A2(n3095), .ZN(n1375) );
  OAI211D4BWP12T U2453 ( .A1(n2951), .A2(n1659), .B(n1376), .C(n1375), .ZN(
        result[31]) );
  CKBD1BWP12T U2454 ( .I(result[31]), .Z(n) );
  OAI22D0BWP12T U2455 ( .A1(n2000), .A2(n2749), .B1(n1999), .B2(n2831), .ZN(
        n1378) );
  OAI22D0BWP12T U2456 ( .A1(n2002), .A2(n2802), .B1(n2001), .B2(n2768), .ZN(
        n1377) );
  NR2D1BWP12T U2457 ( .A1(n1378), .A2(n1377), .ZN(n2014) );
  INR2D1BWP12T U2458 ( .A1(n1379), .B1(n2150), .ZN(n1388) );
  OAI22D0BWP12T U2459 ( .A1(n1414), .A2(n2133), .B1(n1413), .B2(n2095), .ZN(
        n1381) );
  OAI22D0BWP12T U2460 ( .A1(n2205), .A2(n2110), .B1(n2019), .B2(n2150), .ZN(
        n1380) );
  NR2D1BWP12T U2461 ( .A1(n1381), .A2(n1380), .ZN(n2897) );
  NR2D1BWP12T U2462 ( .A1(n2897), .A2(n2431), .ZN(n2214) );
  AOI22D1BWP12T U2463 ( .A1(n2213), .A2(n2459), .B1(n2452), .B2(n2214), .ZN(
        n2103) );
  XNR2D0BWP12T U2464 ( .A1(n1391), .A2(n2262), .ZN(n1792) );
  INR2D0BWP12T U2465 ( .A1(n1382), .B1(n2486), .ZN(n1614) );
  INVD1BWP12T U2466 ( .I(n1384), .ZN(n1386) );
  INVD1BWP12T U2467 ( .I(n1388), .ZN(n2310) );
  INVD1BWP12T U2468 ( .I(n2103), .ZN(n2438) );
  INVD1BWP12T U2469 ( .I(n1392), .ZN(n1590) );
  AOI21D1BWP12T U2470 ( .A1(n1590), .A2(n1589), .B(n1393), .ZN(n1397) );
  ND2D1BWP12T U2471 ( .A1(n1395), .A2(n1394), .ZN(n1396) );
  XOR2XD1BWP12T U2472 ( .A1(n1397), .A2(n1396), .Z(n1622) );
  INVD1BWP12T U2473 ( .I(n1501), .ZN(n1534) );
  INVD1BWP12T U2474 ( .I(n1500), .ZN(n1537) );
  INVD1BWP12T U2475 ( .I(n1401), .ZN(n1803) );
  NR2XD0BWP12T U2476 ( .A1(n1803), .A2(n1804), .ZN(n1806) );
  INVD1BWP12T U2477 ( .I(n1402), .ZN(n1802) );
  OAI21D1BWP12T U2478 ( .A1(n1802), .A2(n1804), .B(n1805), .ZN(n1807) );
  INVD1BWP12T U2479 ( .I(n1679), .ZN(n1683) );
  INVD1BWP12T U2480 ( .I(n1406), .ZN(n1681) );
  CKND2D1BWP12T U2481 ( .A1(n1683), .A2(n1681), .ZN(n1409) );
  INVD0BWP12T U2482 ( .I(n1678), .ZN(n1686) );
  INVD1BWP12T U2483 ( .I(n1680), .ZN(n1407) );
  AOI21D1BWP12T U2484 ( .A1(n1686), .A2(n1681), .B(n1407), .ZN(n1408) );
  OAI21D1BWP12T U2485 ( .A1(n1700), .A2(n1409), .B(n1408), .ZN(n1412) );
  CKND2D1BWP12T U2486 ( .A1(n1902), .A2(n1423), .ZN(n1411) );
  XNR2XD1BWP12T U2487 ( .A1(n1412), .A2(n1411), .ZN(n1682) );
  INVD0BWP12T U2488 ( .I(n2015), .ZN(n1415) );
  TPAOI21D0BWP12T U2489 ( .A1(n1415), .A2(n2089), .B(n2750), .ZN(n1416) );
  TPOAI21D0BWP12T U2490 ( .A1(n2019), .A2(n2095), .B(n1416), .ZN(n1417) );
  AOI21D1BWP12T U2491 ( .A1(n2407), .A2(n2013), .B(n1417), .ZN(n1419) );
  AOI22D0BWP12T U2492 ( .A1(n3098), .A2(n1682), .B1(n2152), .B2(n3091), .ZN(
        n1418) );
  IOA21D1BWP12T U2493 ( .A1(n1758), .A2(n314), .B(n1418), .ZN(n1435) );
  AOI211D0BWP12T U2494 ( .A1(n2750), .A2(n1420), .B(n1419), .C(n2437), .ZN(
        n1421) );
  NR2XD0BWP12T U2495 ( .A1(n1421), .A2(n2101), .ZN(n2024) );
  CKND2D1BWP12T U2496 ( .A1(n1970), .A2(n1960), .ZN(n1422) );
  XOR2XD1BWP12T U2497 ( .A1(n1422), .A2(n2416), .Z(n1969) );
  AOI22D1BWP12T U2498 ( .A1(n3115), .A2(n1969), .B1(n1912), .B2(n3119), .ZN(
        n1433) );
  INVD1BWP12T U2499 ( .I(n2361), .ZN(n1424) );
  MUX2ND0BWP12T U2500 ( .I0(n1424), .I1(n2747), .S(n2407), .ZN(n1425) );
  NR2D1BWP12T U2501 ( .A1(n1425), .A2(n2448), .ZN(n2385) );
  TPNR2D0BWP12T U2502 ( .A1(n2446), .A2(n3038), .ZN(n1431) );
  OAI21D0BWP12T U2503 ( .A1(n2416), .A2(n3066), .B(n3105), .ZN(n1429) );
  MUX2NXD0BWP12T U2504 ( .I0(n3104), .I1(n3103), .S(n2489), .ZN(n1426) );
  ND2XD0BWP12T U2505 ( .A1(n1426), .A2(n3105), .ZN(n1427) );
  MUX2ND0BWP12T U2506 ( .I0(n1427), .I1(n3070), .S(n2281), .ZN(n1428) );
  IOA21D1BWP12T U2507 ( .A1(n2489), .A2(n1429), .B(n1428), .ZN(n1430) );
  AOI211XD0BWP12T U2508 ( .A1(n3040), .A2(n2385), .B(n1431), .C(n1430), .ZN(
        n1432) );
  OAI211D1BWP12T U2509 ( .A1(n2024), .A2(n3044), .B(n1433), .C(n1432), .ZN(
        n1434) );
  AOI211D1BWP12T U2510 ( .A1(n3095), .A2(n1503), .B(n1435), .C(n1434), .ZN(
        n1436) );
  IOA21D1BWP12T U2511 ( .A1(n1622), .A2(n3126), .B(n1436), .ZN(result[12]) );
  ND2D1BWP12T U2512 ( .A1(n1625), .A2(n1438), .ZN(n1439) );
  XNR2D1BWP12T U2513 ( .A1(n1626), .A2(n1439), .ZN(n1634) );
  ND2XD0BWP12T U2514 ( .A1(n1441), .A2(n1440), .ZN(n1442) );
  XNR2D1BWP12T U2515 ( .A1(n1443), .A2(n1442), .ZN(n1759) );
  MUX2XD0BWP12T U2516 ( .I0(n2028), .I1(n2029), .S(n2405), .Z(n1444) );
  AOI21D0BWP12T U2517 ( .A1(n1444), .A2(n2431), .B(n2388), .ZN(n1446) );
  OAI22D0BWP12T U2518 ( .A1(n2113), .A2(n2150), .B1(n2111), .B2(n2095), .ZN(
        n1445) );
  NR2D1BWP12T U2519 ( .A1(n1446), .A2(n1445), .ZN(n1450) );
  NR2D0BWP12T U2520 ( .A1(n1447), .A2(n2431), .ZN(n1448) );
  TPOAI31D0BWP12T U2521 ( .A1(n2090), .A2(n1450), .A3(n1448), .B(n2114), .ZN(
        n2116) );
  MUX2NXD0BWP12T U2522 ( .I0(n2800), .I1(n2169), .S(n2221), .ZN(n1451) );
  AOI21D0BWP12T U2523 ( .A1(n2201), .A2(n2089), .B(n2431), .ZN(n1449) );
  NR2D1BWP12T U2524 ( .A1(n1450), .A2(n1449), .ZN(n2434) );
  TPAOI21D0BWP12T U2525 ( .A1(n2868), .A2(n1451), .B(n2434), .ZN(n2138) );
  CKND2D1BWP12T U2526 ( .A1(n1453), .A2(n1452), .ZN(n1454) );
  XNR2XD1BWP12T U2527 ( .A1(n1455), .A2(n1454), .ZN(n1541) );
  INVD0BWP12T U2528 ( .I(n2808), .ZN(n1457) );
  MUX2ND0BWP12T U2529 ( .I0(n2348), .I1(n1457), .S(n2407), .ZN(n1458) );
  CKND2D1BWP12T U2530 ( .A1(n1458), .A2(n2459), .ZN(n2392) );
  CKND2D1BWP12T U2531 ( .A1(n1460), .A2(n1459), .ZN(n1461) );
  XNR2XD2BWP12T U2532 ( .A1(n1462), .A2(n1461), .ZN(n1721) );
  CKND2D0BWP12T U2533 ( .A1(n1721), .A2(n3098), .ZN(n1471) );
  XNR2XD0BWP12T U2534 ( .A1(n1972), .A2(a[14]), .ZN(n1974) );
  MUX2ND0BWP12T U2535 ( .I0(n2995), .I1(n2994), .S(n2522), .ZN(n1465) );
  NR2D0BWP12T U2536 ( .A1(n1465), .A2(n2996), .ZN(n1466) );
  MUX2NXD0BWP12T U2537 ( .I0(n1466), .I1(n3109), .S(n2280), .ZN(n1469) );
  NR2D0BWP12T U2538 ( .A1(a[14]), .A2(n3066), .ZN(n1467) );
  OA21D0BWP12T U2539 ( .A1(n1467), .A2(n2996), .B(n2522), .Z(n1468) );
  AOI211D1BWP12T U2540 ( .A1(n1974), .A2(n3115), .B(n1469), .C(n1468), .ZN(
        n1470) );
  OAI211D1BWP12T U2541 ( .A1(n2903), .A2(n2392), .B(n1471), .C(n1470), .ZN(
        n1472) );
  AOI211XD0BWP12T U2542 ( .A1(n3130), .A2(n2116), .B(n1473), .C(n1472), .ZN(
        n1474) );
  IOA21D1BWP12T U2543 ( .A1(n314), .A2(n1759), .B(n1474), .ZN(n1475) );
  AO21D2BWP12T U2544 ( .A1(n1634), .A2(n3126), .B(n1475), .Z(result[14]) );
  FA1D1BWP12T U2545 ( .A(n2608), .B(n1734), .CI(n1476), .CO(n1374), .S(n2624)
         );
  FA1D0BWP12T U2546 ( .A(n1736), .B(n2633), .CI(n1477), .CO(n739), .S(n2650)
         );
  FA1D0BWP12T U2547 ( .A(n1821), .B(n2963), .CI(n1478), .CO(n1477), .S(n2988)
         );
  CKND2D0BWP12T U2548 ( .A1(n1480), .A2(n1479), .ZN(n1481) );
  XNR2XD1BWP12T U2549 ( .A1(n1482), .A2(n1481), .ZN(n2946) );
  CKND0BWP12T U2550 ( .I(n1483), .ZN(n1485) );
  CKND2D0BWP12T U2551 ( .A1(n1485), .A2(n1484), .ZN(n1486) );
  XOR2XD1BWP12T U2552 ( .A1(n1487), .A2(n1486), .Z(n2677) );
  CKND2D0BWP12T U2553 ( .A1(n1489), .A2(n1488), .ZN(n1490) );
  XNR2XD1BWP12T U2554 ( .A1(n1491), .A2(n1490), .ZN(n2707) );
  INVD1BWP12T U2555 ( .I(n1492), .ZN(n1495) );
  INVD0BWP12T U2556 ( .I(n1497), .ZN(n1499) );
  CKND0BWP12T U2557 ( .I(n1504), .ZN(n1506) );
  ND2XD0BWP12T U2558 ( .A1(n1506), .A2(n1505), .ZN(n1507) );
  XOR2XD1BWP12T U2559 ( .A1(n1508), .A2(n1507), .Z(n2734) );
  INVD0BWP12T U2560 ( .I(n1514), .ZN(n1510) );
  INVD0BWP12T U2561 ( .I(n1515), .ZN(n1517) );
  INVD1BWP12T U2562 ( .I(n1520), .ZN(n1522) );
  CKND2D1BWP12T U2563 ( .A1(n1522), .A2(n1521), .ZN(n1523) );
  XOR2XD1BWP12T U2564 ( .A1(n1524), .A2(n1523), .Z(n3096) );
  INVD1BWP12T U2565 ( .I(n1527), .ZN(n1528) );
  AOI21D1BWP12T U2566 ( .A1(n1529), .A2(n605), .B(n1528), .ZN(n1533) );
  CKND2D1BWP12T U2567 ( .A1(n1795), .A2(n1531), .ZN(n1532) );
  XOR2XD1BWP12T U2568 ( .A1(n1533), .A2(n1532), .Z(n2739) );
  TPND2D0BWP12T U2569 ( .A1(n1543), .A2(n1542), .ZN(n1544) );
  XNR2XD1BWP12T U2570 ( .A1(n1545), .A2(n1544), .ZN(n2918) );
  FA1D0BWP12T U2571 ( .A(n340), .B(n2993), .CI(n1547), .CO(n1478), .S(n3022)
         );
  OR4D0BWP12T U2572 ( .A1(n2624), .A2(n1554), .A3(n1553), .A4(n1552), .Z(n2482) );
  INVD1BWP12T U2573 ( .I(n1555), .ZN(n1570) );
  CKND2D1BWP12T U2574 ( .A1(n1569), .A2(n1556), .ZN(n1557) );
  XNR2D1BWP12T U2575 ( .A1(n1570), .A2(n1557), .ZN(n2654) );
  CKND2D1BWP12T U2576 ( .A1(n1559), .A2(n1558), .ZN(n1560) );
  XNR2D1BWP12T U2577 ( .A1(n1561), .A2(n1560), .ZN(n3024) );
  INVD1BWP12T U2578 ( .I(n1562), .ZN(n1638) );
  AOI21D1BWP12T U2579 ( .A1(n1638), .A2(n1637), .B(n1563), .ZN(n1567) );
  ND2D1BWP12T U2580 ( .A1(n1565), .A2(n1564), .ZN(n1566) );
  XOR2XD1BWP12T U2581 ( .A1(n1567), .A2(n1566), .Z(n2628) );
  AOI21D1BWP12T U2582 ( .A1(n1570), .A2(n1569), .B(n1568), .ZN(n1574) );
  ND2D1BWP12T U2583 ( .A1(n1572), .A2(n1571), .ZN(n1573) );
  XOR2XD1BWP12T U2584 ( .A1(n1574), .A2(n1573), .Z(n2923) );
  INVD1BWP12T U2585 ( .I(n1577), .ZN(n1579) );
  CKND2D1BWP12T U2586 ( .A1(n1581), .A2(n1580), .ZN(n1582) );
  XOR2XD1BWP12T U2587 ( .A1(n1583), .A2(n1582), .Z(n2889) );
  ND2D1BWP12T U2588 ( .A1(n1585), .A2(n1584), .ZN(n1587) );
  XNR2D1BWP12T U2589 ( .A1(n1587), .A2(n1586), .ZN(n3050) );
  OR2D0BWP12T U2590 ( .A1(n1609), .A2(n1608), .Z(n1612) );
  INVD0BWP12T U2591 ( .I(n1610), .ZN(n1611) );
  AN2XD1BWP12T U2592 ( .A1(n1612), .A2(n1611), .Z(n3127) );
  OR4D1BWP12T U2593 ( .A1(n3127), .A2(n1614), .A3(n2951), .A4(n1613), .Z(n1618) );
  OR4D1BWP12T U2594 ( .A1(n2759), .A2(n1619), .A3(n1618), .A4(n2760), .Z(n1621) );
  OR4D1BWP12T U2595 ( .A1(n2821), .A2(n2791), .A3(n1621), .A4(n1620), .Z(n1623) );
  OR4D1BWP12T U2596 ( .A1(n3087), .A2(n2865), .A3(n1623), .A4(n1622), .Z(n1631) );
  AOI21D1BWP12T U2597 ( .A1(n1626), .A2(n1625), .B(n1624), .ZN(n1630) );
  ND2D1BWP12T U2598 ( .A1(n1628), .A2(n1627), .ZN(n1629) );
  XOR2XD1BWP12T U2599 ( .A1(n1630), .A2(n1629), .Z(n2712) );
  OR4D0BWP12T U2600 ( .A1(n3050), .A2(n2888), .A3(n1631), .A4(n2712), .Z(n1633) );
  OR4D0BWP12T U2601 ( .A1(n2889), .A2(n1634), .A3(n1633), .A4(n1632), .Z(n1635) );
  ND2D1BWP12T U2602 ( .A1(n1637), .A2(n1636), .ZN(n1639) );
  XNR2D1BWP12T U2603 ( .A1(n1639), .A2(n1638), .ZN(n2990) );
  CKND0BWP12T U2604 ( .I(n1642), .ZN(n1643) );
  TPNR2D0BWP12T U2605 ( .A1(n1643), .A2(n1646), .ZN(n1649) );
  CKND1BWP12T U2606 ( .I(n1644), .ZN(n1647) );
  TPOAI21D0BWP12T U2607 ( .A1(n1647), .A2(n1646), .B(n1645), .ZN(n1648) );
  AOI21D1BWP12T U2608 ( .A1(n1650), .A2(n1649), .B(n1648), .ZN(n1655) );
  INVD1BWP12T U2609 ( .I(n1651), .ZN(n1653) );
  ND2D1BWP12T U2610 ( .A1(n1653), .A2(n1652), .ZN(n1654) );
  XOR2XD1BWP12T U2611 ( .A1(n1655), .A2(n1654), .Z(n2601) );
  FA1D2BWP12T U2612 ( .A(n2608), .B(b[29]), .CI(n1661), .CO(n1370), .S(n2602)
         );
  FA1D2BWP12T U2613 ( .A(n2633), .B(b[23]), .CI(n1662), .CO(n704), .S(n2629)
         );
  CKND2D0BWP12T U2614 ( .A1(n1918), .A2(n1917), .ZN(n1664) );
  XNR2XD0BWP12T U2615 ( .A1(n1665), .A2(n1664), .ZN(n2924) );
  INVD0BWP12T U2616 ( .I(n1666), .ZN(n1836) );
  CKND2D0BWP12T U2617 ( .A1(n1836), .A2(n1835), .ZN(n1667) );
  XOR2XD0BWP12T U2618 ( .A1(n1668), .A2(n1667), .Z(n2655) );
  CKND2D0BWP12T U2619 ( .A1(n1840), .A2(n1839), .ZN(n1669) );
  XNR2XD0BWP12T U2620 ( .A1(n1670), .A2(n1669), .ZN(n2683) );
  INVD1BWP12T U2621 ( .I(n1671), .ZN(n1674) );
  CKND2D1BWP12T U2622 ( .A1(n1683), .A2(n1685), .ZN(n1688) );
  AOI21D1BWP12T U2623 ( .A1(n1686), .A2(n1685), .B(n1684), .ZN(n1687) );
  OAI21D1BWP12T U2624 ( .A1(n1700), .A2(n1688), .B(n1687), .ZN(n1692) );
  ND2D1BWP12T U2625 ( .A1(n1690), .A2(n1689), .ZN(n1691) );
  XNR2XD1BWP12T U2626 ( .A1(n1692), .A2(n1691), .ZN(n3026) );
  INVD1BWP12T U2627 ( .I(n1693), .ZN(n1695) );
  CKND2D1BWP12T U2628 ( .A1(n1695), .A2(n1694), .ZN(n1696) );
  XOR2XD0BWP12T U2629 ( .A1(n1697), .A2(n1696), .Z(n2714) );
  ND2XD0BWP12T U2630 ( .A1(n1860), .A2(n1698), .ZN(n1699) );
  INVD1BWP12T U2631 ( .I(n1701), .ZN(n1702) );
  AOI21D1BWP12T U2632 ( .A1(n1718), .A2(n617), .B(n1702), .ZN(n1706) );
  ND2XD0BWP12T U2633 ( .A1(n1876), .A2(n1704), .ZN(n1705) );
  XOR2XD1BWP12T U2634 ( .A1(n1706), .A2(n1705), .Z(n2741) );
  INVD1BWP12T U2635 ( .I(n1707), .ZN(n1709) );
  CKND2D1BWP12T U2636 ( .A1(n1709), .A2(n1708), .ZN(n1710) );
  CKXOR2D1BWP12T U2637 ( .A1(n1711), .A2(n1710), .Z(n3097) );
  INVD1BWP12T U2638 ( .I(n1854), .ZN(n1849) );
  CKND2D0BWP12T U2639 ( .A1(n1844), .A2(n1843), .ZN(n1723) );
  XNR2XD0BWP12T U2640 ( .A1(n1724), .A2(n1723), .ZN(n1725) );
  INVD1BWP12T U2641 ( .I(n1725), .ZN(n2916) );
  FA1D2BWP12T U2642 ( .A(n2993), .B(b[21]), .CI(n1726), .CO(n1663), .S(n3016)
         );
  FA1D1BWP12T U2643 ( .A(n1736), .B(n2633), .CI(n1735), .CO(n702), .S(n2649)
         );
  CKND2D1BWP12T U2644 ( .A1(n1741), .A2(n1740), .ZN(n1742) );
  XNR2D1BWP12T U2645 ( .A1(n1743), .A2(n1742), .ZN(n2947) );
  CKND2D1BWP12T U2646 ( .A1(n1745), .A2(n1744), .ZN(n1746) );
  XNR2D1BWP12T U2647 ( .A1(n1747), .A2(n1746), .ZN(n2708) );
  CKND2D1BWP12T U2648 ( .A1(n1749), .A2(n1748), .ZN(n1750) );
  XNR2D1BWP12T U2649 ( .A1(n1751), .A2(n1750), .ZN(n2919) );
  OAI21D1BWP12T U2650 ( .A1(n1808), .A2(n1753), .B(n1752), .ZN(n1757) );
  CKND2D1BWP12T U2651 ( .A1(n1540), .A2(n1755), .ZN(n1756) );
  XNR2D1BWP12T U2652 ( .A1(n1757), .A2(n1756), .ZN(n3027) );
  NR3D0BWP12T U2653 ( .A1(n1759), .A2(n1758), .A3(n3027), .ZN(n1813) );
  CKND2D1BWP12T U2654 ( .A1(n1506), .A2(n1761), .ZN(n1762) );
  XOR2XD1BWP12T U2655 ( .A1(n1763), .A2(n1762), .Z(n2735) );
  INVD1BWP12T U2656 ( .I(n1764), .ZN(n1796) );
  INVD1BWP12T U2657 ( .I(n1765), .ZN(n1795) );
  AOI21D1BWP12T U2658 ( .A1(n1796), .A2(n1775), .B(n1777), .ZN(n1774) );
  CKND2D1BWP12T U2659 ( .A1(n1517), .A2(n1778), .ZN(n1773) );
  XOR2XD1BWP12T U2660 ( .A1(n1774), .A2(n1773), .Z(n2792) );
  CKND0BWP12T U2661 ( .I(n1775), .ZN(n1776) );
  NR2D0BWP12T U2662 ( .A1(n1776), .A2(n1779), .ZN(n1782) );
  CKND0BWP12T U2663 ( .I(n1777), .ZN(n1780) );
  TPOAI21D0BWP12T U2664 ( .A1(n1780), .A2(n1779), .B(n1778), .ZN(n1781) );
  AOI21D1BWP12T U2665 ( .A1(n1796), .A2(n1782), .B(n1781), .ZN(n1787) );
  INVD0BWP12T U2666 ( .I(n1783), .ZN(n1785) );
  CKND2D1BWP12T U2667 ( .A1(n1785), .A2(n1784), .ZN(n1786) );
  XOR2XD1BWP12T U2668 ( .A1(n1787), .A2(n1786), .Z(n2824) );
  NR2D0BWP12T U2669 ( .A1(n2792), .A2(n2824), .ZN(n1798) );
  ND2D1BWP12T U2670 ( .A1(n1522), .A2(n1789), .ZN(n1791) );
  XOR2XD1BWP12T U2671 ( .A1(n1791), .A2(n1790), .Z(n3099) );
  NR4D0BWP12T U2672 ( .A1(n1793), .A2(n3099), .A3(n1792), .A4(n3020), .ZN(
        n1797) );
  IND4D0BWP12T U2673 ( .A1(n1799), .B1(n1798), .B2(n1797), .B3(n233), .ZN(
        n1800) );
  OR4D0BWP12T U2674 ( .A1(n1801), .A2(n2763), .A3(n2863), .A4(n1800), .Z(n1811) );
  NR4D0BWP12T U2675 ( .A1(n2735), .A2(n1811), .A3(n3085), .A4(n2866), .ZN(
        n1812) );
  IND3D1BWP12T U2676 ( .A1(n2919), .B1(n1813), .B2(n1812), .ZN(n1818) );
  CKND2D1BWP12T U2677 ( .A1(n1485), .A2(n1815), .ZN(n1816) );
  XOR2XD1BWP12T U2678 ( .A1(n1817), .A2(n1816), .Z(n2678) );
  OR4D0BWP12T U2679 ( .A1(n2708), .A2(n1819), .A3(n1818), .A4(n2678), .Z(n1822) );
  FA1D1BWP12T U2680 ( .A(n1821), .B(n2963), .CI(n1820), .CO(n1735), .S(n2961)
         );
  OR4D0BWP12T U2681 ( .A1(n2991), .A2(n2947), .A3(n1822), .A4(n2961), .Z(n1824) );
  OR4D0BWP12T U2682 ( .A1(n1825), .A2(n2649), .A3(n1824), .A4(n1823), .Z(n1827) );
  OR4D1BWP12T U2683 ( .A1(n1829), .A2(n1828), .A3(n1827), .A4(n1826), .Z(n1830) );
  NR4D0BWP12T U2684 ( .A1(n1832), .A2(n1831), .A3(n2623), .A4(n1830), .ZN(
        n2477) );
  FA1D2BWP12T U2685 ( .A(b[22]), .B(n2963), .CI(n1833), .CO(n1922), .S(n2982)
         );
  FA1D0BWP12T U2686 ( .A(n2993), .B(b[21]), .CI(n1834), .CO(n1833), .S(n3015)
         );
  CKND2D0BWP12T U2687 ( .A1(n1836), .A2(n1835), .ZN(n1837) );
  CKXOR2D1BWP12T U2688 ( .A1(n1838), .A2(n1837), .Z(n2656) );
  ND2XD0BWP12T U2689 ( .A1(n1840), .A2(n1839), .ZN(n1841) );
  XNR2XD1BWP12T U2690 ( .A1(n1842), .A2(n1841), .ZN(n2684) );
  ND2XD0BWP12T U2691 ( .A1(n1844), .A2(n1843), .ZN(n1845) );
  XNR2XD1BWP12T U2692 ( .A1(n1846), .A2(n1845), .ZN(n2890) );
  NR2D0BWP12T U2693 ( .A1(n1847), .A2(n2890), .ZN(n1916) );
  INVD1BWP12T U2694 ( .I(n1848), .ZN(n1877) );
  CKND0BWP12T U2695 ( .I(n1850), .ZN(n1851) );
  NR2D1BWP12T U2696 ( .A1(n1851), .A2(n1854), .ZN(n1857) );
  CKND0BWP12T U2697 ( .I(n1852), .ZN(n1855) );
  OAI21D1BWP12T U2698 ( .A1(n1855), .A2(n1854), .B(n1853), .ZN(n1856) );
  AOI21D1BWP12T U2699 ( .A1(n1877), .A2(n1857), .B(n1856), .ZN(n1862) );
  INVD0BWP12T U2700 ( .I(n1858), .ZN(n1860) );
  CKND2D1BWP12T U2701 ( .A1(n1860), .A2(n1859), .ZN(n1861) );
  XOR2XD1BWP12T U2702 ( .A1(n1862), .A2(n1861), .Z(n2839) );
  NR2D0BWP12T U2703 ( .A1(n2794), .A2(n2839), .ZN(n1873) );
  ND2D1BWP12T U2704 ( .A1(n1709), .A2(n1864), .ZN(n1866) );
  XOR2XD1BWP12T U2705 ( .A1(n1866), .A2(n1865), .Z(n3120) );
  NR4D0BWP12T U2706 ( .A1(n1869), .A2(n3120), .A3(n1868), .A4(n1867), .ZN(
        n1872) );
  INVD1BWP12T U2707 ( .I(n1870), .ZN(n1876) );
  CKND0BWP12T U2708 ( .I(n2740), .ZN(n1871) );
  IND4D0BWP12T U2709 ( .A1(n1874), .B1(n1873), .B2(n1872), .B3(n1871), .ZN(
        n1886) );
  INVD0BWP12T U2710 ( .I(n1878), .ZN(n1880) );
  NR4D0BWP12T U2711 ( .A1(n1886), .A2(n1885), .A3(n2777), .A4(n2850), .ZN(
        n1915) );
  INVD1BWP12T U2712 ( .I(n1887), .ZN(n1890) );
  NR2D0BWP12T U2713 ( .A1(n3062), .A2(n2873), .ZN(n1914) );
  TPND2D0BWP12T U2714 ( .A1(n1695), .A2(n1895), .ZN(n1896) );
  XOR2XD1BWP12T U2715 ( .A1(n1897), .A2(n1896), .Z(n2713) );
  CKND0BWP12T U2716 ( .I(n1898), .ZN(n1899) );
  CKND2D1BWP12T U2717 ( .A1(n1899), .A2(n1902), .ZN(n1905) );
  CKND0BWP12T U2718 ( .I(n1900), .ZN(n1903) );
  AOI21D1BWP12T U2719 ( .A1(n1903), .A2(n1902), .B(n1901), .ZN(n1904) );
  OAI21D1BWP12T U2720 ( .A1(n1906), .A2(n1905), .B(n1904), .ZN(n1910) );
  ND2D1BWP12T U2721 ( .A1(n1908), .A2(n1907), .ZN(n1909) );
  XNR2D1BWP12T U2722 ( .A1(n1910), .A2(n1909), .ZN(n3028) );
  NR4D0BWP12T U2723 ( .A1(n1912), .A2(n1911), .A3(n2713), .A4(n3028), .ZN(
        n1913) );
  ND4D1BWP12T U2724 ( .A1(n1916), .A2(n1915), .A3(n1914), .A4(n1913), .ZN(
        n1921) );
  CKND2D0BWP12T U2725 ( .A1(n1918), .A2(n1917), .ZN(n1919) );
  XNR2XD1BWP12T U2726 ( .A1(n1920), .A2(n1919), .ZN(n2925) );
  OR4D0BWP12T U2727 ( .A1(n2656), .A2(n2684), .A3(n1921), .A4(n2925), .Z(n1923) );
  FA1D1BWP12T U2728 ( .A(n2633), .B(b[23]), .CI(n1922), .CO(n705), .S(n2630)
         );
  OR4D0BWP12T U2729 ( .A1(n2982), .A2(n3015), .A3(n1923), .A4(n2630), .Z(n1925) );
  OR4D1BWP12T U2730 ( .A1(n1927), .A2(n1926), .A3(n1925), .A4(n1924), .Z(n1929) );
  FA1D1BWP12T U2731 ( .A(n2608), .B(b[29]), .CI(n1928), .CO(n1324), .S(n2603)
         );
  OR4D1BWP12T U2732 ( .A1(n1931), .A2(n1930), .A3(n1929), .A4(n2603), .Z(n2474) );
  NR4D0BWP12T U2733 ( .A1(n2956), .A2(a[26]), .A3(n2518), .A4(n2403), .ZN(
        n1935) );
  NR4D0BWP12T U2734 ( .A1(n2608), .A2(a[28]), .A3(n2502), .A4(n3067), .ZN(
        n1934) );
  NR4D0BWP12T U2735 ( .A1(a[14]), .A2(n2851), .A3(n2398), .A4(n2874), .ZN(
        n1933) );
  NR4D0BWP12T U2736 ( .A1(n2689), .A2(n2720), .A3(n3033), .A4(n2416), .ZN(
        n1932) );
  ND4D1BWP12T U2737 ( .A1(n1935), .A2(n1934), .A3(n1933), .A4(n1932), .ZN(
        n1991) );
  NR4D0BWP12T U2738 ( .A1(n2993), .A2(a[20]), .A3(n2657), .A4(n2963), .ZN(
        n1940) );
  NR4D0BWP12T U2739 ( .A1(n2764), .A2(n2748), .A3(n2406), .A4(n3110), .ZN(
        n1936) );
  AN4D0BWP12T U2740 ( .A1(n2636), .A2(n1937), .A3(n2996), .A4(n1936), .Z(n1939) );
  NR4D0BWP12T U2741 ( .A1(n2560), .A2(n2891), .A3(n2799), .A4(a[7]), .ZN(n1938) );
  ND4D0BWP12T U2742 ( .A1(n1941), .A2(n1940), .A3(n1939), .A4(n1938), .ZN(
        n1990) );
  HA1D1BWP12T U2743 ( .A(n2607), .B(n1942), .CO(n1323), .S(n2617) );
  HA1D0BWP12T U2744 ( .A(n1944), .B(n1943), .CO(n706), .S(n2644) );
  HA1D0BWP12T U2745 ( .A(n2965), .B(n1945), .CO(n1943), .S(n2962) );
  CKND0BWP12T U2746 ( .I(n1946), .ZN(n1947) );
  NR2D1BWP12T U2747 ( .A1(n1964), .A2(n1947), .ZN(n1948) );
  XNR2XD0BWP12T U2748 ( .A1(n1948), .A2(n2689), .ZN(n2702) );
  NR2XD0BWP12T U2749 ( .A1(n1964), .A2(n1949), .ZN(n1950) );
  XNR2XD0BWP12T U2750 ( .A1(n1950), .A2(n2657), .ZN(n2672) );
  HA1D0BWP12T U2751 ( .A(n1952), .B(n1951), .CO(n1945), .S(n2992) );
  NR4D0BWP12T U2752 ( .A1(n1953), .A2(n2702), .A3(n2672), .A4(n2992), .ZN(
        n1979) );
  HICIND1BWP12T U2753 ( .A(n2928), .CIN(n1954), .CO(n1951), .S(n2940) );
  INVD1BWP12T U2754 ( .I(n1955), .ZN(n1973) );
  CKXOR2D0BWP12T U2755 ( .A1(n1973), .A2(n2748), .Z(n2754) );
  XNR2XD1BWP12T U2756 ( .A1(n3110), .A2(n2486), .ZN(n3116) );
  OR4D0BWP12T U2757 ( .A1(n3116), .A2(n2980), .A3(n1957), .A4(n1956), .Z(n1959) );
  OR4D0BWP12T U2758 ( .A1(n2940), .A2(n2754), .A3(n1959), .A4(n1958), .Z(n1965) );
  CKND0BWP12T U2759 ( .I(n1960), .ZN(n1961) );
  NR2D0BWP12T U2760 ( .A1(n1961), .A2(n2416), .ZN(n1962) );
  CKND2D1BWP12T U2761 ( .A1(n1962), .A2(n1970), .ZN(n1963) );
  XOR2XD1BWP12T U2762 ( .A1(n1963), .A2(n3033), .Z(n3029) );
  CKXOR2D0BWP12T U2763 ( .A1(n1964), .A2(n2891), .Z(n2913) );
  NR3D0BWP12T U2764 ( .A1(n1965), .A2(n3029), .A3(n2913), .ZN(n1978) );
  CKND0BWP12T U2765 ( .I(n1968), .ZN(n1966) );
  CKND2D1BWP12T U2766 ( .A1(n1970), .A2(n1966), .ZN(n1967) );
  XOR2XD1BWP12T U2767 ( .A1(n1967), .A2(n3067), .Z(n3063) );
  OR4D0BWP12T U2768 ( .A1(n2843), .A2(n3063), .A3(n2886), .A4(n1969), .Z(n1976) );
  OR3XD0BWP12T U2769 ( .A1(n1974), .A2(n2716), .A3(n2762), .Z(n1975) );
  NR4D0BWP12T U2770 ( .A1(n1976), .A2(n2845), .A3(n2793), .A4(n1975), .ZN(
        n1977) );
  IND4D1BWP12T U2771 ( .A1(n2962), .B1(n1979), .B2(n1978), .B3(n1977), .ZN(
        n1981) );
  OR4D0BWP12T U2772 ( .A1(n1982), .A2(n2644), .A3(n1981), .A4(n1980), .Z(n1984) );
  OR4D1BWP12T U2773 ( .A1(n1986), .A2(n1985), .A3(n1984), .A4(n1983), .Z(n1987) );
  OR4D1BWP12T U2774 ( .A1(n1988), .A2(n2617), .A3(n1987), .A4(n2596), .Z(n1989) );
  OAI31D0BWP12T U2775 ( .A1(n1991), .A2(n2090), .A3(n1990), .B(n1989), .ZN(
        n2471) );
  CKND0BWP12T U2776 ( .I(n1992), .ZN(n1993) );
  AOI21D0BWP12T U2777 ( .A1(n1993), .A2(n2750), .B(n2359), .ZN(n1994) );
  TPNR2D0BWP12T U2778 ( .A1(n1994), .A2(n2093), .ZN(n2007) );
  CKND1BWP12T U2779 ( .I(n2002), .ZN(n2066) );
  AOI22D1BWP12T U2780 ( .A1(n2066), .A2(n2874), .B1(n2065), .B2(n3067), .ZN(
        n1998) );
  INR2D0BWP12T U2781 ( .A1(n2851), .B1(n2000), .ZN(n1996) );
  TPNR2D0BWP12T U2782 ( .A1(n1999), .A2(n2281), .ZN(n1995) );
  NR2D1BWP12T U2783 ( .A1(n1996), .A2(n1995), .ZN(n1997) );
  ND2D1BWP12T U2784 ( .A1(n1998), .A2(n1997), .ZN(n2069) );
  OAI22D1BWP12T U2785 ( .A1(n2000), .A2(n3031), .B1(n1999), .B2(n2893), .ZN(
        n2004) );
  OAI22D1BWP12T U2786 ( .A1(n2002), .A2(n2722), .B1(n2001), .B2(n2280), .ZN(
        n2003) );
  NR2D1BWP12T U2787 ( .A1(n2004), .A2(n2003), .ZN(n2099) );
  OAI22D0BWP12T U2788 ( .A1(n2098), .A2(n2110), .B1(n2099), .B2(n2095), .ZN(
        n2006) );
  OAI21D0BWP12T U2789 ( .A1(n2096), .A2(n2133), .B(n2431), .ZN(n2005) );
  AOI211D1BWP12T U2790 ( .A1(n2089), .A2(n2069), .B(n2006), .C(n2005), .ZN(
        n2435) );
  TPOAI21D0BWP12T U2791 ( .A1(n2007), .A2(n2435), .B(n2114), .ZN(n2847) );
  CKND2D0BWP12T U2792 ( .A1(n2026), .A2(n2349), .ZN(n2092) );
  AOI21D0BWP12T U2793 ( .A1(n2021), .A2(n2092), .B(n2009), .ZN(n2604) );
  AOI21D0BWP12T U2794 ( .A1(n2033), .A2(n2010), .B(n2009), .ZN(n2012) );
  MUX2NXD0BWP12T U2795 ( .I0(n2044), .I1(n2011), .S(n2405), .ZN(n2080) );
  CKND2D1BWP12T U2796 ( .A1(n2080), .A2(n2349), .ZN(n2196) );
  TPOAI21D0BWP12T U2797 ( .A1(n2040), .A2(n2196), .B(n2021), .ZN(n2632) );
  NR4D0BWP12T U2798 ( .A1(n2847), .A2(n2604), .A3(n2012), .A4(n2632), .ZN(
        n2025) );
  OAI211D0BWP12T U2799 ( .A1(n2297), .A2(n2197), .B(n2936), .C(n2750), .ZN(
        n2020) );
  OA22D1BWP12T U2800 ( .A1(n2015), .A2(n2133), .B1(n2014), .B2(n2150), .Z(
        n2018) );
  AOI21D0BWP12T U2801 ( .A1(n2016), .A2(n2108), .B(n2750), .ZN(n2017) );
  OAI211D1BWP12T U2802 ( .A1(n2019), .A2(n2110), .B(n2018), .C(n2017), .ZN(
        n2136) );
  AOI31D1BWP12T U2803 ( .A1(n2020), .A2(n2452), .A3(n2136), .B(n2101), .ZN(
        n2757) );
  AOI21D0BWP12T U2804 ( .A1(n2297), .A2(n2039), .B(n2021), .ZN(n2023) );
  INVD1BWP12T U2805 ( .I(n2936), .ZN(n2447) );
  OAI21D1BWP12T U2806 ( .A1(n2023), .A2(n2447), .B(n2022), .ZN(n2937) );
  ND4D0BWP12T U2807 ( .A1(n2025), .A2(n2757), .A3(n2024), .A4(n2937), .ZN(
        n2043) );
  OAI22D1BWP12T U2808 ( .A1(n2098), .A2(n2150), .B1(n2097), .B2(n2095), .ZN(
        n2134) );
  AOI21D1BWP12T U2809 ( .A1(n2026), .A2(n2407), .B(n2134), .ZN(n3006) );
  AN4D0BWP12T U2810 ( .A1(n2667), .A2(n2027), .A3(n2897), .A4(n3006), .Z(n2032) );
  OAI22D0BWP12T U2811 ( .A1(n2029), .A2(n2095), .B1(n2028), .B2(n2150), .ZN(
        n2199) );
  AOI21D1BWP12T U2812 ( .A1(n2030), .A2(n2407), .B(n2199), .ZN(n2972) );
  AOI31D0BWP12T U2813 ( .A1(n2032), .A2(n2031), .A3(n2972), .B(n2040), .ZN(
        n2042) );
  INVD1BWP12T U2814 ( .I(n2033), .ZN(n2034) );
  AOI21D1BWP12T U2815 ( .A1(n2034), .A2(n2452), .B(n2459), .ZN(n2038) );
  AOI21D0BWP12T U2816 ( .A1(n2109), .A2(n2089), .B(n2750), .ZN(n2035) );
  OAI21D0BWP12T U2817 ( .A1(n2113), .A2(n2095), .B(n2035), .ZN(n2036) );
  AOI21D1BWP12T U2818 ( .A1(n2407), .A2(n2037), .B(n2036), .ZN(n3082) );
  OAI21D1BWP12T U2819 ( .A1(n2038), .A2(n3082), .B(n2114), .ZN(n3055) );
  OAI21D1BWP12T U2820 ( .A1(n2041), .A2(n2040), .B(n2039), .ZN(n2698) );
  NR4D0BWP12T U2821 ( .A1(n2043), .A2(n2042), .A3(n3055), .A4(n2698), .ZN(
        n2120) );
  CKND0BWP12T U2822 ( .I(n2057), .ZN(n2047) );
  OAI22D0BWP12T U2823 ( .A1(n2044), .A2(n2110), .B1(n2056), .B2(n2133), .ZN(
        n2046) );
  OAI21D0BWP12T U2824 ( .A1(n2058), .A2(n2150), .B(n2431), .ZN(n2045) );
  AO211D1BWP12T U2825 ( .A1(n2108), .A2(n2047), .B(n2046), .C(n2045), .Z(n2139) );
  CKND0BWP12T U2826 ( .I(n2048), .ZN(n2049) );
  OAI21D0BWP12T U2827 ( .A1(n2049), .A2(n2437), .B(n2448), .ZN(n2050) );
  AOI21D0BWP12T U2828 ( .A1(n2139), .A2(n2050), .B(n2101), .ZN(n2884) );
  CKND2D0BWP12T U2829 ( .A1(n2051), .A2(n3130), .ZN(n2052) );
  AOI211D0BWP12T U2830 ( .A1(n2054), .A2(n2207), .B(n2053), .C(n2052), .ZN(
        n2062) );
  OAI21D0BWP12T U2831 ( .A1(n2080), .A2(n2431), .B(n2343), .ZN(n2055) );
  CKND2D0BWP12T U2832 ( .A1(n2055), .A2(n2197), .ZN(n2060) );
  MUX2XD1BWP12T U2833 ( .I0(n2057), .I1(n2056), .S(n2405), .Z(n2081) );
  AOI31D1BWP12T U2834 ( .A1(n2060), .A2(n2452), .A3(n2823), .B(n2101), .ZN(
        n2826) );
  ND4D0BWP12T U2835 ( .A1(n2884), .A2(n2062), .A3(n2826), .A4(n2061), .ZN(
        n2105) );
  AOI22D0BWP12T U2836 ( .A1(n2064), .A2(n2764), .B1(n2063), .B2(n2398), .ZN(
        n2068) );
  AOI22D0BWP12T U2837 ( .A1(n2066), .A2(a[7]), .B1(n2065), .B2(n2799), .ZN(
        n2067) );
  CKND2D1BWP12T U2838 ( .A1(n2068), .A2(n2067), .ZN(n2088) );
  INVD1BWP12T U2839 ( .I(n2069), .ZN(n2085) );
  OAI22D1BWP12T U2840 ( .A1(n2099), .A2(n2110), .B1(n2085), .B2(n2133), .ZN(
        n2077) );
  AOI22D0BWP12T U2841 ( .A1(n2071), .A2(n2404), .B1(n2070), .B2(n3110), .ZN(
        n2075) );
  AOI22D0BWP12T U2842 ( .A1(n2748), .A2(n2073), .B1(n2072), .B2(n2406), .ZN(
        n2074) );
  AOI21D0BWP12T U2843 ( .A1(n2075), .A2(n2074), .B(n2407), .ZN(n2076) );
  AOI211D1BWP12T U2844 ( .A1(n2108), .A2(n2088), .B(n2077), .C(n2076), .ZN(
        n3101) );
  AOI21D1BWP12T U2845 ( .A1(n3101), .A2(n2431), .B(n2090), .ZN(n3092) );
  TPOAI21D0BWP12T U2846 ( .A1(n2078), .A2(n2431), .B(n3092), .ZN(n2079) );
  CKND2D1BWP12T U2847 ( .A1(n2079), .A2(n2114), .ZN(n3129) );
  CKND0BWP12T U2848 ( .I(n2080), .ZN(n2083) );
  OAI22D1BWP12T U2849 ( .A1(n2083), .A2(n2082), .B1(n2081), .B2(n2375), .ZN(
        n2719) );
  AOI21D1BWP12T U2850 ( .A1(n2719), .A2(n2452), .B(n2084), .ZN(n2731) );
  CKND2D0BWP12T U2851 ( .A1(n3006), .A2(n2750), .ZN(n2091) );
  OAI22D0BWP12T U2852 ( .A1(n2096), .A2(n2110), .B1(n2085), .B2(n2095), .ZN(
        n2087) );
  OAI21D0BWP12T U2853 ( .A1(n2099), .A2(n2133), .B(n2431), .ZN(n2086) );
  AOI211D1BWP12T U2854 ( .A1(n2089), .A2(n2088), .B(n2087), .C(n2086), .ZN(
        n2195) );
  NR2D1BWP12T U2855 ( .A1(n2195), .A2(n2090), .ZN(n2441) );
  AOI21D1BWP12T U2856 ( .A1(n2091), .A2(n2441), .B(n2101), .ZN(n2761) );
  CKND0BWP12T U2857 ( .I(n2092), .ZN(n2094) );
  OAI21D1BWP12T U2858 ( .A1(n2094), .A2(n2093), .B(n2452), .ZN(n2100) );
  AOI21D0BWP12T U2859 ( .A1(n2100), .A2(n2448), .B(n2149), .ZN(n2102) );
  NR2D0BWP12T U2860 ( .A1(n2102), .A2(n2101), .ZN(n3045) );
  ND4D0BWP12T U2861 ( .A1(n2103), .A2(n2731), .A3(n2761), .A4(n3045), .ZN(
        n2104) );
  NR4D0BWP12T U2862 ( .A1(n2106), .A2(n2105), .A3(n3129), .A4(n2104), .ZN(
        n2119) );
  CKND0BWP12T U2863 ( .I(n2972), .ZN(n2107) );
  AOI21D1BWP12T U2864 ( .A1(n2107), .A2(n2452), .B(n2459), .ZN(n2115) );
  OAI21D1BWP12T U2865 ( .A1(n2115), .A2(n2812), .B(n2114), .ZN(n2816) );
  NR2D0BWP12T U2866 ( .A1(n2816), .A2(n2116), .ZN(n2117) );
  ND4D0BWP12T U2867 ( .A1(n2120), .A2(n2119), .A3(n2118), .A4(n2117), .ZN(
        n2132) );
  ND4D0BWP12T U2868 ( .A1(n2851), .A2(n2398), .A3(n3067), .A4(n2874), .ZN(
        n2124) );
  ND4D0BWP12T U2869 ( .A1(n2608), .A2(a[28]), .A3(n2502), .A4(n2403), .ZN(
        n2123) );
  ND4D0BWP12T U2870 ( .A1(n2406), .A2(n2404), .A3(n3110), .A4(n2262), .ZN(
        n2122) );
  ND4D0BWP12T U2871 ( .A1(n2633), .A2(n2963), .A3(n2993), .A4(a[20]), .ZN(
        n2121) );
  NR4D0BWP12T U2872 ( .A1(n2124), .A2(n2123), .A3(n2122), .A4(n2121), .ZN(
        n2130) );
  AN4D0BWP12T U2873 ( .A1(n2518), .A2(a[26]), .A3(n2748), .A4(n2764), .Z(n2129) );
  CKND2D0BWP12T U2874 ( .A1(n2720), .A2(n2799), .ZN(n2126) );
  ND4D0BWP12T U2875 ( .A1(n2560), .A2(n2891), .A3(n3033), .A4(n2416), .ZN(
        n2125) );
  NR4D0BWP12T U2876 ( .A1(n2280), .A2(n2126), .A3(n2125), .A4(n3109), .ZN(
        n2128) );
  AN4D0BWP12T U2877 ( .A1(n2689), .A2(n2657), .A3(a[30]), .A4(a[7]), .Z(n2127)
         );
  ND4D1BWP12T U2878 ( .A1(n2130), .A2(n2129), .A3(n2128), .A4(n2127), .ZN(
        n2131) );
  MUX2ND0BWP12T U2879 ( .I0(n2132), .I1(n2131), .S(n2956), .ZN(n2470) );
  INVD1BWP12T U2880 ( .I(n2136), .ZN(n2751) );
  CKND2D0BWP12T U2881 ( .A1(n2936), .A2(n3003), .ZN(n2456) );
  INVD1BWP12T U2882 ( .I(n2234), .ZN(n2835) );
  OAI22D1BWP12T U2883 ( .A1(n2835), .A2(n2170), .B1(n2230), .B2(n2211), .ZN(
        n2715) );
  AOI22D1BWP12T U2884 ( .A1(n2136), .A2(n2447), .B1(n2908), .B2(n2135), .ZN(
        n2744) );
  OAI21D1BWP12T U2885 ( .A1(n2140), .A2(n2431), .B(n2139), .ZN(n2871) );
  TPND2D0BWP12T U2886 ( .A1(n2181), .A2(n2142), .ZN(n2148) );
  AOI22D0BWP12T U2887 ( .A1(n2185), .A2(n2144), .B1(n2183), .B2(n2143), .ZN(
        n2147) );
  TPND2D0BWP12T U2888 ( .A1(n2187), .A2(n2145), .ZN(n2146) );
  ND3D1BWP12T U2889 ( .A1(n2148), .A2(n2147), .A3(n2146), .ZN(n2220) );
  MUX2NXD0BWP12T U2890 ( .I0(n2220), .I1(n2216), .S(n2229), .ZN(n2151) );
  OAI21D1BWP12T U2891 ( .A1(n2151), .A2(n2217), .B(n3037), .ZN(n3025) );
  NR2XD0BWP12T U2892 ( .A1(n2454), .A2(n2431), .ZN(n2153) );
  OAI22D1BWP12T U2893 ( .A1(n2154), .A2(n2217), .B1(n2435), .B2(n2153), .ZN(
        n2864) );
  AOI21D0BWP12T U2894 ( .A1(n2212), .A2(n2431), .B(n2388), .ZN(n2161) );
  AOI22D0BWP12T U2895 ( .A1(n2908), .A2(n2156), .B1(n2155), .B2(n2229), .ZN(
        n2158) );
  NR2D1BWP12T U2896 ( .A1(n2178), .A2(n2157), .ZN(n2232) );
  OAI211D0BWP12T U2897 ( .A1(n2159), .A2(n2868), .B(n2158), .C(n2232), .ZN(
        n2160) );
  OAI21D1BWP12T U2898 ( .A1(n2162), .A2(n2161), .B(n2160), .ZN(n2685) );
  OAI222D1BWP12T U2899 ( .A1(n2170), .A2(n2167), .B1(n2179), .B2(n2166), .C1(
        n2211), .C2(n2165), .ZN(n2926) );
  OAI222D1BWP12T U2900 ( .A1(n2179), .A2(n2800), .B1(n2170), .B2(n2169), .C1(
        n2211), .C2(n2168), .ZN(n2976) );
  AOI22D0BWP12T U2901 ( .A1(n2185), .A2(n2318), .B1(n2183), .B2(n2171), .ZN(
        n2173) );
  CKND2D0BWP12T U2902 ( .A1(n2187), .A2(n2317), .ZN(n2172) );
  CKND2D1BWP12T U2903 ( .A1(n2173), .A2(n2172), .ZN(n2177) );
  NR2D0BWP12T U2904 ( .A1(n2175), .A2(n2174), .ZN(n2176) );
  NR2D1BWP12T U2905 ( .A1(n2177), .A2(n2176), .ZN(n2215) );
  AOI22D0BWP12T U2906 ( .A1(n2178), .A2(n2216), .B1(n2215), .B2(n2904), .ZN(
        n2193) );
  INVD1BWP12T U2907 ( .I(n2179), .ZN(n2906) );
  CKND2D0BWP12T U2908 ( .A1(n2181), .A2(n2180), .ZN(n2190) );
  AOI22D0BWP12T U2909 ( .A1(n2185), .A2(n2184), .B1(n2183), .B2(n2182), .ZN(
        n2189) );
  CKND2D0BWP12T U2910 ( .A1(n2187), .A2(n2186), .ZN(n2188) );
  AOI31D0BWP12T U2911 ( .A1(n2190), .A2(n2189), .A3(n2188), .B(n2211), .ZN(
        n2191) );
  AOI21D0BWP12T U2912 ( .A1(n2220), .A2(n2906), .B(n2191), .ZN(n2192) );
  CKND2D1BWP12T U2913 ( .A1(n2193), .A2(n2192), .ZN(n2616) );
  INVD1BWP12T U2914 ( .I(n2195), .ZN(n2776) );
  CKND2D0BWP12T U2915 ( .A1(n3003), .A2(n2750), .ZN(n2440) );
  CKND0BWP12T U2916 ( .I(n2199), .ZN(n2203) );
  CKND2D0BWP12T U2917 ( .A1(n2201), .A2(n2200), .ZN(n2202) );
  ND2D1BWP12T U2918 ( .A1(n2203), .A2(n2202), .ZN(n2798) );
  ND4D0BWP12T U2919 ( .A1(n2613), .A2(n2205), .A3(n2432), .A4(n2204), .ZN(
        n2206) );
  NR3D0BWP12T U2920 ( .A1(n2798), .A2(n2207), .A3(n2206), .ZN(n2208) );
  CKND2D0BWP12T U2921 ( .A1(n2822), .A2(n2208), .ZN(n2460) );
  OAI22D1BWP12T U2922 ( .A1(n2453), .A2(n2431), .B1(n2211), .B2(n2210), .ZN(
        n3090) );
  INVD1BWP12T U2923 ( .I(n2215), .ZN(n2218) );
  INVD1BWP12T U2924 ( .I(n2216), .ZN(n2772) );
  AOI22D0BWP12T U2925 ( .A1(n2218), .A2(n2908), .B1(n2217), .B2(n2772), .ZN(
        n2219) );
  OAI211D0BWP12T U2926 ( .A1(n2221), .A2(n2220), .B(n2219), .C(n2232), .ZN(
        n3013) );
  AOI22D0BWP12T U2927 ( .A1(n2908), .A2(n2226), .B1(n2225), .B2(n2229), .ZN(
        n2227) );
  OAI211D0BWP12T U2928 ( .A1(n2868), .A2(n2228), .B(n2227), .C(n2232), .ZN(
        n2669) );
  AOI22D0BWP12T U2929 ( .A1(n2231), .A2(n2908), .B1(n2230), .B2(n2229), .ZN(
        n2233) );
  OAI211D0BWP12T U2930 ( .A1(n2868), .A2(n2234), .B(n2233), .C(n2232), .ZN(
        n2631) );
  AOI22D0BWP12T U2931 ( .A1(n2963), .A2(n1821), .B1(n1279), .B2(n2502), .ZN(
        n2245) );
  AOI22D0BWP12T U2932 ( .A1(a[20]), .A2(n2238), .B1(n1736), .B2(n2633), .ZN(
        n2244) );
  AOI22D0BWP12T U2933 ( .A1(n2689), .A2(n2239), .B1(n340), .B2(n2993), .ZN(
        n2243) );
  AOI22D0BWP12T U2934 ( .A1(n2891), .A2(n2241), .B1(n2240), .B2(n2657), .ZN(
        n2242) );
  ND4D1BWP12T U2935 ( .A1(n2245), .A2(n2244), .A3(n2243), .A4(n2242), .ZN(
        n2274) );
  AOI22D0BWP12T U2936 ( .A1(a[14]), .A2(n2247), .B1(n2246), .B2(n2560), .ZN(
        n2257) );
  AOI22D1BWP12T U2937 ( .A1(n2416), .A2(n2249), .B1(n2248), .B2(n2720), .ZN(
        n2256) );
  AOI22D0BWP12T U2938 ( .A1(n3067), .A2(n2251), .B1(n2250), .B2(n3033), .ZN(
        n2255) );
  AOI22D1BWP12T U2939 ( .A1(n2874), .A2(n2253), .B1(n2252), .B2(n2398), .ZN(
        n2254) );
  ND4D1BWP12T U2940 ( .A1(n2257), .A2(n2256), .A3(n2255), .A4(n2254), .ZN(
        n2273) );
  AOI22D1BWP12T U2941 ( .A1(n2799), .A2(n2259), .B1(n2258), .B2(n2851), .ZN(
        n2266) );
  AOI22D0BWP12T U2942 ( .A1(n2748), .A2(n2431), .B1(n2260), .B2(a[7]), .ZN(
        n2265) );
  AOI22D0BWP12T U2943 ( .A1(n2404), .A2(n2297), .B1(n2261), .B2(n2764), .ZN(
        n2264) );
  AOI22D0BWP12T U2944 ( .A1(n2406), .A2(n2349), .B1(n2422), .B2(n2262), .ZN(
        n2263) );
  ND4D1BWP12T U2945 ( .A1(n2266), .A2(n2265), .A3(n2264), .A4(n2263), .ZN(
        n2272) );
  AOI22D0BWP12T U2946 ( .A1(a[28]), .A2(n1205), .B1(n1322), .B2(a[30]), .ZN(
        n2270) );
  AOI22D0BWP12T U2947 ( .A1(a[26]), .A2(n471), .B1(n1734), .B2(n2608), .ZN(
        n2269) );
  AOI22D0BWP12T U2948 ( .A1(n2403), .A2(n703), .B1(n651), .B2(n2518), .ZN(
        n2268) );
  CKND2D0BWP12T U2949 ( .A1(n3111), .A2(n3110), .ZN(n2267) );
  ND4D1BWP12T U2950 ( .A1(n2270), .A2(n2269), .A3(n2268), .A4(n2267), .ZN(
        n2271) );
  NR4D0BWP12T U2951 ( .A1(n2274), .A2(n2273), .A3(n2272), .A4(n2271), .ZN(
        n2430) );
  AOI22D0BWP12T U2952 ( .A1(b[23]), .A2(n2636), .B1(n2965), .B2(b[22]), .ZN(
        n2279) );
  AOI22D0BWP12T U2953 ( .A1(b[20]), .A2(n2928), .B1(n2998), .B2(b[21]), .ZN(
        n2278) );
  AOI22D0BWP12T U2954 ( .A1(b[18]), .A2(n2687), .B1(n2659), .B2(n2663), .ZN(
        n2277) );
  AOI22D0BWP12T U2955 ( .A1(b[16]), .A2(n2893), .B1(n2275), .B2(b[17]), .ZN(
        n2276) );
  ND4D1BWP12T U2956 ( .A1(n2279), .A2(n2278), .A3(n2277), .A4(n2276), .ZN(
        n2309) );
  AOI22D0BWP12T U2957 ( .A1(b[15]), .A2(n2722), .B1(n2280), .B2(n2522), .ZN(
        n2286) );
  AOI22D1BWP12T U2958 ( .A1(n2489), .A2(n2281), .B1(n3031), .B2(b[13]), .ZN(
        n2285) );
  AOI22D0BWP12T U2959 ( .A1(n2880), .A2(n2876), .B1(n3069), .B2(n3074), .ZN(
        n2284) );
  AOI22D0BWP12T U2960 ( .A1(n2501), .A2(n2282), .B1(n2853), .B2(n2857), .ZN(
        n2283) );
  ND4D1BWP12T U2961 ( .A1(n2286), .A2(n2285), .A3(n2284), .A4(n2283), .ZN(
        n2308) );
  AO22XD0BWP12T U2962 ( .A1(b[28]), .A2(n2287), .B1(n2607), .B2(b[29]), .Z(
        n2288) );
  AOI211D0BWP12T U2963 ( .A1(b[30]), .A2(n2289), .B(n2288), .C(n3066), .ZN(
        n2296) );
  AOI22D0BWP12T U2964 ( .A1(b[27]), .A2(n2291), .B1(n2290), .B2(b[26]), .ZN(
        n2295) );
  AOI22D0BWP12T U2965 ( .A1(b[24]), .A2(n2293), .B1(n2292), .B2(b[25]), .ZN(
        n2294) );
  ND4D0BWP12T U2966 ( .A1(n2296), .A2(n2295), .A3(n2294), .A4(n2593), .ZN(
        n2303) );
  AOI22D1BWP12T U2967 ( .A1(n2829), .A2(n2831), .B1(n2802), .B2(n2807), .ZN(
        n2302) );
  AOI22D0BWP12T U2968 ( .A1(n2750), .A2(n2749), .B1(n2768), .B2(n2766), .ZN(
        n2301) );
  OAI22D0BWP12T U2969 ( .A1(n2404), .A2(n2297), .B1(n2349), .B2(n2406), .ZN(
        n2299) );
  AOI211D0BWP12T U2970 ( .A1(n3102), .A2(n3108), .B(n2299), .C(n2298), .ZN(
        n2300) );
  IND4D1BWP12T U2971 ( .A1(n2303), .B1(n2302), .B2(n2301), .B3(n2300), .ZN(
        n2307) );
  OAI21D0BWP12T U2972 ( .A1(n2305), .A2(b[31]), .B(n2304), .ZN(n2306) );
  TPOAI31D0BWP12T U2973 ( .A1(n2309), .A2(n2308), .A3(n2307), .B(n2306), .ZN(
        n2429) );
  MUX2ND0BWP12T U2974 ( .I0(n2387), .I1(n2838), .S(n2407), .ZN(n2316) );
  NR2XD0BWP12T U2975 ( .A1(n2316), .A2(n2448), .ZN(n2728) );
  AOI22D0BWP12T U2976 ( .A1(n2331), .A2(n2318), .B1(n595), .B2(n2317), .ZN(
        n2321) );
  CKND2D0BWP12T U2977 ( .A1(n2319), .A2(n2334), .ZN(n2320) );
  OAI211D0BWP12T U2978 ( .A1(n2323), .A2(n2322), .B(n2321), .C(n2320), .ZN(
        n2357) );
  AOI22D0BWP12T U2979 ( .A1(n595), .A2(n2325), .B1(n2324), .B2(n2331), .ZN(
        n2329) );
  AOI22D0BWP12T U2980 ( .A1(n2336), .A2(n2327), .B1(n2326), .B2(n2334), .ZN(
        n2328) );
  AOI21D0BWP12T U2981 ( .A1(n2329), .A2(n2328), .B(n2375), .ZN(n2330) );
  AOI211D0BWP12T U2982 ( .A1(n2357), .A2(n2381), .B(n2330), .C(n2437), .ZN(
        n2342) );
  AOI22D0BWP12T U2983 ( .A1(n595), .A2(n2333), .B1(n2332), .B2(n2331), .ZN(
        n2339) );
  AOI22D0BWP12T U2984 ( .A1(n2337), .A2(n2336), .B1(n2335), .B2(n2334), .ZN(
        n2338) );
  ND2D1BWP12T U2985 ( .A1(n2339), .A2(n2338), .ZN(n2382) );
  TPND2D0BWP12T U2986 ( .A1(n2382), .A2(n2340), .ZN(n2341) );
  OAI211D0BWP12T U2987 ( .A1(n2774), .A2(n2343), .B(n2342), .C(n2341), .ZN(
        n2605) );
  INVD0BWP12T U2988 ( .I(n2345), .ZN(n2346) );
  OAI22D0BWP12T U2989 ( .A1(n2808), .A2(n2431), .B1(n2346), .B2(n2375), .ZN(
        n2347) );
  AOI211XD0BWP12T U2990 ( .A1(n2407), .A2(n2348), .B(n2347), .C(n2359), .ZN(
        n2975) );
  CKND2D0BWP12T U2991 ( .A1(n2350), .A2(n2349), .ZN(n2373) );
  AOI22D0BWP12T U2992 ( .A1(n2388), .A2(n2352), .B1(n2351), .B2(n2407), .ZN(
        n2353) );
  INVD1BWP12T U2993 ( .I(n2359), .ZN(n2390) );
  OAI211D0BWP12T U2994 ( .A1(n2907), .A2(n2431), .B(n2353), .C(n2390), .ZN(
        n2902) );
  OAI211D0BWP12T U2995 ( .A1(n2373), .A2(n2448), .B(n2902), .C(n3040), .ZN(
        n2354) );
  NR4D0BWP12T U2996 ( .A1(n2356), .A2(n2975), .A3(n2355), .A4(n2354), .ZN(
        n2371) );
  INVD0BWP12T U2997 ( .I(n2357), .ZN(n2358) );
  OAI22D0BWP12T U2998 ( .A1(n2358), .A2(n2375), .B1(n2774), .B2(n2431), .ZN(
        n2360) );
  RCAOI211D0BWP12T U2999 ( .A1(n2407), .A2(n2382), .B(n2360), .C(n2359), .ZN(
        n3009) );
  AOI22D0BWP12T U3000 ( .A1(n2388), .A2(n2362), .B1(n2361), .B2(n2407), .ZN(
        n2363) );
  OA211D0BWP12T U3001 ( .A1(n2747), .A2(n2431), .B(n2363), .C(n2390), .Z(n2933) );
  ND3D1BWP12T U3002 ( .A1(n2364), .A2(n2452), .A3(n2349), .ZN(n2367) );
  AOI222D1BWP12T U3003 ( .A1(n2367), .A2(n2448), .B1(n2366), .B2(n2381), .C1(
        n2365), .C2(n2388), .ZN(n2664) );
  NR4D0BWP12T U3004 ( .A1(n3009), .A2(n2933), .A3(n2368), .A4(n2664), .ZN(
        n2370) );
  IND4D0BWP12T U3005 ( .A1(n2372), .B1(n2371), .B2(n2370), .B3(n2369), .ZN(
        n2397) );
  INVD1BWP12T U3006 ( .I(n2373), .ZN(n2374) );
  AOI21D1BWP12T U3007 ( .A1(n2452), .A2(n2374), .B(n2459), .ZN(n2379) );
  NR3D0BWP12T U3008 ( .A1(n2377), .A2(n2376), .A3(n2375), .ZN(n2378) );
  AOI211D1BWP12T U3009 ( .A1(n2381), .A2(n2380), .B(n2379), .C(n2378), .ZN(
        n2693) );
  INVD1BWP12T U3010 ( .I(n2382), .ZN(n2383) );
  MUX2ND0BWP12T U3011 ( .I0(n2383), .I1(n2774), .S(n2407), .ZN(n2384) );
  NR2XD0BWP12T U3012 ( .A1(n2384), .A2(n2448), .ZN(n3041) );
  NR4D0BWP12T U3013 ( .A1(n2693), .A2(n3041), .A3(n2386), .A4(n2385), .ZN(
        n2393) );
  ND4D0BWP12T U3014 ( .A1(n2393), .A2(n2392), .A3(n2634), .A4(n2391), .ZN(
        n2396) );
  NR4D0BWP12T U3015 ( .A1(n2397), .A2(n2396), .A3(n2395), .A4(n2394), .ZN(
        n2428) );
  AOI22D1BWP12T U3016 ( .A1(n2501), .A2(n2398), .B1(n2807), .B2(n2799), .ZN(
        n2402) );
  AOI22D0BWP12T U3017 ( .A1(n2956), .A2(b[31]), .B1(n2829), .B2(a[7]), .ZN(
        n2401) );
  AOI22D0BWP12T U3018 ( .A1(b[13]), .A2(n3033), .B1(n2522), .B2(a[14]), .ZN(
        n2400) );
  AOI22D0BWP12T U3019 ( .A1(n2880), .A2(n2874), .B1(n3074), .B2(n3067), .ZN(
        n2399) );
  ND4D1BWP12T U3020 ( .A1(n2402), .A2(n2401), .A3(n2400), .A4(n2399), .ZN(
        n2426) );
  AOI22D0BWP12T U3021 ( .A1(b[26]), .A2(a[26]), .B1(n3102), .B2(n3110), .ZN(
        n2411) );
  AOI22D0BWP12T U3022 ( .A1(b[24]), .A2(n2403), .B1(b[25]), .B2(n2502), .ZN(
        n2410) );
  AOI22D0BWP12T U3023 ( .A1(n2766), .A2(n2764), .B1(n2750), .B2(n2748), .ZN(
        n2409) );
  AOI22D0BWP12T U3024 ( .A1(n2407), .A2(n2406), .B1(n2405), .B2(n2404), .ZN(
        n2408) );
  ND4D1BWP12T U3025 ( .A1(n2411), .A2(n2410), .A3(n2409), .A4(n2408), .ZN(
        n2425) );
  AOI22D0BWP12T U3026 ( .A1(b[21]), .A2(n2993), .B1(b[20]), .B2(a[20]), .ZN(
        n2415) );
  AOI22D0BWP12T U3027 ( .A1(b[22]), .A2(n2963), .B1(b[30]), .B2(a[30]), .ZN(
        n2414) );
  AOI22D0BWP12T U3028 ( .A1(b[27]), .A2(n2518), .B1(b[29]), .B2(n2608), .ZN(
        n2413) );
  AOI22D0BWP12T U3029 ( .A1(b[28]), .A2(a[28]), .B1(b[23]), .B2(n2633), .ZN(
        n2412) );
  ND4D1BWP12T U3030 ( .A1(n2415), .A2(n2414), .A3(n2413), .A4(n2412), .ZN(
        n2424) );
  AOI22D0BWP12T U3031 ( .A1(n2489), .A2(n2416), .B1(b[15]), .B2(n2720), .ZN(
        n2419) );
  AOI22D0BWP12T U3032 ( .A1(b[18]), .A2(n2689), .B1(b[16]), .B2(n2891), .ZN(
        n2418) );
  AOI22D0BWP12T U3033 ( .A1(n2663), .A2(n2657), .B1(b[17]), .B2(n2560), .ZN(
        n2417) );
  TPND3D0BWP12T U3034 ( .A1(n2419), .A2(n2418), .A3(n2417), .ZN(n2420) );
  AOI211D0BWP12T U3035 ( .A1(n2857), .A2(n2851), .B(n2994), .C(n2420), .ZN(
        n2421) );
  OAI21D0BWP12T U3036 ( .A1(n2422), .A2(n2486), .B(n2421), .ZN(n2423) );
  NR4D0BWP12T U3037 ( .A1(n2426), .A2(n2425), .A3(n2424), .A4(n2423), .ZN(
        n2427) );
  AOI211XD0BWP12T U3038 ( .A1(n2430), .A2(n2429), .B(n2428), .C(n2427), .ZN(
        n2466) );
  NR2D0BWP12T U3039 ( .A1(n2432), .A2(n2431), .ZN(n2718) );
  OAI31D1BWP12T U3040 ( .A1(n2434), .A2(n2718), .A3(n2433), .B(n2452), .ZN(
        n2464) );
  ND2D1BWP12T U3041 ( .A1(n2454), .A2(n2452), .ZN(n2436) );
  AOI21D0BWP12T U3042 ( .A1(n2436), .A2(n2448), .B(n2435), .ZN(n2849) );
  INVD1BWP12T U3043 ( .I(n2798), .ZN(n2971) );
  AOI211D1BWP12T U3044 ( .A1(n2750), .A2(n2971), .B(n2812), .C(n2437), .ZN(
        n2797) );
  OR4D0BWP12T U3045 ( .A1(n3089), .A2(n2849), .A3(n2797), .A4(n2438), .Z(n2445) );
  ND2D1BWP12T U3046 ( .A1(n3061), .A2(n2452), .ZN(n2439) );
  AOI21D1BWP12T U3047 ( .A1(n2439), .A2(n2448), .B(n3082), .ZN(n3053) );
  INVD1BWP12T U3048 ( .I(n2440), .ZN(n2784) );
  INVD1BWP12T U3049 ( .I(n2441), .ZN(n2783) );
  CKND2D1BWP12T U3050 ( .A1(n2453), .A2(n2750), .ZN(n3088) );
  CKND2D0BWP12T U3051 ( .A1(n3092), .A2(n3088), .ZN(n2443) );
  OAI211D0BWP12T U3052 ( .A1(n2784), .A2(n2783), .B(n2443), .C(n2442), .ZN(
        n2444) );
  NR4D0BWP12T U3053 ( .A1(n2445), .A2(n3053), .A3(n2444), .A4(n2844), .ZN(
        n2463) );
  CKND2D0BWP12T U3054 ( .A1(n2446), .A2(n3037), .ZN(n2451) );
  ND2D1BWP12T U3055 ( .A1(n2447), .A2(n2452), .ZN(n2449) );
  AOI21D1BWP12T U3056 ( .A1(n2449), .A2(n2448), .B(n2751), .ZN(n2746) );
  AOI211D1BWP12T U3057 ( .A1(n2452), .A2(n2451), .B(n2450), .C(n2746), .ZN(
        n2462) );
  INVD1BWP12T U3058 ( .I(n2455), .ZN(n2696) );
  ND4D1BWP12T U3059 ( .A1(n2464), .A2(n2463), .A3(n2462), .A4(n2461), .ZN(
        n2465) );
  OAI211D1BWP12T U3060 ( .A1(n2468), .A2(n2467), .B(n2466), .C(n2465), .ZN(
        n2469) );
  AOI211D1BWP12T U3061 ( .A1(n2471), .A2(n2486), .B(n2470), .C(n2469), .ZN(
        n2472) );
  OAI31D0BWP12T U3062 ( .A1(n2475), .A2(n2474), .A3(n2473), .B(n2472), .ZN(
        n2476) );
  AOI211D1BWP12T U3063 ( .A1(n2479), .A2(n2478), .B(n2477), .C(n2476), .ZN(
        n2480) );
  OAI211D1BWP12T U3064 ( .A1(n2483), .A2(n2482), .B(n2481), .C(n2480), .ZN(z)
         );
  FA1D1BWP12T U3065 ( .A(mult_x_18_n404), .B(mult_x_18_n382), .CI(n2484), .CO(
        n2586), .S(n2587) );
  AO21D0BWP12T U3066 ( .A1(n2487), .A2(n2486), .B(n2485), .Z(n2488) );
  CKXOR2D1BWP12T U3067 ( .A1(mult_x_18_n398), .A2(n2488), .Z(n2510) );
  XNR2XD0BWP12T U3068 ( .A1(n2993), .A2(n2489), .ZN(n2490) );
  OAI22D0BWP12T U3069 ( .A1(n2493), .A2(n2492), .B1(n2491), .B2(n2490), .ZN(
        n2500) );
  XNR2D0BWP12T U3070 ( .A1(n2494), .A2(b[22]), .ZN(n2496) );
  OAI22D0BWP12T U3071 ( .A1(n2498), .A2(n2497), .B1(n2496), .B2(n2495), .ZN(
        n2499) );
  XOR2XD1BWP12T U3072 ( .A1(n2500), .A2(n2499), .Z(n2508) );
  XNR2XD0BWP12T U3073 ( .A1(n2502), .A2(n2501), .ZN(n2503) );
  OAI22D0BWP12T U3074 ( .A1(n2506), .A2(n2505), .B1(n2504), .B2(n2503), .ZN(
        n2507) );
  XOR2XD1BWP12T U3075 ( .A1(n2508), .A2(n2507), .Z(n2509) );
  XOR2XD1BWP12T U3076 ( .A1(n2510), .A2(n2509), .Z(n2511) );
  XOR2XD1BWP12T U3077 ( .A1(mult_x_18_n386), .A2(n2511), .Z(n2527) );
  XOR2XD1BWP12T U3078 ( .A1(n2527), .A2(n2526), .Z(n2528) );
  XOR2XD1BWP12T U3079 ( .A1(mult_x_18_n380), .A2(n2528), .Z(n2583) );
  XOR2XD1BWP12T U3080 ( .A1(mult_x_18_n384), .A2(mult_x_18_n387), .Z(n2581) );
  HA1D0BWP12T U3081 ( .A(n2530), .B(n2529), .CO(n2531), .S(mult_x_18_n402) );
  XOR2XD1BWP12T U3082 ( .A1(mult_x_18_n390), .A2(mult_x_18_n399), .Z(n2577) );
  XNR2XD0BWP12T U3083 ( .A1(n2542), .A2(n2608), .ZN(n2544) );
  OAI22D0BWP12T U3084 ( .A1(n2546), .A2(n2545), .B1(n2544), .B2(n2543), .ZN(
        n2553) );
  XNR2XD0BWP12T U3085 ( .A1(n2547), .A2(n2956), .ZN(n2549) );
  OAI22D0BWP12T U3086 ( .A1(n2551), .A2(n2550), .B1(n2549), .B2(n2548), .ZN(
        n2552) );
  XNR2D1BWP12T U3087 ( .A1(n2553), .A2(n2552), .ZN(n2554) );
  XOR2XD1BWP12T U3088 ( .A1(mult_x_18_n389), .A2(n2554), .Z(n2575) );
  XNR2XD0BWP12T U3089 ( .A1(n2555), .A2(b[26]), .ZN(n2556) );
  OAI22D0BWP12T U3090 ( .A1(n2559), .A2(n2558), .B1(n2557), .B2(n2556), .ZN(
        n2566) );
  XNR2XD0BWP12T U3091 ( .A1(n2560), .A2(b[16]), .ZN(n2562) );
  OAI22D0BWP12T U3092 ( .A1(n2564), .A2(n2563), .B1(n2562), .B2(n2561), .ZN(
        n2565) );
  XOR2XD1BWP12T U3093 ( .A1(n2566), .A2(n2565), .Z(n2573) );
  XNR2XD0BWP12T U3094 ( .A1(n2567), .A2(b[30]), .ZN(n2568) );
  OAI22D0BWP12T U3095 ( .A1(n2571), .A2(n2570), .B1(n2569), .B2(n2568), .ZN(
        n2572) );
  XOR2XD1BWP12T U3096 ( .A1(n2573), .A2(n2572), .Z(n2574) );
  XOR2XD1BWP12T U3097 ( .A1(n2575), .A2(n2574), .Z(n2576) );
  CKXOR2D1BWP12T U3098 ( .A1(n2577), .A2(n2576), .Z(n2578) );
  XOR2XD1BWP12T U3099 ( .A1(n2579), .A2(n2578), .Z(n2580) );
  XOR2XD1BWP12T U3100 ( .A1(n2581), .A2(n2580), .Z(n2582) );
  XOR2XD1BWP12T U3101 ( .A1(n2583), .A2(n2582), .Z(n2584) );
  CKXOR2D1BWP12T U3102 ( .A1(n2584), .A2(mult_x_18_n381), .Z(n2585) );
  XOR2XD1BWP12T U3103 ( .A1(n2586), .A2(n2585), .Z(n2960) );
  CKXOR2D0BWP12T U3104 ( .A1(n2960), .A2(n2587), .Z(n2600) );
  CKND2D0BWP12T U3105 ( .A1(n3020), .A2(n3059), .ZN(n2592) );
  FA1D2BWP12T U3106 ( .A(n2305), .B(b[31]), .CI(n2588), .CO(n2589), .S(n2483)
         );
  FA1D2BWP12T U3107 ( .A(n2305), .B(b[31]), .CI(n2590), .CO(n2591), .S(n1832)
         );
  MUX2NXD0BWP12T U3108 ( .I0(n2592), .I1(n2958), .S(n2956), .ZN(n2594) );
  NR2D1BWP12T U3109 ( .A1(n2594), .A2(n2593), .ZN(n2599) );
  NR2D0BWP12T U3110 ( .A1(n2595), .A2(n2956), .ZN(n2959) );
  XNR2XD1BWP12T U3111 ( .A1(n2959), .A2(n2596), .ZN(n2597) );
  NR2D0BWP12T U3112 ( .A1(n2597), .A2(n2980), .ZN(n2598) );
  AO211D1BWP12T U3113 ( .A1(n2600), .A2(n3126), .B(n2599), .C(n2598), .Z(v) );
  INVD1BWP12T U3114 ( .I(n2601), .ZN(n2627) );
  CKND2D1BWP12T U3115 ( .A1(n2602), .A2(n3098), .ZN(n2621) );
  ND2D1BWP12T U3116 ( .A1(n2603), .A2(n3119), .ZN(n2620) );
  MOAI22D0BWP12T U3117 ( .A1(n2605), .A2(n2903), .B1(n2604), .B2(n3130), .ZN(
        n2615) );
  OAI21D0BWP12T U3118 ( .A1(n2608), .A2(n3066), .B(n3105), .ZN(n2606) );
  AOI22D0BWP12T U3119 ( .A1(n3070), .A2(n2607), .B1(n2606), .B2(b[29]), .ZN(
        n2611) );
  MUX2ND0BWP12T U3120 ( .I0(n2995), .I1(n2994), .S(b[29]), .ZN(n2609) );
  OAI21D0BWP12T U3121 ( .A1(n2609), .A2(n2996), .B(n2608), .ZN(n2610) );
  OAI211D1BWP12T U3122 ( .A1(n2613), .A2(n2612), .B(n2611), .C(n2610), .ZN(
        n2614) );
  RCAOI211D0BWP12T U3123 ( .A1(n3091), .A2(n2616), .B(n2615), .C(n2614), .ZN(
        n2619) );
  ND2D1BWP12T U3124 ( .A1(n2617), .A2(n3115), .ZN(n2618) );
  ND4D1BWP12T U3125 ( .A1(n2621), .A2(n2620), .A3(n2619), .A4(n2618), .ZN(
        n2622) );
  AOI21D1BWP12T U3126 ( .A1(n314), .A2(n2623), .B(n2622), .ZN(n2626) );
  ND2D1BWP12T U3127 ( .A1(n2624), .A2(n3095), .ZN(n2625) );
  OAI211D1BWP12T U3128 ( .A1(n2951), .A2(n2627), .B(n2626), .C(n2625), .ZN(
        result[29]) );
  INVD1BWP12T U3129 ( .I(n2628), .ZN(n2653) );
  INVD1BWP12T U3130 ( .I(n2629), .ZN(n2647) );
  CKND2D1BWP12T U3131 ( .A1(n2630), .A2(n3119), .ZN(n2646) );
  MAOI22D0BWP12T U3132 ( .A1(n3130), .A2(n2632), .B1(n2631), .B2(n3012), .ZN(
        n2642) );
  OAI21D0BWP12T U3133 ( .A1(n2633), .A2(n3066), .B(n3105), .ZN(n2640) );
  NR2D1BWP12T U3134 ( .A1(n2634), .A2(n2903), .ZN(n2639) );
  MUX2ND0BWP12T U3135 ( .I0(n2995), .I1(n2994), .S(b[23]), .ZN(n2635) );
  NR2D0BWP12T U3136 ( .A1(n2635), .A2(n2996), .ZN(n2637) );
  MUX2ND0BWP12T U3137 ( .I0(n2637), .I1(n3109), .S(n2636), .ZN(n2638) );
  AOI211D0BWP12T U3138 ( .A1(b[23]), .A2(n2640), .B(n2639), .C(n2638), .ZN(
        n2641) );
  OAI211D1BWP12T U3139 ( .A1(n2822), .A2(n3004), .B(n2642), .C(n2641), .ZN(
        n2643) );
  AOI21D1BWP12T U3140 ( .A1(n2644), .A2(n3115), .B(n2643), .ZN(n2645) );
  OAI211D1BWP12T U3141 ( .A1(n2647), .A2(n2943), .B(n2646), .C(n2645), .ZN(
        n2648) );
  AOI21D1BWP12T U3142 ( .A1(n314), .A2(n2649), .B(n2648), .ZN(n2652) );
  CKND2D1BWP12T U3143 ( .A1(n2650), .A2(n3095), .ZN(n2651) );
  OAI211D1BWP12T U3144 ( .A1(n2951), .A2(n2653), .B(n2652), .C(n2651), .ZN(
        result[23]) );
  INVD1BWP12T U3145 ( .I(n2654), .ZN(n2681) );
  INVD1BWP12T U3146 ( .I(n2655), .ZN(n2675) );
  CKND2D1BWP12T U3147 ( .A1(n2656), .A2(n3119), .ZN(n2674) );
  OAI21D0BWP12T U3148 ( .A1(n2657), .A2(n3066), .B(n3105), .ZN(n2662) );
  INVD1BWP12T U3149 ( .I(n2970), .ZN(n3001) );
  MUX2ND0BWP12T U3150 ( .I0(n2995), .I1(n2994), .S(n2663), .ZN(n2658) );
  NR2D0BWP12T U3151 ( .A1(n2658), .A2(n2996), .ZN(n2660) );
  MUX2ND0BWP12T U3152 ( .I0(n2660), .I1(n3109), .S(n2659), .ZN(n2661) );
  RCAOI211D0BWP12T U3153 ( .A1(n2663), .A2(n2662), .B(n3001), .C(n2661), .ZN(
        n2666) );
  CKND2D1BWP12T U3154 ( .A1(n2664), .A2(n3040), .ZN(n2665) );
  OAI211D1BWP12T U3155 ( .A1(n3005), .A2(n2667), .B(n2666), .C(n2665), .ZN(
        n2671) );
  OAI22D1BWP12T U3156 ( .A1(n2669), .A2(n3012), .B1(n3004), .B2(n2668), .ZN(
        n2670) );
  AOI211D1BWP12T U3157 ( .A1(n2672), .A2(n3115), .B(n2671), .C(n2670), .ZN(
        n2673) );
  OAI211D1BWP12T U3158 ( .A1(n2675), .A2(n2943), .B(n2674), .C(n2673), .ZN(
        n2676) );
  AOI21D1BWP12T U3159 ( .A1(n3095), .A2(n2677), .B(n2676), .ZN(n2680) );
  CKND2D1BWP12T U3160 ( .A1(n2678), .A2(n314), .ZN(n2679) );
  OAI211D1BWP12T U3161 ( .A1(n2951), .A2(n2681), .B(n2680), .C(n2679), .ZN(
        result[19]) );
  INVD1BWP12T U3162 ( .I(n2682), .ZN(n2711) );
  INVD1BWP12T U3163 ( .I(n2683), .ZN(n2705) );
  CKND2D1BWP12T U3164 ( .A1(n2684), .A2(n3119), .ZN(n2704) );
  ND2D0BWP12T U3165 ( .A1(n2685), .A2(n3091), .ZN(n2695) );
  MUX2ND0BWP12T U3166 ( .I0(n2995), .I1(n2994), .S(b[18]), .ZN(n2686) );
  NR2D0BWP12T U3167 ( .A1(n2686), .A2(n2996), .ZN(n2688) );
  MUX2NXD0BWP12T U3168 ( .I0(n2688), .I1(n3109), .S(n2687), .ZN(n2692) );
  NR2D0BWP12T U3169 ( .A1(n2689), .A2(n3066), .ZN(n2690) );
  OA21XD0BWP12T U3170 ( .A1(n2690), .A2(n2996), .B(b[18]), .Z(n2691) );
  AOI211D1BWP12T U3171 ( .A1(n2693), .A2(n3040), .B(n2692), .C(n2691), .ZN(
        n2694) );
  OAI211D1BWP12T U3172 ( .A1(n2697), .A2(n2696), .B(n2695), .C(n2694), .ZN(
        n2701) );
  INVD1BWP12T U3173 ( .I(n2698), .ZN(n2699) );
  NR2D1BWP12T U3174 ( .A1(n2699), .A2(n3044), .ZN(n2700) );
  RCAOI211D0BWP12T U3175 ( .A1(n2702), .A2(n3115), .B(n2701), .C(n2700), .ZN(
        n2703) );
  OAI211D1BWP12T U3176 ( .A1(n2943), .A2(n2705), .B(n2704), .C(n2703), .ZN(
        n2706) );
  AOI21D1BWP12T U3177 ( .A1(n3095), .A2(n2707), .B(n2706), .ZN(n2710) );
  CKND2D1BWP12T U3178 ( .A1(n2708), .A2(n314), .ZN(n2709) );
  OAI211D1BWP12T U3179 ( .A1(n2951), .A2(n2711), .B(n2710), .C(n2709), .ZN(
        result[18]) );
  INVD1BWP12T U3180 ( .I(n2712), .ZN(n2738) );
  AO22XD1BWP12T U3181 ( .A1(n2714), .A2(n3098), .B1(n2713), .B2(n3119), .Z(
        n2733) );
  AOI22D0BWP12T U3182 ( .A1(n3115), .A2(n2716), .B1(n2715), .B2(n3091), .ZN(
        n2730) );
  OA21D1BWP12T U3183 ( .A1(n2719), .A2(n2718), .B(n2717), .Z(n2727) );
  OAI21D0BWP12T U3184 ( .A1(n2720), .A2(n3066), .B(n3105), .ZN(n2725) );
  MUX2ND0BWP12T U3185 ( .I0(n3104), .I1(n3103), .S(b[15]), .ZN(n2721) );
  ND2XD0BWP12T U3186 ( .A1(n2721), .A2(n3105), .ZN(n2723) );
  MUX2ND0BWP12T U3187 ( .I0(n2723), .I1(n3070), .S(n2722), .ZN(n2724) );
  IOA21D1BWP12T U3188 ( .A1(b[15]), .A2(n2725), .B(n2724), .ZN(n2726) );
  RCAOI211D0BWP12T U3189 ( .A1(n3040), .A2(n2728), .B(n2727), .C(n2726), .ZN(
        n2729) );
  OAI211D1BWP12T U3190 ( .A1(n2731), .A2(n3044), .B(n2730), .C(n2729), .ZN(
        n2732) );
  AOI211D1BWP12T U3191 ( .A1(n3095), .A2(n2734), .B(n2733), .C(n2732), .ZN(
        n2737) );
  CKND2D1BWP12T U3192 ( .A1(n2735), .A2(n314), .ZN(n2736) );
  OAI211D1BWP12T U3193 ( .A1(n2951), .A2(n2738), .B(n2737), .C(n2736), .ZN(
        result[15]) );
  CKND2D0BWP12T U3194 ( .A1(n2739), .A2(n3095), .ZN(n2743) );
  AOI22D0BWP12T U3195 ( .A1(n2741), .A2(n3098), .B1(n2740), .B2(n3119), .ZN(
        n2742) );
  OAI211D1BWP12T U3196 ( .A1(n2744), .A2(n3012), .B(n2743), .C(n2742), .ZN(
        n2745) );
  AOI21D1BWP12T U3197 ( .A1(n3052), .A2(n2746), .B(n2745), .ZN(n2756) );
  NR2D0BWP12T U3198 ( .A1(n233), .A2(n3020), .ZN(n2753) );
  INVD1BWP12T U3199 ( .I(n3060), .ZN(n3100) );
  AOI211D1BWP12T U3200 ( .A1(n2754), .A2(n3115), .B(n2753), .C(n2752), .ZN(
        n2755) );
  OAI211D1BWP12T U3201 ( .A1(n2757), .A2(n3044), .B(n2756), .C(n2755), .ZN(
        n2758) );
  AO21D1BWP12T U3202 ( .A1(n2759), .A2(n3126), .B(n2758), .Z(result[4]) );
  INVD1BWP12T U3203 ( .I(n2760), .ZN(n2790) );
  MAOI22D0BWP12T U3204 ( .A1(n2762), .A2(n3115), .B1(n2761), .B2(n3044), .ZN(
        n2789) );
  INVD1BWP12T U3205 ( .I(n2763), .ZN(n2780) );
  OAI21D0BWP12T U3206 ( .A1(n2764), .A2(n3066), .B(n3105), .ZN(n2765) );
  CKND2D0BWP12T U3207 ( .A1(n2765), .A2(n2766), .ZN(n2771) );
  MUX2ND0BWP12T U3208 ( .I0(n3104), .I1(n3103), .S(n2766), .ZN(n2767) );
  CKND2D0BWP12T U3209 ( .A1(n2767), .A2(n3105), .ZN(n2769) );
  MUX2ND0BWP12T U3210 ( .I0(n2769), .I1(n3070), .S(n2768), .ZN(n2770) );
  OAI211D1BWP12T U3211 ( .A1(n2836), .A2(n2772), .B(n2771), .C(n2770), .ZN(
        n2773) );
  RCAOI21D0BWP12T U3212 ( .A1(n3094), .A2(n2774), .B(n2773), .ZN(n2779) );
  OAI21D0BWP12T U3213 ( .A1(n3003), .A2(n3012), .B(n3100), .ZN(n2775) );
  AOI22D0BWP12T U3214 ( .A1(n2777), .A2(n3119), .B1(n2776), .B2(n2775), .ZN(
        n2778) );
  OAI211D0BWP12T U3215 ( .A1(n3020), .A2(n2780), .B(n2779), .C(n2778), .ZN(
        n2786) );
  CKND2D0BWP12T U3216 ( .A1(n2781), .A2(n3098), .ZN(n2782) );
  TPOAI31D0BWP12T U3217 ( .A1(n2784), .A2(n2783), .A3(n3089), .B(n2782), .ZN(
        n2785) );
  AOI211D1BWP12T U3218 ( .A1(n3095), .A2(n2787), .B(n2786), .C(n2785), .ZN(
        n2788) );
  OAI211D1BWP12T U3219 ( .A1(n2951), .A2(n2790), .B(n2789), .C(n2788), .ZN(
        result[5]) );
  CKND2D1BWP12T U3220 ( .A1(n2791), .A2(n3126), .ZN(n2820) );
  AOI22D0BWP12T U3221 ( .A1(n3115), .A2(n2793), .B1(n2792), .B2(n314), .ZN(
        n2819) );
  AOI22D0BWP12T U3222 ( .A1(n3098), .A2(n2795), .B1(n2794), .B2(n3119), .ZN(
        n2796) );
  IOA21D1BWP12T U3223 ( .A1(n2797), .A2(n3052), .B(n2796), .ZN(n2814) );
  AOI21D0BWP12T U3224 ( .A1(n2798), .A2(n3091), .B(n3060), .ZN(n2811) );
  OAI21D1BWP12T U3225 ( .A1(n2799), .A2(n3066), .B(n3105), .ZN(n2806) );
  NR2D1BWP12T U3226 ( .A1(n2800), .A2(n2836), .ZN(n2805) );
  MUX2ND0BWP12T U3227 ( .I0(n2995), .I1(n2994), .S(n2807), .ZN(n2801) );
  NR2D0BWP12T U3228 ( .A1(n2801), .A2(n2996), .ZN(n2803) );
  MUX2NXD0BWP12T U3229 ( .I0(n2803), .I1(n3109), .S(n2802), .ZN(n2804) );
  AOI211D1BWP12T U3230 ( .A1(n2807), .A2(n2806), .B(n2805), .C(n2804), .ZN(
        n2810) );
  CKND2D1BWP12T U3231 ( .A1(n3094), .A2(n2808), .ZN(n2809) );
  OAI211D1BWP12T U3232 ( .A1(n2812), .A2(n2811), .B(n2810), .C(n2809), .ZN(
        n2813) );
  AOI211D1BWP12T U3233 ( .A1(n3095), .A2(n2815), .B(n2814), .C(n2813), .ZN(
        n2818) );
  ND2XD0BWP12T U3234 ( .A1(n2816), .A2(n3130), .ZN(n2817) );
  ND4D1BWP12T U3235 ( .A1(n2820), .A2(n2819), .A3(n2818), .A4(n2817), .ZN(
        result[6]) );
  INVD1BWP12T U3236 ( .I(n2827), .ZN(n2842) );
  OAI21D0BWP12T U3237 ( .A1(a[7]), .A2(n3066), .B(n3105), .ZN(n2828) );
  CKND2D0BWP12T U3238 ( .A1(n2828), .A2(n2829), .ZN(n2834) );
  MUX2ND0BWP12T U3239 ( .I0(n3104), .I1(n3103), .S(n2829), .ZN(n2830) );
  CKND2D0BWP12T U3240 ( .A1(n2830), .A2(n3105), .ZN(n2832) );
  MUX2NXD0BWP12T U3241 ( .I0(n2832), .I1(n3070), .S(n2831), .ZN(n2833) );
  OAI211D1BWP12T U3242 ( .A1(n2836), .A2(n2835), .B(n2834), .C(n2833), .ZN(
        n2837) );
  AOI21D1BWP12T U3243 ( .A1(n2838), .A2(n3094), .B(n2837), .ZN(n2841) );
  CKND2D0BWP12T U3244 ( .A1(n2839), .A2(n3119), .ZN(n2840) );
  AOI22D0BWP12T U3245 ( .A1(n2850), .A2(n3119), .B1(n3052), .B2(n2849), .ZN(
        n2859) );
  OAI21D0BWP12T U3246 ( .A1(n2851), .A2(n3066), .B(n3105), .ZN(n2856) );
  MUX2ND0BWP12T U3247 ( .I0(n2995), .I1(n2994), .S(n2857), .ZN(n2852) );
  NR2D0BWP12T U3248 ( .A1(n2852), .A2(n2996), .ZN(n2854) );
  MUX2ND0BWP12T U3249 ( .I0(n2854), .I1(n3109), .S(n2853), .ZN(n2855) );
  RCAOI21D0BWP12T U3250 ( .A1(n2857), .A2(n2856), .B(n2855), .ZN(n2858) );
  OAI211D1BWP12T U3251 ( .A1(n2861), .A2(n2860), .B(n2859), .C(n2858), .ZN(
        n2862) );
  CKND2D0BWP12T U3252 ( .A1(n2868), .A2(n3091), .ZN(n3064) );
  OAI22D1BWP12T U3253 ( .A1(n2871), .A2(n2870), .B1(n2869), .B2(n3064), .ZN(
        n2872) );
  OAI21D0BWP12T U3254 ( .A1(n2874), .A2(n3066), .B(n3105), .ZN(n2879) );
  MUX2ND0BWP12T U3255 ( .I0(n2995), .I1(n2994), .S(n2880), .ZN(n2875) );
  NR2D0BWP12T U3256 ( .A1(n2875), .A2(n2996), .ZN(n2877) );
  MUX2NXD0BWP12T U3257 ( .I0(n2877), .I1(n3109), .S(n2876), .ZN(n2878) );
  RCAOI21D0BWP12T U3258 ( .A1(n2880), .A2(n2879), .B(n2878), .ZN(n2883) );
  CKND2D1BWP12T U3259 ( .A1(n2881), .A2(n3078), .ZN(n2882) );
  OAI211D1BWP12T U3260 ( .A1(n3044), .A2(n2884), .B(n2883), .C(n2882), .ZN(
        n2885) );
  INVD1BWP12T U3261 ( .I(n2889), .ZN(n2922) );
  CKND2D1BWP12T U3262 ( .A1(n2890), .A2(n3119), .ZN(n2915) );
  OAI21D0BWP12T U3263 ( .A1(n2891), .A2(n3066), .B(n3105), .ZN(n2896) );
  MUX2ND0BWP12T U3264 ( .I0(n2995), .I1(n2994), .S(b[16]), .ZN(n2892) );
  NR2D0BWP12T U3265 ( .A1(n2892), .A2(n2996), .ZN(n2894) );
  MUX2ND0BWP12T U3266 ( .I0(n2894), .I1(n3109), .S(n2893), .ZN(n2895) );
  RCAOI211D0BWP12T U3267 ( .A1(b[16]), .A2(n2896), .B(n3001), .C(n2895), .ZN(
        n2901) );
  INVD1BWP12T U3268 ( .I(n2897), .ZN(n2898) );
  ND2D1BWP12T U3269 ( .A1(n2899), .A2(n2898), .ZN(n2900) );
  OAI211D1BWP12T U3270 ( .A1(n2903), .A2(n2902), .B(n2901), .C(n2900), .ZN(
        n2912) );
  AOI222D1BWP12T U3271 ( .A1(n2909), .A2(n2908), .B1(n2907), .B2(n2906), .C1(
        n2905), .C2(n2904), .ZN(n2910) );
  NR2D1BWP12T U3272 ( .A1(n2910), .A2(n3012), .ZN(n2911) );
  RCAOI211D0BWP12T U3273 ( .A1(n2913), .A2(n3115), .B(n2912), .C(n2911), .ZN(
        n2914) );
  OAI211D1BWP12T U3274 ( .A1(n2916), .A2(n2943), .B(n2915), .C(n2914), .ZN(
        n2917) );
  AOI21D1BWP12T U3275 ( .A1(n3095), .A2(n2918), .B(n2917), .ZN(n2921) );
  CKND2D1BWP12T U3276 ( .A1(n2919), .A2(n314), .ZN(n2920) );
  OAI211D1BWP12T U3277 ( .A1(n2951), .A2(n2922), .B(n2921), .C(n2920), .ZN(
        result[16]) );
  INVD1BWP12T U3278 ( .I(n2923), .ZN(n2950) );
  INVD1BWP12T U3279 ( .I(n2924), .ZN(n2944) );
  CKND2D1BWP12T U3280 ( .A1(n2925), .A2(n3119), .ZN(n2942) );
  CKND2D0BWP12T U3281 ( .A1(n2926), .A2(n3091), .ZN(n2935) );
  MUX2ND0BWP12T U3282 ( .I0(n2995), .I1(n2994), .S(b[20]), .ZN(n2927) );
  NR2D0BWP12T U3283 ( .A1(n2927), .A2(n2996), .ZN(n2929) );
  MUX2ND0BWP12T U3284 ( .I0(n2929), .I1(n3109), .S(n2928), .ZN(n2932) );
  NR2D0BWP12T U3285 ( .A1(a[20]), .A2(n3066), .ZN(n2930) );
  OA21XD0BWP12T U3286 ( .A1(n2930), .A2(n2996), .B(b[20]), .Z(n2931) );
  RCAOI211D0BWP12T U3287 ( .A1(n2933), .A2(n3040), .B(n2932), .C(n2931), .ZN(
        n2934) );
  OAI211D1BWP12T U3288 ( .A1(n2936), .A2(n3004), .B(n2935), .C(n2934), .ZN(
        n2939) );
  NR2D1BWP12T U3289 ( .A1(n2937), .A2(n3044), .ZN(n2938) );
  AOI211XD0BWP12T U3290 ( .A1(n2940), .A2(n3115), .B(n2939), .C(n2938), .ZN(
        n2941) );
  OAI211D1BWP12T U3291 ( .A1(n2944), .A2(n2943), .B(n2942), .C(n2941), .ZN(
        n2945) );
  AOI21D1BWP12T U3292 ( .A1(n3095), .A2(n2946), .B(n2945), .ZN(n2949) );
  CKND2D1BWP12T U3293 ( .A1(n2947), .A2(n314), .ZN(n2948) );
  OAI211D1BWP12T U3294 ( .A1(n2951), .A2(n2950), .B(n2949), .C(n2948), .ZN(
        result[20]) );
  FA1D2BWP12T U3295 ( .A(n2305), .B(n2953), .CI(n2952), .CO(n2954), .S(n2473)
         );
  FA1D2BWP12T U3296 ( .A(n2956), .B(b[31]), .CI(n2955), .CO(n2957), .S(n1371)
         );
  INVD1BWP12T U3297 ( .I(n2961), .ZN(n2986) );
  INVD1BWP12T U3298 ( .I(n2962), .ZN(n2979) );
  OAI21D0BWP12T U3299 ( .A1(n2963), .A2(n3066), .B(n3105), .ZN(n2968) );
  MUX2ND0BWP12T U3300 ( .I0(n2995), .I1(n2994), .S(b[22]), .ZN(n2964) );
  NR2D0BWP12T U3301 ( .A1(n2964), .A2(n2996), .ZN(n2966) );
  MUX2ND0BWP12T U3302 ( .I0(n2966), .I1(n3109), .S(n2965), .ZN(n2967) );
  AOI21D0BWP12T U3303 ( .A1(b[22]), .A2(n2968), .B(n2967), .ZN(n2969) );
  OAI211D0BWP12T U3304 ( .A1(n2971), .A2(n3004), .B(n2970), .C(n2969), .ZN(
        n2974) );
  NR2D1BWP12T U3305 ( .A1(n2972), .A2(n3005), .ZN(n2973) );
  AOI211XD0BWP12T U3306 ( .A1(n3040), .A2(n2975), .B(n2974), .C(n2973), .ZN(
        n2978) );
  ND2XD0BWP12T U3307 ( .A1(n2976), .A2(n3091), .ZN(n2977) );
  OAI211D1BWP12T U3308 ( .A1(n2980), .A2(n2979), .B(n2978), .C(n2977), .ZN(
        n2981) );
  AOI21D1BWP12T U3309 ( .A1(n2982), .A2(n3119), .B(n2981), .ZN(n2985) );
  TPND2D0BWP12T U3310 ( .A1(n2983), .A2(n3098), .ZN(n2984) );
  OAI211D1BWP12T U3311 ( .A1(n3020), .A2(n2986), .B(n2985), .C(n2984), .ZN(
        n2987) );
  AOI21D1BWP12T U3312 ( .A1(n3095), .A2(n2988), .B(n2987), .ZN(n2989) );
  IOA21D1BWP12T U3313 ( .A1(n2990), .A2(n3126), .B(n2989), .ZN(result[22]) );
  INVD1BWP12T U3314 ( .I(n2991), .ZN(n3019) );
  CKND2D1BWP12T U3315 ( .A1(n2992), .A2(n3115), .ZN(n3011) );
  OAI21D0BWP12T U3316 ( .A1(n2993), .A2(n3066), .B(n3105), .ZN(n3002) );
  MUX2ND0BWP12T U3317 ( .I0(n2995), .I1(n2994), .S(b[21]), .ZN(n2997) );
  NR2D0BWP12T U3318 ( .A1(n2997), .A2(n2996), .ZN(n2999) );
  MUX2ND0BWP12T U3319 ( .I0(n2999), .I1(n3109), .S(n2998), .ZN(n3000) );
  AO211D0BWP12T U3320 ( .A1(b[21]), .A2(n3002), .B(n3001), .C(n3000), .Z(n3008) );
  OAI22D0BWP12T U3321 ( .A1(n3006), .A2(n3005), .B1(n3004), .B2(n3003), .ZN(
        n3007) );
  RCAOI211D0BWP12T U3322 ( .A1(n3040), .A2(n3009), .B(n3008), .C(n3007), .ZN(
        n3010) );
  OAI211D1BWP12T U3323 ( .A1(n3013), .A2(n3012), .B(n3011), .C(n3010), .ZN(
        n3014) );
  AOI21D1BWP12T U3324 ( .A1(n3015), .A2(n3119), .B(n3014), .ZN(n3018) );
  CKND2D1BWP12T U3325 ( .A1(n3016), .A2(n3098), .ZN(n3017) );
  OAI211D1BWP12T U3326 ( .A1(n3020), .A2(n3019), .B(n3018), .C(n3017), .ZN(
        n3021) );
  AOI21D1BWP12T U3327 ( .A1(n3095), .A2(n3022), .B(n3021), .ZN(n3023) );
  IOA21D1BWP12T U3328 ( .A1(n3024), .A2(n3126), .B(n3023), .ZN(result[21]) );
  AOI22D1BWP12T U3329 ( .A1(n3115), .A2(n3029), .B1(n3028), .B2(n3119), .ZN(
        n3043) );
  MUX2ND0BWP12T U3330 ( .I0(n3104), .I1(n3103), .S(b[13]), .ZN(n3030) );
  TPND2D0BWP12T U3331 ( .A1(n3030), .A2(n3105), .ZN(n3032) );
  MUX2ND0BWP12T U3332 ( .I0(n3032), .I1(n3070), .S(n3031), .ZN(n3036) );
  OAI21D0BWP12T U3333 ( .A1(n3033), .A2(n3066), .B(n3105), .ZN(n3034) );
  ND2XD0BWP12T U3334 ( .A1(n3034), .A2(b[13]), .ZN(n3035) );
  OAI211D1BWP12T U3335 ( .A1(n3038), .A2(n3037), .B(n3036), .C(n3035), .ZN(
        n3039) );
  TPAOI21D0BWP12T U3336 ( .A1(n3041), .A2(n3040), .B(n3039), .ZN(n3042) );
  OAI211D1BWP12T U3337 ( .A1(n3045), .A2(n3044), .B(n3043), .C(n3042), .ZN(
        n3046) );
  AOI211XD0BWP12T U3338 ( .A1(n3095), .A2(n3048), .B(n3047), .C(n3046), .ZN(
        n3049) );
  IOA21D1BWP12T U3339 ( .A1(n3050), .A2(n3126), .B(n3049), .ZN(result[13]) );
  INVD1BWP12T U3340 ( .I(n3051), .ZN(n3058) );
  AOI22D0BWP12T U3341 ( .A1(n3054), .A2(n3098), .B1(n3053), .B2(n3052), .ZN(
        n3057) );
  ND2XD0BWP12T U3342 ( .A1(n3055), .A2(n3130), .ZN(n3056) );
  OAI211D1BWP12T U3343 ( .A1(n3059), .A2(n3058), .B(n3057), .C(n3056), .ZN(
        n3084) );
  AOI21D0BWP12T U3344 ( .A1(n3061), .A2(n3091), .B(n3060), .ZN(n3081) );
  AOI22D1BWP12T U3345 ( .A1(n3115), .A2(n3063), .B1(n3062), .B2(n3119), .ZN(
        n3080) );
  NR2D1BWP12T U3346 ( .A1(n3065), .A2(n3064), .ZN(n3076) );
  OAI21D0BWP12T U3347 ( .A1(n3067), .A2(n3066), .B(n3105), .ZN(n3073) );
  MUX2ND0BWP12T U3348 ( .I0(n3104), .I1(n3103), .S(n3074), .ZN(n3068) );
  ND2XD0BWP12T U3349 ( .A1(n3068), .A2(n3105), .ZN(n3071) );
  MUX2ND0BWP12T U3350 ( .I0(n3071), .I1(n3070), .S(n3069), .ZN(n3072) );
  IOA21D1BWP12T U3351 ( .A1(n3074), .A2(n3073), .B(n3072), .ZN(n3075) );
  RCAOI211D0BWP12T U3352 ( .A1(n3078), .A2(n3077), .B(n3076), .C(n3075), .ZN(
        n3079) );
  OAI211D1BWP12T U3353 ( .A1(n3082), .A2(n3081), .B(n3080), .C(n3079), .ZN(
        n3083) );
  AOI211D1BWP12T U3354 ( .A1(n314), .A2(n3085), .B(n3084), .C(n3083), .ZN(
        n3086) );
  IOA21D1BWP12T U3355 ( .A1(n3087), .A2(n3126), .B(n3086), .ZN(result[10]) );
  AOI22D1BWP12T U3356 ( .A1(n3096), .A2(n3095), .B1(n3094), .B2(n3093), .ZN(
        n3123) );
  AOI22D0BWP12T U3357 ( .A1(n3099), .A2(n314), .B1(n3098), .B2(n3097), .ZN(
        n3122) );
  NR2D1BWP12T U3358 ( .A1(n3101), .A2(n3100), .ZN(n3118) );
  MUX2ND0BWP12T U3359 ( .I0(n3104), .I1(n3103), .S(n3102), .ZN(n3106) );
  AOI21D0BWP12T U3360 ( .A1(n3106), .A2(n3105), .B(n3108), .ZN(n3114) );
  AOI21D0BWP12T U3361 ( .A1(n3108), .A2(n3107), .B(n2996), .ZN(n3112) );
  OAI22D0BWP12T U3362 ( .A1(n3112), .A2(n3111), .B1(n3110), .B2(n3109), .ZN(
        n3113) );
  AO211D0BWP12T U3363 ( .A1(n3116), .A2(n3115), .B(n3114), .C(n3113), .Z(n3117) );
  AOI211XD0BWP12T U3364 ( .A1(n3120), .A2(n3119), .B(n3118), .C(n3117), .ZN(
        n3121) );
  ND4D1BWP12T U3365 ( .A1(n3124), .A2(n3123), .A3(n3122), .A4(n3121), .ZN(
        n3125) );
  AOI21D1BWP12T U3366 ( .A1(n3127), .A2(n3126), .B(n3125), .ZN(n3128) );
  IOA21D1BWP12T U3367 ( .A1(n3130), .A2(n3129), .B(n3128), .ZN(result[1]) );
  CMPE42D1BWP12T U3368 ( .A(mult_x_18_n533), .B(mult_x_18_n515), .C(
        mult_x_18_n530), .CIX(mult_x_18_n526), .D(mult_x_18_n512), .CO(
        mult_x_18_n508), .COX(mult_x_18_n507), .S(mult_x_18_n509) );
  CMPE42D1BWP12T U3369 ( .A(mult_x_18_n482), .B(mult_x_18_n457), .C(
        mult_x_18_n476), .CIX(mult_x_18_n454), .D(mult_x_18_n479), .CO(
        mult_x_18_n450), .COX(mult_x_18_n449), .S(mult_x_18_n451) );
  CMPE42D1BWP12T U3370 ( .A(mult_x_18_n499), .B(mult_x_18_n477), .C(
        mult_x_18_n496), .CIX(mult_x_18_n489), .D(mult_x_18_n493), .CO(
        mult_x_18_n470), .COX(mult_x_18_n469), .S(mult_x_18_n471) );
  CMPE42D1BWP12T U3371 ( .A(mult_x_18_n865), .B(mult_x_18_n886), .C(
        mult_x_18_n909), .CIX(mult_x_18_n675), .D(mult_x_18_n934), .CO(
        mult_x_18_n667), .COX(mult_x_18_n666), .S(mult_x_18_n668) );
  CMPE42D1BWP12T U3372 ( .A(mult_x_18_n551), .B(mult_x_18_n570), .C(
        mult_x_18_n567), .CIX(mult_x_18_n560), .D(mult_x_18_n564), .CO(
        mult_x_18_n544), .COX(mult_x_18_n543), .S(mult_x_18_n545) );
  CMPE42D1BWP12T U3373 ( .A(mult_x_18_n862), .B(mult_x_18_n843), .C(
        mult_x_18_n650), .CIX(mult_x_18_n647), .D(mult_x_18_n638), .CO(
        mult_x_18_n632), .COX(mult_x_18_n631), .S(mult_x_18_n633) );
  CMPE42D1BWP12T U3374 ( .A(mult_x_18_n601), .B(mult_x_18_n955), .C(
        mult_x_18_n605), .CIX(mult_x_18_n596), .D(mult_x_18_n599), .CO(
        mult_x_18_n592), .COX(mult_x_18_n591), .S(mult_x_18_n593) );
  CMPE42D1BWP12T U3375 ( .A(mult_x_18_n957), .B(mult_x_18_n882), .C(
        mult_x_18_n842), .CIX(mult_x_18_n627), .D(mult_x_18_n631), .CO(
        mult_x_18_n620), .COX(mult_x_18_n619), .S(mult_x_18_n621) );
  CMPE42D1BWP12T U3376 ( .A(mult_x_18_n800), .B(mult_x_18_n776), .C(
        mult_x_18_n832), .CIX(mult_x_18_n478), .D(mult_x_18_n851), .CO(
        mult_x_18_n459), .COX(mult_x_18_n458), .S(mult_x_18_n460) );
  CMPE42D1BWP12T U3377 ( .A(mult_x_18_n949), .B(mult_x_18_n778), .C(
        mult_x_18_n802), .CIX(mult_x_18_n513), .D(mult_x_18_n834), .CO(
        mult_x_18_n496), .COX(mult_x_18_n495), .S(mult_x_18_n497) );
  CMPE42D1BWP12T U3378 ( .A(mult_x_18_n791), .B(mult_x_18_n876), .C(
        mult_x_18_n951), .CIX(mult_x_18_n552), .D(mult_x_18_n539), .CO(
        mult_x_18_n530), .COX(mult_x_18_n529), .S(mult_x_18_n531) );
  CMPE42D1BWP12T U3379 ( .A(mult_x_18_n804), .B(mult_x_18_n780), .C(
        mult_x_18_n836), .CIX(mult_x_18_n549), .D(mult_x_18_n855), .CO(
        mult_x_18_n533), .COX(mult_x_18_n532), .S(mult_x_18_n534) );
  CMPE42D1BWP12T U3380 ( .A(mult_x_18_n921), .B(mult_x_18_n777), .C(
        mult_x_18_n977), .CIX(mult_x_18_n492), .D(mult_x_18_n485), .CO(
        mult_x_18_n482), .COX(mult_x_18_n481), .S(mult_x_18_n483) );
  CMPE42D1BWP12T U3381 ( .A(mult_x_18_n394), .B(mult_x_18_n397), .C(
        mult_x_18_n391), .CIX(mult_x_18_n406), .D(mult_x_18_n419), .CO(
        mult_x_18_n384), .COX(mult_x_18_n383), .S(mult_x_18_n385) );
  CMPE42D1BWP12T U3382 ( .A(mult_x_18_n437), .B(mult_x_18_n440), .C(
        mult_x_18_n434), .CIX(mult_x_18_n427), .D(mult_x_18_n430), .CO(
        mult_x_18_n407), .COX(mult_x_18_n406), .S(mult_x_18_n408) );
  CMPE42D1BWP12T U3383 ( .A(mult_x_18_n462), .B(mult_x_18_n435), .C(
        mult_x_18_n459), .CIX(mult_x_18_n453), .D(mult_x_18_n452), .CO(
        mult_x_18_n428), .COX(mult_x_18_n427), .S(mult_x_18_n429) );
  CMPE42D1BWP12T U3384 ( .A(mult_x_18_n514), .B(mult_x_18_n500), .C(
        mult_x_18_n517), .CIX(mult_x_18_n507), .D(mult_x_18_n494), .CO(
        mult_x_18_n490), .COX(mult_x_18_n489), .S(mult_x_18_n491) );
  CMPE42D1BWP12T U3385 ( .A(mult_x_18_n571), .B(mult_x_18_n793), .C(
        mult_x_18_n568), .CIX(mult_x_18_n582), .D(mult_x_18_n565), .CO(
        mult_x_18_n561), .COX(mult_x_18_n560), .S(mult_x_18_n562) );
  CMPE42D1BWP12T U3386 ( .A(mult_x_18_n740), .B(mult_x_18_n845), .C(
        mult_x_18_n864), .CIX(mult_x_18_n669), .D(mult_x_18_n908), .CO(
        mult_x_18_n656), .COX(mult_x_18_n655), .S(mult_x_18_n657) );
  CMPE42D1BWP12T U3387 ( .A(mult_x_18_n894), .B(mult_x_18_n814), .C(
        mult_x_18_n919), .CIX(mult_x_18_n455), .D(mult_x_18_n445), .CO(
        mult_x_18_n440), .COX(mult_x_18_n439), .S(mult_x_18_n441) );
  CMPE42D1BWP12T U3388 ( .A(mult_x_18_n902), .B(mult_x_18_n794), .C(
        mult_x_18_n927), .CIX(mult_x_18_n594), .D(mult_x_18_n587), .CO(
        mult_x_18_n582), .COX(mult_x_18_n581), .S(mult_x_18_n583) );
  CMPE42D1BWP12T U3389 ( .A(mult_x_18_n757), .B(mult_x_18_n773), .C(
        mult_x_18_n869), .CIX(mult_x_18_n421), .D(mult_x_18_n764), .CO(
        mult_x_18_n390), .COX(mult_x_18_n389), .S(mult_x_18_n391) );
  CMPE42D1BWP12T U3390 ( .A(mult_x_18_n849), .B(mult_x_18_n753), .C(
        mult_x_18_n893), .CIX(mult_x_18_n433), .D(mult_x_18_n918), .CO(
        mult_x_18_n419), .COX(mult_x_18_n418), .S(mult_x_18_n420) );
  CMPE42D1BWP12T U3391 ( .A(mult_x_18_n465), .B(mult_x_18_n872), .C(
        mult_x_18_n472), .CIX(mult_x_18_n460), .D(mult_x_18_n463), .CO(
        mult_x_18_n453), .COX(mult_x_18_n452), .S(mult_x_18_n454) );
  CMPE42D1BWP12T U3392 ( .A(mult_x_18_n1025), .B(mult_x_18_n890), .C(
        mult_x_18_n913), .CIX(mult_x_18_n707), .D(mult_x_18_n709), .CO(
        mult_x_18_n702), .COX(mult_x_18_n701), .S(mult_x_18_n703) );
  CMPE42D1BWP12T U3393 ( .A(mult_x_18_n937), .B(mult_x_18_n889), .C(
        mult_x_18_n993), .CIX(mult_x_18_n698), .D(mult_x_18_n697), .CO(
        mult_x_18_n694), .COX(mult_x_18_n693), .S(mult_x_18_n695) );
  CMPE42D1BWP12T U3394 ( .A(mult_x_18_n929), .B(mult_x_18_n881), .C(
        mult_x_18_n985), .CIX(mult_x_18_n619), .D(mult_x_18_n615), .CO(
        mult_x_18_n612), .COX(mult_x_18_n611), .S(mult_x_18_n613) );
  CMPE42D1BWP12T U3395 ( .A(mult_x_18_n1009), .B(mult_x_18_n762), .C(
        mult_x_18_n978), .CIX(mult_x_18_n519), .D(mult_x_18_n521), .CO(
        mult_x_18_n502), .COX(mult_x_18_n501), .S(mult_x_18_n503) );
  CMPE42D1BWP12T U3396 ( .A(mult_x_18_n833), .B(mult_x_18_n761), .C(
        mult_x_18_n852), .CIX(mult_x_18_n495), .D(mult_x_18_n896), .CO(
        mult_x_18_n479), .COX(mult_x_18_n478), .S(mult_x_18_n480) );
  CMPE42D1BWP12T U3397 ( .A(mult_x_18_n585), .B(mult_x_18_n600), .C(
        mult_x_18_n583), .CIX(mult_x_18_n591), .D(mult_x_18_n580), .CO(
        mult_x_18_n576), .COX(mult_x_18_n575), .S(mult_x_18_n577) );
  CMPE42D1BWP12T U3398 ( .A(mult_x_18_n1017), .B(mult_x_18_n810), .C(
        mult_x_18_n986), .CIX(mult_x_18_n637), .D(mult_x_18_n639), .CO(
        mult_x_18_n626), .COX(mult_x_18_n625), .S(mult_x_18_n627) );
  CMPE42D1BWP12T U3399 ( .A(mult_x_18_n738), .B(mult_x_18_n809), .C(
        mult_x_18_n625), .CIX(mult_x_18_n613), .D(mult_x_18_n626), .CO(
        mult_x_18_n606), .COX(mult_x_18_n605), .S(mult_x_18_n607) );
  CMPE42D1BWP12T U3400 ( .A(mult_x_18_n550), .B(mult_x_18_n537), .C(
        mult_x_18_n547), .CIX(mult_x_18_n543), .D(mult_x_18_n531), .CO(
        mult_x_18_n527), .COX(mult_x_18_n526), .S(mult_x_18_n528) );
  CMPE42D1BWP12T U3401 ( .A(mult_x_18_n925), .B(mult_x_18_n736), .C(
        mult_x_18_n981), .CIX(mult_x_18_n563), .D(mult_x_18_n556), .CO(
        mult_x_18_n553), .COX(mult_x_18_n552), .S(mult_x_18_n554) );
  CMPE42D1BWP12T U3402 ( .A(mult_x_18_n898), .B(mult_x_18_n770), .C(
        mult_x_18_n923), .CIX(mult_x_18_n529), .D(mult_x_18_n522), .CO(
        mult_x_18_n517), .COX(mult_x_18_n516), .S(mult_x_18_n518) );
  CMPE42D1BWP12T U3403 ( .A(mult_x_18_n768), .B(mult_x_18_n873), .C(
        mult_x_18_n501), .CIX(mult_x_18_n483), .D(mult_x_18_n502), .CO(
        mult_x_18_n473), .COX(mult_x_18_n472), .S(mult_x_18_n474) );
  CMPE42D1BWP12T U3404 ( .A(mult_x_18_n910), .B(mult_x_18_n866), .C(
        mult_x_18_n935), .CIX(mult_x_18_n685), .D(mult_x_18_n681), .CO(
        mult_x_18_n676), .COX(mult_x_18_n675), .S(mult_x_18_n677) );
  CMPE42D1BWP12T U3405 ( .A(mult_x_18_n870), .B(mult_x_18_n774), .C(
        mult_x_18_n765), .CIX(mult_x_18_n439), .D(mult_x_18_n785), .CO(
        mult_x_18_n413), .COX(mult_x_18_n412), .S(mult_x_18_n414) );
  CMPE42D1BWP12T U3406 ( .A(mult_x_18_n808), .B(mult_x_18_n880), .C(
        mult_x_18_n840), .CIX(mult_x_18_n611), .D(mult_x_18_n859), .CO(
        mult_x_18_n595), .COX(mult_x_18_n594), .S(mult_x_18_n596) );
  CMPE42D1BWP12T U3407 ( .A(mult_x_18_n792), .B(mult_x_18_n877), .C(
        mult_x_18_n952), .CIX(mult_x_18_n569), .D(mult_x_18_n805), .CO(
        mult_x_18_n547), .COX(mult_x_18_n546), .S(mult_x_18_n548) );
  CMPE42D1BWP12T U3408 ( .A(mult_x_18_n841), .B(mult_x_18_n956), .C(
        mult_x_18_n860), .CIX(mult_x_18_n622), .D(mult_x_18_n904), .CO(
        mult_x_18_n609), .COX(mult_x_18_n608), .S(mult_x_18_n610) );
  CMPE42D1BWP12T U3409 ( .A(mult_x_18_n844), .B(mult_x_18_n959), .C(
        mult_x_18_n863), .CIX(mult_x_18_n658), .D(mult_x_18_n651), .CO(
        mult_x_18_n645), .COX(mult_x_18_n644), .S(mult_x_18_n646) );
  CMPE42D1BWP12T U3410 ( .A(mult_x_18_n807), .B(mult_x_18_n954), .C(
        mult_x_18_n839), .CIX(mult_x_18_n597), .D(mult_x_18_n858), .CO(
        mult_x_18_n579), .COX(mult_x_18_n578), .S(mult_x_18_n580) );
  CMPE42D1BWP12T U3411 ( .A(mult_x_18_n400), .B(mult_x_18_n422), .C(
        mult_x_18_n416), .CIX(mult_x_18_n409), .D(mult_x_18_n413), .CO(
        mult_x_18_n387), .COX(mult_x_18_n386), .S(mult_x_18_n388) );
  CMPE42D1BWP12T U3412 ( .A(mult_x_18_n443), .B(mult_x_18_n464), .C(
        mult_x_18_n441), .CIX(mult_x_18_n456), .D(mult_x_18_n438), .CO(
        mult_x_18_n431), .COX(mult_x_18_n430), .S(mult_x_18_n432) );
  CMPE42D1BWP12T U3413 ( .A(mult_x_18_n892), .B(mult_x_18_n749), .C(
        mult_x_18_n973), .CIX(mult_x_18_n412), .D(mult_x_18_n402), .CO(
        mult_x_18_n399), .COX(mult_x_18_n398), .S(mult_x_18_n400) );
  CMPE42D1BWP12T U3414 ( .A(mult_x_18_n1005), .B(mult_x_18_n750), .C(
        mult_x_18_n974), .CIX(mult_x_18_n442), .D(mult_x_18_n444), .CO(
        mult_x_18_n422), .COX(mult_x_18_n421), .S(mult_x_18_n423) );
  CMPE42D1BWP12T U3415 ( .A(mult_x_18_n1021), .B(mult_x_18_n846), .C(
        mult_x_18_n990), .CIX(mult_x_18_n678), .D(mult_x_18_n680), .CO(
        mult_x_18_n670), .COX(mult_x_18_n669), .S(mult_x_18_n671) );
  CMPE42D1BWP12T U3416 ( .A(mult_x_18_n784), .B(mult_x_18_n812), .C(
        mult_x_18_n944), .CIX(mult_x_18_n418), .D(mult_x_18_n797), .CO(
        mult_x_18_n393), .COX(mult_x_18_n392), .S(mult_x_18_n394) );
  CMPE42D1BWP12T U3417 ( .A(mult_x_18_n423), .B(mult_x_18_n758), .C(
        mult_x_18_n420), .CIX(mult_x_18_n414), .D(mult_x_18_n417), .CO(
        mult_x_18_n410), .COX(mult_x_18_n409), .S(mult_x_18_n411) );
  CMPE42D1BWP12T U3418 ( .A(mult_x_18_n829), .B(mult_x_18_n752), .C(
        mult_x_18_n848), .CIX(mult_x_18_n415), .D(mult_x_18_n917), .CO(
        mult_x_18_n396), .COX(mult_x_18_n395), .S(mult_x_18_n397) );
  CMPE42D1BWP12T U3419 ( .A(mult_x_18_n766), .B(mult_x_18_n871), .C(
        mult_x_18_n786), .CIX(mult_x_18_n461), .D(mult_x_18_n946), .CO(
        mult_x_18_n434), .COX(mult_x_18_n433), .S(mult_x_18_n435) );
  CMPE42D1BWP12T U3420 ( .A(mult_x_18_n899), .B(mult_x_18_n819), .C(
        mult_x_18_n924), .CIX(mult_x_18_n546), .D(mult_x_18_n555), .CO(
        mult_x_18_n536), .COX(mult_x_18_n535), .S(mult_x_18_n537) );
  CMPE42D1BWP12T U3421 ( .A(mult_x_18_n861), .B(mult_x_18_n825), .C(
        mult_x_18_n905), .CIX(mult_x_18_n634), .D(mult_x_18_n930), .CO(
        mult_x_18_n623), .COX(mult_x_18_n622), .S(mult_x_18_n624) );
  CMPE42D1BWP12T U3422 ( .A(mult_x_18_n788), .B(mult_x_18_n734), .C(
        mult_x_18_n948), .CIX(mult_x_18_n498), .D(mult_x_18_n801), .CO(
        mult_x_18_n476), .COX(mult_x_18_n475), .S(mult_x_18_n477) );
  CMPE42D1BWP12T U3423 ( .A(mult_x_18_n388), .B(mult_x_18_n410), .C(
        mult_x_18_n385), .CIX(mult_x_18_n403), .D(mult_x_18_n407), .CO(
        mult_x_18_n381), .COX(mult_x_18_n380), .S(mult_x_18_n382) );
  CMPE42D1BWP12T U3424 ( .A(mult_x_18_n431), .B(mult_x_18_n411), .C(
        mult_x_18_n408), .CIX(mult_x_18_n424), .D(mult_x_18_n428), .CO(
        mult_x_18_n404), .COX(mult_x_18_n403), .S(mult_x_18_n405) );
  CMPE42D1BWP12T U3425 ( .A(mult_x_18_n945), .B(mult_x_18_n813), .C(
        mult_x_18_n798), .CIX(mult_x_18_n436), .D(mult_x_18_n830), .CO(
        mult_x_18_n416), .COX(mult_x_18_n415), .S(mult_x_18_n417) );
  CMPE42D1BWP12T U3426 ( .A(mult_x_18_n799), .B(mult_x_18_n759), .C(
        mult_x_18_n831), .CIX(mult_x_18_n458), .D(mult_x_18_n850), .CO(
        mult_x_18_n437), .COX(mult_x_18_n436), .S(mult_x_18_n438) );
  CMPE42D1BWP12T U3427 ( .A(mult_x_18_n769), .B(mult_x_18_n874), .C(
        mult_x_18_n789), .CIX(mult_x_18_n503), .D(mult_x_18_n510), .CO(
        mult_x_18_n493), .COX(mult_x_18_n492), .S(mult_x_18_n494) );
  CMPE42D1BWP12T U3428 ( .A(mult_x_18_n953), .B(mult_x_18_n878), .C(
        mult_x_18_n806), .CIX(mult_x_18_n581), .D(mult_x_18_n838), .CO(
        mult_x_18_n564), .COX(mult_x_18_n563), .S(mult_x_18_n565) );
  CMPE42D1BWP12T U3429 ( .A(mult_x_18_n903), .B(mult_x_18_n823), .C(
        mult_x_18_n928), .CIX(mult_x_18_n608), .D(mult_x_18_n614), .CO(
        mult_x_18_n598), .COX(mult_x_18_n597), .S(mult_x_18_n599) );
  CMPE42D1BWP12T U3430 ( .A(mult_x_18_n895), .B(mult_x_18_n815), .C(
        mult_x_18_n920), .CIX(mult_x_18_n475), .D(mult_x_18_n484), .CO(
        mult_x_18_n462), .COX(mult_x_18_n461), .S(mult_x_18_n463) );
  CMPE42D1BWP12T U3431 ( .A(mult_x_18_n609), .B(mult_x_18_n612), .C(
        mult_x_18_n606), .CIX(mult_x_18_n593), .D(mult_x_18_n602), .CO(
        mult_x_18_n589), .COX(mult_x_18_n588), .S(mult_x_18_n590) );
  CMPE42D1BWP12T U3432 ( .A(mult_x_18_n912), .B(mult_x_18_n964), .C(
        mult_x_18_n701), .CIX(mult_x_18_n695), .D(mult_x_18_n702), .CO(
        mult_x_18_n691), .COX(mult_x_18_n690), .S(mult_x_18_n692) );
  CMPE42D1BWP12T U3433 ( .A(mult_x_18_n595), .B(mult_x_18_n598), .C(
        mult_x_18_n592), .CIX(mult_x_18_n577), .D(mult_x_18_n588), .CO(
        mult_x_18_n573), .COX(mult_x_18_n572), .S(mult_x_18_n574) );
  CMPE42D1BWP12T U3434 ( .A(mult_x_18_n575), .B(mult_x_18_n579), .C(
        mult_x_18_n562), .CIX(mult_x_18_n572), .D(mult_x_18_n576), .CO(
        mult_x_18_n558), .COX(mult_x_18_n557), .S(mult_x_18_n559) );
  CMPE42D1BWP12T U3435 ( .A(mult_x_18_n469), .B(mult_x_18_n473), .C(
        mult_x_18_n451), .CIX(mult_x_18_n466), .D(mult_x_18_n470), .CO(
        mult_x_18_n447), .COX(mult_x_18_n446), .S(mult_x_18_n448) );
  CMPE42D1BWP12T U3436 ( .A(mult_x_18_n553), .B(mult_x_18_n534), .C(
        mult_x_18_n544), .CIX(mult_x_18_n540), .D(mult_x_18_n528), .CO(
        mult_x_18_n524), .COX(mult_x_18_n523), .S(mult_x_18_n525) );
  CMPE42D1BWP12T U3437 ( .A(mult_x_18_n933), .B(mult_x_18_n960), .C(
        mult_x_18_n989), .CIX(mult_x_18_n666), .D(mult_x_18_n662), .CO(
        mult_x_18_n659), .COX(mult_x_18_n658), .S(mult_x_18_n660) );
  CMPE42D1BWP12T U3438 ( .A(mult_x_18_n689), .B(mult_x_18_n963), .C(
        mult_x_18_n690), .CIX(mult_x_18_n694), .D(mult_x_18_n687), .CO(
        mult_x_18_n683), .COX(mult_x_18_n682), .S(mult_x_18_n684) );
endmodule


module top7 ( clk, reset, MEM_MEMCTRL_from_mem_data, 
        MEMCTRL_MEM_to_mem_read_enable, MEMCTRL_MEM_to_mem_write_enable, 
        MEMCTRL_MEM_to_mem_mem_enable, MEMCTRL_MEM_to_mem_address, 
        MEMCTRL_MEM_to_mem_data );
  input [15:0] MEM_MEMCTRL_from_mem_data;
  output [11:0] MEMCTRL_MEM_to_mem_address;
  output [15:0] MEMCTRL_MEM_to_mem_data;
  input clk, reset;
  output MEMCTRL_MEM_to_mem_read_enable, MEMCTRL_MEM_to_mem_write_enable,
         MEMCTRL_MEM_to_mem_mem_enable;
  wire   DEC_CPSR_update_flag_n, new_n, ALU_OUT_n, RF_OUT_n,
         DEC_CPSR_update_flag_c, new_c, ALU_OUT_c, RF_OUT_c,
         DEC_CPSR_update_flag_z, new_z, ALU_OUT_z, RF_OUT_z,
         DEC_CPSR_update_flag_v, new_v, ALU_OUT_v, RF_OUT_v,
         DEC_RF_alu_write_to_reg_enable, DEC_RF_memory_write_to_reg_enable,
         DEC_MISC_OUT_memory_address_source_is_reg,
         DEC_MEMCTRL_memorycontroller_sign_extend,
         DEC_MEMCTRL_memory_load_request, DEC_MEMCTRL_memory_store_request,
         DEC_IF_stall_to_instructionfetch, ALU_IN_c, irdecode_inst1_N1022,
         irdecode_inst1_N1021, irdecode_inst1_N1020, irdecode_inst1_N1019,
         irdecode_inst1_N1018, irdecode_inst1_N1017, irdecode_inst1_N1016,
         irdecode_inst1_N1015, irdecode_inst1_N1014, irdecode_inst1_N1013,
         irdecode_inst1_N1012, irdecode_inst1_N1011, irdecode_inst1_N1010,
         irdecode_inst1_N1009, irdecode_inst1_N1008, irdecode_inst1_N1007,
         irdecode_inst1_N1006, irdecode_inst1_N1005, irdecode_inst1_N1004,
         irdecode_inst1_N1003, irdecode_inst1_N1002, irdecode_inst1_N1001,
         irdecode_inst1_N1000, irdecode_inst1_N999, irdecode_inst1_N998,
         irdecode_inst1_N997, irdecode_inst1_N996, irdecode_inst1_N995,
         irdecode_inst1_N994, irdecode_inst1_N993, irdecode_inst1_N992,
         irdecode_inst1_N991, irdecode_inst1_N990, irdecode_inst1_N988,
         irdecode_inst1_N987, irdecode_inst1_N986, irdecode_inst1_N985,
         irdecode_inst1_N984, irdecode_inst1_N983, irdecode_inst1_N982,
         irdecode_inst1_N981, irdecode_inst1_N980, irdecode_inst1_N979,
         irdecode_inst1_N978, irdecode_inst1_N977, irdecode_inst1_N976,
         irdecode_inst1_N975, irdecode_inst1_N974, irdecode_inst1_N973,
         irdecode_inst1_N972, irdecode_inst1_N971, irdecode_inst1_N970,
         irdecode_inst1_N969, irdecode_inst1_N968, irdecode_inst1_N967,
         irdecode_inst1_N966, irdecode_inst1_N965, irdecode_inst1_N964,
         irdecode_inst1_N755, irdecode_inst1_N754, irdecode_inst1_N753,
         irdecode_inst1_N751, irdecode_inst1_next_split_instruction,
         irdecode_inst1_split_instruction, irdecode_inst1_next_step_0_,
         irdecode_inst1_next_step_1_, irdecode_inst1_next_step_2_,
         irdecode_inst1_next_step_3_, irdecode_inst1_next_step_4_,
         irdecode_inst1_next_step_5_, irdecode_inst1_next_step_6_,
         irdecode_inst1_next_step_7_, irdecode_inst1_itstate_0_,
         irdecode_inst1_itstate_1_, irdecode_inst1_itstate_2_,
         irdecode_inst1_itstate_3_, irdecode_inst1_itstate_4_,
         irdecode_inst1_itstate_5_, irdecode_inst1_itstate_6_,
         irdecode_inst1_itstate_7_,
         irdecode_inst1_next_stall_to_instructionfetch,
         irdecode_inst1_next_alu_write_to_reg_enable,
         irdecode_inst1_next_update_flag_v, irdecode_inst1_next_update_flag_c,
         irdecode_inst1_next_update_flag_n,
         memory_interface_inst1_delayed_is_signed, Instruction_Fetch_inst1_N99,
         Instruction_Fetch_inst1_N98, Instruction_Fetch_inst1_N97,
         Instruction_Fetch_inst1_N96, Instruction_Fetch_inst1_N95,
         Instruction_Fetch_inst1_N94, Instruction_Fetch_inst1_N93,
         Instruction_Fetch_inst1_N92, Instruction_Fetch_inst1_N91,
         Instruction_Fetch_inst1_N90, Instruction_Fetch_inst1_N89,
         Instruction_Fetch_inst1_N88, Instruction_Fetch_inst1_N87,
         Instruction_Fetch_inst1_N86, Instruction_Fetch_inst1_N85,
         Instruction_Fetch_inst1_N84, Instruction_Fetch_inst1_N80,
         Instruction_Fetch_inst1_N79,
         Instruction_Fetch_inst1_first_instruction_fetched,
         Instruction_Fetch_inst1_fetched_instruction_reg_0_,
         Instruction_Fetch_inst1_fetched_instruction_reg_1_,
         Instruction_Fetch_inst1_fetched_instruction_reg_2_,
         Instruction_Fetch_inst1_fetched_instruction_reg_3_,
         Instruction_Fetch_inst1_fetched_instruction_reg_4_,
         Instruction_Fetch_inst1_fetched_instruction_reg_5_,
         Instruction_Fetch_inst1_fetched_instruction_reg_6_,
         Instruction_Fetch_inst1_fetched_instruction_reg_7_,
         Instruction_Fetch_inst1_fetched_instruction_reg_8_,
         Instruction_Fetch_inst1_fetched_instruction_reg_9_,
         Instruction_Fetch_inst1_fetched_instruction_reg_10_,
         Instruction_Fetch_inst1_fetched_instruction_reg_11_,
         Instruction_Fetch_inst1_fetched_instruction_reg_12_,
         Instruction_Fetch_inst1_fetched_instruction_reg_13_,
         Instruction_Fetch_inst1_fetched_instruction_reg_14_,
         Instruction_Fetch_inst1_fetched_instruction_reg_15_,
         Instruction_Fetch_inst1_currentState_0_,
         Instruction_Fetch_inst1_currentState_1_,
         memory_interface_inst1_fsm_N35, memory_interface_inst1_fsm_N34,
         memory_interface_inst1_fsm_N33, memory_interface_inst1_fsm_N32,
         memory_interface_inst1_fsm_state_0_,
         memory_interface_inst1_fsm_state_1_,
         memory_interface_inst1_fsm_state_2_,
         memory_interface_inst1_fsm_state_3_, n755, n779, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41,
         SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43,
         SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45,
         SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47,
         SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49,
         SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51,
         SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53;
  wire   [4:0] DEC_RF_operand_a;
  wire   [4:0] DEC_RF_operand_b;
  wire   [31:0] DEC_RF_offset_b;
  wire   [4:0] DEC_ALU_alu_opcode;
  wire   [4:0] DEC_RF_alu_write_to_reg;
  wire   [4:0] DEC_RF_memory_write_to_reg;
  wire   [4:0] DEC_RF_memory_store_data_reg;
  wire   [4:0] DEC_RF_memory_store_address_reg;
  wire   [1:0] DEC_MEMCTRL_load_store_width;
  wire   [31:0] ALU_MISC_OUT_result;
  wire   [31:0] MEMCTRL_RF_IF_data_in;
  wire   [31:0] IF_RF_incremented_pc_out;
  wire   [31:0] RF_ALU_operand_a;
  wire   [31:0] RF_ALU_operand_b;
  wire   [31:0] RF_MEMCTRL_data_reg;
  wire   [12:2] RF_MEMCTRL_address_reg;
  wire   [31:0] RF_pc_out;
  wire   [11:0] MEMCTRL_IN_address;
  wire   [7:0] irdecode_inst1_step;
  wire   [4:0] irdecode_inst1_next_alu_write_to_reg;
  wire   [4:0] irdecode_inst1_next_alu_opcode;
  wire   [31:0] irdecode_inst1_next_offset_b;
  wire   [4:0] irdecode_inst1_next_operand_a;
  wire   [15:0] memory_interface_inst1_delay_first_two_bytes_out;
  wire   [31:0] memory_interface_inst1_delay_data_in32;
  wire   [11:0] memory_interface_inst1_delay_addr_for_adder;

  register_file register_file_inst1 ( .readA_sel(DEC_RF_operand_a), 
        .readB_sel(DEC_RF_operand_b), .readC_sel(DEC_RF_memory_store_data_reg), 
        .readD_sel(DEC_RF_memory_store_address_reg), .write1_sel(
        DEC_RF_alu_write_to_reg), .write2_sel(DEC_RF_memory_write_to_reg), 
        .write1_en(DEC_RF_alu_write_to_reg_enable), .write2_en(
        DEC_RF_memory_write_to_reg_enable), .write1_in(ALU_MISC_OUT_result), 
        .write2_in(MEMCTRL_RF_IF_data_in), .immediate1_in({n819, n819, n819, 
        n819, n819, n819, n819, n819, n819, n819, n819, n819, n819, n819, n819, 
        n819, n819, n819, n819, n819, n819, n819, n819, n819, n819, n819, n819, 
        n819, n819, n819, n819, n819}), .immediate2_in(DEC_RF_offset_b), 
        .next_pc_in({IF_RF_incremented_pc_out[31:2], MEMCTRL_IN_address[0], 
        IF_RF_incremented_pc_out[0]}), .next_cpsr_in({new_n, new_c, new_z, 
        new_v}), .next_sp_in({n819, n819, n819, n819, n819, n819, n819, n819, 
        n819, n819, n819, n819, n819, n819, n819, n819, n819, n819, n819, n819, 
        n819, n819, n819, n819, n819, n819, n819, n819, n819, n819, n819, n819}), .clk(clk), .reset(reset), .regA_out(RF_ALU_operand_a), .regB_out(
        RF_ALU_operand_b), .regC_out(RF_MEMCTRL_data_reg), .regD_out({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        RF_MEMCTRL_address_reg, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21}), .pc_out(RF_pc_out), .cpsr_out({RF_OUT_n, 
        RF_OUT_c, RF_OUT_z, RF_OUT_v}), .sp_out({SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53}), .next_pc_en_BAR(n755) );
  ALU_VARIABLE ALU_VARIABLE_inst1 ( .a(RF_ALU_operand_a), .b(RF_ALU_operand_b), 
        .op(DEC_ALU_alu_opcode[3:0]), .c_in(ALU_IN_c), .result(
        ALU_MISC_OUT_result), .c_out(ALU_OUT_c), .z(ALU_OUT_z), .n(ALU_OUT_n), 
        .v(ALU_OUT_v) );
  CKAN2D2BWP12T irdecode_inst1_C2448 ( .A1(irdecode_inst1_next_step_2_), .A2(
        n817), .Z(irdecode_inst1_N753) );
  OR3XD4BWP12T irdecode_inst1_C4464 ( .A1(irdecode_inst1_next_step_0_), .A2(
        irdecode_inst1_N751), .A3(irdecode_inst1_N754), .Z(irdecode_inst1_N755) );
  CKAN2D2BWP12T irdecode_inst1_C2445 ( .A1(irdecode_inst1_next_step_1_), .A2(
        n816), .Z(irdecode_inst1_N751) );
  CKAN2D2BWP12T irdecode_inst1_C2449 ( .A1(irdecode_inst1_N753), .A2(n816), 
        .Z(irdecode_inst1_N754) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_0_ ( .D(
        MEM_MEMCTRL_from_mem_data[8]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[0]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_1_ ( .D(
        MEM_MEMCTRL_from_mem_data[9]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[1]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_2_ ( .D(
        MEM_MEMCTRL_from_mem_data[10]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_3_ ( .D(
        MEM_MEMCTRL_from_mem_data[11]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_4_ ( .D(
        MEM_MEMCTRL_from_mem_data[12]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[4]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_5_ ( .D(
        MEM_MEMCTRL_from_mem_data[13]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[5]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_6_ ( .D(
        MEM_MEMCTRL_from_mem_data[14]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_7_ ( .D(
        MEM_MEMCTRL_from_mem_data[15]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_8_ ( .D(
        MEM_MEMCTRL_from_mem_data[0]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_9_ ( .D(
        MEM_MEMCTRL_from_mem_data[1]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_10_ ( .D(
        MEM_MEMCTRL_from_mem_data[2]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_11_ ( .D(
        MEM_MEMCTRL_from_mem_data[3]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[11]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_12_ ( .D(
        MEM_MEMCTRL_from_mem_data[4]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[12]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_13_ ( .D(
        MEM_MEMCTRL_from_mem_data[5]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[13]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_14_ ( .D(
        MEM_MEMCTRL_from_mem_data[6]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[14]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_15_ ( .D(
        MEM_MEMCTRL_from_mem_data[7]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[15]) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_3_ ( .D(
        memory_interface_inst1_fsm_N35), .CP(clk), .Q(
        memory_interface_inst1_fsm_state_3_) );
  DFQD1BWP12T Instruction_Fetch_inst1_first_instruction_fetched_reg ( .D(n815), 
        .CP(clk), .Q(Instruction_Fetch_inst1_first_instruction_fetched) );
  DFQD1BWP12T irdecode_inst1_memorycontroller_sign_extend_reg ( .D(n785), .CP(
        clk), .Q(DEC_MEMCTRL_memorycontroller_sign_extend) );
  DFQD1BWP12T memory_interface_inst1_delayed_is_signed_reg ( .D(
        DEC_MEMCTRL_memorycontroller_sign_extend), .CP(clk), .Q(
        memory_interface_inst1_delayed_is_signed) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_14_ ( .D(
        Instruction_Fetch_inst1_N98), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_14_) );
  DFQD1BWP12T irdecode_inst1_load_store_width_reg_1_ ( .D(n787), .CP(clk), .Q(
        DEC_MEMCTRL_load_store_width[1]) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_1_ ( .D(
        memory_interface_inst1_fsm_N33), .CP(clk), .Q(
        memory_interface_inst1_fsm_state_1_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_1_ ( .D(
        Instruction_Fetch_inst1_N85), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_1_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_2_ ( .D(
        Instruction_Fetch_inst1_N86), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_2_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_0_ ( .D(
        Instruction_Fetch_inst1_N84), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_0_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_3_ ( .D(
        Instruction_Fetch_inst1_N87), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_3_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_4_ ( .D(
        Instruction_Fetch_inst1_N88), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_4_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_7_ ( .D(
        Instruction_Fetch_inst1_N91), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_7_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_5_ ( .D(
        Instruction_Fetch_inst1_N89), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_5_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_6_ ( .D(
        Instruction_Fetch_inst1_N90), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_6_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_15_ ( .D(
        Instruction_Fetch_inst1_N99), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_15_) );
  DFQD1BWP12T irdecode_inst1_step_reg_7_ ( .D(irdecode_inst1_next_step_7_), 
        .CP(clk), .Q(irdecode_inst1_step[7]) );
  DFQD1BWP12T irdecode_inst1_memory_store_request_reg ( .D(n814), .CP(clk), 
        .Q(DEC_MEMCTRL_memory_store_request) );
  DFQD1BWP12T irdecode_inst1_step_reg_6_ ( .D(irdecode_inst1_next_step_6_), 
        .CP(clk), .Q(irdecode_inst1_step[6]) );
  DFQD1BWP12T irdecode_inst1_step_reg_5_ ( .D(irdecode_inst1_next_step_5_), 
        .CP(clk), .Q(irdecode_inst1_step[5]) );
  DFQD1BWP12T irdecode_inst1_memory_load_request_reg ( .D(n805), .CP(clk), .Q(
        DEC_MEMCTRL_memory_load_request) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_2_ ( .D(
        memory_interface_inst1_fsm_N34), .CP(clk), .Q(
        memory_interface_inst1_fsm_state_2_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_8_ ( .D(
        Instruction_Fetch_inst1_N92), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_8_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_9_ ( .D(
        Instruction_Fetch_inst1_N93), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_9_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_11_ ( .D(
        Instruction_Fetch_inst1_N95), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_11_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_12_ ( .D(
        Instruction_Fetch_inst1_N96), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_12_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_10_ ( .D(
        Instruction_Fetch_inst1_N94), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_10_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_13_ ( .D(
        Instruction_Fetch_inst1_N97), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_13_) );
  DFQD1BWP12T irdecode_inst1_stall_to_instructionfetch_reg ( .D(
        irdecode_inst1_next_stall_to_instructionfetch), .CP(clk), .Q(
        DEC_IF_stall_to_instructionfetch) );
  DFQD1BWP12T Instruction_Fetch_inst1_currentState_reg_1_ ( .D(
        Instruction_Fetch_inst1_N80), .CP(clk), .Q(
        Instruction_Fetch_inst1_currentState_1_) );
  DFQD1BWP12T Instruction_Fetch_inst1_currentState_reg_0_ ( .D(
        Instruction_Fetch_inst1_N79), .CP(clk), .Q(
        Instruction_Fetch_inst1_currentState_0_) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_0_ ( .D(
        MEMCTRL_IN_address[0]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[0]) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_1_ ( .D(n790), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[1]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_23_ ( .D(
        irdecode_inst1_next_offset_b[23]), .CP(clk), .Q(DEC_RF_offset_b[23])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_24_ ( .D(
        irdecode_inst1_next_offset_b[24]), .CP(clk), .Q(DEC_RF_offset_b[24])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_25_ ( .D(
        irdecode_inst1_next_offset_b[25]), .CP(clk), .Q(DEC_RF_offset_b[25])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_26_ ( .D(
        irdecode_inst1_next_offset_b[26]), .CP(clk), .Q(DEC_RF_offset_b[26])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_27_ ( .D(
        irdecode_inst1_next_offset_b[27]), .CP(clk), .Q(DEC_RF_offset_b[27])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_28_ ( .D(
        irdecode_inst1_next_offset_b[28]), .CP(clk), .Q(DEC_RF_offset_b[28])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_29_ ( .D(
        irdecode_inst1_next_offset_b[29]), .CP(clk), .Q(DEC_RF_offset_b[29])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_30_ ( .D(
        irdecode_inst1_next_offset_b[30]), .CP(clk), .Q(DEC_RF_offset_b[30])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_31_ ( .D(
        irdecode_inst1_next_offset_b[31]), .CP(clk), .Q(DEC_RF_offset_b[31])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_12_ ( .D(
        irdecode_inst1_next_offset_b[12]), .CP(clk), .Q(DEC_RF_offset_b[12])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_13_ ( .D(
        irdecode_inst1_next_offset_b[13]), .CP(clk), .Q(DEC_RF_offset_b[13])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_14_ ( .D(
        irdecode_inst1_next_offset_b[14]), .CP(clk), .Q(DEC_RF_offset_b[14])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_15_ ( .D(
        irdecode_inst1_next_offset_b[15]), .CP(clk), .Q(DEC_RF_offset_b[15])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_16_ ( .D(
        irdecode_inst1_next_offset_b[16]), .CP(clk), .Q(DEC_RF_offset_b[16])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_17_ ( .D(
        irdecode_inst1_next_offset_b[17]), .CP(clk), .Q(DEC_RF_offset_b[17])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_18_ ( .D(
        irdecode_inst1_next_offset_b[18]), .CP(clk), .Q(DEC_RF_offset_b[18])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_19_ ( .D(
        irdecode_inst1_next_offset_b[19]), .CP(clk), .Q(DEC_RF_offset_b[19])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_20_ ( .D(
        irdecode_inst1_next_offset_b[20]), .CP(clk), .Q(DEC_RF_offset_b[20])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_21_ ( .D(
        irdecode_inst1_next_offset_b[21]), .CP(clk), .Q(DEC_RF_offset_b[21])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_22_ ( .D(
        irdecode_inst1_next_offset_b[22]), .CP(clk), .Q(DEC_RF_offset_b[22])
         );
  DFQD1BWP12T irdecode_inst1_itstate_reg_0_ ( .D(n813), .CP(clk), .Q(
        irdecode_inst1_itstate_0_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_1_ ( .D(n812), .CP(clk), .Q(
        irdecode_inst1_itstate_1_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_2_ ( .D(n811), .CP(clk), .Q(
        irdecode_inst1_itstate_2_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_3_ ( .D(n810), .CP(clk), .Q(
        irdecode_inst1_itstate_3_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_4_ ( .D(n809), .CP(clk), .Q(
        irdecode_inst1_itstate_4_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_5_ ( .D(n808), .CP(clk), .Q(
        irdecode_inst1_itstate_5_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_6_ ( .D(n807), .CP(clk), .Q(
        irdecode_inst1_itstate_6_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_7_ ( .D(n806), .CP(clk), .Q(
        irdecode_inst1_itstate_7_) );
  DFQD1BWP12T irdecode_inst1_update_flag_v_reg ( .D(
        irdecode_inst1_next_update_flag_v), .CP(clk), .Q(
        DEC_CPSR_update_flag_v) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_1_ ( .D(
        irdecode_inst1_next_alu_write_to_reg[1]), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[1]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_enable_reg ( .D(
        irdecode_inst1_next_alu_write_to_reg_enable), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg_enable) );
  DFQD1BWP12T irdecode_inst1_step_reg_2_ ( .D(irdecode_inst1_next_step_2_), 
        .CP(clk), .Q(irdecode_inst1_step[2]) );
  DFQD1BWP12T irdecode_inst1_step_reg_3_ ( .D(irdecode_inst1_next_step_3_), 
        .CP(clk), .Q(irdecode_inst1_step[3]) );
  DFQD1BWP12T irdecode_inst1_step_reg_4_ ( .D(irdecode_inst1_next_step_4_), 
        .CP(clk), .Q(irdecode_inst1_step[4]) );
  DFQD1BWP12T irdecode_inst1_step_reg_0_ ( .D(irdecode_inst1_next_step_0_), 
        .CP(clk), .Q(irdecode_inst1_step[0]) );
  DFQD1BWP12T irdecode_inst1_step_reg_1_ ( .D(irdecode_inst1_next_step_1_), 
        .CP(clk), .Q(irdecode_inst1_step[1]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_9_ ( .D(
        irdecode_inst1_next_offset_b[9]), .CP(clk), .Q(DEC_RF_offset_b[9]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_10_ ( .D(
        irdecode_inst1_next_offset_b[10]), .CP(clk), .Q(DEC_RF_offset_b[10])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_11_ ( .D(
        irdecode_inst1_next_offset_b[11]), .CP(clk), .Q(DEC_RF_offset_b[11])
         );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_6_ ( .D(
        irdecode_inst1_next_offset_b[6]), .CP(clk), .Q(DEC_RF_offset_b[6]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_7_ ( .D(
        irdecode_inst1_next_offset_b[7]), .CP(clk), .Q(DEC_RF_offset_b[7]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_8_ ( .D(
        irdecode_inst1_next_offset_b[8]), .CP(clk), .Q(DEC_RF_offset_b[8]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_1_ ( .D(n801), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[1]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_4_ ( .D(n804), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[4]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_5_ ( .D(
        irdecode_inst1_next_offset_b[5]), .CP(clk), .Q(DEC_RF_offset_b[5]) );
  DFQD1BWP12T irdecode_inst1_load_store_width_reg_0_ ( .D(n786), .CP(clk), .Q(
        DEC_MEMCTRL_load_store_width[0]) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_0_ ( .D(
        memory_interface_inst1_fsm_N32), .CP(clk), .Q(
        memory_interface_inst1_fsm_state_0_) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_enable_reg ( .D(n799), .CP(
        clk), .Q(DEC_RF_memory_write_to_reg_enable) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_4_ ( .D(n798), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[4]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_1_ ( .D(n795), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[1]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_4_ ( .D(
        irdecode_inst1_next_alu_opcode[4]), .CP(clk), .Q(DEC_ALU_alu_opcode[4]) );
  DFQD1BWP12T irdecode_inst1_split_instruction_reg ( .D(
        irdecode_inst1_next_split_instruction), .CP(clk), .Q(
        irdecode_inst1_split_instruction) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_3_ ( .D(n803), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[3]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_3_ ( .D(n797), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[3]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_2_ ( .D(n802), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[2]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_2_ ( .D(n796), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[2]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_0_ ( .D(n800), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[0]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_0_ ( .D(n794), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[0]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_0_ ( .D(
        irdecode_inst1_next_alu_write_to_reg[0]), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[0]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_2_ ( .D(
        irdecode_inst1_next_alu_write_to_reg[2]), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[2]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_4_ ( .D(
        irdecode_inst1_next_alu_write_to_reg[4]), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[4]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_3_ ( .D(
        irdecode_inst1_next_alu_opcode[3]), .CP(clk), .Q(DEC_ALU_alu_opcode[3]) );
  DFQD1BWP12T irdecode_inst1_memory_address_source_is_reg_reg ( .D(n788), .CP(
        clk), .Q(DEC_MISC_OUT_memory_address_source_is_reg) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_3_ ( .D(
        irdecode_inst1_next_offset_b[3]), .CP(clk), .Q(DEC_RF_offset_b[3]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_4_ ( .D(
        irdecode_inst1_next_offset_b[4]), .CP(clk), .Q(DEC_RF_offset_b[4]) );
  DFQD1BWP12T irdecode_inst1_update_flag_c_reg ( .D(
        irdecode_inst1_next_update_flag_c), .CP(clk), .Q(
        DEC_CPSR_update_flag_c) );
  DFQD1BWP12T irdecode_inst1_update_flag_n_reg ( .D(
        irdecode_inst1_next_update_flag_n), .CP(clk), .Q(
        DEC_CPSR_update_flag_n) );
  DFQD1BWP12T irdecode_inst1_update_flag_z_reg ( .D(
        irdecode_inst1_next_update_flag_n), .CP(clk), .Q(
        DEC_CPSR_update_flag_z) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_2_ ( .D(
        irdecode_inst1_next_alu_opcode[2]), .CP(clk), .Q(DEC_ALU_alu_opcode[2]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_0_ ( .D(
        irdecode_inst1_next_alu_opcode[0]), .CP(clk), .Q(DEC_ALU_alu_opcode[0]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_1_ ( .D(
        irdecode_inst1_next_alu_opcode[1]), .CP(clk), .Q(DEC_ALU_alu_opcode[1]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_0_ ( .D(
        irdecode_inst1_next_offset_b[0]), .CP(clk), .Q(DEC_RF_offset_b[0]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_1_ ( .D(
        irdecode_inst1_next_offset_b[1]), .CP(clk), .Q(DEC_RF_offset_b[1]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_2_ ( .D(
        irdecode_inst1_next_offset_b[2]), .CP(clk), .Q(DEC_RF_offset_b[2]) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_4_ ( .D(n793), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[4]) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_3_ ( .D(n792), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[3]) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_2_ ( .D(n791), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[2]) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_0_ ( .D(n789), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[0]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_3_ ( .D(
        irdecode_inst1_next_alu_write_to_reg[3]), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_0_ ( .D(
        RF_MEMCTRL_data_reg[0]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[0]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_1_ ( .D(
        RF_MEMCTRL_data_reg[1]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[1]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_2_ ( .D(
        RF_MEMCTRL_data_reg[2]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_3_ ( .D(
        RF_MEMCTRL_data_reg[3]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_4_ ( .D(
        RF_MEMCTRL_data_reg[4]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[4]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_5_ ( .D(
        RF_MEMCTRL_data_reg[5]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[5]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_6_ ( .D(
        RF_MEMCTRL_data_reg[6]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_7_ ( .D(
        RF_MEMCTRL_data_reg[7]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_8_ ( .D(
        RF_MEMCTRL_data_reg[8]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_9_ ( .D(
        RF_MEMCTRL_data_reg[9]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_10_ ( .D(
        RF_MEMCTRL_data_reg[10]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_11_ ( .D(
        RF_MEMCTRL_data_reg[11]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[11]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_12_ ( .D(
        RF_MEMCTRL_data_reg[12]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[12]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_13_ ( .D(
        RF_MEMCTRL_data_reg[13]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[13]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_14_ ( .D(
        RF_MEMCTRL_data_reg[14]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[14]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_15_ ( .D(
        RF_MEMCTRL_data_reg[15]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[15]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_16_ ( .D(
        RF_MEMCTRL_data_reg[16]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[16]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_17_ ( .D(
        RF_MEMCTRL_data_reg[17]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[17]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_18_ ( .D(
        RF_MEMCTRL_data_reg[18]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[18]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_19_ ( .D(
        RF_MEMCTRL_data_reg[19]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[19]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_20_ ( .D(
        RF_MEMCTRL_data_reg[20]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[20]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_21_ ( .D(
        RF_MEMCTRL_data_reg[21]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[21]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_22_ ( .D(
        RF_MEMCTRL_data_reg[22]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[22]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_23_ ( .D(
        RF_MEMCTRL_data_reg[23]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[23]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_24_ ( .D(
        RF_MEMCTRL_data_reg[24]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[24]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_25_ ( .D(
        RF_MEMCTRL_data_reg[25]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[25]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_26_ ( .D(
        RF_MEMCTRL_data_reg[26]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[26]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_27_ ( .D(
        RF_MEMCTRL_data_reg[27]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[27]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_28_ ( .D(
        RF_MEMCTRL_data_reg[28]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[28]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_29_ ( .D(
        RF_MEMCTRL_data_reg[29]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[29]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_30_ ( .D(
        RF_MEMCTRL_data_reg[30]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[30]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_31_ ( .D(
        RF_MEMCTRL_data_reg[31]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[31]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_1_ ( .D(
        MEMCTRL_IN_address[1]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[1]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_2_ ( .D(
        MEMCTRL_IN_address[2]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_3_ ( .D(
        MEMCTRL_IN_address[3]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_4_ ( .D(
        MEMCTRL_IN_address[4]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[4]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_5_ ( .D(
        MEMCTRL_IN_address[5]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[5]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_6_ ( .D(
        MEMCTRL_IN_address[6]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_7_ ( .D(
        MEMCTRL_IN_address[7]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_8_ ( .D(
        MEMCTRL_IN_address[8]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_9_ ( .D(
        MEMCTRL_IN_address[9]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_10_ ( .D(
        MEMCTRL_IN_address[10]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_11_ ( .D(
        MEMCTRL_IN_address[11]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[11]) );
  LHQD1BWP12T irdecode_inst1_next_step_reg_7_ ( .E(irdecode_inst1_N969), .D(
        irdecode_inst1_N988), .Q(irdecode_inst1_next_step_7_) );
  LHQD1BWP12T irdecode_inst1_next_step_reg_6_ ( .E(irdecode_inst1_N969), .D(
        irdecode_inst1_N987), .Q(irdecode_inst1_next_step_6_) );
  LHQD1BWP12T irdecode_inst1_next_step_reg_5_ ( .E(irdecode_inst1_N969), .D(
        irdecode_inst1_N986), .Q(irdecode_inst1_next_step_5_) );
  LHQD1BWP12T irdecode_inst1_next_stall_to_instructionfetch_reg ( .E(
        irdecode_inst1_N969), .D(irdecode_inst1_N980), .Q(
        irdecode_inst1_next_stall_to_instructionfetch) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_23_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1014), .Q(irdecode_inst1_next_offset_b[23]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_24_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1015), .Q(irdecode_inst1_next_offset_b[24]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_25_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1016), .Q(irdecode_inst1_next_offset_b[25]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_26_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1017), .Q(irdecode_inst1_next_offset_b[26]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_27_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1018), .Q(irdecode_inst1_next_offset_b[27]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_28_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1019), .Q(irdecode_inst1_next_offset_b[28]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_29_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1020), .Q(irdecode_inst1_next_offset_b[29]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_30_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1021), .Q(irdecode_inst1_next_offset_b[30]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_31_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1022), .Q(irdecode_inst1_next_offset_b[31]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_12_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1003), .Q(irdecode_inst1_next_offset_b[12]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_13_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1004), .Q(irdecode_inst1_next_offset_b[13]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_14_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1005), .Q(irdecode_inst1_next_offset_b[14]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_15_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1006), .Q(irdecode_inst1_next_offset_b[15]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_16_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1007), .Q(irdecode_inst1_next_offset_b[16]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_17_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1008), .Q(irdecode_inst1_next_offset_b[17]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_18_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1009), .Q(irdecode_inst1_next_offset_b[18]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_19_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1010), .Q(irdecode_inst1_next_offset_b[19]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_20_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1011), .Q(irdecode_inst1_next_offset_b[20]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_21_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1012), .Q(irdecode_inst1_next_offset_b[21]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_22_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1013), .Q(irdecode_inst1_next_offset_b[22]) );
  LHQD1BWP12T irdecode_inst1_next_operand_a_reg_1_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N971), .Q(irdecode_inst1_next_operand_a[1]) );
  LHQD1BWP12T irdecode_inst1_next_alu_write_to_reg_reg_1_ ( .E(
        irdecode_inst1_N969), .D(irdecode_inst1_N976), .Q(
        irdecode_inst1_next_alu_write_to_reg[1]) );
  LHQD1BWP12T irdecode_inst1_next_step_reg_2_ ( .E(irdecode_inst1_N969), .D(
        irdecode_inst1_N983), .Q(irdecode_inst1_next_step_2_) );
  LHQD1BWP12T irdecode_inst1_next_step_reg_3_ ( .E(irdecode_inst1_N969), .D(
        irdecode_inst1_N984), .Q(irdecode_inst1_next_step_3_) );
  LHQD1BWP12T irdecode_inst1_next_step_reg_4_ ( .E(irdecode_inst1_N969), .D(
        irdecode_inst1_N985), .Q(irdecode_inst1_next_step_4_) );
  LHQD1BWP12T irdecode_inst1_next_step_reg_0_ ( .E(irdecode_inst1_N969), .D(
        irdecode_inst1_N981), .Q(irdecode_inst1_next_step_0_) );
  LHQD1BWP12T irdecode_inst1_next_step_reg_1_ ( .E(irdecode_inst1_N969), .D(
        irdecode_inst1_N982), .Q(irdecode_inst1_next_step_1_) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_9_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1000), .Q(irdecode_inst1_next_offset_b[9]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_10_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1001), .Q(irdecode_inst1_next_offset_b[10]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_11_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N1002), .Q(irdecode_inst1_next_offset_b[11]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_6_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N997), .Q(irdecode_inst1_next_offset_b[6]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_7_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N998), .Q(irdecode_inst1_next_offset_b[7]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_8_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N999), .Q(irdecode_inst1_next_offset_b[8]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_5_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N996), .Q(irdecode_inst1_next_offset_b[5]) );
  LHQD1BWP12T irdecode_inst1_next_alu_opcode_reg_4_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N968), .Q(irdecode_inst1_next_alu_opcode[4]) );
  LHQD1BWP12T irdecode_inst1_next_split_instruction_reg ( .E(
        irdecode_inst1_N969), .D(irdecode_inst1_N990), .Q(
        irdecode_inst1_next_split_instruction) );
  LHQD1BWP12T irdecode_inst1_next_alu_write_to_reg_reg_0_ ( .E(
        irdecode_inst1_N969), .D(irdecode_inst1_N975), .Q(
        irdecode_inst1_next_alu_write_to_reg[0]) );
  LHQD1BWP12T irdecode_inst1_next_alu_write_to_reg_reg_2_ ( .E(
        irdecode_inst1_N969), .D(irdecode_inst1_N977), .Q(
        irdecode_inst1_next_alu_write_to_reg[2]) );
  LHQD1BWP12T irdecode_inst1_next_alu_write_to_reg_reg_4_ ( .E(
        irdecode_inst1_N969), .D(irdecode_inst1_N979), .Q(
        irdecode_inst1_next_alu_write_to_reg[4]) );
  LHQD1BWP12T irdecode_inst1_next_operand_a_reg_0_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N970), .Q(irdecode_inst1_next_operand_a[0]) );
  LHQD1BWP12T irdecode_inst1_next_operand_a_reg_2_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N972), .Q(irdecode_inst1_next_operand_a[2]) );
  LHQD1BWP12T irdecode_inst1_next_operand_a_reg_3_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N973), .Q(irdecode_inst1_next_operand_a[3]) );
  LHQD1BWP12T irdecode_inst1_next_operand_a_reg_4_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N974), .Q(irdecode_inst1_next_operand_a[4]) );
  LHQD1BWP12T irdecode_inst1_next_alu_opcode_reg_3_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N967), .Q(irdecode_inst1_next_alu_opcode[3]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_3_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N994), .Q(irdecode_inst1_next_offset_b[3]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_4_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N995), .Q(irdecode_inst1_next_offset_b[4]) );
  LHQD1BWP12T irdecode_inst1_next_alu_opcode_reg_2_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N966), .Q(irdecode_inst1_next_alu_opcode[2]) );
  LHQD1BWP12T irdecode_inst1_next_alu_opcode_reg_0_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N964), .Q(irdecode_inst1_next_alu_opcode[0]) );
  LHQD1BWP12T irdecode_inst1_next_alu_opcode_reg_1_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N965), .Q(irdecode_inst1_next_alu_opcode[1]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_0_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N991), .Q(irdecode_inst1_next_offset_b[0]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_1_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N992), .Q(irdecode_inst1_next_offset_b[1]) );
  LHQD1BWP12T irdecode_inst1_next_offset_b_reg_2_ ( .E(irdecode_inst1_N969), 
        .D(irdecode_inst1_N993), .Q(irdecode_inst1_next_offset_b[2]) );
  LHQD1BWP12T irdecode_inst1_next_alu_write_to_reg_reg_3_ ( .E(
        irdecode_inst1_N969), .D(irdecode_inst1_N978), .Q(
        irdecode_inst1_next_alu_write_to_reg[3]) );
  DFQD4BWP12T irdecode_inst1_operand_a_reg_3_ ( .D(
        irdecode_inst1_next_operand_a[3]), .CP(clk), .Q(DEC_RF_operand_a[3])
         );
  DFQD4BWP12T irdecode_inst1_operand_b_reg_0_ ( .D(n784), .CP(clk), .Q(
        DEC_RF_operand_b[0]) );
  DFQD4BWP12T irdecode_inst1_operand_a_reg_1_ ( .D(
        irdecode_inst1_next_operand_a[1]), .CP(clk), .Q(DEC_RF_operand_a[1])
         );
  DFQD4BWP12T irdecode_inst1_operand_a_reg_2_ ( .D(
        irdecode_inst1_next_operand_a[2]), .CP(clk), .Q(DEC_RF_operand_a[2])
         );
  DFQD4BWP12T irdecode_inst1_operand_b_reg_2_ ( .D(n782), .CP(clk), .Q(
        DEC_RF_operand_b[2]) );
  DFQD4BWP12T irdecode_inst1_operand_b_reg_3_ ( .D(n781), .CP(clk), .Q(
        DEC_RF_operand_b[3]) );
  DFQD4BWP12T irdecode_inst1_operand_a_reg_0_ ( .D(
        irdecode_inst1_next_operand_a[0]), .CP(clk), .Q(DEC_RF_operand_a[0])
         );
  DFQD4BWP12T irdecode_inst1_operand_a_reg_4_ ( .D(
        irdecode_inst1_next_operand_a[4]), .CP(clk), .Q(DEC_RF_operand_a[4])
         );
  DFQD4BWP12T irdecode_inst1_operand_b_reg_1_ ( .D(n783), .CP(clk), .Q(
        DEC_RF_operand_b[1]) );
  DFQD4BWP12T irdecode_inst1_operand_b_reg_4_ ( .D(n779), .CP(clk), .Q(
        DEC_RF_operand_b[4]) );
  TIELBWP12T U1017 ( .ZN(n819) );
  INVD1BWP12T U1018 ( .I(n819), .ZN(MEMCTRL_MEM_to_mem_mem_enable) );
  MUX2ND0BWP12T U1019 ( .I0(MEM_MEMCTRL_from_mem_data[15]), .I1(n1564), .S(
        n1563), .ZN(n1580) );
  INVD1BWP12T U1020 ( .I(n1187), .ZN(n1185) );
  MAOI22D0BWP12T U1021 ( .A1(RF_pc_out[11]), .A2(n1064), .B1(RF_pc_out[11]), 
        .B2(n1064), .ZN(n1137) );
  MAOI22D0BWP12T U1022 ( .A1(RF_pc_out[9]), .A2(n1067), .B1(RF_pc_out[9]), 
        .B2(n1067), .ZN(n1144) );
  MAOI22D0BWP12T U1023 ( .A1(RF_pc_out[7]), .A2(n1071), .B1(RF_pc_out[7]), 
        .B2(n1071), .ZN(n1145) );
  MAOI22D0BWP12T U1024 ( .A1(RF_pc_out[5]), .A2(n1073), .B1(RF_pc_out[5]), 
        .B2(n1073), .ZN(n1140) );
  MAOI22D0BWP12T U1025 ( .A1(RF_pc_out[4]), .A2(n1077), .B1(RF_pc_out[4]), 
        .B2(n1077), .ZN(n1139) );
  MAOI22D0BWP12T U1026 ( .A1(RF_pc_out[2]), .A2(n1188), .B1(RF_pc_out[2]), 
        .B2(n1188), .ZN(n1135) );
  INVD1BWP12T U1027 ( .I(n1476), .ZN(n1593) );
  MAOI22D0BWP12T U1028 ( .A1(n1428), .A2(
        memory_interface_inst1_delay_data_in32[24]), .B1(n1570), .B2(n1409), 
        .ZN(n1402) );
  MAOI22D0BWP12T U1029 ( .A1(n1428), .A2(
        memory_interface_inst1_delay_data_in32[25]), .B1(n1572), .B2(n1409), 
        .ZN(n1405) );
  MAOI22D0BWP12T U1030 ( .A1(n1498), .A2(n1335), .B1(n1337), .B2(n1625), .ZN(
        n1331) );
  MAOI22D0BWP12T U1031 ( .A1(n1103), .A2(n1592), .B1(n1103), .B2(n1592), .ZN(
        n1109) );
  MAOI22D0BWP12T U1032 ( .A1(n1452), .A2(n1106), .B1(n1452), .B2(n1106), .ZN(
        n1107) );
  MAOI22D0BWP12T U1033 ( .A1(n1278), .A2(n1095), .B1(n1095), .B2(n1549), .ZN(
        n1102) );
  MOAI22D0BWP12T U1034 ( .A1(n1096), .A2(n1549), .B1(n1096), .B2(n1278), .ZN(
        n1101) );
  AO22D0BWP12T U1035 ( .A1(MEMCTRL_RF_IF_data_in[7]), .A2(n1610), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_7_), .B2(n1155), .Z(
        n1348) );
  NR2D0BWP12T U1036 ( .A1(RF_pc_out[2]), .A2(RF_pc_out[1]), .ZN(n820) );
  MAOI22D0BWP12T U1037 ( .A1(RF_pc_out[3]), .A2(n820), .B1(RF_pc_out[3]), .B2(
        n820), .ZN(n1141) );
  CKND0BWP12T U1038 ( .I(RF_MEMCTRL_data_reg[10]), .ZN(n821) );
  MAOI22D0BWP12T U1039 ( .A1(n1428), .A2(
        memory_interface_inst1_delay_data_in32[26]), .B1(n1409), .B2(n1582), 
        .ZN(n822) );
  CKND2D0BWP12T U1040 ( .A1(n1410), .A2(
        memory_interface_inst1_delay_data_in32[10]), .ZN(n823) );
  OAI211D0BWP12T U1041 ( .A1(n1414), .A2(n821), .B(n822), .C(n823), .ZN(
        MEMCTRL_MEM_to_mem_data[2]) );
  MAOI22D0BWP12T U1042 ( .A1(n1155), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_3_), .B1(n1615), .B2(
        n755), .ZN(n1329) );
  CKND0BWP12T U1043 ( .I(RF_MEMCTRL_data_reg[11]), .ZN(n824) );
  MAOI22D0BWP12T U1044 ( .A1(n1428), .A2(
        memory_interface_inst1_delay_data_in32[27]), .B1(n1409), .B2(n1569), 
        .ZN(n825) );
  CKND2D0BWP12T U1045 ( .A1(n1410), .A2(
        memory_interface_inst1_delay_data_in32[11]), .ZN(n826) );
  OAI211D0BWP12T U1046 ( .A1(n1414), .A2(n824), .B(n825), .C(n826), .ZN(
        MEMCTRL_MEM_to_mem_data[3]) );
  INR2D0BWP12T U1047 ( .A1(n1162), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[13]) );
  AOI31D0BWP12T U1048 ( .A1(n1513), .A2(n1515), .A3(n1514), .B(n1594), .ZN(
        n827) );
  NR3D0BWP12T U1049 ( .A1(n1510), .A2(n1509), .A3(n1511), .ZN(n828) );
  AOI31D0BWP12T U1050 ( .A1(n1514), .A2(n1512), .A3(n828), .B(n1626), .ZN(n829) );
  AOI211D0BWP12T U1051 ( .A1(n1516), .A2(n1523), .B(n827), .C(n829), .ZN(n1527) );
  CKND0BWP12T U1052 ( .I(RF_MEMCTRL_data_reg[12]), .ZN(n830) );
  MAOI22D0BWP12T U1053 ( .A1(n1428), .A2(
        memory_interface_inst1_delay_data_in32[28]), .B1(n1409), .B2(n1568), 
        .ZN(n831) );
  CKND2D0BWP12T U1054 ( .A1(n1410), .A2(
        memory_interface_inst1_delay_data_in32[12]), .ZN(n832) );
  OAI211D0BWP12T U1055 ( .A1(n1414), .A2(n830), .B(n831), .C(n832), .ZN(
        MEMCTRL_MEM_to_mem_data[4]) );
  INR2D0BWP12T U1056 ( .A1(n1160), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[14]) );
  MAOI22D0BWP12T U1057 ( .A1(n1155), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_2_), .B1(n1617), .B2(
        n755), .ZN(n1328) );
  CKND0BWP12T U1058 ( .I(RF_MEMCTRL_data_reg[13]), .ZN(n833) );
  MAOI22D0BWP12T U1059 ( .A1(n1428), .A2(
        memory_interface_inst1_delay_data_in32[29]), .B1(n1409), .B2(n1567), 
        .ZN(n834) );
  CKND2D0BWP12T U1060 ( .A1(n1410), .A2(
        memory_interface_inst1_delay_data_in32[13]), .ZN(n835) );
  OAI211D0BWP12T U1061 ( .A1(n1414), .A2(n833), .B(n834), .C(n835), .ZN(
        MEMCTRL_MEM_to_mem_data[5]) );
  INR2D0BWP12T U1062 ( .A1(n1133), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[15]) );
  IOA21D0BWP12T U1063 ( .A1(Instruction_Fetch_inst1_fetched_instruction_reg_8_), .A2(n1155), .B(n1158), .ZN(n836) );
  AO21D0BWP12T U1064 ( .A1(n1187), .A2(MEMCTRL_RF_IF_data_in[8]), .B(n836), 
        .Z(n1592) );
  CKND0BWP12T U1065 ( .I(RF_MEMCTRL_data_reg[14]), .ZN(n837) );
  MAOI22D0BWP12T U1066 ( .A1(n1428), .A2(
        memory_interface_inst1_delay_data_in32[30]), .B1(n1409), .B2(n1565), 
        .ZN(n838) );
  CKND2D0BWP12T U1067 ( .A1(n1410), .A2(
        memory_interface_inst1_delay_data_in32[14]), .ZN(n839) );
  OAI211D0BWP12T U1068 ( .A1(n1414), .A2(n837), .B(n838), .C(n839), .ZN(
        MEMCTRL_MEM_to_mem_data[6]) );
  INR2D0BWP12T U1069 ( .A1(n1131), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[16]) );
  CKND0BWP12T U1070 ( .I(MEMCTRL_RF_IF_data_in[6]), .ZN(n840) );
  MOAI22D0BWP12T U1071 ( .A1(n755), .A2(n840), .B1(n1155), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_6_), .ZN(n1545) );
  AN2D0BWP12T U1072 ( .A1(memory_interface_inst1_fsm_state_0_), .A2(n922), .Z(
        n1430) );
  CKND0BWP12T U1073 ( .I(RF_MEMCTRL_data_reg[15]), .ZN(n841) );
  MAOI22D0BWP12T U1074 ( .A1(n1428), .A2(
        memory_interface_inst1_delay_data_in32[31]), .B1(n1409), .B2(n1566), 
        .ZN(n842) );
  CKND2D0BWP12T U1075 ( .A1(n1410), .A2(
        memory_interface_inst1_delay_data_in32[15]), .ZN(n843) );
  OAI211D0BWP12T U1076 ( .A1(n1414), .A2(n841), .B(n842), .C(n843), .ZN(
        MEMCTRL_MEM_to_mem_data[7]) );
  INR2D0BWP12T U1077 ( .A1(n1129), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[17]) );
  INR2D0BWP12T U1078 ( .A1(n981), .B1(n1013), .ZN(n1232) );
  AOI31D0BWP12T U1079 ( .A1(memory_interface_inst1_fsm_state_0_), .A2(n917), 
        .A3(n1371), .B(n919), .ZN(n927) );
  IND2D0BWP12T U1080 ( .A1(n1215), .B1(n1216), .ZN(n1307) );
  CKND2D0BWP12T U1081 ( .A1(n1053), .A2(n1246), .ZN(n844) );
  NR3D0BWP12T U1082 ( .A1(n844), .A2(n1054), .A3(n1532), .ZN(n845) );
  AOI32D0BWP12T U1083 ( .A1(n1515), .A2(n1533), .A3(n845), .B1(n1508), .B2(
        n1533), .ZN(n1458) );
  CKND0BWP12T U1084 ( .I(n1476), .ZN(n846) );
  OR4D0BWP12T U1085 ( .A1(n963), .A2(n1025), .A3(n1097), .A4(n846), .Z(n1623)
         );
  CKND0BWP12T U1086 ( .I(n1414), .ZN(n847) );
  AOI222D0BWP12T U1087 ( .A1(n847), .A2(RF_MEMCTRL_data_reg[0]), .B1(n1412), 
        .B2(memory_interface_inst1_delay_data_in32[0]), .C1(n1428), .C2(
        memory_interface_inst1_delay_data_in32[16]), .ZN(n848) );
  IOA21D0BWP12T U1088 ( .A1(n1413), .A2(RF_MEMCTRL_data_reg[16]), .B(n848), 
        .ZN(MEMCTRL_MEM_to_mem_data[8]) );
  INR2D0BWP12T U1089 ( .A1(n1127), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[18]) );
  INR3D0BWP12T U1090 ( .A1(n972), .B1(n1012), .B2(n973), .ZN(n1510) );
  CKND0BWP12T U1091 ( .I(n1414), .ZN(n849) );
  AOI222D0BWP12T U1092 ( .A1(n849), .A2(RF_MEMCTRL_data_reg[1]), .B1(n1412), 
        .B2(memory_interface_inst1_delay_data_in32[1]), .C1(n1428), .C2(
        memory_interface_inst1_delay_data_in32[17]), .ZN(n850) );
  IOA21D0BWP12T U1093 ( .A1(RF_MEMCTRL_data_reg[17]), .A2(n1413), .B(n850), 
        .ZN(MEMCTRL_MEM_to_mem_data[9]) );
  CKND2D0BWP12T U1094 ( .A1(memory_interface_inst1_delay_addr_for_adder[0]), 
        .A2(memory_interface_inst1_delay_addr_for_adder[1]), .ZN(n851) );
  CKND0BWP12T U1095 ( .I(memory_interface_inst1_delay_addr_for_adder[1]), .ZN(
        n852) );
  AO21D0BWP12T U1096 ( .A1(n1393), .A2(n852), .B(n1400), .Z(n853) );
  AOI22D0BWP12T U1097 ( .A1(n1605), .A2(MEMCTRL_IN_address[2]), .B1(
        memory_interface_inst1_delay_addr_for_adder[2]), .B2(n853), .ZN(n854)
         );
  OAI31D0BWP12T U1098 ( .A1(n1416), .A2(
        memory_interface_inst1_delay_addr_for_adder[2]), .A3(n851), .B(n854), 
        .ZN(MEMCTRL_MEM_to_mem_address[2]) );
  INR2D0BWP12T U1099 ( .A1(n1122), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[19]) );
  CKND0BWP12T U1100 ( .I(n1334), .ZN(n855) );
  AOI222D0BWP12T U1101 ( .A1(n855), .A2(n1546), .B1(n1498), .B2(n1336), .C1(
        DEC_RF_offset_b[2]), .C2(n1627), .ZN(n856) );
  OAI222D0BWP12T U1102 ( .A1(n1624), .A2(n1315), .B1(n1328), .B2(n1358), .C1(
        n1452), .C2(n1366), .ZN(n857) );
  CKND2D0BWP12T U1103 ( .A1(n1364), .A2(n857), .ZN(n858) );
  OAI211D0BWP12T U1104 ( .A1(n1544), .A2(n1340), .B(n856), .C(n858), .ZN(
        irdecode_inst1_N993) );
  INR2D0BWP12T U1105 ( .A1(n968), .B1(n1281), .ZN(n1011) );
  IOA21D0BWP12T U1106 ( .A1(n1032), .A2(n1510), .B(n1206), .ZN(n1483) );
  ND3D0BWP12T U1107 ( .A1(n1594), .A2(n1315), .A3(n1318), .ZN(n859) );
  AOI21D0BWP12T U1108 ( .A1(n1476), .A2(n859), .B(n1521), .ZN(n1314) );
  AO22D0BWP12T U1109 ( .A1(MEMCTRL_RF_IF_data_in[4]), .A2(n1610), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_4_), .B2(n1155), .Z(
        n1338) );
  CKND0BWP12T U1110 ( .I(n1414), .ZN(n860) );
  AOI222D0BWP12T U1111 ( .A1(n860), .A2(RF_MEMCTRL_data_reg[2]), .B1(n1412), 
        .B2(memory_interface_inst1_delay_data_in32[2]), .C1(n1428), .C2(
        memory_interface_inst1_delay_data_in32[18]), .ZN(n861) );
  IOA21D0BWP12T U1112 ( .A1(RF_MEMCTRL_data_reg[18]), .A2(n1413), .B(n861), 
        .ZN(MEMCTRL_MEM_to_mem_data[10]) );
  CKND0BWP12T U1113 ( .I(memory_interface_inst1_delay_addr_for_adder[3]), .ZN(
        n862) );
  AO21D0BWP12T U1114 ( .A1(n1393), .A2(n862), .B(n1382), .Z(n863) );
  AOI22D0BWP12T U1115 ( .A1(n1605), .A2(MEMCTRL_IN_address[4]), .B1(
        memory_interface_inst1_delay_addr_for_adder[4]), .B2(n863), .ZN(n864)
         );
  OAI31D0BWP12T U1116 ( .A1(n1416), .A2(n1383), .A3(
        memory_interface_inst1_delay_addr_for_adder[4]), .B(n864), .ZN(
        MEMCTRL_MEM_to_mem_address[4]) );
  INR2D0BWP12T U1117 ( .A1(n1118), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[21]) );
  OAI211D0BWP12T U1118 ( .A1(n1323), .A2(n1500), .B(n1322), .C(n1537), .ZN(
        n865) );
  AOI31D0BWP12T U1119 ( .A1(n1324), .A2(n1361), .A3(n865), .B(n1540), .ZN(n866) );
  AOI211D0BWP12T U1120 ( .A1(DEC_ALU_alu_opcode[1]), .A2(n1627), .B(n1325), 
        .C(n866), .ZN(n867) );
  OAI31D0BWP12T U1121 ( .A1(n1326), .A2(n1625), .A3(n1346), .B(n867), .ZN(n868) );
  AO211D0BWP12T U1122 ( .A1(n1590), .A2(n1330), .B(n1327), .C(n868), .Z(
        irdecode_inst1_N965) );
  NR2D0BWP12T U1123 ( .A1(n1011), .A2(n1031), .ZN(n869) );
  OAI31D0BWP12T U1124 ( .A1(n1014), .A2(n1008), .A3(n869), .B(n1049), .ZN(n870) );
  NR3D0BWP12T U1125 ( .A1(n1486), .A2(n1485), .A3(n870), .ZN(n1036) );
  MOAI22D0BWP12T U1126 ( .A1(n919), .A2(n1578), .B1(n919), .B2(
        memory_interface_inst1_delay_first_two_bytes_out[0]), .ZN(
        MEMCTRL_RF_IF_data_in[0]) );
  MAOI22D0BWP12T U1127 ( .A1(n1155), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_5_), .B1(n1614), .B2(
        n755), .ZN(n1442) );
  CKND0BWP12T U1128 ( .I(n1414), .ZN(n871) );
  AOI222D0BWP12T U1129 ( .A1(n871), .A2(RF_MEMCTRL_data_reg[3]), .B1(n1412), 
        .B2(memory_interface_inst1_delay_data_in32[3]), .C1(n1428), .C2(
        memory_interface_inst1_delay_data_in32[19]), .ZN(n872) );
  IOA21D0BWP12T U1130 ( .A1(RF_MEMCTRL_data_reg[19]), .A2(n1413), .B(n872), 
        .ZN(MEMCTRL_MEM_to_mem_data[11]) );
  CKND0BWP12T U1131 ( .I(memory_interface_inst1_delay_addr_for_adder[7]), .ZN(
        n873) );
  AO21D0BWP12T U1132 ( .A1(n1393), .A2(n873), .B(n1392), .Z(n874) );
  AOI22D0BWP12T U1133 ( .A1(n1605), .A2(MEMCTRL_IN_address[8]), .B1(
        memory_interface_inst1_delay_addr_for_adder[8]), .B2(n874), .ZN(n875)
         );
  OAI31D0BWP12T U1134 ( .A1(n1416), .A2(n1394), .A3(
        memory_interface_inst1_delay_addr_for_adder[8]), .B(n875), .ZN(
        MEMCTRL_MEM_to_mem_address[8]) );
  INR2D0BWP12T U1135 ( .A1(n1116), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[22]) );
  CKND0BWP12T U1136 ( .I(DEC_RF_offset_b[4]), .ZN(n876) );
  AOI22D0BWP12T U1137 ( .A1(n1454), .A2(n1335), .B1(n1438), .B2(n1336), .ZN(
        n877) );
  MAOI22D0BWP12T U1138 ( .A1(n1338), .A2(n1339), .B1(n1452), .B2(n1334), .ZN(
        n878) );
  OA211D0BWP12T U1139 ( .A1(n1449), .A2(n1337), .B(n877), .C(n878), .Z(n879)
         );
  OAI222D0BWP12T U1140 ( .A1(n876), .A2(n1482), .B1(n1540), .B2(n879), .C1(
        n1625), .C2(n1340), .ZN(irdecode_inst1_N995) );
  OAI21D0BWP12T U1141 ( .A1(n1554), .A2(n1321), .B(n1320), .ZN(n880) );
  AOI22D0BWP12T U1142 ( .A1(DEC_ALU_alu_opcode[3]), .A2(n1627), .B1(n1476), 
        .B2(n880), .ZN(n881) );
  ND3D0BWP12T U1143 ( .A1(n1467), .A2(n1599), .A3(n881), .ZN(
        irdecode_inst1_N967) );
  MOAI22D0BWP12T U1144 ( .A1(n919), .A2(n1576), .B1(n919), .B2(
        memory_interface_inst1_delay_first_two_bytes_out[2]), .ZN(
        MEMCTRL_RF_IF_data_in[2]) );
  CKND0BWP12T U1145 ( .I(n1414), .ZN(n882) );
  AOI222D0BWP12T U1146 ( .A1(n882), .A2(RF_MEMCTRL_data_reg[4]), .B1(n1412), 
        .B2(memory_interface_inst1_delay_data_in32[4]), .C1(n1428), .C2(
        memory_interface_inst1_delay_data_in32[20]), .ZN(n883) );
  IOA21D0BWP12T U1147 ( .A1(RF_MEMCTRL_data_reg[20]), .A2(n1413), .B(n883), 
        .ZN(MEMCTRL_MEM_to_mem_data[12]) );
  INR2D0BWP12T U1148 ( .A1(n1091), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[23]) );
  OAI22D0BWP12T U1149 ( .A1(n1624), .A2(n1296), .B1(n1452), .B2(n1303), .ZN(
        n884) );
  CKND0BWP12T U1150 ( .I(n1300), .ZN(n885) );
  AO211D0BWP12T U1151 ( .A1(n1438), .A2(n1307), .B(n1297), .C(n885), .Z(n886)
         );
  NR4D0BWP12T U1152 ( .A1(n1298), .A2(n1299), .A3(n884), .A4(n886), .ZN(n887)
         );
  CKND2D0BWP12T U1153 ( .A1(DEC_RF_operand_a[0]), .A2(n1627), .ZN(n888) );
  OAI211D0BWP12T U1154 ( .A1(n1593), .A2(n887), .B(n1314), .C(n888), .ZN(
        irdecode_inst1_N970) );
  MOAI22D0BWP12T U1155 ( .A1(n919), .A2(n1575), .B1(n919), .B2(
        memory_interface_inst1_delay_first_two_bytes_out[3]), .ZN(
        MEMCTRL_RF_IF_data_in[3]) );
  OA21D0BWP12T U1156 ( .A1(n1593), .A2(n1016), .B(n1533), .Z(n1344) );
  CKND0BWP12T U1157 ( .I(n1320), .ZN(n889) );
  AOI21D0BWP12T U1158 ( .A1(n1536), .A2(n1094), .B(n889), .ZN(n1541) );
  MAOI22D0BWP12T U1159 ( .A1(n1155), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_1_), .B1(n1616), .B2(
        n755), .ZN(n1491) );
  IOA21D0BWP12T U1160 ( .A1(n919), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[8]), .B(n966), .ZN(
        n890) );
  AO21D0BWP12T U1161 ( .A1(MEM_MEMCTRL_from_mem_data[0]), .A2(n965), .B(n890), 
        .Z(MEMCTRL_RF_IF_data_in[8]) );
  MOAI22D0BWP12T U1162 ( .A1(n919), .A2(n1571), .B1(n919), .B2(
        memory_interface_inst1_delay_first_two_bytes_out[7]), .ZN(
        MEMCTRL_RF_IF_data_in[7]) );
  CKND0BWP12T U1163 ( .I(n1414), .ZN(n891) );
  AOI222D0BWP12T U1164 ( .A1(n891), .A2(RF_MEMCTRL_data_reg[5]), .B1(n1412), 
        .B2(memory_interface_inst1_delay_data_in32[5]), .C1(n1428), .C2(
        memory_interface_inst1_delay_data_in32[21]), .ZN(n892) );
  IOA21D0BWP12T U1165 ( .A1(RF_MEMCTRL_data_reg[21]), .A2(n1413), .B(n892), 
        .ZN(MEMCTRL_MEM_to_mem_data[13]) );
  INR2D0BWP12T U1166 ( .A1(n1186), .B1(n1185), .ZN(IF_RF_incremented_pc_out[2]) );
  INR2D0BWP12T U1167 ( .A1(n1089), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[24]) );
  OR4D0BWP12T U1168 ( .A1(n1590), .A2(n1279), .A3(n1299), .A4(n1351), .Z(n893)
         );
  AOI22D0BWP12T U1169 ( .A1(n1364), .A2(n893), .B1(DEC_ALU_alu_opcode[4]), 
        .B2(n1627), .ZN(n894) );
  AOI32D0BWP12T U1170 ( .A1(n1271), .A2(n894), .A3(n1280), .B1(n1496), .B2(
        n894), .ZN(irdecode_inst1_N968) );
  AO22D0BWP12T U1171 ( .A1(n1509), .A2(n970), .B1(n1054), .B2(n969), .Z(n1010)
         );
  OAI21D0BWP12T U1172 ( .A1(n1462), .A2(n1626), .B(n1520), .ZN(n895) );
  AOI21D0BWP12T U1173 ( .A1(n1476), .A2(n895), .B(n1521), .ZN(n1468) );
  MAOI22D0BWP12T U1174 ( .A1(n1155), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_0_), .B1(n1618), .B2(
        n755), .ZN(n1624) );
  MOAI22D0BWP12T U1175 ( .A1(n919), .A2(n1579), .B1(n919), .B2(
        memory_interface_inst1_delay_first_two_bytes_out[4]), .ZN(
        MEMCTRL_RF_IF_data_in[4]) );
  CKND0BWP12T U1176 ( .I(n1414), .ZN(n896) );
  AOI222D0BWP12T U1177 ( .A1(n896), .A2(RF_MEMCTRL_data_reg[6]), .B1(n1412), 
        .B2(memory_interface_inst1_delay_data_in32[6]), .C1(n1428), .C2(
        memory_interface_inst1_delay_data_in32[22]), .ZN(n897) );
  IOA21D0BWP12T U1178 ( .A1(RF_MEMCTRL_data_reg[22]), .A2(n1413), .B(n897), 
        .ZN(MEMCTRL_MEM_to_mem_data[14]) );
  AO222D0BWP12T U1179 ( .A1(memory_interface_inst1_delay_addr_for_adder[9]), 
        .A2(n1608), .B1(n1607), .B2(n1606), .C1(MEMCTRL_IN_address[9]), .C2(
        n1605), .Z(MEMCTRL_MEM_to_mem_address[9]) );
  CKND0BWP12T U1180 ( .I(RF_OUT_c), .ZN(n898) );
  MOAI22D0BWP12T U1181 ( .A1(DEC_CPSR_update_flag_c), .A2(n898), .B1(
        DEC_CPSR_update_flag_c), .B2(ALU_OUT_c), .ZN(new_c) );
  INR2D0BWP12T U1182 ( .A1(n1182), .B1(n1185), .ZN(IF_RF_incremented_pc_out[3]) );
  INR2D0BWP12T U1183 ( .A1(n1176), .B1(n1185), .ZN(IF_RF_incremented_pc_out[7]) );
  INR2D0BWP12T U1184 ( .A1(n1170), .B1(n1185), .ZN(IF_RF_incremented_pc_out[9]) );
  INR2D0BWP12T U1185 ( .A1(n1076), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[27]) );
  CKND0BWP12T U1186 ( .I(n1588), .ZN(n899) );
  CKND2D0BWP12T U1187 ( .A1(n1292), .A2(n1287), .ZN(n900) );
  AOI222D0BWP12T U1188 ( .A1(n899), .A2(n1498), .B1(DEC_RF_alu_write_to_reg[1]), .B2(n1627), .C1(n900), .C2(n1267), .ZN(n901) );
  IOA21D0BWP12T U1189 ( .A1(n1221), .A2(n1364), .B(n901), .ZN(
        irdecode_inst1_N976) );
  MOAI22D0BWP12T U1190 ( .A1(n919), .A2(n1577), .B1(n919), .B2(
        memory_interface_inst1_delay_first_two_bytes_out[1]), .ZN(
        MEMCTRL_RF_IF_data_in[1]) );
  MOAI22D0BWP12T U1191 ( .A1(n919), .A2(n1574), .B1(n919), .B2(
        memory_interface_inst1_delay_first_two_bytes_out[5]), .ZN(
        MEMCTRL_RF_IF_data_in[5]) );
  MOAI22D0BWP12T U1192 ( .A1(n919), .A2(n1573), .B1(n919), .B2(
        memory_interface_inst1_delay_first_two_bytes_out[6]), .ZN(
        MEMCTRL_RF_IF_data_in[6]) );
  CKND0BWP12T U1193 ( .I(n1414), .ZN(n902) );
  AOI222D0BWP12T U1194 ( .A1(n902), .A2(RF_MEMCTRL_data_reg[7]), .B1(n1412), 
        .B2(memory_interface_inst1_delay_data_in32[7]), .C1(n1428), .C2(
        memory_interface_inst1_delay_data_in32[23]), .ZN(n903) );
  IOA21D0BWP12T U1195 ( .A1(RF_MEMCTRL_data_reg[23]), .A2(n1413), .B(n903), 
        .ZN(MEMCTRL_MEM_to_mem_data[15]) );
  CKND0BWP12T U1196 ( .I(memory_interface_inst1_delay_addr_for_adder[5]), .ZN(
        n904) );
  AO21D0BWP12T U1197 ( .A1(n1393), .A2(n904), .B(n1387), .Z(n905) );
  AOI22D0BWP12T U1198 ( .A1(n1605), .A2(MEMCTRL_IN_address[6]), .B1(
        memory_interface_inst1_delay_addr_for_adder[6]), .B2(n905), .ZN(n906)
         );
  OAI31D0BWP12T U1199 ( .A1(n1416), .A2(n1388), .A3(
        memory_interface_inst1_delay_addr_for_adder[6]), .B(n906), .ZN(
        MEMCTRL_MEM_to_mem_address[6]) );
  INR2D0BWP12T U1200 ( .A1(RF_pc_out[0]), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[0]) );
  INR2D0BWP12T U1201 ( .A1(n1184), .B1(n1185), .ZN(IF_RF_incremented_pc_out[4]) );
  INR2D0BWP12T U1202 ( .A1(n1172), .B1(n1185), .ZN(IF_RF_incremented_pc_out[8]) );
  INR2D0BWP12T U1203 ( .A1(n1168), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[10]) );
  INR2D0BWP12T U1204 ( .A1(n1066), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[28]) );
  OAI21D0BWP12T U1205 ( .A1(n1516), .A2(n1525), .B(n963), .ZN(n907) );
  AOI32D0BWP12T U1206 ( .A1(n1046), .A2(n907), .A3(n1490), .B1(n1328), .B2(
        n907), .ZN(n908) );
  AOI211D0BWP12T U1207 ( .A1(n1530), .A2(n1108), .B(n1517), .C(n908), .ZN(n909) );
  AOI31D0BWP12T U1208 ( .A1(n909), .A2(n1461), .A3(n1456), .B(n1593), .ZN(n910) );
  AO211D0BWP12T U1209 ( .A1(DEC_RF_memory_write_to_reg[2]), .A2(n1627), .B(
        n910), .C(n1458), .Z(n802) );
  MUX2ND0BWP12T U1210 ( .I0(MEMCTRL_RF_IF_data_in[8]), .I1(
        Instruction_Fetch_inst1_fetched_instruction_reg_8_), .S(n755), .ZN(
        n911) );
  CKND2D0BWP12T U1211 ( .A1(n1609), .A2(n911), .ZN(Instruction_Fetch_inst1_N92) );
  INVD1BWP12T U1212 ( .I(n919), .ZN(n1581) );
  INVD1BWP12T U1213 ( .I(memory_interface_inst1_fsm_state_0_), .ZN(n916) );
  INR2D1BWP12T U1214 ( .A1(memory_interface_inst1_fsm_state_1_), .B1(
        memory_interface_inst1_fsm_state_2_), .ZN(n922) );
  INR2D0BWP12T U1215 ( .A1(n916), .B1(n922), .ZN(n913) );
  INVD1BWP12T U1216 ( .I(memory_interface_inst1_fsm_state_1_), .ZN(n917) );
  ND2D1BWP12T U1217 ( .A1(n917), .A2(memory_interface_inst1_fsm_state_2_), 
        .ZN(n918) );
  AOI21D0BWP12T U1218 ( .A1(memory_interface_inst1_fsm_state_1_), .A2(
        memory_interface_inst1_fsm_state_2_), .B(n916), .ZN(n912) );
  INVD0BWP12T U1219 ( .I(memory_interface_inst1_fsm_state_3_), .ZN(n1429) );
  AOI211D1BWP12T U1220 ( .A1(n913), .A2(n918), .B(n912), .C(n1429), .ZN(n1374)
         );
  CKND2D0BWP12T U1221 ( .A1(memory_interface_inst1_fsm_state_3_), .A2(
        memory_interface_inst1_fsm_state_0_), .ZN(n914) );
  NR2D1BWP12T U1222 ( .A1(n918), .A2(n914), .ZN(n1428) );
  NR3D1BWP12T U1223 ( .A1(n1374), .A2(n1430), .A3(n1428), .ZN(n1370) );
  NR2D1BWP12T U1224 ( .A1(memory_interface_inst1_fsm_state_2_), .A2(
        memory_interface_inst1_fsm_state_3_), .ZN(n1371) );
  INVD1BWP12T U1225 ( .I(n1371), .ZN(n915) );
  INR2D1BWP12T U1226 ( .A1(n917), .B1(n915), .ZN(n1559) );
  ND2D1BWP12T U1227 ( .A1(n1559), .A2(n916), .ZN(n1414) );
  ND2D1BWP12T U1228 ( .A1(n1370), .A2(n1414), .ZN(n1562) );
  NR2D1BWP12T U1229 ( .A1(memory_interface_inst1_fsm_state_3_), .A2(
        memory_interface_inst1_fsm_state_0_), .ZN(n921) );
  INR2D1BWP12T U1230 ( .A1(n921), .B1(n918), .ZN(n919) );
  INVD0BWP12T U1231 ( .I(n927), .ZN(n920) );
  NR2D1BWP12T U1232 ( .A1(n1562), .A2(n920), .ZN(n925) );
  NR2D1BWP12T U1233 ( .A1(n925), .A2(n919), .ZN(n965) );
  ND2D1BWP12T U1234 ( .A1(n922), .A2(n921), .ZN(n1560) );
  TPNR2D0BWP12T U1235 ( .A1(n1560), .A2(
        memory_interface_inst1_delayed_is_signed), .ZN(n923) );
  NR2D1BWP12T U1236 ( .A1(n923), .A2(MEM_MEMCTRL_from_mem_data[15]), .ZN(n924)
         );
  ND2D1BWP12T U1237 ( .A1(n925), .A2(n924), .ZN(n966) );
  IOA21D0BWP12T U1238 ( .A1(n919), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[14]), .B(n966), .ZN(
        n926) );
  AOI21D1BWP12T U1239 ( .A1(n965), .A2(MEM_MEMCTRL_from_mem_data[6]), .B(n926), 
        .ZN(n1621) );
  INVD1BWP12T U1240 ( .I(n1621), .ZN(MEMCTRL_RF_IF_data_in[14]) );
  INVD1BWP12T U1241 ( .I(Instruction_Fetch_inst1_currentState_0_), .ZN(n928)
         );
  AN2XD1BWP12T U1242 ( .A1(n928), .A2(Instruction_Fetch_inst1_currentState_1_), 
        .Z(n1187) );
  ND2D1BWP12T U1243 ( .A1(n927), .A2(n1560), .ZN(n1433) );
  IND2D1BWP12T U1244 ( .A1(n1185), .B1(n1433), .ZN(n755) );
  INVD1BWP12T U1245 ( .I(n755), .ZN(n1610) );
  NR2D1BWP12T U1246 ( .A1(Instruction_Fetch_inst1_currentState_1_), .A2(n928), 
        .ZN(n1155) );
  AOI22D1BWP12T U1247 ( .A1(MEMCTRL_RF_IF_data_in[14]), .A2(n1610), .B1(n1155), 
        .B2(Instruction_Fetch_inst1_fetched_instruction_reg_14_), .ZN(n990) );
  INVD1BWP12T U1248 ( .I(n990), .ZN(n987) );
  INVD1BWP12T U1249 ( .I(n965), .ZN(n960) );
  TPND2D0BWP12T U1250 ( .A1(n919), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[15]), .ZN(n929) );
  OAI211D1BWP12T U1251 ( .A1(n1566), .A2(n960), .B(n966), .C(n929), .ZN(
        MEMCTRL_RF_IF_data_in[15]) );
  INR2D0BWP12T U1252 ( .A1(MEMCTRL_RF_IF_data_in[15]), .B1(n1185), .ZN(n930)
         );
  NR2D1BWP12T U1253 ( .A1(n1610), .A2(n1155), .ZN(n961) );
  AOI211D1BWP12T U1254 ( .A1(n1155), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_15_), .B(n930), .C(
        n961), .ZN(n1021) );
  INVD1BWP12T U1255 ( .I(n1021), .ZN(n994) );
  TPND2D0BWP12T U1256 ( .A1(n919), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[12]), .ZN(n931) );
  OAI211D1BWP12T U1257 ( .A1(n1568), .A2(n960), .B(n966), .C(n931), .ZN(
        MEMCTRL_RF_IF_data_in[12]) );
  INR2D0BWP12T U1258 ( .A1(MEMCTRL_RF_IF_data_in[12]), .B1(n1185), .ZN(n932)
         );
  AOI211D1BWP12T U1259 ( .A1(n1155), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_12_), .B(n932), .C(
        n961), .ZN(n1472) );
  INVD1BWP12T U1260 ( .I(n1472), .ZN(n1347) );
  TPND2D0BWP12T U1261 ( .A1(n919), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[13]), .ZN(n933) );
  OAI211D1BWP12T U1262 ( .A1(n1567), .A2(n960), .B(n966), .C(n933), .ZN(
        MEMCTRL_RF_IF_data_in[13]) );
  AOI22D0BWP12T U1263 ( .A1(n1187), .A2(MEMCTRL_RF_IF_data_in[13]), .B1(n1155), 
        .B2(Instruction_Fetch_inst1_fetched_instruction_reg_13_), .ZN(n934) );
  INVD1BWP12T U1264 ( .I(n961), .ZN(n1158) );
  ND2D1BWP12T U1265 ( .A1(n934), .A2(n1158), .ZN(n988) );
  NR2XD0BWP12T U1266 ( .A1(n1347), .A2(n988), .ZN(n993) );
  ND3D1BWP12T U1267 ( .A1(n987), .A2(n994), .A3(n993), .ZN(n1626) );
  INVD1BWP12T U1268 ( .I(irdecode_inst1_itstate_6_), .ZN(n1444) );
  INVD1BWP12T U1269 ( .I(irdecode_inst1_itstate_7_), .ZN(n1443) );
  CKND2D1BWP12T U1270 ( .A1(n1444), .A2(n1443), .ZN(n936) );
  OR4XD1BWP12T U1271 ( .A1(irdecode_inst1_itstate_2_), .A2(
        irdecode_inst1_itstate_1_), .A3(irdecode_inst1_itstate_0_), .A4(
        irdecode_inst1_itstate_3_), .Z(n935) );
  NR4D0BWP12T U1272 ( .A1(irdecode_inst1_itstate_4_), .A2(
        irdecode_inst1_itstate_5_), .A3(n936), .A4(n935), .ZN(n1550) );
  INVD0BWP12T U1273 ( .I(irdecode_inst1_itstate_4_), .ZN(n950) );
  AOI32D0BWP12T U1274 ( .A1(RF_OUT_c), .A2(n1444), .A3(n1443), .B1(RF_OUT_v), 
        .B2(irdecode_inst1_itstate_6_), .ZN(n938) );
  INVD0BWP12T U1275 ( .I(RF_OUT_v), .ZN(n1098) );
  CKND1BWP12T U1276 ( .I(RF_OUT_n), .ZN(n1095) );
  AOI22D1BWP12T U1277 ( .A1(RF_OUT_v), .A2(RF_OUT_n), .B1(n1098), .B2(n1095), 
        .ZN(n1104) );
  IOA21D0BWP12T U1278 ( .A1(n1444), .A2(n1104), .B(irdecode_inst1_itstate_7_), 
        .ZN(n937) );
  INVD1BWP12T U1279 ( .I(irdecode_inst1_itstate_5_), .ZN(n1441) );
  AOI21D1BWP12T U1280 ( .A1(n938), .A2(n937), .B(n1441), .ZN(n949) );
  NR2D1BWP12T U1281 ( .A1(n1104), .A2(RF_OUT_z), .ZN(n1096) );
  NR2D0BWP12T U1282 ( .A1(n1096), .A2(n1444), .ZN(n942) );
  INVD1BWP12T U1283 ( .I(RF_OUT_c), .ZN(n1556) );
  TPNR2D0BWP12T U1284 ( .A1(n1556), .A2(RF_OUT_z), .ZN(n943) );
  INVD0BWP12T U1285 ( .I(n943), .ZN(n1105) );
  CKND0BWP12T U1286 ( .I(RF_OUT_z), .ZN(n939) );
  AOI22D0BWP12T U1287 ( .A1(irdecode_inst1_itstate_7_), .A2(n1105), .B1(n939), 
        .B2(n1443), .ZN(n940) );
  OAI32D0BWP12T U1288 ( .A1(n1444), .A2(RF_OUT_n), .A3(
        irdecode_inst1_itstate_7_), .B1(irdecode_inst1_itstate_6_), .B2(n940), 
        .ZN(n941) );
  AOI211XD0BWP12T U1289 ( .A1(irdecode_inst1_itstate_7_), .A2(n942), .B(
        irdecode_inst1_itstate_5_), .C(n941), .ZN(n948) );
  AOI22D0BWP12T U1290 ( .A1(irdecode_inst1_itstate_6_), .A2(RF_OUT_n), .B1(
        RF_OUT_z), .B2(n1444), .ZN(n945) );
  AOI32D0BWP12T U1291 ( .A1(n943), .A2(n1444), .A3(n1441), .B1(
        irdecode_inst1_itstate_6_), .B2(n1096), .ZN(n944) );
  OAI32D0BWP12T U1292 ( .A1(irdecode_inst1_itstate_7_), .A2(
        irdecode_inst1_itstate_5_), .A3(n945), .B1(n944), .B2(n1443), .ZN(n946) );
  NR2D1BWP12T U1293 ( .A1(n949), .A2(n946), .ZN(n947) );
  OAI32D1BWP12T U1294 ( .A1(n950), .A2(n949), .A3(n948), .B1(n947), .B2(
        irdecode_inst1_itstate_4_), .ZN(n951) );
  NR2D1BWP12T U1295 ( .A1(n1550), .A2(n951), .ZN(n1302) );
  ND2D1BWP12T U1296 ( .A1(irdecode_inst1_split_instruction), .A2(
        DEC_IF_stall_to_instructionfetch), .ZN(n953) );
  INVD1BWP12T U1297 ( .I(DEC_MEMCTRL_memory_load_request), .ZN(n952) );
  INVD1BWP12T U1298 ( .I(DEC_MEMCTRL_memory_store_request), .ZN(n1421) );
  OAI22D1BWP12T U1299 ( .A1(n1433), .A2(n952), .B1(n1374), .B2(n1421), .ZN(
        n954) );
  AOI211D1BWP12T U1300 ( .A1(n755), .A2(n953), .B(n954), .C(reset), .ZN(n1476)
         );
  IND2D1BWP12T U1301 ( .A1(n1302), .B1(n1476), .ZN(n1540) );
  INR2D2BWP12T U1302 ( .A1(n954), .B1(reset), .ZN(n1627) );
  NR2D1BWP12T U1303 ( .A1(n1021), .A2(n987), .ZN(n992) );
  CKND2D1BWP12T U1304 ( .A1(n992), .A2(n988), .ZN(n991) );
  OR2XD1BWP12T U1305 ( .A1(n991), .A2(n1472), .Z(n998) );
  TPND2D0BWP12T U1306 ( .A1(n919), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[10]), .ZN(n955) );
  OAI211D1BWP12T U1307 ( .A1(n1582), .A2(n960), .B(n966), .C(n955), .ZN(
        MEMCTRL_RF_IF_data_in[10]) );
  AOI22D0BWP12T U1308 ( .A1(n1187), .A2(MEMCTRL_RF_IF_data_in[10]), .B1(n1155), 
        .B2(Instruction_Fetch_inst1_fetched_instruction_reg_10_), .ZN(n956) );
  ND2D1BWP12T U1309 ( .A1(n956), .A2(n1158), .ZN(n1475) );
  IND2XD1BWP12T U1310 ( .A1(n998), .B1(n1475), .ZN(n1025) );
  TPND2D0BWP12T U1311 ( .A1(n919), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[9]), .ZN(n957) );
  OAI211D1BWP12T U1312 ( .A1(n1572), .A2(n960), .B(n966), .C(n957), .ZN(
        MEMCTRL_RF_IF_data_in[9]) );
  AOI22D0BWP12T U1313 ( .A1(n1187), .A2(MEMCTRL_RF_IF_data_in[9]), .B1(n1155), 
        .B2(Instruction_Fetch_inst1_fetched_instruction_reg_9_), .ZN(n958) );
  ND2D1BWP12T U1314 ( .A1(n958), .A2(n1158), .ZN(n1489) );
  NR2D1BWP12T U1315 ( .A1(n1025), .A2(n1489), .ZN(n1479) );
  INVD1BWP12T U1316 ( .I(n1540), .ZN(n1364) );
  ND2D1BWP12T U1317 ( .A1(n1479), .A2(n1364), .ZN(n1496) );
  TPND2D0BWP12T U1318 ( .A1(n919), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[11]), .ZN(n959) );
  OAI211D1BWP12T U1319 ( .A1(n1569), .A2(n960), .B(n966), .C(n959), .ZN(
        MEMCTRL_RF_IF_data_in[11]) );
  INR2D0BWP12T U1320 ( .A1(MEMCTRL_RF_IF_data_in[11]), .B1(n1185), .ZN(n962)
         );
  RCAOI211D0BWP12T U1321 ( .A1(n1155), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_11_), .B(n962), .C(
        n961), .ZN(n963) );
  INVD1BWP12T U1322 ( .I(MEM_MEMCTRL_from_mem_data[9]), .ZN(n1577) );
  INVD1BWP12T U1323 ( .I(MEMCTRL_RF_IF_data_in[1]), .ZN(n1616) );
  INVD1BWP12T U1324 ( .I(irdecode_inst1_next_step_1_), .ZN(n817) );
  OR2XD1BWP12T U1325 ( .A1(n1491), .A2(n817), .Z(n968) );
  INVD1BWP12T U1326 ( .I(irdecode_inst1_next_step_0_), .ZN(n816) );
  INVD1BWP12T U1327 ( .I(MEM_MEMCTRL_from_mem_data[8]), .ZN(n1578) );
  INVD1BWP12T U1328 ( .I(MEMCTRL_RF_IF_data_in[0]), .ZN(n1618) );
  NR2D1BWP12T U1329 ( .A1(n816), .A2(n1624), .ZN(n1226) );
  NR2D1BWP12T U1330 ( .A1(n968), .A2(n1226), .ZN(n1031) );
  INVD0BWP12T U1331 ( .I(n1031), .ZN(n1514) );
  INVD1BWP12T U1332 ( .I(MEM_MEMCTRL_from_mem_data[12]), .ZN(n1579) );
  ND2D1BWP12T U1333 ( .A1(n1338), .A2(irdecode_inst1_next_step_4_), .ZN(n967)
         );
  IND2D1BWP12T U1334 ( .A1(n1226), .B1(n968), .ZN(n1012) );
  INVD1BWP12T U1335 ( .I(MEM_MEMCTRL_from_mem_data[10]), .ZN(n1576) );
  INVD0BWP12T U1336 ( .I(MEMCTRL_RF_IF_data_in[2]), .ZN(n1617) );
  INVD1BWP12T U1337 ( .I(n1328), .ZN(n1454) );
  ND2D1BWP12T U1338 ( .A1(n1454), .A2(irdecode_inst1_next_step_2_), .ZN(n972)
         );
  INVD1BWP12T U1339 ( .I(MEM_MEMCTRL_from_mem_data[11]), .ZN(n1575) );
  INVD0BWP12T U1340 ( .I(MEMCTRL_RF_IF_data_in[3]), .ZN(n1615) );
  INVD1BWP12T U1341 ( .I(n1329), .ZN(n1438) );
  ND2D1BWP12T U1342 ( .A1(n1438), .A2(irdecode_inst1_next_step_3_), .ZN(n973)
         );
  ND2D1BWP12T U1343 ( .A1(n972), .A2(n973), .ZN(n1008) );
  NR2D1BWP12T U1344 ( .A1(n1012), .A2(n1008), .ZN(n964) );
  IND2D1BWP12T U1345 ( .A1(n967), .B1(n964), .ZN(n1200) );
  INVD1BWP12T U1346 ( .I(MEM_MEMCTRL_from_mem_data[13]), .ZN(n1574) );
  INVD0BWP12T U1347 ( .I(MEMCTRL_RF_IF_data_in[5]), .ZN(n1614) );
  INVD1BWP12T U1348 ( .I(n1442), .ZN(n1308) );
  ND2D1BWP12T U1349 ( .A1(n1308), .A2(irdecode_inst1_next_step_5_), .ZN(n974)
         );
  ND2D1BWP12T U1350 ( .A1(n964), .A2(n967), .ZN(n975) );
  NR2D1BWP12T U1351 ( .A1(n974), .A2(n975), .ZN(n1509) );
  INVD0BWP12T U1352 ( .I(n1509), .ZN(n1035) );
  INVD1BWP12T U1353 ( .I(n1592), .ZN(n1452) );
  INVD1BWP12T U1354 ( .I(MEM_MEMCTRL_from_mem_data[14]), .ZN(n1573) );
  ND2D1BWP12T U1355 ( .A1(n1545), .A2(irdecode_inst1_next_step_6_), .ZN(n977)
         );
  INVD1BWP12T U1356 ( .I(MEM_MEMCTRL_from_mem_data[15]), .ZN(n1571) );
  ND2D1BWP12T U1357 ( .A1(n1348), .A2(irdecode_inst1_next_step_7_), .ZN(n978)
         );
  AN2XD1BWP12T U1358 ( .A1(n977), .A2(n978), .Z(n970) );
  ND2D1BWP12T U1359 ( .A1(n970), .A2(n974), .ZN(n1018) );
  NR3D1BWP12T U1360 ( .A1(n1452), .A2(n1018), .A3(n975), .ZN(n1532) );
  INVD1BWP12T U1361 ( .I(n1018), .ZN(n969) );
  ND2D1BWP12T U1362 ( .A1(n967), .A2(n969), .ZN(n1014) );
  INVD1BWP12T U1363 ( .I(n1014), .ZN(n980) );
  INVD0BWP12T U1364 ( .I(n1226), .ZN(n1281) );
  IAO21D0BWP12T U1365 ( .A1(n1031), .A2(n1011), .B(n1008), .ZN(n971) );
  INVD1BWP12T U1366 ( .I(n1200), .ZN(n1054) );
  AOI32D1BWP12T U1367 ( .A1(n980), .A2(n1452), .A3(n971), .B1(n1010), .B2(
        n1452), .ZN(n985) );
  INVD1BWP12T U1368 ( .I(n1510), .ZN(n1513) );
  NR2D1BWP12T U1369 ( .A1(n1012), .A2(n972), .ZN(n1204) );
  ND2D0BWP12T U1370 ( .A1(n1204), .A2(n973), .ZN(n1009) );
  CKND2D1BWP12T U1371 ( .A1(n1513), .A2(n1009), .ZN(n979) );
  IND2XD1BWP12T U1372 ( .A1(n975), .B1(n974), .ZN(n976) );
  INR3XD0BWP12T U1373 ( .A1(n977), .B1(n978), .B2(n976), .ZN(n1052) );
  INVD1BWP12T U1374 ( .I(n1052), .ZN(n1512) );
  NR2D1BWP12T U1375 ( .A1(n977), .A2(n976), .ZN(n1033) );
  ND2D1BWP12T U1376 ( .A1(n1033), .A2(n978), .ZN(n1053) );
  ND2D1BWP12T U1377 ( .A1(n1512), .A2(n1053), .ZN(n1484) );
  AOI32D1BWP12T U1378 ( .A1(n980), .A2(n1452), .A3(n979), .B1(n1484), .B2(
        n1452), .ZN(n984) );
  ND2D1BWP12T U1379 ( .A1(n985), .A2(n984), .ZN(n1282) );
  NR3D1BWP12T U1380 ( .A1(n1226), .A2(n1532), .A3(n1282), .ZN(n1271) );
  INVD1BWP12T U1381 ( .I(n1271), .ZN(n1196) );
  AOI31D1BWP12T U1382 ( .A1(n1514), .A2(n1200), .A3(n1035), .B(n1196), .ZN(
        n1270) );
  NR2D1BWP12T U1383 ( .A1(n1196), .A2(n1031), .ZN(n981) );
  NR2D1BWP12T U1384 ( .A1(n1510), .A2(n1204), .ZN(n1013) );
  ND3D1BWP12T U1385 ( .A1(n981), .A2(n1013), .A3(n1200), .ZN(n1017) );
  INVD1BWP12T U1386 ( .I(n1017), .ZN(n982) );
  AOI21D1BWP12T U1387 ( .A1(n1052), .A2(n982), .B(n1232), .ZN(n983) );
  ND2D1BWP12T U1388 ( .A1(n1033), .A2(n982), .ZN(n1246) );
  ND2D1BWP12T U1389 ( .A1(n983), .A2(n1246), .ZN(n1269) );
  INR3XD0BWP12T U1390 ( .A1(n984), .B1(n1532), .B2(n1269), .ZN(n1497) );
  IND4D1BWP12T U1391 ( .A1(n1270), .B1(n985), .B2(n1497), .B3(n1281), .ZN(
        n1044) );
  CKND2D1BWP12T U1392 ( .A1(n963), .A2(n1044), .ZN(n1507) );
  NR2D1BWP12T U1393 ( .A1(n1496), .A2(n1507), .ZN(n1327) );
  AOI21D1BWP12T U1394 ( .A1(n1627), .A2(
        DEC_MISC_OUT_memory_address_source_is_reg), .B(n1327), .ZN(n986) );
  OAI21D1BWP12T U1395 ( .A1(n1626), .A2(n1540), .B(n986), .ZN(n788) );
  INVD1BWP12T U1396 ( .I(n988), .ZN(n1323) );
  ND2D0BWP12T U1397 ( .A1(n1323), .A2(n1347), .ZN(n1322) );
  OR2XD1BWP12T U1398 ( .A1(n1322), .A2(n1021), .Z(n989) );
  NR2D1BWP12T U1399 ( .A1(n987), .A2(n989), .ZN(n1518) );
  ND3D1BWP12T U1400 ( .A1(n1021), .A2(n1323), .A3(n987), .ZN(n1001) );
  NR2D1BWP12T U1401 ( .A1(n1347), .A2(n1001), .ZN(n1043) );
  INVD1BWP12T U1402 ( .I(n963), .ZN(n1500) );
  ND2XD0BWP12T U1403 ( .A1(n1043), .A2(n1500), .ZN(n1503) );
  INVD1BWP12T U1404 ( .I(n1503), .ZN(n1218) );
  NR2D1BWP12T U1405 ( .A1(n1518), .A2(n1218), .ZN(n1255) );
  TPND2D0BWP12T U1406 ( .A1(n1347), .A2(n1500), .ZN(n1326) );
  CKND2D1BWP12T U1407 ( .A1(n990), .A2(n1021), .ZN(n1015) );
  TPNR2D0BWP12T U1408 ( .A1(n988), .A2(n1015), .ZN(n1093) );
  TPOAI21D0BWP12T U1409 ( .A1(n1475), .A2(n1326), .B(n1093), .ZN(n1366) );
  CKND1BWP12T U1410 ( .I(n1489), .ZN(n1321) );
  TPND2D0BWP12T U1411 ( .A1(n1452), .A2(n1321), .ZN(n1278) );
  INVD1BWP12T U1412 ( .I(n1475), .ZN(n1449) );
  ND2D1BWP12T U1413 ( .A1(n1449), .A2(n963), .ZN(n1453) );
  NR3D1BWP12T U1414 ( .A1(n998), .A2(n1278), .A3(n1453), .ZN(n1590) );
  TPNR2D0BWP12T U1415 ( .A1(n990), .A2(n989), .ZN(n1194) );
  TPNR2D0BWP12T U1416 ( .A1(n990), .A2(n1323), .ZN(n1020) );
  ND2D1BWP12T U1417 ( .A1(n1020), .A2(n994), .ZN(n997) );
  CKND2D0BWP12T U1418 ( .A1(n1472), .A2(n963), .ZN(n1217) );
  NR2D1BWP12T U1419 ( .A1(n997), .A2(n1217), .ZN(n1239) );
  NR2D1BWP12T U1420 ( .A1(n1194), .A2(n1239), .ZN(n1300) );
  NR2D1BWP12T U1421 ( .A1(n997), .A2(n1472), .ZN(n1274) );
  INVD1BWP12T U1422 ( .I(n1274), .ZN(n1237) );
  ND2D1BWP12T U1423 ( .A1(n1300), .A2(n1237), .ZN(n1221) );
  NR2D1BWP12T U1424 ( .A1(n1347), .A2(n991), .ZN(n1219) );
  INVD1BWP12T U1425 ( .I(n1219), .ZN(n1256) );
  TPND2D0BWP12T U1426 ( .A1(n1626), .A2(n1256), .ZN(n1478) );
  CKND0BWP12T U1427 ( .I(n1478), .ZN(n1191) );
  CKND2D1BWP12T U1428 ( .A1(n993), .A2(n992), .ZN(n1340) );
  OAI211D0BWP12T U1429 ( .A1(n1323), .A2(n994), .B(n1191), .C(n1340), .ZN(n995) );
  NR4D0BWP12T U1430 ( .A1(n1479), .A2(n1590), .A3(n1221), .A4(n995), .ZN(n996)
         );
  ND3D1BWP12T U1431 ( .A1(n1255), .A2(n1366), .A3(n996), .ZN(n1082) );
  CKND2D1BWP12T U1432 ( .A1(n1500), .A2(n1449), .ZN(n1108) );
  INVD1BWP12T U1433 ( .I(n1108), .ZN(n1125) );
  AOI211D0BWP12T U1434 ( .A1(n1449), .A2(n1592), .B(n1125), .C(n1489), .ZN(
        n999) );
  TPND2D0BWP12T U1435 ( .A1(n1472), .A2(n1500), .ZN(n1092) );
  OAI22D1BWP12T U1436 ( .A1(n999), .A2(n998), .B1(n997), .B2(n1092), .ZN(n1297) );
  OAI21D0BWP12T U1437 ( .A1(n1082), .A2(n1297), .B(n1476), .ZN(n1000) );
  OR2XD1BWP12T U1438 ( .A1(n1476), .A2(n1627), .Z(n1533) );
  INVD1BWP12T U1439 ( .I(n1302), .ZN(n1016) );
  ND2D1BWP12T U1440 ( .A1(n1000), .A2(n1344), .ZN(n1190) );
  INVD1BWP12T U1441 ( .I(n1190), .ZN(n1070) );
  NR2D1BWP12T U1442 ( .A1(n1472), .A2(n1001), .ZN(n1123) );
  NR2D1BWP12T U1443 ( .A1(n1123), .A2(n1093), .ZN(n1216) );
  INVD1BWP12T U1444 ( .I(n1545), .ZN(n1447) );
  CKND2D1BWP12T U1445 ( .A1(n1043), .A2(n963), .ZN(n1296) );
  OAI22D0BWP12T U1446 ( .A1(n1216), .A2(n1447), .B1(n1329), .B2(n1296), .ZN(
        n1002) );
  AOI22D1BWP12T U1447 ( .A1(n1002), .A2(n1476), .B1(n1627), .B2(
        DEC_RF_operand_b[0]), .ZN(n1003) );
  ND2D1BWP12T U1448 ( .A1(n1070), .A2(n1003), .ZN(n784) );
  IND2XD1BWP12T U1449 ( .A1(n1453), .B1(n1043), .ZN(n1554) );
  INVD1BWP12T U1450 ( .I(n1348), .ZN(n1543) );
  OR2XD1BWP12T U1451 ( .A1(n1540), .A2(n1543), .Z(n1544) );
  NR2D1BWP12T U1452 ( .A1(n1554), .A2(n1544), .ZN(n1325) );
  TPND2D0BWP12T U1453 ( .A1(n1093), .A2(n1326), .ZN(n1337) );
  NR2D1BWP12T U1454 ( .A1(n1015), .A2(n1323), .ZN(n1339) );
  INVD1BWP12T U1455 ( .I(n1339), .ZN(n1358) );
  INVD1BWP12T U1456 ( .I(n1296), .ZN(n1305) );
  CKND2D1BWP12T U1457 ( .A1(n1475), .A2(n1305), .ZN(n1277) );
  INVD1BWP12T U1458 ( .I(n1277), .ZN(n1312) );
  NR2D1BWP12T U1459 ( .A1(n1452), .A2(n1489), .ZN(n1549) );
  ND2D1BWP12T U1460 ( .A1(n1312), .A2(n1549), .ZN(n1324) );
  OA21D1BWP12T U1461 ( .A1(n1092), .A2(n1358), .B(n1324), .Z(n1320) );
  TPND2D0BWP12T U1462 ( .A1(n1489), .A2(n1452), .ZN(n1099) );
  INVD1BWP12T U1463 ( .I(n1099), .ZN(n1547) );
  MOAI22D0BWP12T U1464 ( .A1(n1320), .A2(n1540), .B1(n1325), .B2(n1547), .ZN(
        n1005) );
  NR3D0BWP12T U1465 ( .A1(n1472), .A2(n1500), .A3(n1358), .ZN(n1272) );
  TPNR2D0BWP12T U1466 ( .A1(n1015), .A2(n1326), .ZN(n1279) );
  CKND2D0BWP12T U1467 ( .A1(n1550), .A2(n1476), .ZN(n1538) );
  CKND0BWP12T U1468 ( .I(n1538), .ZN(n1004) );
  OAI32D1BWP12T U1469 ( .A1(n1005), .A2(n1272), .A3(n1279), .B1(n1004), .B2(
        n1005), .ZN(n1551) );
  INVD1BWP12T U1470 ( .I(n1554), .ZN(n1536) );
  AOI32D0BWP12T U1471 ( .A1(n1452), .A2(n1536), .A3(n1545), .B1(n1549), .B2(
        n1536), .ZN(n1006) );
  AOI32D0BWP12T U1472 ( .A1(n1337), .A2(n1551), .A3(n1006), .B1(n1538), .B2(
        n1551), .ZN(n1007) );
  AO31D1BWP12T U1473 ( .A1(n1325), .A2(n1550), .A3(n1321), .B(n1007), .Z(
        irdecode_inst1_next_update_flag_c) );
  CKND2D0BWP12T U1474 ( .A1(n1430), .A2(memory_interface_inst1_fsm_state_3_), 
        .ZN(n1373) );
  INVD1BWP12T U1475 ( .I(n1373), .ZN(n1423) );
  NR2D0BWP12T U1476 ( .A1(n1423), .A2(n1428), .ZN(n1411) );
  AOI211D0BWP12T U1477 ( .A1(DEC_MEMCTRL_load_store_width[0]), .A2(
        DEC_MEMCTRL_load_store_width[1]), .B(n1414), .C(reset), .ZN(n1173) );
  NR2D0BWP12T U1478 ( .A1(Instruction_Fetch_inst1_currentState_1_), .A2(
        DEC_MEMCTRL_memory_load_request), .ZN(n1422) );
  ND3XD0BWP12T U1479 ( .A1(n1173), .A2(DEC_MEMCTRL_memory_store_request), .A3(
        n1422), .ZN(n1432) );
  OAI21D0BWP12T U1480 ( .A1(reset), .A2(n1411), .B(n1432), .ZN(
        memory_interface_inst1_fsm_N35) );
  INVD1BWP12T U1481 ( .I(n1533), .ZN(n1521) );
  TPNR2D0BWP12T U1482 ( .A1(n1014), .A2(n1009), .ZN(n1486) );
  INVD0BWP12T U1483 ( .I(n1010), .ZN(n1049) );
  TPNR2D0BWP12T U1484 ( .A1(n1014), .A2(n1513), .ZN(n1485) );
  CKND2D1BWP12T U1485 ( .A1(n1036), .A2(n1053), .ZN(n1029) );
  NR2D1BWP12T U1486 ( .A1(n1012), .A2(n1029), .ZN(n1032) );
  CKND2D1BWP12T U1487 ( .A1(n1013), .A2(n1032), .ZN(n1034) );
  NR2D1BWP12T U1488 ( .A1(n1014), .A2(n1034), .ZN(n1511) );
  INVD1BWP12T U1489 ( .I(n1511), .ZN(n1462) );
  ND3D1BWP12T U1490 ( .A1(n1123), .A2(n1489), .A3(n1453), .ZN(n1046) );
  INVD1BWP12T U1491 ( .I(n1046), .ZN(n1524) );
  INVD1BWP12T U1492 ( .I(n1015), .ZN(n1537) );
  TPNR3D0BWP12T U1493 ( .A1(n1043), .A2(n1590), .A3(n1537), .ZN(n1022) );
  NR2D1BWP12T U1494 ( .A1(n1221), .A2(n1297), .ZN(n1290) );
  TPND3D0BWP12T U1495 ( .A1(n1022), .A2(n1290), .A3(n1016), .ZN(n1470) );
  NR4D0BWP12T U1496 ( .A1(n1524), .A2(n1219), .A3(n1500), .A4(n1470), .ZN(
        n1520) );
  CKND2D1BWP12T U1497 ( .A1(n1476), .A2(n1479), .ZN(n1508) );
  INVD1BWP12T U1498 ( .I(n1508), .ZN(n1531) );
  NR2D1BWP12T U1499 ( .A1(n1018), .A2(n1017), .ZN(n1504) );
  OR2XD1BWP12T U1500 ( .A1(n1532), .A2(n1504), .Z(n1464) );
  TPAOI22D0BWP12T U1501 ( .A1(n1627), .A2(DEC_RF_memory_store_data_reg[3]), 
        .B1(n1531), .B2(n1464), .ZN(n1019) );
  ND2D1BWP12T U1502 ( .A1(n1468), .A2(n1019), .ZN(n797) );
  TPND2D0BWP12T U1503 ( .A1(n1021), .A2(n1020), .ZN(n1334) );
  ND2D1BWP12T U1504 ( .A1(n1340), .A2(n1334), .ZN(n1215) );
  TPNR2D0BWP12T U1505 ( .A1(n1123), .A2(n1215), .ZN(n1057) );
  INVD1BWP12T U1506 ( .I(n1518), .ZN(n1028) );
  ND3D1BWP12T U1507 ( .A1(n1022), .A2(n1057), .A3(n1028), .ZN(n1192) );
  CKND2D1BWP12T U1508 ( .A1(n1290), .A2(n1256), .ZN(n1048) );
  NR2D1BWP12T U1509 ( .A1(n1192), .A2(n1048), .ZN(n1235) );
  ND2XD0BWP12T U1510 ( .A1(n1627), .A2(DEC_RF_memory_store_address_reg[4]), 
        .ZN(n1023) );
  OAI211D0BWP12T U1511 ( .A1(n1235), .A2(n1593), .B(n1344), .C(n1023), .ZN(
        n793) );
  ND4D1BWP12T U1512 ( .A1(n1491), .A2(n1624), .A3(n1329), .A4(n1328), .ZN(
        n1024) );
  TPND2D0BWP12T U1513 ( .A1(n1592), .A2(n1489), .ZN(n1097) );
  INR2D1BWP12T U1514 ( .A1(n1024), .B1(n1623), .ZN(n1439) );
  OAI22D1BWP12T U1515 ( .A1(n1623), .A2(n1024), .B1(reset), .B2(n1476), .ZN(
        n1622) );
  TPNR3D0BWP12T U1516 ( .A1(irdecode_inst1_itstate_2_), .A2(
        irdecode_inst1_itstate_1_), .A3(irdecode_inst1_itstate_0_), .ZN(n1027)
         );
  TPNR3D0BWP12T U1517 ( .A1(n963), .A2(n1025), .A3(n1097), .ZN(n1026) );
  AOI211D1BWP12T U1518 ( .A1(irdecode_inst1_itstate_3_), .A2(n1027), .B(n1593), 
        .C(n1026), .ZN(n1440) );
  AO222D1BWP12T U1519 ( .A1(n1338), .A2(n1439), .B1(n1622), .B2(
        irdecode_inst1_itstate_4_), .C1(irdecode_inst1_itstate_3_), .C2(n1440), 
        .Z(n809) );
  AOI21D1BWP12T U1520 ( .A1(n1321), .A2(n1123), .B(n1215), .ZN(n1490) );
  CKND2D1BWP12T U1521 ( .A1(n1490), .A2(n1028), .ZN(n1041) );
  INVD1BWP12T U1522 ( .I(n1123), .ZN(n1474) );
  NR2D1BWP12T U1523 ( .A1(n1453), .A2(n1474), .ZN(n1517) );
  RCAOI21D0BWP12T U1524 ( .A1(n963), .A2(n1041), .B(n1517), .ZN(n1460) );
  CKND0BWP12T U1525 ( .I(n1029), .ZN(n1030) );
  OAI21D0BWP12T U1526 ( .A1(n1226), .A2(n1031), .B(n1030), .ZN(n1197) );
  CKND2D0BWP12T U1527 ( .A1(n1204), .A2(n1032), .ZN(n1206) );
  CKND0BWP12T U1528 ( .I(n1033), .ZN(n1487) );
  AOI31D0BWP12T U1529 ( .A1(n1035), .A2(n1487), .A3(n1200), .B(n1034), .ZN(
        n1051) );
  INR3D0BWP12T U1530 ( .A1(n1197), .B1(n1483), .B2(n1051), .ZN(n1040) );
  NR3XD0BWP12T U1531 ( .A1(n1040), .A2(n1626), .A3(n1540), .ZN(n1284) );
  AOI211D1BWP12T U1532 ( .A1(n1627), .A2(DEC_MEMCTRL_memory_store_request), 
        .B(n1284), .C(n1327), .ZN(n1038) );
  INVD1BWP12T U1533 ( .I(n1626), .ZN(n1493) );
  INVD0BWP12T U1534 ( .I(n1036), .ZN(n1039) );
  AOI32D0BWP12T U1535 ( .A1(n963), .A2(n1493), .A3(n1039), .B1(n1484), .B2(
        n1493), .ZN(n1037) );
  AOI32D0BWP12T U1536 ( .A1(n1460), .A2(n1038), .A3(n1037), .B1(n1540), .B2(
        n1038), .ZN(n814) );
  TPNR2D0BWP12T U1537 ( .A1(n1484), .A2(n1039), .ZN(n1211) );
  AOI21D0BWP12T U1538 ( .A1(n1211), .A2(n1040), .B(n1626), .ZN(n1042) );
  TPOAI31D0BWP12T U1539 ( .A1(n1043), .A2(n1042), .A3(n1041), .B(n1500), .ZN(
        n1045) );
  IND3D1BWP12T U1540 ( .A1(n1496), .B1(n1500), .B2(n1044), .ZN(n1354) );
  AOI31D1BWP12T U1541 ( .A1(n1045), .A2(n1046), .A3(n1354), .B(n1540), .ZN(
        n1542) );
  AO21D0BWP12T U1542 ( .A1(n1627), .A2(DEC_RF_memory_write_to_reg_enable), .B(
        n1542), .Z(n799) );
  INVD0BWP12T U1543 ( .I(n1255), .ZN(n1530) );
  INVD1BWP12T U1544 ( .I(n1490), .ZN(n1516) );
  INVD1BWP12T U1545 ( .I(n1479), .ZN(n1594) );
  CKND2D0BWP12T U1546 ( .A1(n1626), .A2(n1594), .ZN(n1525) );
  INVD1BWP12T U1547 ( .I(n1590), .ZN(n1349) );
  ND2D0BWP12T U1548 ( .A1(n1349), .A2(n1296), .ZN(n1047) );
  NR4D0BWP12T U1549 ( .A1(n1302), .A2(n1537), .A3(n1048), .A4(n1047), .ZN(
        n1461) );
  CKND2D0BWP12T U1550 ( .A1(n1049), .A2(n1462), .ZN(n1050) );
  TPOAI31D0BWP12T U1551 ( .A1(n1484), .A2(n1051), .A3(n1050), .B(n1493), .ZN(
        n1456) );
  NR3D1BWP12T U1552 ( .A1(n1052), .A2(n1509), .A3(n1504), .ZN(n1515) );
  RCIAO22D1BWP12T U1553 ( .B1(n1055), .B2(RF_pc_out[31]), .A1(n1055), .A2(
        RF_pc_out[31]), .ZN(n1056) );
  INR2XD0BWP12T U1554 ( .A1(n1056), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[31]) );
  ND2D1BWP12T U1555 ( .A1(n1057), .A2(n1255), .ZN(n1291) );
  NR2D1BWP12T U1556 ( .A1(n1297), .A2(n1291), .ZN(n1587) );
  NR2D1BWP12T U1557 ( .A1(n816), .A2(n1237), .ZN(n1299) );
  ND2D1BWP12T U1558 ( .A1(n1299), .A2(n1500), .ZN(n1361) );
  AOI21D0BWP12T U1559 ( .A1(n1545), .A2(n1543), .B(n1099), .ZN(n1094) );
  AOI31D1BWP12T U1560 ( .A1(n1587), .A2(n1361), .A3(n1541), .B(n1593), .ZN(
        n1058) );
  INVD1BWP12T U1561 ( .I(n1344), .ZN(n1288) );
  AO211D0BWP12T U1562 ( .A1(n1627), .A2(DEC_RF_alu_write_to_reg[4]), .B(n1058), 
        .C(n1288), .Z(irdecode_inst1_N979) );
  HA1D0BWP12T U1563 ( .A(n1059), .B(RF_pc_out[30]), .CO(n1055), .S(n1060) );
  INR2XD0BWP12T U1564 ( .A1(n1060), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[30]) );
  NR4D0BWP12T U1565 ( .A1(RF_pc_out[4]), .A2(RF_pc_out[3]), .A3(RF_pc_out[2]), 
        .A4(RF_pc_out[1]), .ZN(n1073) );
  IND2XD1BWP12T U1566 ( .A1(RF_pc_out[5]), .B1(n1073), .ZN(n1085) );
  NR2XD0BWP12T U1567 ( .A1(RF_pc_out[6]), .A2(n1085), .ZN(n1071) );
  IND2D1BWP12T U1568 ( .A1(RF_pc_out[7]), .B1(n1071), .ZN(n1074) );
  NR2XD0BWP12T U1569 ( .A1(RF_pc_out[8]), .A2(n1074), .ZN(n1067) );
  IND2D1BWP12T U1570 ( .A1(RF_pc_out[9]), .B1(n1067), .ZN(n1072) );
  TPNR2D0BWP12T U1571 ( .A1(RF_pc_out[10]), .A2(n1072), .ZN(n1064) );
  IND2XD0BWP12T U1572 ( .A1(RF_pc_out[11]), .B1(n1064), .ZN(n1061) );
  MOAI22D0BWP12T U1573 ( .A1(RF_pc_out[12]), .A2(n1061), .B1(RF_pc_out[12]), 
        .B2(n1061), .ZN(n1138) );
  NR2D1BWP12T U1574 ( .A1(Instruction_Fetch_inst1_currentState_1_), .A2(
        DEC_MISC_OUT_memory_address_source_is_reg), .ZN(n1086) );
  INR2XD0BWP12T U1575 ( .A1(DEC_MISC_OUT_memory_address_source_is_reg), .B1(
        Instruction_Fetch_inst1_currentState_1_), .ZN(n1087) );
  AO222D0BWP12T U1576 ( .A1(n1187), .A2(n1138), .B1(ALU_MISC_OUT_result[12]), 
        .B2(n1086), .C1(n1087), .C2(RF_MEMCTRL_address_reg[12]), .Z(
        MEMCTRL_IN_address[11]) );
  HA1D0BWP12T U1577 ( .A(n1062), .B(RF_pc_out[29]), .CO(n1059), .S(n1063) );
  INR2D0BWP12T U1578 ( .A1(n1063), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[29]) );
  AO222D0BWP12T U1579 ( .A1(n1187), .A2(n1137), .B1(n1087), .B2(
        RF_MEMCTRL_address_reg[11]), .C1(ALU_MISC_OUT_result[11]), .C2(n1086), 
        .Z(MEMCTRL_IN_address[10]) );
  HA1D0BWP12T U1580 ( .A(n1065), .B(RF_pc_out[28]), .CO(n1062), .S(n1066) );
  AO222D0BWP12T U1581 ( .A1(n1187), .A2(n1144), .B1(n1087), .B2(
        RF_MEMCTRL_address_reg[9]), .C1(ALU_MISC_OUT_result[9]), .C2(n1086), 
        .Z(MEMCTRL_IN_address[8]) );
  OAI22D0BWP12T U1582 ( .A1(n1216), .A2(n1452), .B1(n1296), .B2(n1442), .ZN(
        n1068) );
  AOI22D0BWP12T U1583 ( .A1(n1068), .A2(n1476), .B1(n1627), .B2(
        DEC_RF_operand_b[2]), .ZN(n1069) );
  CKND2D1BWP12T U1584 ( .A1(n1070), .A2(n1069), .ZN(n782) );
  AO222D0BWP12T U1585 ( .A1(n1187), .A2(n1145), .B1(n1087), .B2(
        RF_MEMCTRL_address_reg[7]), .C1(ALU_MISC_OUT_result[7]), .C2(n1086), 
        .Z(MEMCTRL_IN_address[6]) );
  INVD0BWP12T U1586 ( .I(RF_pc_out[1]), .ZN(n1188) );
  AO222D0BWP12T U1587 ( .A1(n1187), .A2(n1135), .B1(n1087), .B2(
        RF_MEMCTRL_address_reg[2]), .C1(ALU_MISC_OUT_result[2]), .C2(n1086), 
        .Z(MEMCTRL_IN_address[1]) );
  MOAI22D0BWP12T U1588 ( .A1(RF_pc_out[10]), .A2(n1072), .B1(RF_pc_out[10]), 
        .B2(n1072), .ZN(n1136) );
  AO222D0BWP12T U1589 ( .A1(n1187), .A2(n1136), .B1(n1087), .B2(
        RF_MEMCTRL_address_reg[10]), .C1(ALU_MISC_OUT_result[10]), .C2(n1086), 
        .Z(MEMCTRL_IN_address[9]) );
  AO222D0BWP12T U1590 ( .A1(n1187), .A2(n1140), .B1(n1087), .B2(
        RF_MEMCTRL_address_reg[5]), .C1(ALU_MISC_OUT_result[5]), .C2(n1086), 
        .Z(MEMCTRL_IN_address[4]) );
  MOAI22D0BWP12T U1591 ( .A1(RF_pc_out[8]), .A2(n1074), .B1(RF_pc_out[8]), 
        .B2(n1074), .ZN(n1142) );
  AO222D0BWP12T U1592 ( .A1(n1187), .A2(n1142), .B1(n1087), .B2(
        RF_MEMCTRL_address_reg[8]), .C1(ALU_MISC_OUT_result[8]), .C2(n1086), 
        .Z(MEMCTRL_IN_address[7]) );
  HA1D0BWP12T U1593 ( .A(n1075), .B(RF_pc_out[27]), .CO(n1065), .S(n1076) );
  AO21D0BWP12T U1594 ( .A1(n1627), .A2(DEC_RF_operand_b[4]), .B(n1190), .Z(
        n779) );
  AO222D0BWP12T U1595 ( .A1(n1187), .A2(n1141), .B1(n1087), .B2(
        RF_MEMCTRL_address_reg[3]), .C1(ALU_MISC_OUT_result[3]), .C2(n1086), 
        .Z(MEMCTRL_IN_address[2]) );
  NR3D0BWP12T U1596 ( .A1(RF_pc_out[3]), .A2(RF_pc_out[2]), .A3(RF_pc_out[1]), 
        .ZN(n1077) );
  AO222D0BWP12T U1597 ( .A1(n1187), .A2(n1139), .B1(n1087), .B2(
        RF_MEMCTRL_address_reg[4]), .C1(ALU_MISC_OUT_result[4]), .C2(n1086), 
        .Z(MEMCTRL_IN_address[3]) );
  HA1D0BWP12T U1598 ( .A(n1078), .B(RF_pc_out[26]), .CO(n1075), .S(n1079) );
  INR2D0BWP12T U1599 ( .A1(n1079), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[26]) );
  HA1D0BWP12T U1600 ( .A(n1080), .B(RF_pc_out[25]), .CO(n1078), .S(n1081) );
  INR2D0BWP12T U1601 ( .A1(n1081), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[25]) );
  INVD1BWP12T U1602 ( .I(DEC_RF_operand_b[1]), .ZN(n1084) );
  INVD1BWP12T U1603 ( .I(n1627), .ZN(n1482) );
  AOI21D0BWP12T U1604 ( .A1(n1305), .A2(n1338), .B(n1082), .ZN(n1083) );
  OAI222D0BWP12T U1605 ( .A1(n1084), .A2(n1482), .B1(n1540), .B2(n1083), .C1(
        n1544), .C2(n1216), .ZN(n783) );
  MOAI22D0BWP12T U1606 ( .A1(RF_pc_out[6]), .A2(n1085), .B1(RF_pc_out[6]), 
        .B2(n1085), .ZN(n1143) );
  AO222D0BWP12T U1607 ( .A1(n1187), .A2(n1143), .B1(n1087), .B2(
        RF_MEMCTRL_address_reg[6]), .C1(ALU_MISC_OUT_result[6]), .C2(n1086), 
        .Z(MEMCTRL_IN_address[5]) );
  HA1D0BWP12T U1608 ( .A(n1088), .B(RF_pc_out[24]), .CO(n1080), .S(n1089) );
  INVD0BWP12T U1609 ( .I(n1297), .ZN(n1317) );
  IND4D1BWP12T U1610 ( .A1(n1192), .B1(n1300), .B2(n1317), .B3(n1256), .ZN(
        n1210) );
  NR2D1BWP12T U1611 ( .A1(n1274), .A2(n1210), .ZN(n1242) );
  AOI32D1BWP12T U1612 ( .A1(n1242), .A2(n1344), .A3(n1594), .B1(n1593), .B2(
        n1344), .ZN(n1450) );
  AO21D0BWP12T U1613 ( .A1(n1627), .A2(DEC_RF_memory_store_address_reg[3]), 
        .B(n1450), .Z(n792) );
  HA1D0BWP12T U1614 ( .A(n1090), .B(RF_pc_out[23]), .CO(n1088), .S(n1091) );
  AOI21D0BWP12T U1615 ( .A1(n1092), .A2(n1339), .B(n1478), .ZN(n1292) );
  OAI21D0BWP12T U1616 ( .A1(n1549), .A2(n1277), .B(n1292), .ZN(n1342) );
  CKND0BWP12T U1617 ( .I(n1093), .ZN(n1346) );
  OAI21D0BWP12T U1618 ( .A1(n1094), .A2(n1554), .B(n1346), .ZN(n1207) );
  OAI221D0BWP12T U1619 ( .A1(RF_OUT_v), .A2(n1099), .B1(n1098), .B2(n1097), 
        .C(n1475), .ZN(n1100) );
  AOI221D0BWP12T U1620 ( .A1(n963), .A2(n1102), .B1(n1500), .B2(n1101), .C(
        n1100), .ZN(n1111) );
  AOI22D0BWP12T U1621 ( .A1(n1321), .A2(RF_OUT_z), .B1(RF_OUT_c), .B2(n1489), 
        .ZN(n1103) );
  AOI22D0BWP12T U1622 ( .A1(n1321), .A2(n1105), .B1(n1104), .B2(n1489), .ZN(
        n1106) );
  OAI22D0BWP12T U1623 ( .A1(n1453), .A2(n1109), .B1(n1108), .B2(n1107), .ZN(
        n1110) );
  OA21D0BWP12T U1624 ( .A1(n1111), .A2(n1110), .B(n1194), .Z(n1112) );
  OR4D1BWP12T U1625 ( .A1(n1207), .A2(n1239), .A3(n1274), .A4(n1112), .Z(n1113) );
  TPOAI31D0BWP12T U1626 ( .A1(n1590), .A2(n1342), .A3(n1113), .B(n1364), .ZN(
        n1114) );
  CKND2D1BWP12T U1627 ( .A1(n1114), .A2(n1496), .ZN(
        irdecode_inst1_next_alu_write_to_reg_enable) );
  HA1D0BWP12T U1628 ( .A(n1115), .B(RF_pc_out[22]), .CO(n1090), .S(n1116) );
  HA1D0BWP12T U1629 ( .A(n1117), .B(RF_pc_out[21]), .CO(n1115), .S(n1118) );
  HA1D1BWP12T U1630 ( .A(n1119), .B(RF_pc_out[20]), .CO(n1117), .S(n1120) );
  INR2D0BWP12T U1631 ( .A1(n1120), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[20]) );
  HA1D1BWP12T U1632 ( .A(n1121), .B(RF_pc_out[19]), .CO(n1119), .S(n1122) );
  INR2XD0BWP12T U1633 ( .A1(n1489), .B1(n1540), .ZN(n1267) );
  TPND2D0BWP12T U1634 ( .A1(n1123), .A2(n1267), .ZN(n1628) );
  INVD0BWP12T U1635 ( .I(DEC_MEMCTRL_load_store_width[0]), .ZN(n1124) );
  OAI222D0BWP12T U1636 ( .A1(n1540), .A2(n1340), .B1(n1628), .B2(n1125), .C1(
        n1482), .C2(n1124), .ZN(n786) );
  HA1D1BWP12T U1637 ( .A(n1126), .B(RF_pc_out[18]), .CO(n1121), .S(n1127) );
  HA1D0BWP12T U1638 ( .A(n1128), .B(RF_pc_out[17]), .CO(n1126), .S(n1129) );
  HA1D0BWP12T U1639 ( .A(n1130), .B(RF_pc_out[16]), .CO(n1128), .S(n1131) );
  HA1D0BWP12T U1640 ( .A(n1132), .B(RF_pc_out[15]), .CO(n1130), .S(n1133) );
  OR4D0BWP12T U1641 ( .A1(RF_pc_out[15]), .A2(RF_pc_out[18]), .A3(
        RF_pc_out[20]), .A4(RF_pc_out[19]), .Z(n1134) );
  NR4D0BWP12T U1642 ( .A1(n1135), .A2(RF_pc_out[17]), .A3(RF_pc_out[16]), .A4(
        n1134), .ZN(n1153) );
  NR4D0BWP12T U1643 ( .A1(RF_pc_out[14]), .A2(RF_pc_out[13]), .A3(
        RF_pc_out[27]), .A4(RF_pc_out[26]), .ZN(n1152) );
  NR4D0BWP12T U1644 ( .A1(RF_pc_out[25]), .A2(RF_pc_out[24]), .A3(
        RF_pc_out[23]), .A4(RF_pc_out[22]), .ZN(n1151) );
  NR4D0BWP12T U1645 ( .A1(n1138), .A2(n1137), .A3(n1136), .A4(RF_pc_out[28]), 
        .ZN(n1149) );
  NR4D0BWP12T U1646 ( .A1(RF_pc_out[31]), .A2(RF_pc_out[30]), .A3(
        RF_pc_out[21]), .A4(RF_pc_out[29]), .ZN(n1148) );
  NR4D0BWP12T U1647 ( .A1(n1141), .A2(n1140), .A3(n1139), .A4(n1188), .ZN(
        n1147) );
  NR4D0BWP12T U1648 ( .A1(n1145), .A2(n1144), .A3(n1143), .A4(n1142), .ZN(
        n1146) );
  AN4XD1BWP12T U1649 ( .A1(n1149), .A2(n1148), .A3(n1147), .A4(n1146), .Z(
        n1150) );
  AN4XD1BWP12T U1650 ( .A1(n1153), .A2(n1152), .A3(n1151), .A4(n1150), .Z(
        n1434) );
  TPND3D0BWP12T U1651 ( .A1(n1187), .A2(
        Instruction_Fetch_inst1_first_instruction_fetched), .A3(n1434), .ZN(
        n1157) );
  OAI21D0BWP12T U1652 ( .A1(Instruction_Fetch_inst1_currentState_1_), .A2(
        DEC_IF_stall_to_instructionfetch), .B(
        Instruction_Fetch_inst1_currentState_0_), .ZN(n1154) );
  AOI31D0BWP12T U1653 ( .A1(n1157), .A2(n755), .A3(n1154), .B(reset), .ZN(
        Instruction_Fetch_inst1_N79) );
  CKND0BWP12T U1654 ( .I(DEC_IF_stall_to_instructionfetch), .ZN(n1261) );
  CKND2D0BWP12T U1655 ( .A1(n1155), .A2(n1261), .ZN(n1156) );
  TPAOI31D0BWP12T U1656 ( .A1(n1158), .A2(n1157), .A3(n1156), .B(reset), .ZN(
        Instruction_Fetch_inst1_N80) );
  HA1D0BWP12T U1657 ( .A(n1159), .B(RF_pc_out[14]), .CO(n1132), .S(n1160) );
  HA1D1BWP12T U1658 ( .A(n1161), .B(RF_pc_out[13]), .CO(n1159), .S(n1162) );
  INVD1BWP12T U1659 ( .I(reset), .ZN(n1609) );
  AO221D0BWP12T U1660 ( .A1(n1610), .A2(MEMCTRL_RF_IF_data_in[13]), .B1(n755), 
        .B2(Instruction_Fetch_inst1_fetched_instruction_reg_13_), .C(reset), 
        .Z(Instruction_Fetch_inst1_N97) );
  AO221D0BWP12T U1661 ( .A1(n1610), .A2(MEMCTRL_RF_IF_data_in[10]), .B1(n755), 
        .B2(Instruction_Fetch_inst1_fetched_instruction_reg_10_), .C(reset), 
        .Z(Instruction_Fetch_inst1_N94) );
  HA1D1BWP12T U1662 ( .A(n1163), .B(RF_pc_out[12]), .CO(n1161), .S(n1164) );
  INR2D0BWP12T U1663 ( .A1(n1164), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[12]) );
  AO221D0BWP12T U1664 ( .A1(n755), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_12_), .B1(n1610), .B2(
        MEMCTRL_RF_IF_data_in[12]), .C(reset), .Z(Instruction_Fetch_inst1_N96)
         );
  AO221D0BWP12T U1665 ( .A1(n755), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_11_), .B1(n1610), .B2(
        MEMCTRL_RF_IF_data_in[11]), .C(reset), .Z(Instruction_Fetch_inst1_N95)
         );
  AO221D0BWP12T U1666 ( .A1(n1610), .A2(MEMCTRL_RF_IF_data_in[9]), .B1(n755), 
        .B2(Instruction_Fetch_inst1_fetched_instruction_reg_9_), .C(reset), 
        .Z(Instruction_Fetch_inst1_N93) );
  AO221D0BWP12T U1667 ( .A1(n755), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_15_), .B1(n1610), .B2(
        MEMCTRL_RF_IF_data_in[15]), .C(reset), .Z(Instruction_Fetch_inst1_N99)
         );
  HA1D1BWP12T U1668 ( .A(n1165), .B(RF_pc_out[11]), .CO(n1163), .S(n1166) );
  INR2D0BWP12T U1669 ( .A1(n1166), .B1(n1185), .ZN(
        IF_RF_incremented_pc_out[11]) );
  HA1D1BWP12T U1670 ( .A(n1167), .B(RF_pc_out[10]), .CO(n1165), .S(n1168) );
  HA1D1BWP12T U1671 ( .A(n1169), .B(RF_pc_out[9]), .CO(n1167), .S(n1170) );
  HA1D1BWP12T U1672 ( .A(n1171), .B(RF_pc_out[8]), .CO(n1169), .S(n1172) );
  NR2D1BWP12T U1673 ( .A1(DEC_MEMCTRL_load_store_width[0]), .A2(
        DEC_MEMCTRL_load_store_width[1]), .ZN(n1601) );
  CKND0BWP12T U1674 ( .I(n1173), .ZN(n1174) );
  OAI31D0BWP12T U1675 ( .A1(n1601), .A2(n1422), .A3(n1174), .B(n1432), .ZN(
        memory_interface_inst1_fsm_N32) );
  HA1D1BWP12T U1676 ( .A(n1175), .B(RF_pc_out[7]), .CO(n1171), .S(n1176) );
  HA1D0BWP12T U1677 ( .A(n1177), .B(RF_pc_out[6]), .CO(n1175), .S(n1178) );
  INR2D0BWP12T U1678 ( .A1(n1178), .B1(n1185), .ZN(IF_RF_incremented_pc_out[6]) );
  HA1D0BWP12T U1679 ( .A(n1179), .B(RF_pc_out[5]), .CO(n1177), .S(n1180) );
  INR2D0BWP12T U1680 ( .A1(n1180), .B1(n1185), .ZN(IF_RF_incremented_pc_out[5]) );
  HA1D0BWP12T U1681 ( .A(n1181), .B(RF_pc_out[3]), .CO(n1183), .S(n1182) );
  HA1D0BWP12T U1682 ( .A(n1183), .B(RF_pc_out[4]), .CO(n1179), .S(n1184) );
  HA1D0BWP12T U1683 ( .A(RF_pc_out[1]), .B(RF_pc_out[2]), .CO(n1181), .S(n1186) );
  AN2XD0BWP12T U1684 ( .A1(n1188), .A2(n1187), .Z(MEMCTRL_IN_address[0]) );
  NR3D0BWP12T U1685 ( .A1(n1447), .A2(n1277), .A3(n1593), .ZN(n1189) );
  AO211D0BWP12T U1686 ( .A1(n1627), .A2(DEC_RF_operand_b[3]), .B(n1190), .C(
        n1189), .Z(n781) );
  NR2D0BWP12T U1687 ( .A1(n1500), .A2(n1237), .ZN(n1298) );
  CKND2D0BWP12T U1688 ( .A1(n1300), .A2(n1191), .ZN(n1273) );
  OR3XD0BWP12T U1689 ( .A1(n1479), .A2(n1192), .A3(n1273), .Z(n1259) );
  NR4D0BWP12T U1690 ( .A1(irdecode_inst1_N755), .A2(n1298), .A3(n1259), .A4(
        n1540), .ZN(n1193) );
  ND2D1BWP12T U1691 ( .A1(n1193), .A2(n1317), .ZN(irdecode_inst1_N969) );
  ND2D1BWP12T U1692 ( .A1(n1364), .A2(n1298), .ZN(n1254) );
  INVD1BWP12T U1693 ( .I(n1254), .ZN(n1230) );
  AOI22D1BWP12T U1694 ( .A1(n1627), .A2(DEC_RF_offset_b[22]), .B1(n1475), .B2(
        n1230), .ZN(n1195) );
  INVD1BWP12T U1695 ( .I(n1544), .ZN(n1330) );
  ND2D1BWP12T U1696 ( .A1(n1330), .A2(n1194), .ZN(n1585) );
  ND2D1BWP12T U1697 ( .A1(n1195), .A2(n1585), .ZN(irdecode_inst1_N1013) );
  OAI32D1BWP12T U1698 ( .A1(n1302), .A2(n1504), .A3(n1196), .B1(n1479), .B2(
        n1302), .ZN(n1233) );
  ND2D1BWP12T U1699 ( .A1(n1211), .A2(n1197), .ZN(n1198) );
  OAI21D1BWP12T U1700 ( .A1(n1511), .A2(n1198), .B(n1493), .ZN(n1234) );
  ND4D1BWP12T U1701 ( .A1(n1233), .A2(n1235), .A3(n1234), .A4(n1514), .ZN(
        n1203) );
  OAI32D0BWP12T U1702 ( .A1(n1521), .A2(n1232), .A3(n1203), .B1(n1476), .B2(
        n1521), .ZN(n1584) );
  CKND2D0BWP12T U1703 ( .A1(irdecode_inst1_step[5]), .A2(n1627), .ZN(n1199) );
  OAI211D1BWP12T U1704 ( .A1(n1593), .A2(n1200), .B(n1584), .C(n1199), .ZN(
        irdecode_inst1_N986) );
  AOI22D1BWP12T U1705 ( .A1(n1627), .A2(DEC_RF_offset_b[18]), .B1(n1230), .B2(
        n1545), .ZN(n1201) );
  ND2D1BWP12T U1706 ( .A1(n1201), .A2(n1585), .ZN(irdecode_inst1_N1009) );
  AOI22D1BWP12T U1707 ( .A1(n1627), .A2(DEC_RF_offset_b[16]), .B1(n1230), .B2(
        n1338), .ZN(n1202) );
  ND2D1BWP12T U1708 ( .A1(n1202), .A2(n1585), .ZN(irdecode_inst1_N1007) );
  AOI21D0BWP12T U1709 ( .A1(n1476), .A2(n1203), .B(n1521), .ZN(n1583) );
  AOI22D1BWP12T U1710 ( .A1(n1627), .A2(irdecode_inst1_step[3]), .B1(n1204), 
        .B2(n1531), .ZN(n1205) );
  OAI211D1BWP12T U1711 ( .A1(n1593), .A2(n1206), .B(n1583), .C(n1205), .ZN(
        irdecode_inst1_N984) );
  AOI21D1BWP12T U1712 ( .A1(n1312), .A2(n1452), .B(n1207), .ZN(n1588) );
  NR2D1BWP12T U1713 ( .A1(n1540), .A2(n1491), .ZN(n1498) );
  ND2D1BWP12T U1714 ( .A1(n1312), .A2(n1592), .ZN(n1287) );
  AOI22D1BWP12T U1715 ( .A1(n1627), .A2(DEC_RF_offset_b[20]), .B1(n1230), .B2(
        n1592), .ZN(n1208) );
  ND2D1BWP12T U1716 ( .A1(n1208), .A2(n1585), .ZN(irdecode_inst1_N1011) );
  ND2D1BWP12T U1717 ( .A1(n1627), .A2(DEC_RF_offset_b[13]), .ZN(n1209) );
  OAI211D1BWP12T U1718 ( .A1(n1491), .A2(n1254), .B(n1209), .C(n1585), .ZN(
        irdecode_inst1_N1004) );
  NR2D1BWP12T U1719 ( .A1(n1282), .A2(n1464), .ZN(n1214) );
  AOI211D1BWP12T U1720 ( .A1(n1274), .A2(irdecode_inst1_N754), .B(n1298), .C(
        n1210), .ZN(n1212) );
  AOI32D1BWP12T U1721 ( .A1(n1462), .A2(n1212), .A3(n1211), .B1(n1626), .B2(
        n1212), .ZN(n1227) );
  AOI22D0BWP12T U1722 ( .A1(n1627), .A2(irdecode_inst1_step[0]), .B1(n1476), 
        .B2(n1227), .ZN(n1213) );
  OAI211D1BWP12T U1723 ( .A1(n1214), .A2(n1508), .B(n1344), .C(n1213), .ZN(
        irdecode_inst1_N981) );
  OAI22D1BWP12T U1724 ( .A1(n1321), .A2(n1277), .B1(n1358), .B2(n1217), .ZN(
        n1301) );
  AO211D1BWP12T U1725 ( .A1(n1219), .A2(n963), .B(n1218), .C(n1301), .Z(n1220)
         );
  AOI211D1BWP12T U1726 ( .A1(n1338), .A2(n1307), .B(n1221), .C(n1220), .ZN(
        n1224) );
  NR2D1BWP12T U1727 ( .A1(n1493), .A2(n1339), .ZN(n1303) );
  INVD1BWP12T U1728 ( .I(n1267), .ZN(n1625) );
  MAOI22D0BWP12T U1729 ( .A1(n1627), .A2(DEC_RF_operand_a[1]), .B1(n1303), 
        .B2(n1625), .ZN(n1223) );
  ND2D1BWP12T U1730 ( .A1(n1498), .A2(n1305), .ZN(n1222) );
  OAI211D1BWP12T U1731 ( .A1(n1224), .A2(n1540), .B(n1223), .C(n1222), .ZN(
        irdecode_inst1_N971) );
  AOI22D1BWP12T U1732 ( .A1(n1489), .A2(n1230), .B1(n1627), .B2(
        DEC_RF_offset_b[21]), .ZN(n1225) );
  ND2D1BWP12T U1733 ( .A1(n1225), .A2(n1585), .ZN(irdecode_inst1_N1012) );
  NR3D1BWP12T U1734 ( .A1(n1227), .A2(n1226), .A3(n1299), .ZN(n1228) );
  AOI21D1BWP12T U1735 ( .A1(n1233), .A2(n1228), .B(n1593), .ZN(n1229) );
  AO211D1BWP12T U1736 ( .A1(n1627), .A2(irdecode_inst1_step[1]), .B(n1521), 
        .C(n1229), .Z(irdecode_inst1_N982) );
  AOI22D1BWP12T U1737 ( .A1(DEC_RF_offset_b[19]), .A2(n1627), .B1(n1230), .B2(
        n1348), .ZN(n1231) );
  ND2D1BWP12T U1738 ( .A1(n1231), .A2(n1585), .ZN(irdecode_inst1_N1010) );
  INR3D0BWP12T U1739 ( .A1(n1233), .B1(n1232), .B2(n1270), .ZN(n1243) );
  AOI31D1BWP12T U1740 ( .A1(n1243), .A2(n1235), .A3(n1234), .B(n1593), .ZN(
        n1236) );
  AO211D1BWP12T U1741 ( .A1(n1627), .A2(irdecode_inst1_step[6]), .B(n1236), 
        .C(n1521), .Z(irdecode_inst1_N987) );
  NR2D1BWP12T U1742 ( .A1(n963), .A2(n1237), .ZN(n1316) );
  ND2D1BWP12T U1743 ( .A1(irdecode_inst1_N751), .A2(n1316), .ZN(n1285) );
  INVD1BWP12T U1744 ( .I(n1285), .ZN(n1238) );
  OAI21D1BWP12T U1745 ( .A1(n1239), .A2(n1238), .B(n1364), .ZN(n1252) );
  ND2D1BWP12T U1746 ( .A1(n1255), .A2(n1256), .ZN(n1240) );
  AOI22D1BWP12T U1747 ( .A1(n1330), .A2(n1240), .B1(n1627), .B2(
        DEC_RF_offset_b[9]), .ZN(n1241) );
  OAI211D1BWP12T U1748 ( .A1(n1452), .A2(n1252), .B(n1241), .C(n1585), .ZN(
        irdecode_inst1_N1000) );
  AOI31D1BWP12T U1749 ( .A1(n1243), .A2(n1242), .A3(n1626), .B(n1593), .ZN(
        n1244) );
  AOI211D1BWP12T U1750 ( .A1(n1627), .A2(irdecode_inst1_step[7]), .B(n1521), 
        .C(n1244), .ZN(n1245) );
  OAI21D1BWP12T U1751 ( .A1(n1508), .A2(n1246), .B(n1245), .ZN(
        irdecode_inst1_N988) );
  ND2D1BWP12T U1752 ( .A1(n1627), .A2(DEC_RF_offset_b[17]), .ZN(n1247) );
  OAI211D1BWP12T U1753 ( .A1(n1442), .A2(n1254), .B(n1247), .C(n1585), .ZN(
        irdecode_inst1_N1008) );
  ND2D1BWP12T U1754 ( .A1(n1627), .A2(DEC_RF_offset_b[10]), .ZN(n1248) );
  OAI211D1BWP12T U1755 ( .A1(n1321), .A2(n1252), .B(n1585), .C(n1248), .ZN(
        irdecode_inst1_N1001) );
  ND2D1BWP12T U1756 ( .A1(n1627), .A2(DEC_RF_offset_b[15]), .ZN(n1249) );
  OAI211D1BWP12T U1757 ( .A1(n1329), .A2(n1254), .B(n1249), .C(n1585), .ZN(
        irdecode_inst1_N1006) );
  ND2D1BWP12T U1758 ( .A1(n1627), .A2(DEC_RF_offset_b[14]), .ZN(n1250) );
  OAI211D1BWP12T U1759 ( .A1(n1328), .A2(n1254), .B(n1250), .C(n1585), .ZN(
        irdecode_inst1_N1005) );
  ND2D1BWP12T U1760 ( .A1(n1627), .A2(DEC_RF_offset_b[11]), .ZN(n1251) );
  OAI211D1BWP12T U1761 ( .A1(n1449), .A2(n1252), .B(n1585), .C(n1251), .ZN(
        irdecode_inst1_N1002) );
  ND2D1BWP12T U1762 ( .A1(n1627), .A2(DEC_RF_offset_b[12]), .ZN(n1253) );
  OAI211D1BWP12T U1763 ( .A1(n1624), .A2(n1254), .B(n1253), .C(n1585), .ZN(
        irdecode_inst1_N1003) );
  ND2D1BWP12T U1764 ( .A1(n1285), .A2(n1300), .ZN(n1336) );
  INVD1BWP12T U1765 ( .I(n1336), .ZN(n1586) );
  ND3D1BWP12T U1766 ( .A1(n1349), .A2(n1256), .A3(n1255), .ZN(n1335) );
  INVD1BWP12T U1767 ( .I(n1335), .ZN(n1315) );
  INVD1BWP12T U1768 ( .I(n1338), .ZN(n1257) );
  OAI222D1BWP12T U1769 ( .A1(n1449), .A2(n1334), .B1(n1442), .B2(n1586), .C1(
        n1315), .C2(n1257), .ZN(n1258) );
  NR2D1BWP12T U1770 ( .A1(n1540), .A2(n1447), .ZN(n1546) );
  AO222D1BWP12T U1771 ( .A1(n1258), .A2(n1364), .B1(n1339), .B2(n1546), .C1(
        n1627), .C2(DEC_RF_offset_b[6]), .Z(irdecode_inst1_N997) );
  OAI31D0BWP12T U1772 ( .A1(n1302), .A2(n1316), .A3(n1259), .B(n1476), .ZN(
        n1260) );
  OAI21D1BWP12T U1773 ( .A1(n1261), .A2(n1482), .B(n1260), .ZN(
        irdecode_inst1_N980) );
  ND2D1BWP12T U1774 ( .A1(n1335), .A2(n1308), .ZN(n1262) );
  MAOI22D0BWP12T U1775 ( .A1(n1627), .A2(DEC_RF_offset_b[7]), .B1(n1540), .B2(
        n1262), .ZN(n1264) );
  ND2D1BWP12T U1776 ( .A1(n1546), .A2(n1336), .ZN(n1263) );
  OAI211D1BWP12T U1777 ( .A1(n1358), .A2(n1544), .B(n1264), .C(n1263), .ZN(
        irdecode_inst1_N998) );
  AO222D1BWP12T U1778 ( .A1(n1330), .A2(n1336), .B1(n1546), .B2(n1335), .C1(
        n1627), .C2(DEC_RF_offset_b[8]), .Z(irdecode_inst1_N999) );
  AOI22D1BWP12T U1779 ( .A1(n1336), .A2(n1338), .B1(n1335), .B2(n1438), .ZN(
        n1266) );
  INVD1BWP12T U1780 ( .I(n1340), .ZN(n1360) );
  ND2D1BWP12T U1781 ( .A1(n1475), .A2(n1360), .ZN(n1265) );
  OAI211D1BWP12T U1782 ( .A1(n1442), .A2(n1358), .B(n1266), .C(n1265), .ZN(
        n1268) );
  INVD0BWP12T U1783 ( .I(n1334), .ZN(n1471) );
  AO222D1BWP12T U1784 ( .A1(n1268), .A2(n1364), .B1(n1627), .B2(
        DEC_RF_offset_b[5]), .C1(n1267), .C2(n1471), .Z(irdecode_inst1_N996)
         );
  NR2D1BWP12T U1785 ( .A1(n1270), .A2(n1269), .ZN(n1280) );
  NR2D1BWP12T U1786 ( .A1(n1298), .A2(n1272), .ZN(n1276) );
  AOI211D1BWP12T U1787 ( .A1(n1274), .A2(irdecode_inst1_N751), .B(n1291), .C(
        n1273), .ZN(n1275) );
  OAI211D1BWP12T U1788 ( .A1(n1278), .A2(n1277), .B(n1276), .C(n1275), .ZN(
        n1351) );
  OAI32D1BWP12T U1789 ( .A1(n1496), .A2(n1282), .A3(n1281), .B1(n1280), .B2(
        n1496), .ZN(n1283) );
  AOI211D1BWP12T U1790 ( .A1(irdecode_inst1_split_instruction), .A2(n1627), 
        .B(n1284), .C(n1283), .ZN(n1286) );
  AOI32D1BWP12T U1791 ( .A1(n1361), .A2(n1286), .A3(n1285), .B1(n1540), .B2(
        n1286), .ZN(irdecode_inst1_N990) );
  ND2D1BWP12T U1792 ( .A1(n1541), .A2(n1287), .ZN(n1289) );
  AOI21D0BWP12T U1793 ( .A1(n1476), .A2(n1289), .B(n1288), .ZN(n1596) );
  INVD1BWP12T U1794 ( .I(n1290), .ZN(n1311) );
  NR4D0BWP12T U1795 ( .A1(n1479), .A2(n1590), .A3(n1311), .A4(n1291), .ZN(
        n1367) );
  INVD1BWP12T U1796 ( .I(n1292), .ZN(n1591) );
  ND2D1BWP12T U1797 ( .A1(n1475), .A2(n1591), .ZN(n1293) );
  OAI211D1BWP12T U1798 ( .A1(n1328), .A2(n1588), .B(n1367), .C(n1293), .ZN(
        n1294) );
  AOI22D0BWP12T U1799 ( .A1(n1476), .A2(n1294), .B1(n1627), .B2(
        DEC_RF_alu_write_to_reg[2]), .ZN(n1295) );
  ND2D1BWP12T U1800 ( .A1(n1596), .A2(n1295), .ZN(irdecode_inst1_N977) );
  NR2D1BWP12T U1801 ( .A1(n1302), .A2(n1301), .ZN(n1318) );
  NR2D1BWP12T U1802 ( .A1(n1303), .A2(n1449), .ZN(n1304) );
  AO211D1BWP12T U1803 ( .A1(n1305), .A2(n1454), .B(n1304), .C(n1311), .Z(n1306) );
  AOI21D1BWP12T U1804 ( .A1(n1308), .A2(n1307), .B(n1306), .ZN(n1310) );
  CKND2D0BWP12T U1805 ( .A1(n1627), .A2(DEC_RF_operand_a[2]), .ZN(n1309) );
  OAI211D1BWP12T U1806 ( .A1(n1310), .A2(n1593), .B(n1314), .C(n1309), .ZN(
        irdecode_inst1_N972) );
  AOI22D0BWP12T U1807 ( .A1(n1476), .A2(n1311), .B1(n1627), .B2(
        DEC_RF_operand_a[3]), .ZN(n1313) );
  ND3D0BWP12T U1808 ( .A1(n1476), .A2(n1312), .A3(n1348), .ZN(n1368) );
  ND3D1BWP12T U1809 ( .A1(n1314), .A2(n1313), .A3(n1368), .ZN(
        irdecode_inst1_N973) );
  CKND2D1BWP12T U1810 ( .A1(n1504), .A2(n1531), .ZN(n1467) );
  ND2D1BWP12T U1811 ( .A1(n1316), .A2(irdecode_inst1_N754), .ZN(n1355) );
  AOI31D1BWP12T U1812 ( .A1(n1318), .A2(n1317), .A3(n1355), .B(n1593), .ZN(
        n1319) );
  NR2D1BWP12T U1813 ( .A1(n1521), .A2(n1319), .ZN(n1599) );
  OA222D1BWP12T U1814 ( .A1(n1358), .A2(n1329), .B1(n1452), .B2(n1340), .C1(
        n1586), .C2(n1328), .Z(n1333) );
  AOI22D1BWP12T U1815 ( .A1(n1330), .A2(n1471), .B1(n1627), .B2(
        DEC_RF_offset_b[3]), .ZN(n1332) );
  OAI211D1BWP12T U1816 ( .A1(n1333), .A2(n1540), .B(n1332), .C(n1331), .ZN(
        irdecode_inst1_N994) );
  CKND0BWP12T U1817 ( .I(DEC_ALU_alu_opcode[2]), .ZN(n1345) );
  OAI21D1BWP12T U1818 ( .A1(n1452), .A2(n1554), .B(n1367), .ZN(n1341) );
  OAI31D0BWP12T U1819 ( .A1(n1342), .A2(n1347), .A3(n1341), .B(n1476), .ZN(
        n1343) );
  OAI211D1BWP12T U1820 ( .A1(n1482), .A2(n1345), .B(n1344), .C(n1343), .ZN(
        irdecode_inst1_N966) );
  CKND0BWP12T U1821 ( .I(DEC_ALU_alu_opcode[0]), .ZN(n1555) );
  AOI211D1BWP12T U1822 ( .A1(n1347), .A2(n1489), .B(n963), .C(n1346), .ZN(
        n1352) );
  OAI22D1BWP12T U1823 ( .A1(n1447), .A2(n1554), .B1(n1349), .B2(n1348), .ZN(
        n1350) );
  OAI31D1BWP12T U1824 ( .A1(n1352), .A2(n1351), .A3(n1350), .B(n1364), .ZN(
        n1353) );
  OAI211D1BWP12T U1825 ( .A1(n1482), .A2(n1555), .B(n1354), .C(n1353), .ZN(
        irdecode_inst1_N964) );
  OAI21D1BWP12T U1826 ( .A1(n1624), .A2(n1358), .B(n1355), .ZN(n1357) );
  INVD1BWP12T U1827 ( .I(n1366), .ZN(n1356) );
  AO222D1BWP12T U1828 ( .A1(n1357), .A2(n1364), .B1(n1356), .B2(n1546), .C1(
        DEC_RF_offset_b[0]), .C2(n1627), .Z(irdecode_inst1_N991) );
  OAI22D1BWP12T U1829 ( .A1(n1624), .A2(n1586), .B1(n1491), .B2(n1358), .ZN(
        n1359) );
  AOI211D1BWP12T U1830 ( .A1(n1360), .A2(n1545), .B(n1493), .C(n1359), .ZN(
        n1362) );
  ND2D1BWP12T U1831 ( .A1(n1362), .A2(n1361), .ZN(n1363) );
  AOI22D1BWP12T U1832 ( .A1(n1364), .A2(n1363), .B1(n1627), .B2(
        DEC_RF_offset_b[1]), .ZN(n1365) );
  OAI211D1BWP12T U1833 ( .A1(n1366), .A2(n1544), .B(n1365), .C(n1496), .ZN(
        irdecode_inst1_N992) );
  MAOI22D0BWP12T U1834 ( .A1(n1627), .A2(DEC_RF_alu_write_to_reg[3]), .B1(
        n1367), .B2(n1593), .ZN(n1369) );
  ND3D1BWP12T U1835 ( .A1(n1596), .A2(n1369), .A3(n1368), .ZN(
        irdecode_inst1_N978) );
  CKND0BWP12T U1836 ( .I(n1433), .ZN(n1376) );
  CKND2D0BWP12T U1837 ( .A1(n1376), .A2(n1370), .ZN(n1602) );
  CKND0BWP12T U1838 ( .I(n1374), .ZN(n1372) );
  NR2D0BWP12T U1839 ( .A1(n919), .A2(n1371), .ZN(n1603) );
  ND2D1BWP12T U1840 ( .A1(n1372), .A2(n1603), .ZN(n1377) );
  ND2D1BWP12T U1841 ( .A1(n1602), .A2(n1377), .ZN(n1398) );
  ND2D1BWP12T U1842 ( .A1(n1373), .A2(n1398), .ZN(n1412) );
  NR2D1BWP12T U1843 ( .A1(n1602), .A2(n1377), .ZN(n1413) );
  CKND0BWP12T U1844 ( .I(n1414), .ZN(n1426) );
  NR2D0BWP12T U1845 ( .A1(n1426), .A2(n1374), .ZN(n1375) );
  ND2D1BWP12T U1846 ( .A1(n1376), .A2(n1375), .ZN(n1605) );
  INVD1BWP12T U1847 ( .I(n1428), .ZN(n1378) );
  INR2D1BWP12T U1848 ( .A1(n1378), .B1(n1377), .ZN(n1407) );
  NR2D1BWP12T U1849 ( .A1(n1605), .A2(n1407), .ZN(n1396) );
  INVD1BWP12T U1850 ( .I(n1396), .ZN(n1416) );
  INVD1BWP12T U1851 ( .I(n1605), .ZN(n1393) );
  INVD1BWP12T U1852 ( .I(n1407), .ZN(n1409) );
  OAI21D1BWP12T U1853 ( .A1(memory_interface_inst1_delay_addr_for_adder[0]), 
        .A2(n1605), .B(n1409), .ZN(n1400) );
  ND3D1BWP12T U1854 ( .A1(memory_interface_inst1_delay_addr_for_adder[0]), 
        .A2(memory_interface_inst1_delay_addr_for_adder[1]), .A3(
        memory_interface_inst1_delay_addr_for_adder[2]), .ZN(n1380) );
  INVD1BWP12T U1855 ( .I(n1380), .ZN(n1381) );
  OAI21D1BWP12T U1856 ( .A1(n1381), .A2(n1605), .B(n1409), .ZN(n1382) );
  AOI22D1BWP12T U1857 ( .A1(memory_interface_inst1_delay_addr_for_adder[3]), 
        .A2(n1382), .B1(n1605), .B2(MEMCTRL_IN_address[3]), .ZN(n1379) );
  OAI31D1BWP12T U1858 ( .A1(memory_interface_inst1_delay_addr_for_adder[3]), 
        .A2(n1416), .A3(n1380), .B(n1379), .ZN(MEMCTRL_MEM_to_mem_address[3])
         );
  ND2D1BWP12T U1859 ( .A1(n1381), .A2(
        memory_interface_inst1_delay_addr_for_adder[3]), .ZN(n1383) );
  INR2D1BWP12T U1860 ( .A1(memory_interface_inst1_delay_addr_for_adder[4]), 
        .B1(n1383), .ZN(n1386) );
  INVD1BWP12T U1861 ( .I(n1386), .ZN(n1385) );
  OAI21D1BWP12T U1862 ( .A1(n1386), .A2(n1605), .B(n1409), .ZN(n1387) );
  AOI22D1BWP12T U1863 ( .A1(memory_interface_inst1_delay_addr_for_adder[5]), 
        .A2(n1387), .B1(n1605), .B2(MEMCTRL_IN_address[5]), .ZN(n1384) );
  OAI31D1BWP12T U1864 ( .A1(memory_interface_inst1_delay_addr_for_adder[5]), 
        .A2(n1416), .A3(n1385), .B(n1384), .ZN(MEMCTRL_MEM_to_mem_address[5])
         );
  ND2D1BWP12T U1865 ( .A1(n1386), .A2(
        memory_interface_inst1_delay_addr_for_adder[5]), .ZN(n1388) );
  INR2D1BWP12T U1866 ( .A1(memory_interface_inst1_delay_addr_for_adder[6]), 
        .B1(n1388), .ZN(n1391) );
  INVD1BWP12T U1867 ( .I(n1391), .ZN(n1390) );
  OAI21D1BWP12T U1868 ( .A1(n1391), .A2(n1605), .B(n1409), .ZN(n1392) );
  AOI22D1BWP12T U1869 ( .A1(memory_interface_inst1_delay_addr_for_adder[7]), 
        .A2(n1392), .B1(n1605), .B2(MEMCTRL_IN_address[7]), .ZN(n1389) );
  OAI31D1BWP12T U1870 ( .A1(memory_interface_inst1_delay_addr_for_adder[7]), 
        .A2(n1416), .A3(n1390), .B(n1389), .ZN(MEMCTRL_MEM_to_mem_address[7])
         );
  ND2D1BWP12T U1871 ( .A1(n1391), .A2(
        memory_interface_inst1_delay_addr_for_adder[7]), .ZN(n1394) );
  INR2D1BWP12T U1872 ( .A1(memory_interface_inst1_delay_addr_for_adder[8]), 
        .B1(n1394), .ZN(n1395) );
  AN2XD0BWP12T U1873 ( .A1(n1395), .A2(n1396), .Z(n1607) );
  ND2D1BWP12T U1874 ( .A1(memory_interface_inst1_delay_addr_for_adder[9]), 
        .A2(n1607), .ZN(n1419) );
  INVD1BWP12T U1875 ( .I(memory_interface_inst1_delay_addr_for_adder[10]), 
        .ZN(n1420) );
  INVD1BWP12T U1876 ( .I(memory_interface_inst1_delay_addr_for_adder[9]), .ZN(
        n1606) );
  OAI21D1BWP12T U1877 ( .A1(n1395), .A2(n1605), .B(n1409), .ZN(n1608) );
  AOI21D1BWP12T U1878 ( .A1(n1396), .A2(n1606), .B(n1608), .ZN(n1415) );
  ND2D1BWP12T U1879 ( .A1(n1605), .A2(MEMCTRL_IN_address[10]), .ZN(n1397) );
  OAI221D1BWP12T U1880 ( .A1(memory_interface_inst1_delay_addr_for_adder[10]), 
        .A2(n1419), .B1(n1420), .B2(n1415), .C(n1397), .ZN(
        MEMCTRL_MEM_to_mem_address[10]) );
  INVD1BWP12T U1881 ( .I(MEM_MEMCTRL_from_mem_data[2]), .ZN(n1582) );
  INVD1BWP12T U1882 ( .I(n1398), .ZN(n1410) );
  NR2D1BWP12T U1883 ( .A1(memory_interface_inst1_delay_addr_for_adder[1]), 
        .A2(n1416), .ZN(n1399) );
  AO222D1BWP12T U1884 ( .A1(n1400), .A2(
        memory_interface_inst1_delay_addr_for_adder[1]), .B1(n1605), .B2(
        MEMCTRL_IN_address[1]), .C1(
        memory_interface_inst1_delay_addr_for_adder[0]), .C2(n1399), .Z(
        MEMCTRL_MEM_to_mem_address[1]) );
  INVD1BWP12T U1885 ( .I(RF_MEMCTRL_data_reg[8]), .ZN(n1403) );
  INVD1BWP12T U1886 ( .I(MEM_MEMCTRL_from_mem_data[0]), .ZN(n1570) );
  ND2D1BWP12T U1887 ( .A1(n1410), .A2(
        memory_interface_inst1_delay_data_in32[8]), .ZN(n1401) );
  OAI211D1BWP12T U1888 ( .A1(n1403), .A2(n1414), .B(n1402), .C(n1401), .ZN(
        MEMCTRL_MEM_to_mem_data[0]) );
  INVD1BWP12T U1889 ( .I(RF_MEMCTRL_data_reg[9]), .ZN(n1406) );
  INVD1BWP12T U1890 ( .I(MEM_MEMCTRL_from_mem_data[1]), .ZN(n1572) );
  ND2D1BWP12T U1891 ( .A1(n1410), .A2(
        memory_interface_inst1_delay_data_in32[9]), .ZN(n1404) );
  OAI211D1BWP12T U1892 ( .A1(n1406), .A2(n1414), .B(n1405), .C(n1404), .ZN(
        MEMCTRL_MEM_to_mem_data[1]) );
  AOI22D1BWP12T U1893 ( .A1(n1407), .A2(
        memory_interface_inst1_delay_addr_for_adder[0]), .B1(
        MEMCTRL_IN_address[0]), .B2(n1605), .ZN(n1408) );
  OAI21D1BWP12T U1894 ( .A1(memory_interface_inst1_delay_addr_for_adder[0]), 
        .A2(n1416), .B(n1408), .ZN(MEMCTRL_MEM_to_mem_address[0]) );
  INVD1BWP12T U1895 ( .I(MEM_MEMCTRL_from_mem_data[3]), .ZN(n1569) );
  INVD1BWP12T U1896 ( .I(MEM_MEMCTRL_from_mem_data[4]), .ZN(n1568) );
  INVD1BWP12T U1897 ( .I(MEM_MEMCTRL_from_mem_data[5]), .ZN(n1567) );
  INVD1BWP12T U1898 ( .I(MEM_MEMCTRL_from_mem_data[6]), .ZN(n1565) );
  INVD1BWP12T U1899 ( .I(MEM_MEMCTRL_from_mem_data[7]), .ZN(n1566) );
  OAI31D1BWP12T U1900 ( .A1(n1601), .A2(n1421), .A3(n1602), .B(n1411), .ZN(
        MEMCTRL_MEM_to_mem_write_enable) );
  OAI21D1BWP12T U1901 ( .A1(memory_interface_inst1_delay_addr_for_adder[10]), 
        .A2(n1416), .B(n1415), .ZN(n1417) );
  AOI22D1BWP12T U1902 ( .A1(memory_interface_inst1_delay_addr_for_adder[11]), 
        .A2(n1417), .B1(n1605), .B2(MEMCTRL_IN_address[11]), .ZN(n1418) );
  OAI31D1BWP12T U1903 ( .A1(memory_interface_inst1_delay_addr_for_adder[11]), 
        .A2(n1420), .A3(n1419), .B(n1418), .ZN(MEMCTRL_MEM_to_mem_address[11])
         );
  OAI21D0BWP12T U1904 ( .A1(DEC_MEMCTRL_load_store_width[1]), .A2(n1421), .B(
        n1422), .ZN(n1425) );
  CKND0BWP12T U1905 ( .I(n1422), .ZN(n1600) );
  ND2D0BWP12T U1906 ( .A1(n1600), .A2(DEC_MEMCTRL_load_store_width[0]), .ZN(
        n1424) );
  TPAOI31D0BWP12T U1907 ( .A1(n1426), .A2(n1425), .A3(n1424), .B(n1423), .ZN(
        n1427) );
  NR2D1BWP12T U1908 ( .A1(n1427), .A2(reset), .ZN(
        memory_interface_inst1_fsm_N33) );
  AOI21D0BWP12T U1909 ( .A1(n1430), .A2(n1429), .B(n1428), .ZN(n1431) );
  OAI22D1BWP12T U1910 ( .A1(n1432), .A2(n1601), .B1(reset), .B2(n1431), .ZN(
        memory_interface_inst1_fsm_N34) );
  AOI21D0BWP12T U1911 ( .A1(n1434), .A2(n1433), .B(
        Instruction_Fetch_inst1_first_instruction_fetched), .ZN(n1435) );
  NR2D1BWP12T U1912 ( .A1(reset), .A2(n1435), .ZN(n815) );
  CKND0BWP12T U1913 ( .I(n1491), .ZN(n1436) );
  INVD1BWP12T U1914 ( .I(n1623), .ZN(n1437) );
  AO222D1BWP12T U1915 ( .A1(n1436), .A2(n1437), .B1(n1622), .B2(
        irdecode_inst1_itstate_1_), .C1(n1440), .C2(irdecode_inst1_itstate_0_), 
        .Z(n812) );
  AO222D1BWP12T U1916 ( .A1(n1454), .A2(n1437), .B1(n1622), .B2(
        irdecode_inst1_itstate_2_), .C1(n1440), .C2(irdecode_inst1_itstate_1_), 
        .Z(n811) );
  AO222D1BWP12T U1917 ( .A1(n1438), .A2(n1437), .B1(n1622), .B2(
        irdecode_inst1_itstate_3_), .C1(n1440), .C2(irdecode_inst1_itstate_2_), 
        .Z(n810) );
  INVD1BWP12T U1918 ( .I(n1439), .ZN(n1446) );
  NR2D1BWP12T U1919 ( .A1(n1440), .A2(n1622), .ZN(n1445) );
  OAI22D1BWP12T U1920 ( .A1(n1446), .A2(n1442), .B1(n1445), .B2(n1441), .ZN(
        n808) );
  OAI22D1BWP12T U1921 ( .A1(n1543), .A2(n1446), .B1(n1445), .B2(n1443), .ZN(
        n806) );
  OAI22D1BWP12T U1922 ( .A1(n1447), .A2(n1446), .B1(n1445), .B2(n1444), .ZN(
        n807) );
  AOI21D0BWP12T U1923 ( .A1(n1627), .A2(DEC_RF_memory_store_address_reg[2]), 
        .B(n1450), .ZN(n1448) );
  OAI21D1BWP12T U1924 ( .A1(n1449), .A2(n1593), .B(n1448), .ZN(n791) );
  AOI21D0BWP12T U1925 ( .A1(n1627), .A2(DEC_RF_memory_store_address_reg[0]), 
        .B(n1450), .ZN(n1451) );
  OAI21D1BWP12T U1926 ( .A1(n1452), .A2(n1593), .B(n1451), .ZN(n789) );
  OR2XD0BWP12T U1927 ( .A1(n1517), .A2(n1516), .Z(n1455) );
  AOI22D0BWP12T U1928 ( .A1(n1455), .A2(n1454), .B1(n1518), .B2(n1453), .ZN(
        n1457) );
  TPAOI31D0BWP12T U1929 ( .A1(n1457), .A2(n1520), .A3(n1456), .B(n1593), .ZN(
        n1459) );
  AO211D1BWP12T U1930 ( .A1(n1627), .A2(DEC_RF_memory_store_data_reg[2]), .B(
        n1459), .C(n1458), .Z(n796) );
  CKND0BWP12T U1931 ( .I(DEC_RF_memory_write_to_reg[3]), .ZN(n1466) );
  CKND2D1BWP12T U1932 ( .A1(n1461), .A2(n1460), .ZN(n1529) );
  AOI21D0BWP12T U1933 ( .A1(n1462), .A2(n1500), .B(n1626), .ZN(n1463) );
  OAI32D0BWP12T U1934 ( .A1(n1521), .A2(n1529), .A3(n1463), .B1(n1476), .B2(
        n1521), .ZN(n1506) );
  TPOAI21D0BWP12T U1935 ( .A1(n963), .A2(n1464), .B(n1531), .ZN(n1465) );
  OAI211D1BWP12T U1936 ( .A1(n1482), .A2(n1466), .B(n1506), .C(n1465), .ZN(
        n803) );
  CKND0BWP12T U1937 ( .I(DEC_RF_memory_store_data_reg[4]), .ZN(n1469) );
  OAI211D1BWP12T U1938 ( .A1(n1482), .A2(n1469), .B(n1468), .C(n1467), .ZN(
        n798) );
  INVD1BWP12T U1939 ( .I(DEC_MEMCTRL_load_store_width[1]), .ZN(n1481) );
  AOI211D0BWP12T U1940 ( .A1(n1472), .A2(n1471), .B(n1518), .C(n1470), .ZN(
        n1473) );
  OAI31D0BWP12T U1941 ( .A1(n1475), .A2(n1489), .A3(n1474), .B(n1473), .ZN(
        n1477) );
  OAI31D0BWP12T U1942 ( .A1(n1479), .A2(n1478), .A3(n1477), .B(n1476), .ZN(
        n1480) );
  OAI211D1BWP12T U1943 ( .A1(n1482), .A2(n1481), .B(n1480), .C(n1533), .ZN(
        n787) );
  NR4D0BWP12T U1944 ( .A1(n1486), .A2(n1485), .A3(n1484), .A4(n1483), .ZN(
        n1488) );
  CKND2D1BWP12T U1945 ( .A1(n1488), .A2(n1487), .ZN(n1494) );
  MOAI22D0BWP12T U1946 ( .A1(n1491), .A2(n1490), .B1(n1518), .B2(n1489), .ZN(
        n1492) );
  AOI21D1BWP12T U1947 ( .A1(n1494), .A2(n1493), .B(n1492), .ZN(n1495) );
  OAI22D1BWP12T U1948 ( .A1(n1497), .A2(n1496), .B1(n1495), .B2(n1540), .ZN(
        n1499) );
  AO222D1BWP12T U1949 ( .A1(n1499), .A2(n963), .B1(n1517), .B2(n1498), .C1(
        n1627), .C2(DEC_RF_memory_store_data_reg[1]), .Z(n795) );
  AOI22D0BWP12T U1950 ( .A1(n1627), .A2(DEC_RF_memory_write_to_reg[1]), .B1(
        n1524), .B2(n1498), .ZN(n1502) );
  CKND2D1BWP12T U1951 ( .A1(n1500), .A2(n1499), .ZN(n1501) );
  OAI211D1BWP12T U1952 ( .A1(n1625), .A2(n1503), .B(n1502), .C(n1501), .ZN(
        n801) );
  AOI22D0BWP12T U1953 ( .A1(n1627), .A2(DEC_RF_memory_write_to_reg[4]), .B1(
        n1504), .B2(n1531), .ZN(n1505) );
  OAI211D1BWP12T U1954 ( .A1(n1508), .A2(n1507), .B(n1506), .C(n1505), .ZN(
        n804) );
  CKND0BWP12T U1955 ( .I(n1624), .ZN(n1523) );
  AOI22D0BWP12T U1956 ( .A1(n1518), .A2(n1592), .B1(n1517), .B2(n1523), .ZN(
        n1519) );
  AOI31D1BWP12T U1957 ( .A1(n1520), .A2(n1527), .A3(n1519), .B(n1593), .ZN(
        n1522) );
  AO211D1BWP12T U1958 ( .A1(n1627), .A2(DEC_RF_memory_store_data_reg[0]), .B(
        n1522), .C(n1521), .Z(n794) );
  AOI22D0BWP12T U1959 ( .A1(n963), .A2(n1525), .B1(n1524), .B2(n1523), .ZN(
        n1526) );
  CKND2D1BWP12T U1960 ( .A1(n1527), .A2(n1526), .ZN(n1528) );
  RCAOI211D0BWP12T U1961 ( .A1(n1592), .A2(n1530), .B(n1529), .C(n1528), .ZN(
        n1535) );
  AOI22D0BWP12T U1962 ( .A1(n1627), .A2(DEC_RF_memory_write_to_reg[0]), .B1(
        n1532), .B2(n1531), .ZN(n1534) );
  OAI211D1BWP12T U1963 ( .A1(n1535), .A2(n1593), .B(n1534), .C(n1533), .ZN(
        n800) );
  NR2D1BWP12T U1964 ( .A1(n1537), .A2(n1536), .ZN(n1539) );
  OAI22D1BWP12T U1965 ( .A1(n1541), .A2(n1540), .B1(n1539), .B2(n1538), .ZN(
        irdecode_inst1_next_update_flag_n) );
  AO21D1BWP12T U1966 ( .A1(DEC_MEMCTRL_memory_load_request), .A2(n1627), .B(
        n1542), .Z(n805) );
  MOAI22D0BWP12T U1967 ( .A1(n1545), .A2(n1544), .B1(n1543), .B2(n1546), .ZN(
        n1548) );
  TPAOI22D0BWP12T U1968 ( .A1(n1549), .A2(n1548), .B1(n1547), .B2(n1546), .ZN(
        n1553) );
  CKND0BWP12T U1969 ( .I(n1550), .ZN(n1552) );
  OAI31D1BWP12T U1970 ( .A1(n1554), .A2(n1553), .A3(n1552), .B(n1551), .ZN(
        irdecode_inst1_next_update_flag_v) );
  MUX2D1BWP12T U1971 ( .I0(RF_OUT_z), .I1(ALU_OUT_z), .S(
        DEC_CPSR_update_flag_z), .Z(new_z) );
  MUX2D1BWP12T U1972 ( .I0(RF_OUT_v), .I1(ALU_OUT_v), .S(
        DEC_CPSR_update_flag_v), .Z(new_v) );
  MUX2D1BWP12T U1973 ( .I0(RF_OUT_n), .I1(ALU_OUT_n), .S(
        DEC_CPSR_update_flag_n), .Z(new_n) );
  IND3D0BWP12T U1974 ( .A1(DEC_ALU_alu_opcode[3]), .B1(DEC_ALU_alu_opcode[4]), 
        .B2(DEC_ALU_alu_opcode[2]), .ZN(n1558) );
  CKND2D0BWP12T U1975 ( .A1(n1555), .A2(DEC_ALU_alu_opcode[1]), .ZN(n1557) );
  OAI22D1BWP12T U1976 ( .A1(n1558), .A2(n1557), .B1(DEC_ALU_alu_opcode[4]), 
        .B2(n1556), .ZN(ALU_IN_c) );
  AN3XD1BWP12T U1977 ( .A1(n1559), .A2(MEM_MEMCTRL_from_mem_data[7]), .A3(
        memory_interface_inst1_delayed_is_signed), .Z(n1564) );
  INR2D1BWP12T U1978 ( .A1(memory_interface_inst1_delayed_is_signed), .B1(
        n1560), .ZN(n1561) );
  NR2D1BWP12T U1979 ( .A1(n1562), .A2(n1561), .ZN(n1563) );
  OAI21D1BWP12T U1980 ( .A1(n1565), .A2(n1581), .B(n1580), .ZN(
        MEMCTRL_RF_IF_data_in[30]) );
  OAI21D1BWP12T U1981 ( .A1(n1566), .A2(n1581), .B(n1580), .ZN(
        MEMCTRL_RF_IF_data_in[31]) );
  OAI21D1BWP12T U1982 ( .A1(n1567), .A2(n1581), .B(n1580), .ZN(
        MEMCTRL_RF_IF_data_in[29]) );
  OAI21D1BWP12T U1983 ( .A1(n1568), .A2(n1581), .B(n1580), .ZN(
        MEMCTRL_RF_IF_data_in[28]) );
  OAI21D1BWP12T U1984 ( .A1(n1569), .A2(n1581), .B(n1580), .ZN(
        MEMCTRL_RF_IF_data_in[27]) );
  OAI21D1BWP12T U1985 ( .A1(n1570), .A2(n1581), .B(n1580), .ZN(
        MEMCTRL_RF_IF_data_in[24]) );
  OAI21D1BWP12T U1986 ( .A1(n1581), .A2(n1571), .B(n1580), .ZN(
        MEMCTRL_RF_IF_data_in[23]) );
  OAI21D1BWP12T U1987 ( .A1(n1572), .A2(n1581), .B(n1580), .ZN(
        MEMCTRL_RF_IF_data_in[25]) );
  OAI21D1BWP12T U1988 ( .A1(n1581), .A2(n1573), .B(n1580), .ZN(
        MEMCTRL_RF_IF_data_in[22]) );
  OAI21D1BWP12T U1989 ( .A1(n1581), .A2(n1574), .B(n1580), .ZN(
        MEMCTRL_RF_IF_data_in[21]) );
  OAI21D1BWP12T U1990 ( .A1(n1581), .A2(n1575), .B(n1580), .ZN(
        MEMCTRL_RF_IF_data_in[19]) );
  OAI21D1BWP12T U1991 ( .A1(n1581), .A2(n1576), .B(n1580), .ZN(
        MEMCTRL_RF_IF_data_in[18]) );
  OAI21D1BWP12T U1992 ( .A1(n1581), .A2(n1577), .B(n1580), .ZN(
        MEMCTRL_RF_IF_data_in[17]) );
  OAI21D1BWP12T U1993 ( .A1(n1581), .A2(n1578), .B(n1580), .ZN(
        MEMCTRL_RF_IF_data_in[16]) );
  OAI21D1BWP12T U1994 ( .A1(n1581), .A2(n1579), .B(n1580), .ZN(
        MEMCTRL_RF_IF_data_in[20]) );
  OAI21D1BWP12T U1995 ( .A1(n1582), .A2(n1581), .B(n1580), .ZN(
        MEMCTRL_RF_IF_data_in[26]) );
  IOA21D1BWP12T U1996 ( .A1(n1627), .A2(irdecode_inst1_step[2]), .B(n1583), 
        .ZN(irdecode_inst1_N983) );
  IOA21D1BWP12T U1997 ( .A1(n1627), .A2(DEC_RF_offset_b[31]), .B(n1585), .ZN(
        irdecode_inst1_N1022) );
  IOA21D1BWP12T U1998 ( .A1(n1627), .A2(DEC_RF_offset_b[29]), .B(n1585), .ZN(
        irdecode_inst1_N1020) );
  IOA21D1BWP12T U1999 ( .A1(n1627), .A2(irdecode_inst1_step[4]), .B(n1584), 
        .ZN(irdecode_inst1_N985) );
  IOA21D1BWP12T U2000 ( .A1(n1627), .A2(DEC_RF_offset_b[28]), .B(n1585), .ZN(
        irdecode_inst1_N1019) );
  IOA21D1BWP12T U2001 ( .A1(n1627), .A2(DEC_RF_offset_b[27]), .B(n1585), .ZN(
        irdecode_inst1_N1018) );
  IOA21D1BWP12T U2002 ( .A1(n1627), .A2(DEC_RF_offset_b[26]), .B(n1585), .ZN(
        irdecode_inst1_N1017) );
  IOA21D1BWP12T U2003 ( .A1(n1627), .A2(DEC_RF_offset_b[25]), .B(n1585), .ZN(
        irdecode_inst1_N1016) );
  IOA21D1BWP12T U2004 ( .A1(n1627), .A2(DEC_RF_offset_b[24]), .B(n1585), .ZN(
        irdecode_inst1_N1015) );
  IOA21D1BWP12T U2005 ( .A1(n1627), .A2(DEC_RF_offset_b[23]), .B(n1585), .ZN(
        irdecode_inst1_N1014) );
  IOA21D1BWP12T U2006 ( .A1(n1627), .A2(DEC_RF_offset_b[30]), .B(n1585), .ZN(
        irdecode_inst1_N1021) );
  OAI211D1BWP12T U2007 ( .A1(n1624), .A2(n1588), .B(n1587), .C(n1586), .ZN(
        n1589) );
  AOI211D1BWP12T U2008 ( .A1(n1592), .A2(n1591), .B(n1590), .C(n1589), .ZN(
        n1595) );
  AOI21D1BWP12T U2009 ( .A1(n1595), .A2(n1594), .B(n1593), .ZN(n1598) );
  INVD1BWP12T U2010 ( .I(n1596), .ZN(n1597) );
  AO211D0BWP12T U2011 ( .A1(n1627), .A2(DEC_RF_alu_write_to_reg[0]), .B(n1598), 
        .C(n1597), .Z(irdecode_inst1_N975) );
  IOA21D1BWP12T U2012 ( .A1(n1627), .A2(DEC_RF_operand_a[4]), .B(n1599), .ZN(
        irdecode_inst1_N974) );
  NR2D1BWP12T U2013 ( .A1(n1601), .A2(n1600), .ZN(n1604) );
  MUX2ND0BWP12T U2014 ( .I0(n1604), .I1(n1603), .S(n1602), .ZN(
        MEMCTRL_MEM_to_mem_read_enable) );
  CKND0BWP12T U2015 ( .I(MEMCTRL_RF_IF_data_in[7]), .ZN(n1611) );
  CKND2D1BWP12T U2016 ( .A1(n1610), .A2(n1609), .ZN(n1620) );
  NR2D1BWP12T U2017 ( .A1(reset), .A2(n1610), .ZN(n1619) );
  MOAI22D0BWP12T U2018 ( .A1(n1611), .A2(n1620), .B1(n1619), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_7_), .ZN(
        Instruction_Fetch_inst1_N91) );
  CKND0BWP12T U2019 ( .I(MEMCTRL_RF_IF_data_in[4]), .ZN(n1612) );
  MOAI22D0BWP12T U2020 ( .A1(n1612), .A2(n1620), .B1(n1619), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_4_), .ZN(
        Instruction_Fetch_inst1_N88) );
  CKND0BWP12T U2021 ( .I(MEMCTRL_RF_IF_data_in[6]), .ZN(n1613) );
  MOAI22D0BWP12T U2022 ( .A1(n1613), .A2(n1620), .B1(n1619), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_6_), .ZN(
        Instruction_Fetch_inst1_N90) );
  MOAI22D0BWP12T U2023 ( .A1(n1614), .A2(n1620), .B1(n1619), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_5_), .ZN(
        Instruction_Fetch_inst1_N89) );
  MOAI22D0BWP12T U2024 ( .A1(n1615), .A2(n1620), .B1(n1619), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_3_), .ZN(
        Instruction_Fetch_inst1_N87) );
  MOAI22D0BWP12T U2025 ( .A1(n1616), .A2(n1620), .B1(n1619), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_1_), .ZN(
        Instruction_Fetch_inst1_N85) );
  MOAI22D0BWP12T U2026 ( .A1(n1617), .A2(n1620), .B1(n1619), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_2_), .ZN(
        Instruction_Fetch_inst1_N86) );
  MOAI22D0BWP12T U2027 ( .A1(n1618), .A2(n1620), .B1(n1619), .B2(
        Instruction_Fetch_inst1_fetched_instruction_reg_0_), .ZN(
        Instruction_Fetch_inst1_N84) );
  MOAI22D0BWP12T U2028 ( .A1(n1621), .A2(n1620), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_14_), .B2(n1619), .ZN(
        Instruction_Fetch_inst1_N98) );
  MOAI22D0BWP12T U2029 ( .A1(n1624), .A2(n1623), .B1(irdecode_inst1_itstate_0_), .B2(n1622), .ZN(n813) );
  MOAI22D0BWP12T U2030 ( .A1(n1626), .A2(n1625), .B1(n1627), .B2(
        DEC_RF_memory_store_address_reg[1]), .ZN(n790) );
  MOAI22D0BWP12T U2031 ( .A1(n963), .A2(n1628), .B1(n1627), .B2(
        DEC_MEMCTRL_memorycontroller_sign_extend), .ZN(n785) );
endmodule

