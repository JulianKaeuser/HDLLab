module Instruction_Fetch(

input clk, reset, stall_decoder_in, stall_memory, 
input[31:0] pc_in, 
input[15:0] instruction_in, 

output reg read_enable, pc_en, valid, /*stall_decoder_out,*/  
output reg[11:0] address, 
output reg [31:0] pc_out, 
output reg[15:0] instruction_out

);


localparam[1:0]
RESET = 2'b01,
WAIT = 2'b00,
READ = 2'b10;
//D = 2'b11;

reg[1:0] currentState, nextState;


always@(currentState or stall_decoder_in or stall_memory or pc_in or instruction_in) begin
pc_out = pc_in + 1;

case(currentState)
		
	RESET: begin
		nextState = (reset == 1) ? RESET:WAIT;
		pc_out = 32'b00000000000000000000000000000100;
		read_enable = 1'b1;
		pc_en = 1'b1;
		address = 12'b0;
		instruction_out = 16'b0001110000000000;
		valid = 1'b1;
		//stall_decoder_out = 1'b0;
	end
	WAIT: begin
		nextState = (stall_memory == 1 || stall_decoder_in == 1) ? WAIT:READ;
		read_enable = (stall_decoder_in == 0) ? 1'b1: 1'b0;
		pc_en = 1'b0;
		//stall_decoder_out = 1'b0;
		address = pc_in;
		instruction_out = 16'bx;
		valid = 1'b0;
	end
	/*C: begin
		nextState = (stall_memory == 0) ? C:D;
		read_enable = (stall_memory == 1) ? 1'b0:1'b1;
		pc_en = 1'b1;
		address = pc_in - 4;
		//stall_decoder_out = 1'b1;
		instruction = instruction_out;
	end
	D: begin
		nextState = (stall_memory == 1)? D: (stall_decoder_in == 1)? B: C;
		read_enable = 1'b0;
		//stall_decoder_out = 1'b1;
		instruction= (stall_memory == 1) ? instruction_out: instruction_in ;
		pc_en = 1'b1;
		address = 12'bx;
	end*/
	READ: begin
		nextState = (stall_memory == 1 || stall_decoder_in == 1) ? WAIT : READ;
		read_enable = 1'b0;
		//stall_decoder_out = 1'b1;
		instruction_out =  instruction_in ;
		address = pc_in;
		read_enable = (stall_decoder_in == 0 && stall_memory == 0) ? 1'b1: 1'b0;
		valid = 1'b1;
		pc_en = 1'b1;
	end
	default: begin
		read_enable = 1'bx;
		instruction_out = 16'bx;
		address = 12'bx;
		pc_en = 1'bx;
		nextState = WAIT;
		pc_out = 32'bx;
		valid = 0;
		//stall_decoder_out = 1'bx;
	end
endcase
end

always@(posedge clk or posedge reset) begin
	if(reset) begin
	currentState <= RESET;
	end
	
	else begin
	currentState <= nextState;
	end 
end
endmodule
