
module register_file ( readA_sel, readB_sel, readC_sel, readD_sel, write1_sel, 
        write2_sel, write1_en, write2_en, write1_in, write2_in, immediate1_in, 
        immediate2_in, next_pc_in, next_cpsr_in, next_sp_in, clk, reset, 
        regA_out, regB_out, regC_out, regD_out, pc_out, cpsr_out, sp_out, 
        next_pc_en_BAR );
  input [4:0] readA_sel;
  input [4:0] readB_sel;
  input [4:0] readC_sel;
  input [4:0] readD_sel;
  input [4:0] write1_sel;
  input [4:0] write2_sel;
  input [31:0] write1_in;
  input [31:0] write2_in;
  input [31:0] immediate1_in;
  input [31:0] immediate2_in;
  input [31:0] next_pc_in;
  input [3:0] next_cpsr_in;
  input [31:0] next_sp_in;
  output [31:0] regA_out;
  output [31:0] regB_out;
  output [31:0] regC_out;
  output [31:0] regD_out;
  output [31:0] pc_out;
  output [3:0] cpsr_out;
  output [31:0] sp_out;
  input write1_en, write2_en, clk, reset, next_pc_en_BAR;
  wire   n2136, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2137, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935;
  wire   [2937:2968] n;
  wire   [31:0] r0;
  wire   [31:0] r1;
  wire   [31:0] r2;
  wire   [31:0] r3;
  wire   [31:0] r4;
  wire   [31:0] r5;
  wire   [31:0] r6;
  wire   [31:0] r7;
  wire   [31:0] r8;
  wire   [31:0] r9;
  wire   [31:0] r10;
  wire   [31:0] r11;
  wire   [31:0] r12;
  wire   [31:0] lr;
  wire   [31:0] tmp1;
  wire   [31:0] spin;
  wire   [3:0] cpsrin;

  DFQD1BWP12T r0_reg_31_ ( .D(n2648), .CP(clk), .Q(r0[31]) );
  DFQD1BWP12T r0_reg_30_ ( .D(n2647), .CP(clk), .Q(r0[30]) );
  DFQD1BWP12T r0_reg_29_ ( .D(n2646), .CP(clk), .Q(r0[29]) );
  DFQD1BWP12T r0_reg_28_ ( .D(n2645), .CP(clk), .Q(r0[28]) );
  DFQD1BWP12T r0_reg_27_ ( .D(n2644), .CP(clk), .Q(r0[27]) );
  DFQD1BWP12T r0_reg_26_ ( .D(n2643), .CP(clk), .Q(r0[26]) );
  DFQD1BWP12T r0_reg_25_ ( .D(n2642), .CP(clk), .Q(r0[25]) );
  DFQD1BWP12T r0_reg_24_ ( .D(n2641), .CP(clk), .Q(r0[24]) );
  DFQD1BWP12T r0_reg_23_ ( .D(n2640), .CP(clk), .Q(r0[23]) );
  DFQD1BWP12T r0_reg_22_ ( .D(n2639), .CP(clk), .Q(r0[22]) );
  DFQD1BWP12T r0_reg_21_ ( .D(n2638), .CP(clk), .Q(r0[21]) );
  DFQD1BWP12T r0_reg_20_ ( .D(n2637), .CP(clk), .Q(r0[20]) );
  DFQD1BWP12T r0_reg_19_ ( .D(n2636), .CP(clk), .Q(r0[19]) );
  DFQD1BWP12T r0_reg_18_ ( .D(n2635), .CP(clk), .Q(r0[18]) );
  DFQD1BWP12T r0_reg_17_ ( .D(n2634), .CP(clk), .Q(r0[17]) );
  DFQD1BWP12T r0_reg_16_ ( .D(n2633), .CP(clk), .Q(r0[16]) );
  DFQD1BWP12T r0_reg_15_ ( .D(n2632), .CP(clk), .Q(r0[15]) );
  DFQD1BWP12T r0_reg_14_ ( .D(n2631), .CP(clk), .Q(r0[14]) );
  DFQD1BWP12T r0_reg_13_ ( .D(n2630), .CP(clk), .Q(r0[13]) );
  DFQD1BWP12T r0_reg_12_ ( .D(n2629), .CP(clk), .Q(r0[12]) );
  DFQD1BWP12T r0_reg_11_ ( .D(n2628), .CP(clk), .Q(r0[11]) );
  DFQD1BWP12T r0_reg_10_ ( .D(n2627), .CP(clk), .Q(r0[10]) );
  DFQD1BWP12T r0_reg_9_ ( .D(n2626), .CP(clk), .Q(r0[9]) );
  DFQD1BWP12T r0_reg_8_ ( .D(n2625), .CP(clk), .Q(r0[8]) );
  DFQD1BWP12T r0_reg_7_ ( .D(n2624), .CP(clk), .Q(r0[7]) );
  DFQD1BWP12T r0_reg_6_ ( .D(n2623), .CP(clk), .Q(r0[6]) );
  DFQD1BWP12T r0_reg_5_ ( .D(n2622), .CP(clk), .Q(r0[5]) );
  DFQD1BWP12T r0_reg_4_ ( .D(n2621), .CP(clk), .Q(r0[4]) );
  DFQD1BWP12T r0_reg_3_ ( .D(n2620), .CP(clk), .Q(r0[3]) );
  DFQD1BWP12T r0_reg_2_ ( .D(n2619), .CP(clk), .Q(r0[2]) );
  DFQD1BWP12T r0_reg_1_ ( .D(n2618), .CP(clk), .Q(r0[1]) );
  DFQD1BWP12T r0_reg_0_ ( .D(n2617), .CP(clk), .Q(r0[0]) );
  DFQD1BWP12T r1_reg_31_ ( .D(n2616), .CP(clk), .Q(r1[31]) );
  DFQD1BWP12T r1_reg_30_ ( .D(n2615), .CP(clk), .Q(r1[30]) );
  DFQD1BWP12T r1_reg_29_ ( .D(n2614), .CP(clk), .Q(r1[29]) );
  DFQD1BWP12T r1_reg_28_ ( .D(n2613), .CP(clk), .Q(r1[28]) );
  DFQD1BWP12T r1_reg_27_ ( .D(n2612), .CP(clk), .Q(r1[27]) );
  DFQD1BWP12T r1_reg_26_ ( .D(n2611), .CP(clk), .Q(r1[26]) );
  DFQD1BWP12T r1_reg_25_ ( .D(n2610), .CP(clk), .Q(r1[25]) );
  DFQD1BWP12T r1_reg_24_ ( .D(n2609), .CP(clk), .Q(r1[24]) );
  DFQD1BWP12T r1_reg_23_ ( .D(n2608), .CP(clk), .Q(r1[23]) );
  DFQD1BWP12T r1_reg_22_ ( .D(n2607), .CP(clk), .Q(r1[22]) );
  DFQD1BWP12T r1_reg_21_ ( .D(n2606), .CP(clk), .Q(r1[21]) );
  DFQD1BWP12T r1_reg_20_ ( .D(n2605), .CP(clk), .Q(r1[20]) );
  DFQD1BWP12T r1_reg_19_ ( .D(n2604), .CP(clk), .Q(r1[19]) );
  DFQD1BWP12T r1_reg_18_ ( .D(n2603), .CP(clk), .Q(r1[18]) );
  DFQD1BWP12T r1_reg_17_ ( .D(n2602), .CP(clk), .Q(r1[17]) );
  DFQD1BWP12T r1_reg_16_ ( .D(n2601), .CP(clk), .Q(r1[16]) );
  DFQD1BWP12T r1_reg_15_ ( .D(n2600), .CP(clk), .Q(r1[15]) );
  DFQD1BWP12T r1_reg_14_ ( .D(n2599), .CP(clk), .Q(r1[14]) );
  DFQD1BWP12T r1_reg_13_ ( .D(n2598), .CP(clk), .Q(r1[13]) );
  DFQD1BWP12T r1_reg_12_ ( .D(n2597), .CP(clk), .Q(r1[12]) );
  DFQD1BWP12T r1_reg_11_ ( .D(n2596), .CP(clk), .Q(r1[11]) );
  DFQD1BWP12T r1_reg_10_ ( .D(n2595), .CP(clk), .Q(r1[10]) );
  DFQD1BWP12T r1_reg_9_ ( .D(n2594), .CP(clk), .Q(r1[9]) );
  DFQD1BWP12T r1_reg_8_ ( .D(n2593), .CP(clk), .Q(r1[8]) );
  DFQD1BWP12T r1_reg_7_ ( .D(n2592), .CP(clk), .Q(r1[7]) );
  DFQD1BWP12T r1_reg_6_ ( .D(n2591), .CP(clk), .Q(r1[6]) );
  DFQD1BWP12T r1_reg_5_ ( .D(n2590), .CP(clk), .Q(r1[5]) );
  DFQD1BWP12T r1_reg_4_ ( .D(n2589), .CP(clk), .Q(r1[4]) );
  DFQD1BWP12T r1_reg_3_ ( .D(n2588), .CP(clk), .Q(r1[3]) );
  DFQD1BWP12T r1_reg_2_ ( .D(n2587), .CP(clk), .Q(r1[2]) );
  DFQD1BWP12T r1_reg_1_ ( .D(n2586), .CP(clk), .Q(r1[1]) );
  DFQD1BWP12T r1_reg_0_ ( .D(n2585), .CP(clk), .Q(r1[0]) );
  DFQD1BWP12T r2_reg_31_ ( .D(n2584), .CP(clk), .Q(r2[31]) );
  DFQD1BWP12T r2_reg_30_ ( .D(n2583), .CP(clk), .Q(r2[30]) );
  DFQD1BWP12T r2_reg_29_ ( .D(n2582), .CP(clk), .Q(r2[29]) );
  DFQD1BWP12T r2_reg_28_ ( .D(n2581), .CP(clk), .Q(r2[28]) );
  DFQD1BWP12T r2_reg_27_ ( .D(n2580), .CP(clk), .Q(r2[27]) );
  DFQD1BWP12T r2_reg_26_ ( .D(n2579), .CP(clk), .Q(r2[26]) );
  DFQD1BWP12T r2_reg_25_ ( .D(n2578), .CP(clk), .Q(r2[25]) );
  DFQD1BWP12T r2_reg_24_ ( .D(n2577), .CP(clk), .Q(r2[24]) );
  DFQD1BWP12T r2_reg_23_ ( .D(n2576), .CP(clk), .Q(r2[23]) );
  DFQD1BWP12T r2_reg_22_ ( .D(n2575), .CP(clk), .Q(r2[22]) );
  DFQD1BWP12T r2_reg_21_ ( .D(n2574), .CP(clk), .Q(r2[21]) );
  DFQD1BWP12T r2_reg_20_ ( .D(n2573), .CP(clk), .Q(r2[20]) );
  DFQD1BWP12T r2_reg_19_ ( .D(n2572), .CP(clk), .Q(r2[19]) );
  DFQD1BWP12T r2_reg_18_ ( .D(n2571), .CP(clk), .Q(r2[18]) );
  DFQD1BWP12T r2_reg_17_ ( .D(n2570), .CP(clk), .Q(r2[17]) );
  DFQD1BWP12T r2_reg_16_ ( .D(n2569), .CP(clk), .Q(r2[16]) );
  DFQD1BWP12T r2_reg_15_ ( .D(n2568), .CP(clk), .Q(r2[15]) );
  DFQD1BWP12T r2_reg_14_ ( .D(n2567), .CP(clk), .Q(r2[14]) );
  DFQD1BWP12T r2_reg_13_ ( .D(n2566), .CP(clk), .Q(r2[13]) );
  DFQD1BWP12T r2_reg_12_ ( .D(n2565), .CP(clk), .Q(r2[12]) );
  DFQD1BWP12T r2_reg_11_ ( .D(n2564), .CP(clk), .Q(r2[11]) );
  DFQD1BWP12T r2_reg_10_ ( .D(n2563), .CP(clk), .Q(r2[10]) );
  DFQD1BWP12T r2_reg_9_ ( .D(n2562), .CP(clk), .Q(r2[9]) );
  DFQD1BWP12T r2_reg_8_ ( .D(n2561), .CP(clk), .Q(r2[8]) );
  DFQD1BWP12T r2_reg_7_ ( .D(n2560), .CP(clk), .Q(r2[7]) );
  DFQD1BWP12T r2_reg_6_ ( .D(n2559), .CP(clk), .Q(r2[6]) );
  DFQD1BWP12T r2_reg_5_ ( .D(n2558), .CP(clk), .Q(r2[5]) );
  DFQD1BWP12T r2_reg_4_ ( .D(n2557), .CP(clk), .Q(r2[4]) );
  DFQD1BWP12T r2_reg_3_ ( .D(n2556), .CP(clk), .Q(r2[3]) );
  DFQD1BWP12T r2_reg_2_ ( .D(n2555), .CP(clk), .Q(r2[2]) );
  DFQD1BWP12T r2_reg_1_ ( .D(n2554), .CP(clk), .Q(r2[1]) );
  DFQD1BWP12T r2_reg_0_ ( .D(n2553), .CP(clk), .Q(r2[0]) );
  DFQD1BWP12T r3_reg_31_ ( .D(n2552), .CP(clk), .Q(r3[31]) );
  DFQD1BWP12T r3_reg_30_ ( .D(n2551), .CP(clk), .Q(r3[30]) );
  DFQD1BWP12T r3_reg_29_ ( .D(n2550), .CP(clk), .Q(r3[29]) );
  DFQD1BWP12T r3_reg_28_ ( .D(n2549), .CP(clk), .Q(r3[28]) );
  DFQD1BWP12T r3_reg_27_ ( .D(n2548), .CP(clk), .Q(r3[27]) );
  DFQD1BWP12T r3_reg_26_ ( .D(n2547), .CP(clk), .Q(r3[26]) );
  DFQD1BWP12T r3_reg_25_ ( .D(n2546), .CP(clk), .Q(r3[25]) );
  DFQD1BWP12T r3_reg_24_ ( .D(n2545), .CP(clk), .Q(r3[24]) );
  DFQD1BWP12T r3_reg_23_ ( .D(n2544), .CP(clk), .Q(r3[23]) );
  DFQD1BWP12T r3_reg_22_ ( .D(n2543), .CP(clk), .Q(r3[22]) );
  DFQD1BWP12T r3_reg_21_ ( .D(n2542), .CP(clk), .Q(r3[21]) );
  DFQD1BWP12T r3_reg_20_ ( .D(n2541), .CP(clk), .Q(r3[20]) );
  DFQD1BWP12T r3_reg_19_ ( .D(n2540), .CP(clk), .Q(r3[19]) );
  DFQD1BWP12T r3_reg_18_ ( .D(n2539), .CP(clk), .Q(r3[18]) );
  DFQD1BWP12T r3_reg_17_ ( .D(n2538), .CP(clk), .Q(r3[17]) );
  DFQD1BWP12T r3_reg_16_ ( .D(n2537), .CP(clk), .Q(r3[16]) );
  DFQD1BWP12T r3_reg_15_ ( .D(n2536), .CP(clk), .Q(r3[15]) );
  DFQD1BWP12T r3_reg_14_ ( .D(n2535), .CP(clk), .Q(r3[14]) );
  DFQD1BWP12T r3_reg_13_ ( .D(n2534), .CP(clk), .Q(r3[13]) );
  DFQD1BWP12T r3_reg_12_ ( .D(n2533), .CP(clk), .Q(r3[12]) );
  DFQD1BWP12T r3_reg_11_ ( .D(n2532), .CP(clk), .Q(r3[11]) );
  DFQD1BWP12T r3_reg_10_ ( .D(n2531), .CP(clk), .Q(r3[10]) );
  DFQD1BWP12T r3_reg_9_ ( .D(n2530), .CP(clk), .Q(r3[9]) );
  DFQD1BWP12T r3_reg_8_ ( .D(n2529), .CP(clk), .Q(r3[8]) );
  DFQD1BWP12T r3_reg_7_ ( .D(n2528), .CP(clk), .Q(r3[7]) );
  DFQD1BWP12T r3_reg_6_ ( .D(n2527), .CP(clk), .Q(r3[6]) );
  DFQD1BWP12T r3_reg_5_ ( .D(n2526), .CP(clk), .Q(r3[5]) );
  DFQD1BWP12T r3_reg_4_ ( .D(n2525), .CP(clk), .Q(r3[4]) );
  DFQD1BWP12T r3_reg_3_ ( .D(n2524), .CP(clk), .Q(r3[3]) );
  DFQD1BWP12T r3_reg_2_ ( .D(n2523), .CP(clk), .Q(r3[2]) );
  DFQD1BWP12T r3_reg_1_ ( .D(n2522), .CP(clk), .Q(r3[1]) );
  DFQD1BWP12T r3_reg_0_ ( .D(n2521), .CP(clk), .Q(r3[0]) );
  DFQD1BWP12T r4_reg_31_ ( .D(n2520), .CP(clk), .Q(r4[31]) );
  DFQD1BWP12T r4_reg_30_ ( .D(n2519), .CP(clk), .Q(r4[30]) );
  DFQD1BWP12T r4_reg_29_ ( .D(n2518), .CP(clk), .Q(r4[29]) );
  DFQD1BWP12T r4_reg_28_ ( .D(n2517), .CP(clk), .Q(r4[28]) );
  DFQD1BWP12T r4_reg_27_ ( .D(n2516), .CP(clk), .Q(r4[27]) );
  DFQD1BWP12T r4_reg_26_ ( .D(n2515), .CP(clk), .Q(r4[26]) );
  DFQD1BWP12T r4_reg_25_ ( .D(n2514), .CP(clk), .Q(r4[25]) );
  DFQD1BWP12T r4_reg_24_ ( .D(n2513), .CP(clk), .Q(r4[24]) );
  DFQD1BWP12T r4_reg_23_ ( .D(n2512), .CP(clk), .Q(r4[23]) );
  DFQD1BWP12T r4_reg_22_ ( .D(n2511), .CP(clk), .Q(r4[22]) );
  DFQD1BWP12T r4_reg_21_ ( .D(n2510), .CP(clk), .Q(r4[21]) );
  DFQD1BWP12T r4_reg_20_ ( .D(n2509), .CP(clk), .Q(r4[20]) );
  DFQD1BWP12T r4_reg_19_ ( .D(n2508), .CP(clk), .Q(r4[19]) );
  DFQD1BWP12T r4_reg_18_ ( .D(n2507), .CP(clk), .Q(r4[18]) );
  DFQD1BWP12T r4_reg_17_ ( .D(n2506), .CP(clk), .Q(r4[17]) );
  DFQD1BWP12T r4_reg_16_ ( .D(n2505), .CP(clk), .Q(r4[16]) );
  DFQD1BWP12T r4_reg_15_ ( .D(n2504), .CP(clk), .Q(r4[15]) );
  DFQD1BWP12T r4_reg_14_ ( .D(n2503), .CP(clk), .Q(r4[14]) );
  DFQD1BWP12T r4_reg_13_ ( .D(n2502), .CP(clk), .Q(r4[13]) );
  DFQD1BWP12T r4_reg_12_ ( .D(n2501), .CP(clk), .Q(r4[12]) );
  DFQD1BWP12T r4_reg_11_ ( .D(n2500), .CP(clk), .Q(r4[11]) );
  DFQD1BWP12T r4_reg_10_ ( .D(n2499), .CP(clk), .Q(r4[10]) );
  DFQD1BWP12T r4_reg_9_ ( .D(n2498), .CP(clk), .Q(r4[9]) );
  DFQD1BWP12T r4_reg_8_ ( .D(n2497), .CP(clk), .Q(r4[8]) );
  DFQD1BWP12T r4_reg_7_ ( .D(n2496), .CP(clk), .Q(r4[7]) );
  DFQD1BWP12T r4_reg_6_ ( .D(n2495), .CP(clk), .Q(r4[6]) );
  DFQD1BWP12T r4_reg_5_ ( .D(n2494), .CP(clk), .Q(r4[5]) );
  DFQD1BWP12T r4_reg_4_ ( .D(n2493), .CP(clk), .Q(r4[4]) );
  DFQD1BWP12T r4_reg_3_ ( .D(n2492), .CP(clk), .Q(r4[3]) );
  DFQD1BWP12T r4_reg_2_ ( .D(n2491), .CP(clk), .Q(r4[2]) );
  DFQD1BWP12T r4_reg_1_ ( .D(n2490), .CP(clk), .Q(r4[1]) );
  DFQD1BWP12T r4_reg_0_ ( .D(n2489), .CP(clk), .Q(r4[0]) );
  DFQD1BWP12T r5_reg_31_ ( .D(n2488), .CP(clk), .Q(r5[31]) );
  DFQD1BWP12T r5_reg_30_ ( .D(n2487), .CP(clk), .Q(r5[30]) );
  DFQD1BWP12T r5_reg_29_ ( .D(n2486), .CP(clk), .Q(r5[29]) );
  DFQD1BWP12T r5_reg_28_ ( .D(n2485), .CP(clk), .Q(r5[28]) );
  DFQD1BWP12T r5_reg_27_ ( .D(n2484), .CP(clk), .Q(r5[27]) );
  DFQD1BWP12T r5_reg_26_ ( .D(n2483), .CP(clk), .Q(r5[26]) );
  DFQD1BWP12T r5_reg_25_ ( .D(n2482), .CP(clk), .Q(r5[25]) );
  DFQD1BWP12T r5_reg_24_ ( .D(n2481), .CP(clk), .Q(r5[24]) );
  DFQD1BWP12T r5_reg_23_ ( .D(n2480), .CP(clk), .Q(r5[23]) );
  DFQD1BWP12T r5_reg_22_ ( .D(n2479), .CP(clk), .Q(r5[22]) );
  DFQD1BWP12T r5_reg_21_ ( .D(n2478), .CP(clk), .Q(r5[21]) );
  DFQD1BWP12T r5_reg_20_ ( .D(n2477), .CP(clk), .Q(r5[20]) );
  DFQD1BWP12T r5_reg_19_ ( .D(n2476), .CP(clk), .Q(r5[19]) );
  DFQD1BWP12T r5_reg_18_ ( .D(n2475), .CP(clk), .Q(r5[18]) );
  DFQD1BWP12T r5_reg_17_ ( .D(n2474), .CP(clk), .Q(r5[17]) );
  DFQD1BWP12T r5_reg_16_ ( .D(n2473), .CP(clk), .Q(r5[16]) );
  DFQD1BWP12T r5_reg_15_ ( .D(n2472), .CP(clk), .Q(r5[15]) );
  DFQD1BWP12T r5_reg_14_ ( .D(n2471), .CP(clk), .Q(r5[14]) );
  DFQD1BWP12T r5_reg_13_ ( .D(n2470), .CP(clk), .Q(r5[13]) );
  DFQD1BWP12T r5_reg_12_ ( .D(n2469), .CP(clk), .Q(r5[12]) );
  DFQD1BWP12T r5_reg_11_ ( .D(n2468), .CP(clk), .Q(r5[11]) );
  DFQD1BWP12T r5_reg_10_ ( .D(n2467), .CP(clk), .Q(r5[10]) );
  DFQD1BWP12T r5_reg_9_ ( .D(n2466), .CP(clk), .Q(r5[9]) );
  DFQD1BWP12T r5_reg_8_ ( .D(n2465), .CP(clk), .Q(r5[8]) );
  DFQD1BWP12T r5_reg_7_ ( .D(n2464), .CP(clk), .Q(r5[7]) );
  DFQD1BWP12T r5_reg_6_ ( .D(n2463), .CP(clk), .Q(r5[6]) );
  DFQD1BWP12T r5_reg_5_ ( .D(n2462), .CP(clk), .Q(r5[5]) );
  DFQD1BWP12T r5_reg_3_ ( .D(n2460), .CP(clk), .Q(r5[3]) );
  DFQD1BWP12T r5_reg_2_ ( .D(n2459), .CP(clk), .Q(r5[2]) );
  DFQD1BWP12T r5_reg_1_ ( .D(n2458), .CP(clk), .Q(r5[1]) );
  DFQD1BWP12T r5_reg_0_ ( .D(n2457), .CP(clk), .Q(r5[0]) );
  DFQD1BWP12T r6_reg_31_ ( .D(n2456), .CP(clk), .Q(r6[31]) );
  DFQD1BWP12T r6_reg_30_ ( .D(n2455), .CP(clk), .Q(r6[30]) );
  DFQD1BWP12T r6_reg_29_ ( .D(n2454), .CP(clk), .Q(r6[29]) );
  DFQD1BWP12T r6_reg_28_ ( .D(n2453), .CP(clk), .Q(r6[28]) );
  DFQD1BWP12T r6_reg_27_ ( .D(n2452), .CP(clk), .Q(r6[27]) );
  DFQD1BWP12T r6_reg_26_ ( .D(n2451), .CP(clk), .Q(r6[26]) );
  DFQD1BWP12T r6_reg_25_ ( .D(n2450), .CP(clk), .Q(r6[25]) );
  DFQD1BWP12T r6_reg_24_ ( .D(n2449), .CP(clk), .Q(r6[24]) );
  DFQD1BWP12T r6_reg_23_ ( .D(n2448), .CP(clk), .Q(r6[23]) );
  DFQD1BWP12T r6_reg_22_ ( .D(n2447), .CP(clk), .Q(r6[22]) );
  DFQD1BWP12T r6_reg_21_ ( .D(n2446), .CP(clk), .Q(r6[21]) );
  DFQD1BWP12T r6_reg_20_ ( .D(n2445), .CP(clk), .Q(r6[20]) );
  DFQD1BWP12T r6_reg_19_ ( .D(n2444), .CP(clk), .Q(r6[19]) );
  DFQD1BWP12T r6_reg_18_ ( .D(n2443), .CP(clk), .Q(r6[18]) );
  DFQD1BWP12T r6_reg_17_ ( .D(n2442), .CP(clk), .Q(r6[17]) );
  DFQD1BWP12T r6_reg_16_ ( .D(n2441), .CP(clk), .Q(r6[16]) );
  DFQD1BWP12T r6_reg_15_ ( .D(n2440), .CP(clk), .Q(r6[15]) );
  DFQD1BWP12T r6_reg_14_ ( .D(n2439), .CP(clk), .Q(r6[14]) );
  DFQD1BWP12T r6_reg_13_ ( .D(n2438), .CP(clk), .Q(r6[13]) );
  DFQD1BWP12T r6_reg_12_ ( .D(n2437), .CP(clk), .Q(r6[12]) );
  DFQD1BWP12T r6_reg_11_ ( .D(n2436), .CP(clk), .Q(r6[11]) );
  DFQD1BWP12T r6_reg_10_ ( .D(n2435), .CP(clk), .Q(r6[10]) );
  DFQD1BWP12T r6_reg_9_ ( .D(n2434), .CP(clk), .Q(r6[9]) );
  DFQD1BWP12T r6_reg_8_ ( .D(n2433), .CP(clk), .Q(r6[8]) );
  DFQD1BWP12T r6_reg_7_ ( .D(n2432), .CP(clk), .Q(r6[7]) );
  DFQD1BWP12T r6_reg_6_ ( .D(n2431), .CP(clk), .Q(r6[6]) );
  DFQD1BWP12T r6_reg_5_ ( .D(n2430), .CP(clk), .Q(r6[5]) );
  DFQD1BWP12T r6_reg_4_ ( .D(n2429), .CP(clk), .Q(r6[4]) );
  DFQD1BWP12T r6_reg_3_ ( .D(n2428), .CP(clk), .Q(r6[3]) );
  DFQD1BWP12T r6_reg_2_ ( .D(n2427), .CP(clk), .Q(r6[2]) );
  DFQD1BWP12T r6_reg_1_ ( .D(n2426), .CP(clk), .Q(r6[1]) );
  DFQD1BWP12T r6_reg_0_ ( .D(n2425), .CP(clk), .Q(r6[0]) );
  DFQD1BWP12T r7_reg_31_ ( .D(n2424), .CP(clk), .Q(r7[31]) );
  DFQD1BWP12T r7_reg_30_ ( .D(n2423), .CP(clk), .Q(r7[30]) );
  DFQD1BWP12T r7_reg_29_ ( .D(n2422), .CP(clk), .Q(r7[29]) );
  DFQD1BWP12T r7_reg_28_ ( .D(n2421), .CP(clk), .Q(r7[28]) );
  DFQD1BWP12T r7_reg_27_ ( .D(n2420), .CP(clk), .Q(r7[27]) );
  DFQD1BWP12T r7_reg_26_ ( .D(n2419), .CP(clk), .Q(r7[26]) );
  DFQD1BWP12T r7_reg_25_ ( .D(n2418), .CP(clk), .Q(r7[25]) );
  DFQD1BWP12T r7_reg_24_ ( .D(n2417), .CP(clk), .Q(r7[24]) );
  DFQD1BWP12T r7_reg_23_ ( .D(n2416), .CP(clk), .Q(r7[23]) );
  DFQD1BWP12T r7_reg_22_ ( .D(n2415), .CP(clk), .Q(r7[22]) );
  DFQD1BWP12T r7_reg_21_ ( .D(n2414), .CP(clk), .Q(r7[21]) );
  DFQD1BWP12T r7_reg_20_ ( .D(n2413), .CP(clk), .Q(r7[20]) );
  DFQD1BWP12T r7_reg_19_ ( .D(n2412), .CP(clk), .Q(r7[19]) );
  DFQD1BWP12T r7_reg_18_ ( .D(n2411), .CP(clk), .Q(r7[18]) );
  DFQD1BWP12T r7_reg_17_ ( .D(n2410), .CP(clk), .Q(r7[17]) );
  DFQD1BWP12T r7_reg_16_ ( .D(n2409), .CP(clk), .Q(r7[16]) );
  DFQD1BWP12T r7_reg_15_ ( .D(n2408), .CP(clk), .Q(r7[15]) );
  DFQD1BWP12T r7_reg_14_ ( .D(n2407), .CP(clk), .Q(r7[14]) );
  DFQD1BWP12T r7_reg_13_ ( .D(n2406), .CP(clk), .Q(r7[13]) );
  DFQD1BWP12T r7_reg_12_ ( .D(n2405), .CP(clk), .Q(r7[12]) );
  DFQD1BWP12T r7_reg_11_ ( .D(n2404), .CP(clk), .Q(r7[11]) );
  DFQD1BWP12T r7_reg_10_ ( .D(n2403), .CP(clk), .Q(r7[10]) );
  DFQD1BWP12T r7_reg_9_ ( .D(n2402), .CP(clk), .Q(r7[9]) );
  DFQD1BWP12T r7_reg_8_ ( .D(n2401), .CP(clk), .Q(r7[8]) );
  DFQD1BWP12T r7_reg_7_ ( .D(n2400), .CP(clk), .Q(r7[7]) );
  DFQD1BWP12T r7_reg_6_ ( .D(n2399), .CP(clk), .Q(r7[6]) );
  DFQD1BWP12T r7_reg_5_ ( .D(n2398), .CP(clk), .Q(r7[5]) );
  DFQD1BWP12T r7_reg_4_ ( .D(n2397), .CP(clk), .Q(r7[4]) );
  DFQD1BWP12T r7_reg_3_ ( .D(n2396), .CP(clk), .Q(r7[3]) );
  DFQD1BWP12T r7_reg_2_ ( .D(n2395), .CP(clk), .Q(r7[2]) );
  DFQD1BWP12T r7_reg_1_ ( .D(n2394), .CP(clk), .Q(r7[1]) );
  DFQD1BWP12T r7_reg_0_ ( .D(n2393), .CP(clk), .Q(r7[0]) );
  DFQD1BWP12T r8_reg_31_ ( .D(n2392), .CP(clk), .Q(r8[31]) );
  DFQD1BWP12T r8_reg_30_ ( .D(n2391), .CP(clk), .Q(r8[30]) );
  DFQD1BWP12T r8_reg_29_ ( .D(n2390), .CP(clk), .Q(r8[29]) );
  DFQD1BWP12T r8_reg_28_ ( .D(n2389), .CP(clk), .Q(r8[28]) );
  DFQD1BWP12T r8_reg_27_ ( .D(n2388), .CP(clk), .Q(r8[27]) );
  DFQD1BWP12T r8_reg_26_ ( .D(n2387), .CP(clk), .Q(r8[26]) );
  DFQD1BWP12T r8_reg_25_ ( .D(n2386), .CP(clk), .Q(r8[25]) );
  DFQD1BWP12T r8_reg_24_ ( .D(n2385), .CP(clk), .Q(r8[24]) );
  DFQD1BWP12T r8_reg_23_ ( .D(n2384), .CP(clk), .Q(r8[23]) );
  DFQD1BWP12T r8_reg_22_ ( .D(n2383), .CP(clk), .Q(r8[22]) );
  DFQD1BWP12T r8_reg_21_ ( .D(n2382), .CP(clk), .Q(r8[21]) );
  DFQD1BWP12T r8_reg_20_ ( .D(n2381), .CP(clk), .Q(r8[20]) );
  DFQD1BWP12T r8_reg_19_ ( .D(n2380), .CP(clk), .Q(r8[19]) );
  DFQD1BWP12T r8_reg_18_ ( .D(n2379), .CP(clk), .Q(r8[18]) );
  DFQD1BWP12T r8_reg_17_ ( .D(n2378), .CP(clk), .Q(r8[17]) );
  DFQD1BWP12T r8_reg_16_ ( .D(n2377), .CP(clk), .Q(r8[16]) );
  DFQD1BWP12T r8_reg_15_ ( .D(n2376), .CP(clk), .Q(r8[15]) );
  DFQD1BWP12T r8_reg_14_ ( .D(n2375), .CP(clk), .Q(r8[14]) );
  DFQD1BWP12T r8_reg_13_ ( .D(n2374), .CP(clk), .Q(r8[13]) );
  DFQD1BWP12T r8_reg_12_ ( .D(n2373), .CP(clk), .Q(r8[12]) );
  DFQD1BWP12T r8_reg_11_ ( .D(n2372), .CP(clk), .Q(r8[11]) );
  DFQD1BWP12T r8_reg_10_ ( .D(n2371), .CP(clk), .Q(r8[10]) );
  DFQD1BWP12T r8_reg_9_ ( .D(n2370), .CP(clk), .Q(r8[9]) );
  DFQD1BWP12T r8_reg_8_ ( .D(n2369), .CP(clk), .Q(r8[8]) );
  DFQD1BWP12T r8_reg_7_ ( .D(n2368), .CP(clk), .Q(r8[7]) );
  DFQD1BWP12T r8_reg_6_ ( .D(n2367), .CP(clk), .Q(r8[6]) );
  DFQD1BWP12T r8_reg_5_ ( .D(n2366), .CP(clk), .Q(r8[5]) );
  DFQD1BWP12T r8_reg_4_ ( .D(n2365), .CP(clk), .Q(r8[4]) );
  DFQD1BWP12T r8_reg_3_ ( .D(n2364), .CP(clk), .Q(r8[3]) );
  DFQD1BWP12T r8_reg_2_ ( .D(n2363), .CP(clk), .Q(r8[2]) );
  DFQD1BWP12T r8_reg_1_ ( .D(n2362), .CP(clk), .Q(r8[1]) );
  DFQD1BWP12T r8_reg_0_ ( .D(n2361), .CP(clk), .Q(r8[0]) );
  DFQD1BWP12T r9_reg_31_ ( .D(n2360), .CP(clk), .Q(r9[31]) );
  DFQD1BWP12T r9_reg_30_ ( .D(n2359), .CP(clk), .Q(r9[30]) );
  DFQD1BWP12T r9_reg_29_ ( .D(n2358), .CP(clk), .Q(r9[29]) );
  DFQD1BWP12T r9_reg_28_ ( .D(n2357), .CP(clk), .Q(r9[28]) );
  DFQD1BWP12T r9_reg_27_ ( .D(n2356), .CP(clk), .Q(r9[27]) );
  DFQD1BWP12T r9_reg_26_ ( .D(n2355), .CP(clk), .Q(r9[26]) );
  DFQD1BWP12T r9_reg_25_ ( .D(n2354), .CP(clk), .Q(r9[25]) );
  DFQD1BWP12T r9_reg_24_ ( .D(n2353), .CP(clk), .Q(r9[24]) );
  DFQD1BWP12T r9_reg_23_ ( .D(n2352), .CP(clk), .Q(r9[23]) );
  DFQD1BWP12T r9_reg_22_ ( .D(n2351), .CP(clk), .Q(r9[22]) );
  DFQD1BWP12T r9_reg_21_ ( .D(n2350), .CP(clk), .Q(r9[21]) );
  DFQD1BWP12T r9_reg_20_ ( .D(n2349), .CP(clk), .Q(r9[20]) );
  DFQD1BWP12T r9_reg_19_ ( .D(n2348), .CP(clk), .Q(r9[19]) );
  DFQD1BWP12T r9_reg_18_ ( .D(n2347), .CP(clk), .Q(r9[18]) );
  DFQD1BWP12T r9_reg_17_ ( .D(n2346), .CP(clk), .Q(r9[17]) );
  DFQD1BWP12T r9_reg_16_ ( .D(n2345), .CP(clk), .Q(r9[16]) );
  DFQD1BWP12T r9_reg_15_ ( .D(n2344), .CP(clk), .Q(r9[15]) );
  DFQD1BWP12T r9_reg_14_ ( .D(n2343), .CP(clk), .Q(r9[14]) );
  DFQD1BWP12T r9_reg_13_ ( .D(n2342), .CP(clk), .Q(r9[13]) );
  DFQD1BWP12T r9_reg_12_ ( .D(n2341), .CP(clk), .Q(r9[12]) );
  DFQD1BWP12T r9_reg_11_ ( .D(n2340), .CP(clk), .Q(r9[11]) );
  DFQD1BWP12T r9_reg_10_ ( .D(n2339), .CP(clk), .Q(r9[10]) );
  DFQD1BWP12T r9_reg_9_ ( .D(n2338), .CP(clk), .Q(r9[9]) );
  DFQD1BWP12T r9_reg_8_ ( .D(n2337), .CP(clk), .Q(r9[8]) );
  DFQD1BWP12T r9_reg_7_ ( .D(n2336), .CP(clk), .Q(r9[7]) );
  DFQD1BWP12T r9_reg_6_ ( .D(n2335), .CP(clk), .Q(r9[6]) );
  DFQD1BWP12T r9_reg_5_ ( .D(n2334), .CP(clk), .Q(r9[5]) );
  DFQD1BWP12T r9_reg_4_ ( .D(n2333), .CP(clk), .Q(r9[4]) );
  DFQD1BWP12T r9_reg_3_ ( .D(n2332), .CP(clk), .Q(r9[3]) );
  DFQD1BWP12T r9_reg_2_ ( .D(n2331), .CP(clk), .Q(r9[2]) );
  DFQD1BWP12T r9_reg_0_ ( .D(n2329), .CP(clk), .Q(r9[0]) );
  DFQD1BWP12T r10_reg_31_ ( .D(n2328), .CP(clk), .Q(r10[31]) );
  DFQD1BWP12T r10_reg_30_ ( .D(n2327), .CP(clk), .Q(r10[30]) );
  DFQD1BWP12T r10_reg_29_ ( .D(n2326), .CP(clk), .Q(r10[29]) );
  DFQD1BWP12T r10_reg_28_ ( .D(n2325), .CP(clk), .Q(r10[28]) );
  DFQD1BWP12T r10_reg_27_ ( .D(n2324), .CP(clk), .Q(r10[27]) );
  DFQD1BWP12T r10_reg_26_ ( .D(n2323), .CP(clk), .Q(r10[26]) );
  DFQD1BWP12T r10_reg_25_ ( .D(n2322), .CP(clk), .Q(r10[25]) );
  DFQD1BWP12T r10_reg_24_ ( .D(n2321), .CP(clk), .Q(r10[24]) );
  DFQD1BWP12T r10_reg_23_ ( .D(n2320), .CP(clk), .Q(r10[23]) );
  DFQD1BWP12T r10_reg_22_ ( .D(n2319), .CP(clk), .Q(r10[22]) );
  DFQD1BWP12T r10_reg_21_ ( .D(n2318), .CP(clk), .Q(r10[21]) );
  DFQD1BWP12T r10_reg_20_ ( .D(n2317), .CP(clk), .Q(r10[20]) );
  DFQD1BWP12T r10_reg_19_ ( .D(n2316), .CP(clk), .Q(r10[19]) );
  DFQD1BWP12T r10_reg_18_ ( .D(n2315), .CP(clk), .Q(r10[18]) );
  DFQD1BWP12T r10_reg_17_ ( .D(n2314), .CP(clk), .Q(r10[17]) );
  DFQD1BWP12T r10_reg_16_ ( .D(n2313), .CP(clk), .Q(r10[16]) );
  DFQD1BWP12T r10_reg_15_ ( .D(n2312), .CP(clk), .Q(r10[15]) );
  DFQD1BWP12T r10_reg_14_ ( .D(n2311), .CP(clk), .Q(r10[14]) );
  DFQD1BWP12T r10_reg_13_ ( .D(n2310), .CP(clk), .Q(r10[13]) );
  DFQD1BWP12T r10_reg_12_ ( .D(n2309), .CP(clk), .Q(r10[12]) );
  DFQD1BWP12T r10_reg_11_ ( .D(n2308), .CP(clk), .Q(r10[11]) );
  DFQD1BWP12T r10_reg_10_ ( .D(n2307), .CP(clk), .Q(r10[10]) );
  DFQD1BWP12T r10_reg_9_ ( .D(n2306), .CP(clk), .Q(r10[9]) );
  DFQD1BWP12T r10_reg_8_ ( .D(n2305), .CP(clk), .Q(r10[8]) );
  DFQD1BWP12T r10_reg_7_ ( .D(n2304), .CP(clk), .Q(r10[7]) );
  DFQD1BWP12T r10_reg_6_ ( .D(n2303), .CP(clk), .Q(r10[6]) );
  DFQD1BWP12T r10_reg_5_ ( .D(n2302), .CP(clk), .Q(r10[5]) );
  DFQD1BWP12T r10_reg_4_ ( .D(n2301), .CP(clk), .Q(r10[4]) );
  DFQD1BWP12T r10_reg_3_ ( .D(n2300), .CP(clk), .Q(r10[3]) );
  DFQD1BWP12T r10_reg_2_ ( .D(n2299), .CP(clk), .Q(r10[2]) );
  DFQD1BWP12T r10_reg_1_ ( .D(n2298), .CP(clk), .Q(r10[1]) );
  DFQD1BWP12T r10_reg_0_ ( .D(n2297), .CP(clk), .Q(r10[0]) );
  DFQD1BWP12T r11_reg_31_ ( .D(n2296), .CP(clk), .Q(r11[31]) );
  DFQD1BWP12T r11_reg_30_ ( .D(n2295), .CP(clk), .Q(r11[30]) );
  DFQD1BWP12T r11_reg_29_ ( .D(n2294), .CP(clk), .Q(r11[29]) );
  DFQD1BWP12T r11_reg_28_ ( .D(n2293), .CP(clk), .Q(r11[28]) );
  DFQD1BWP12T r11_reg_27_ ( .D(n2292), .CP(clk), .Q(r11[27]) );
  DFQD1BWP12T r11_reg_26_ ( .D(n2291), .CP(clk), .Q(r11[26]) );
  DFQD1BWP12T r11_reg_25_ ( .D(n2290), .CP(clk), .Q(r11[25]) );
  DFQD1BWP12T r11_reg_24_ ( .D(n2289), .CP(clk), .Q(r11[24]) );
  DFQD1BWP12T r11_reg_23_ ( .D(n2288), .CP(clk), .Q(r11[23]) );
  DFQD1BWP12T r11_reg_22_ ( .D(n2287), .CP(clk), .Q(r11[22]) );
  DFQD1BWP12T r11_reg_21_ ( .D(n2286), .CP(clk), .Q(r11[21]) );
  DFQD1BWP12T r11_reg_20_ ( .D(n2285), .CP(clk), .Q(r11[20]) );
  DFQD1BWP12T r11_reg_19_ ( .D(n2284), .CP(clk), .Q(r11[19]) );
  DFQD1BWP12T r11_reg_18_ ( .D(n2283), .CP(clk), .Q(r11[18]) );
  DFQD1BWP12T r11_reg_17_ ( .D(n2282), .CP(clk), .Q(r11[17]) );
  DFQD1BWP12T r11_reg_16_ ( .D(n2281), .CP(clk), .Q(r11[16]) );
  DFQD1BWP12T r11_reg_15_ ( .D(n2280), .CP(clk), .Q(r11[15]) );
  DFQD1BWP12T r11_reg_14_ ( .D(n2279), .CP(clk), .Q(r11[14]) );
  DFQD1BWP12T r11_reg_13_ ( .D(n2278), .CP(clk), .Q(r11[13]) );
  DFQD1BWP12T r11_reg_12_ ( .D(n2277), .CP(clk), .Q(r11[12]) );
  DFQD1BWP12T r11_reg_11_ ( .D(n2276), .CP(clk), .Q(r11[11]) );
  DFQD1BWP12T r11_reg_10_ ( .D(n2275), .CP(clk), .Q(r11[10]) );
  DFQD1BWP12T r11_reg_9_ ( .D(n2274), .CP(clk), .Q(r11[9]) );
  DFQD1BWP12T r11_reg_8_ ( .D(n2273), .CP(clk), .Q(r11[8]) );
  DFQD1BWP12T r11_reg_7_ ( .D(n2272), .CP(clk), .Q(r11[7]) );
  DFQD1BWP12T r11_reg_6_ ( .D(n2271), .CP(clk), .Q(r11[6]) );
  DFQD1BWP12T r11_reg_5_ ( .D(n2270), .CP(clk), .Q(r11[5]) );
  DFQD1BWP12T r11_reg_4_ ( .D(n2269), .CP(clk), .Q(r11[4]) );
  DFQD1BWP12T r11_reg_3_ ( .D(n2268), .CP(clk), .Q(r11[3]) );
  DFQD1BWP12T r11_reg_2_ ( .D(n2267), .CP(clk), .Q(r11[2]) );
  DFQD1BWP12T r11_reg_1_ ( .D(n2266), .CP(clk), .Q(r11[1]) );
  DFQD1BWP12T r11_reg_0_ ( .D(n2265), .CP(clk), .Q(r11[0]) );
  DFQD1BWP12T r12_reg_31_ ( .D(n2264), .CP(clk), .Q(r12[31]) );
  DFQD1BWP12T r12_reg_30_ ( .D(n2263), .CP(clk), .Q(r12[30]) );
  DFQD1BWP12T r12_reg_29_ ( .D(n2262), .CP(clk), .Q(r12[29]) );
  DFQD1BWP12T r12_reg_28_ ( .D(n2261), .CP(clk), .Q(r12[28]) );
  DFQD1BWP12T r12_reg_27_ ( .D(n2260), .CP(clk), .Q(r12[27]) );
  DFQD1BWP12T r12_reg_26_ ( .D(n2259), .CP(clk), .Q(r12[26]) );
  DFQD1BWP12T r12_reg_25_ ( .D(n2258), .CP(clk), .Q(r12[25]) );
  DFQD1BWP12T r12_reg_24_ ( .D(n2257), .CP(clk), .Q(r12[24]) );
  DFQD1BWP12T r12_reg_23_ ( .D(n2256), .CP(clk), .Q(r12[23]) );
  DFQD1BWP12T r12_reg_22_ ( .D(n2255), .CP(clk), .Q(r12[22]) );
  DFQD1BWP12T r12_reg_21_ ( .D(n2254), .CP(clk), .Q(r12[21]) );
  DFQD1BWP12T r12_reg_20_ ( .D(n2253), .CP(clk), .Q(r12[20]) );
  DFQD1BWP12T r12_reg_19_ ( .D(n2252), .CP(clk), .Q(r12[19]) );
  DFQD1BWP12T r12_reg_18_ ( .D(n2251), .CP(clk), .Q(r12[18]) );
  DFQD1BWP12T r12_reg_17_ ( .D(n2250), .CP(clk), .Q(r12[17]) );
  DFQD1BWP12T r12_reg_16_ ( .D(n2249), .CP(clk), .Q(r12[16]) );
  DFQD1BWP12T r12_reg_15_ ( .D(n2248), .CP(clk), .Q(r12[15]) );
  DFQD1BWP12T r12_reg_14_ ( .D(n2247), .CP(clk), .Q(r12[14]) );
  DFQD1BWP12T r12_reg_13_ ( .D(n2246), .CP(clk), .Q(r12[13]) );
  DFQD1BWP12T r12_reg_12_ ( .D(n2245), .CP(clk), .Q(r12[12]) );
  DFQD1BWP12T r12_reg_11_ ( .D(n2244), .CP(clk), .Q(r12[11]) );
  DFQD1BWP12T r12_reg_10_ ( .D(n2243), .CP(clk), .Q(r12[10]) );
  DFQD1BWP12T r12_reg_9_ ( .D(n2242), .CP(clk), .Q(r12[9]) );
  DFQD1BWP12T r12_reg_8_ ( .D(n2241), .CP(clk), .Q(r12[8]) );
  DFQD1BWP12T r12_reg_7_ ( .D(n2240), .CP(clk), .Q(r12[7]) );
  DFQD1BWP12T r12_reg_6_ ( .D(n2239), .CP(clk), .Q(r12[6]) );
  DFQD1BWP12T r12_reg_5_ ( .D(n2238), .CP(clk), .Q(r12[5]) );
  DFQD1BWP12T r12_reg_4_ ( .D(n2237), .CP(clk), .Q(r12[4]) );
  DFQD1BWP12T r12_reg_3_ ( .D(n2236), .CP(clk), .Q(r12[3]) );
  DFQD1BWP12T r12_reg_2_ ( .D(n2235), .CP(clk), .Q(r12[2]) );
  DFQD1BWP12T r12_reg_1_ ( .D(n2234), .CP(clk), .Q(r12[1]) );
  DFQD1BWP12T r12_reg_0_ ( .D(n2233), .CP(clk), .Q(r12[0]) );
  DFQD1BWP12T lr_reg_31_ ( .D(n2232), .CP(clk), .Q(lr[31]) );
  DFQD1BWP12T lr_reg_30_ ( .D(n2231), .CP(clk), .Q(lr[30]) );
  DFQD1BWP12T lr_reg_29_ ( .D(n2230), .CP(clk), .Q(lr[29]) );
  DFQD1BWP12T lr_reg_28_ ( .D(n2229), .CP(clk), .Q(lr[28]) );
  DFQD1BWP12T lr_reg_27_ ( .D(n2228), .CP(clk), .Q(lr[27]) );
  DFQD1BWP12T lr_reg_26_ ( .D(n2227), .CP(clk), .Q(lr[26]) );
  DFQD1BWP12T lr_reg_25_ ( .D(n2226), .CP(clk), .Q(lr[25]) );
  DFQD1BWP12T lr_reg_24_ ( .D(n2225), .CP(clk), .Q(lr[24]) );
  DFQD1BWP12T lr_reg_23_ ( .D(n2224), .CP(clk), .Q(lr[23]) );
  DFQD1BWP12T lr_reg_22_ ( .D(n2223), .CP(clk), .Q(lr[22]) );
  DFQD1BWP12T lr_reg_21_ ( .D(n2222), .CP(clk), .Q(lr[21]) );
  DFQD1BWP12T lr_reg_20_ ( .D(n2221), .CP(clk), .Q(lr[20]) );
  DFQD1BWP12T lr_reg_19_ ( .D(n2220), .CP(clk), .Q(lr[19]) );
  DFQD1BWP12T lr_reg_18_ ( .D(n2219), .CP(clk), .Q(lr[18]) );
  DFQD1BWP12T lr_reg_17_ ( .D(n2218), .CP(clk), .Q(lr[17]) );
  DFQD1BWP12T lr_reg_16_ ( .D(n2217), .CP(clk), .Q(lr[16]) );
  DFQD1BWP12T lr_reg_15_ ( .D(n2216), .CP(clk), .Q(lr[15]) );
  DFQD1BWP12T lr_reg_14_ ( .D(n2215), .CP(clk), .Q(lr[14]) );
  DFQD1BWP12T lr_reg_13_ ( .D(n2214), .CP(clk), .Q(lr[13]) );
  DFQD1BWP12T lr_reg_12_ ( .D(n2213), .CP(clk), .Q(lr[12]) );
  DFQD1BWP12T lr_reg_11_ ( .D(n2212), .CP(clk), .Q(lr[11]) );
  DFQD1BWP12T lr_reg_10_ ( .D(n2211), .CP(clk), .Q(lr[10]) );
  DFQD1BWP12T lr_reg_9_ ( .D(n2210), .CP(clk), .Q(lr[9]) );
  DFQD1BWP12T lr_reg_8_ ( .D(n2209), .CP(clk), .Q(lr[8]) );
  DFQD1BWP12T lr_reg_7_ ( .D(n2208), .CP(clk), .Q(lr[7]) );
  DFQD1BWP12T lr_reg_6_ ( .D(n2207), .CP(clk), .Q(lr[6]) );
  DFQD1BWP12T lr_reg_5_ ( .D(n2206), .CP(clk), .Q(lr[5]) );
  DFQD1BWP12T lr_reg_4_ ( .D(n2205), .CP(clk), .Q(lr[4]) );
  DFQD1BWP12T lr_reg_3_ ( .D(n2204), .CP(clk), .Q(lr[3]) );
  DFQD1BWP12T lr_reg_2_ ( .D(n2203), .CP(clk), .Q(lr[2]) );
  DFQD1BWP12T lr_reg_1_ ( .D(n2202), .CP(clk), .Q(lr[1]) );
  DFQD1BWP12T lr_reg_0_ ( .D(n2201), .CP(clk), .Q(lr[0]) );
  DFQD1BWP12T sp_reg_31_ ( .D(spin[31]), .CP(clk), .Q(n[2937]) );
  DFQD1BWP12T sp_reg_30_ ( .D(spin[30]), .CP(clk), .Q(n[2938]) );
  DFQD1BWP12T sp_reg_29_ ( .D(spin[29]), .CP(clk), .Q(n[2939]) );
  DFQD1BWP12T sp_reg_28_ ( .D(spin[28]), .CP(clk), .Q(n[2940]) );
  DFQD1BWP12T sp_reg_27_ ( .D(spin[27]), .CP(clk), .Q(n[2941]) );
  DFQD1BWP12T sp_reg_26_ ( .D(spin[26]), .CP(clk), .Q(n[2942]) );
  DFQD1BWP12T sp_reg_25_ ( .D(spin[25]), .CP(clk), .Q(n[2943]) );
  DFQD1BWP12T sp_reg_24_ ( .D(spin[24]), .CP(clk), .Q(n[2944]) );
  DFQD1BWP12T sp_reg_23_ ( .D(spin[23]), .CP(clk), .Q(n[2945]) );
  DFQD1BWP12T sp_reg_22_ ( .D(spin[22]), .CP(clk), .Q(n[2946]) );
  DFQD1BWP12T sp_reg_21_ ( .D(spin[21]), .CP(clk), .Q(n[2947]) );
  DFQD1BWP12T sp_reg_20_ ( .D(spin[20]), .CP(clk), .Q(n[2948]) );
  DFQD1BWP12T sp_reg_19_ ( .D(spin[19]), .CP(clk), .Q(n[2949]) );
  DFQD1BWP12T sp_reg_18_ ( .D(spin[18]), .CP(clk), .Q(n[2950]) );
  DFQD1BWP12T sp_reg_17_ ( .D(spin[17]), .CP(clk), .Q(n[2951]) );
  DFQD1BWP12T sp_reg_16_ ( .D(spin[16]), .CP(clk), .Q(n[2952]) );
  DFQD1BWP12T sp_reg_15_ ( .D(spin[15]), .CP(clk), .Q(n[2953]) );
  DFQD1BWP12T sp_reg_14_ ( .D(spin[14]), .CP(clk), .Q(n[2954]) );
  DFQD1BWP12T sp_reg_13_ ( .D(spin[13]), .CP(clk), .Q(n[2955]) );
  DFQD1BWP12T sp_reg_12_ ( .D(spin[12]), .CP(clk), .Q(n[2956]) );
  DFQD1BWP12T sp_reg_11_ ( .D(spin[11]), .CP(clk), .Q(n[2957]) );
  DFQD1BWP12T sp_reg_10_ ( .D(spin[10]), .CP(clk), .Q(n[2958]) );
  DFQD1BWP12T sp_reg_9_ ( .D(spin[9]), .CP(clk), .Q(n[2959]) );
  DFQD1BWP12T sp_reg_8_ ( .D(spin[8]), .CP(clk), .Q(n[2960]) );
  DFQD1BWP12T sp_reg_7_ ( .D(spin[7]), .CP(clk), .Q(n[2961]) );
  DFQD1BWP12T sp_reg_6_ ( .D(spin[6]), .CP(clk), .Q(n[2962]) );
  DFQD1BWP12T sp_reg_5_ ( .D(spin[5]), .CP(clk), .Q(n[2963]) );
  DFQD1BWP12T sp_reg_3_ ( .D(spin[3]), .CP(clk), .Q(n[2965]) );
  DFQD1BWP12T sp_reg_2_ ( .D(spin[2]), .CP(clk), .Q(n[2966]) );
  DFQD1BWP12T sp_reg_1_ ( .D(spin[1]), .CP(clk), .Q(n[2967]) );
  DFQD1BWP12T sp_reg_0_ ( .D(spin[0]), .CP(clk), .Q(n[2968]) );
  DFQD1BWP12T pc_reg_31_ ( .D(n2200), .CP(clk), .Q(pc_out[31]) );
  DFQD1BWP12T pc_reg_30_ ( .D(n2199), .CP(clk), .Q(pc_out[30]) );
  DFQD1BWP12T pc_reg_29_ ( .D(n2198), .CP(clk), .Q(pc_out[29]) );
  DFQD1BWP12T pc_reg_28_ ( .D(n2197), .CP(clk), .Q(pc_out[28]) );
  DFQD1BWP12T pc_reg_27_ ( .D(n2196), .CP(clk), .Q(pc_out[27]) );
  DFQD1BWP12T pc_reg_26_ ( .D(n2195), .CP(clk), .Q(pc_out[26]) );
  DFQD1BWP12T pc_reg_25_ ( .D(n2194), .CP(clk), .Q(pc_out[25]) );
  DFQD1BWP12T pc_reg_24_ ( .D(n2193), .CP(clk), .Q(pc_out[24]) );
  DFQD1BWP12T pc_reg_23_ ( .D(n2192), .CP(clk), .Q(pc_out[23]) );
  DFQD1BWP12T pc_reg_22_ ( .D(n2191), .CP(clk), .Q(pc_out[22]) );
  DFQD1BWP12T pc_reg_21_ ( .D(n2190), .CP(clk), .Q(pc_out[21]) );
  DFQD1BWP12T pc_reg_20_ ( .D(n2189), .CP(clk), .Q(pc_out[20]) );
  DFQD1BWP12T pc_reg_19_ ( .D(n2188), .CP(clk), .Q(pc_out[19]) );
  DFQD1BWP12T pc_reg_18_ ( .D(n2187), .CP(clk), .Q(pc_out[18]) );
  DFQD1BWP12T pc_reg_17_ ( .D(n2186), .CP(clk), .Q(pc_out[17]) );
  DFQD1BWP12T pc_reg_16_ ( .D(n2185), .CP(clk), .Q(pc_out[16]) );
  DFQD1BWP12T pc_reg_15_ ( .D(n2184), .CP(clk), .Q(pc_out[15]) );
  DFQD1BWP12T pc_reg_14_ ( .D(n2183), .CP(clk), .Q(pc_out[14]) );
  DFQD1BWP12T pc_reg_13_ ( .D(n2182), .CP(clk), .Q(pc_out[13]) );
  DFQD1BWP12T pc_reg_12_ ( .D(n2181), .CP(clk), .Q(pc_out[12]) );
  DFQD1BWP12T pc_reg_11_ ( .D(n2180), .CP(clk), .Q(pc_out[11]) );
  DFQD1BWP12T pc_reg_10_ ( .D(n2179), .CP(clk), .Q(pc_out[10]) );
  DFQD1BWP12T pc_reg_9_ ( .D(n2178), .CP(clk), .Q(pc_out[9]) );
  DFQD1BWP12T pc_reg_8_ ( .D(n2177), .CP(clk), .Q(pc_out[8]) );
  DFQD1BWP12T pc_reg_7_ ( .D(n2176), .CP(clk), .Q(pc_out[7]) );
  DFQD1BWP12T pc_reg_6_ ( .D(n2175), .CP(clk), .Q(pc_out[6]) );
  DFQD1BWP12T pc_reg_5_ ( .D(n2174), .CP(clk), .Q(pc_out[5]) );
  DFQD1BWP12T pc_reg_4_ ( .D(n2173), .CP(clk), .Q(pc_out[4]) );
  DFQD1BWP12T pc_reg_3_ ( .D(n2172), .CP(clk), .Q(pc_out[3]) );
  DFQD1BWP12T pc_reg_0_ ( .D(n2169), .CP(clk), .Q(pc_out[0]) );
  DFQD1BWP12T cpsr_reg_3_ ( .D(cpsrin[3]), .CP(clk), .Q(cpsr_out[3]) );
  DFQD1BWP12T cpsr_reg_2_ ( .D(cpsrin[2]), .CP(clk), .Q(cpsr_out[2]) );
  DFQD1BWP12T cpsr_reg_1_ ( .D(cpsrin[1]), .CP(clk), .Q(cpsr_out[1]) );
  DFQD1BWP12T cpsr_reg_0_ ( .D(cpsrin[0]), .CP(clk), .Q(cpsr_out[0]) );
  DFQD1BWP12T tmp1_reg_31_ ( .D(n2168), .CP(clk), .Q(tmp1[31]) );
  DFQD1BWP12T tmp1_reg_30_ ( .D(n2167), .CP(clk), .Q(tmp1[30]) );
  DFQD1BWP12T tmp1_reg_29_ ( .D(n2166), .CP(clk), .Q(tmp1[29]) );
  DFQD1BWP12T tmp1_reg_28_ ( .D(n2165), .CP(clk), .Q(tmp1[28]) );
  DFQD1BWP12T tmp1_reg_27_ ( .D(n2164), .CP(clk), .Q(tmp1[27]) );
  DFQD1BWP12T tmp1_reg_26_ ( .D(n2163), .CP(clk), .Q(tmp1[26]) );
  DFQD1BWP12T tmp1_reg_25_ ( .D(n2162), .CP(clk), .Q(tmp1[25]) );
  DFQD1BWP12T tmp1_reg_24_ ( .D(n2161), .CP(clk), .Q(tmp1[24]) );
  DFQD1BWP12T tmp1_reg_23_ ( .D(n2160), .CP(clk), .Q(tmp1[23]) );
  DFQD1BWP12T tmp1_reg_22_ ( .D(n2159), .CP(clk), .Q(tmp1[22]) );
  DFQD1BWP12T tmp1_reg_21_ ( .D(n2158), .CP(clk), .Q(tmp1[21]) );
  DFQD1BWP12T tmp1_reg_20_ ( .D(n2157), .CP(clk), .Q(tmp1[20]) );
  DFQD1BWP12T tmp1_reg_19_ ( .D(n2156), .CP(clk), .Q(tmp1[19]) );
  DFQD1BWP12T tmp1_reg_18_ ( .D(n2155), .CP(clk), .Q(tmp1[18]) );
  DFQD1BWP12T tmp1_reg_17_ ( .D(n2154), .CP(clk), .Q(tmp1[17]) );
  DFQD1BWP12T tmp1_reg_16_ ( .D(n2153), .CP(clk), .Q(tmp1[16]) );
  DFQD1BWP12T tmp1_reg_15_ ( .D(n2152), .CP(clk), .Q(tmp1[15]) );
  DFQD1BWP12T tmp1_reg_14_ ( .D(n2151), .CP(clk), .Q(tmp1[14]) );
  DFQD1BWP12T tmp1_reg_13_ ( .D(n2150), .CP(clk), .Q(tmp1[13]) );
  DFQD1BWP12T tmp1_reg_12_ ( .D(n2149), .CP(clk), .Q(tmp1[12]) );
  DFQD1BWP12T tmp1_reg_11_ ( .D(n2148), .CP(clk), .Q(tmp1[11]) );
  DFQD1BWP12T tmp1_reg_10_ ( .D(n2147), .CP(clk), .Q(tmp1[10]) );
  DFQD1BWP12T tmp1_reg_9_ ( .D(n2146), .CP(clk), .Q(tmp1[9]) );
  DFQD1BWP12T tmp1_reg_8_ ( .D(n2145), .CP(clk), .Q(tmp1[8]) );
  DFQD1BWP12T tmp1_reg_7_ ( .D(n2144), .CP(clk), .Q(tmp1[7]) );
  DFQD1BWP12T tmp1_reg_6_ ( .D(n2143), .CP(clk), .Q(tmp1[6]) );
  DFQD1BWP12T tmp1_reg_5_ ( .D(n2142), .CP(clk), .Q(tmp1[5]) );
  DFQD1BWP12T tmp1_reg_4_ ( .D(n2141), .CP(clk), .Q(tmp1[4]) );
  DFQD1BWP12T tmp1_reg_3_ ( .D(n2140), .CP(clk), .Q(tmp1[3]) );
  DFQD1BWP12T tmp1_reg_2_ ( .D(n2139), .CP(clk), .Q(tmp1[2]) );
  DFQD1BWP12T tmp1_reg_1_ ( .D(n2138), .CP(clk), .Q(tmp1[1]) );
  DFQD1BWP12T tmp1_reg_0_ ( .D(n2136), .CP(clk), .Q(tmp1[0]) );
  DFQD1BWP12T r9_reg_1_ ( .D(n2330), .CP(clk), .Q(r9[1]) );
  DFQD1BWP12T r5_reg_4_ ( .D(n2461), .CP(clk), .Q(r5[4]) );
  DFQD1BWP12T sp_reg_4_ ( .D(spin[4]), .CP(clk), .Q(n[2964]) );
  DFQD2BWP12T pc_reg_2_ ( .D(n2171), .CP(clk), .Q(pc_out[2]) );
  DFQD1BWP12T pc_reg_1_ ( .D(n2170), .CP(clk), .Q(pc_out[1]) );
  ND4D2BWP12T U3 ( .A1(n391), .A2(n390), .A3(n389), .A4(n388), .ZN(
        regB_out[25]) );
  INVD1BWP12T U4 ( .I(n1720), .ZN(n1725) );
  AN3XD1BWP12T U5 ( .A1(n376), .A2(n375), .A3(n374), .Z(n379) );
  OAI22D1BWP12T U6 ( .A1(n842), .A2(n2680), .B1(n2679), .B2(n1139), .ZN(n138)
         );
  NR2D1BWP12T U7 ( .A1(n2860), .A2(n840), .ZN(n841) );
  ND2D1BWP12T U8 ( .A1(write1_in[23]), .A2(n2920), .ZN(n1645) );
  ND3D1BWP12T U9 ( .A1(n790), .A2(n789), .A3(n788), .ZN(regA_out[27]) );
  AOI22D1BWP12T U10 ( .A1(r9[1]), .A2(n105), .B1(n2753), .B2(r4[1]), .ZN(n111)
         );
  ND4D1BWP12T U11 ( .A1(n836), .A2(n835), .A3(n834), .A4(n833), .ZN(
        regA_out[19]) );
  ND3D1BWP12T U12 ( .A1(n589), .A2(n588), .A3(n587), .ZN(n590) );
  AOI21D1BWP12T U13 ( .A1(n2819), .A2(r9[7]), .B(n618), .ZN(n619) );
  NR2D1BWP12T U14 ( .A1(n2880), .A2(n685), .ZN(n618) );
  ND2D1BWP12T U15 ( .A1(n461), .A2(n460), .ZN(n463) );
  MOAI22D0BWP12T U16 ( .A1(n1875), .A2(n2666), .B1(n2745), .B2(
        immediate2_in[2]), .ZN(n464) );
  ND2D1BWP12T U17 ( .A1(write1_in[22]), .A2(n2920), .ZN(n1700) );
  INR3D0BWP12T U18 ( .A1(n902), .B1(write1_sel[2]), .B2(write1_sel[1]), .ZN(
        n191) );
  AOI22D1BWP12T U19 ( .A1(n2814), .A2(r1[13]), .B1(n2813), .B2(r12[13]), .ZN(
        n720) );
  ND3D1BWP12T U20 ( .A1(n369), .A2(n368), .A3(n367), .ZN(regA_out[16]) );
  INVD2BWP12T U21 ( .I(n104), .ZN(n309) );
  INVD3BWP12T U22 ( .I(readA_sel[2]), .ZN(n1856) );
  AOI21D1BWP12T U23 ( .A1(write1_in[2]), .A2(n2920), .B(n433), .ZN(n434) );
  NR2D1BWP12T U24 ( .A1(n303), .A2(n302), .ZN(n1622) );
  NR2D1BWP12T U25 ( .A1(n303), .A2(n301), .ZN(n1625) );
  INVD1BWP12T U26 ( .I(n2924), .ZN(n1690) );
  INVD1BWP12T U27 ( .I(n1740), .ZN(n1735) );
  OAI21D1BWP12T U28 ( .A1(n1679), .A2(n2916), .B(n2915), .ZN(n2927) );
  INVD1BWP12T U29 ( .I(write1_in[29]), .ZN(n1679) );
  AOI21D1BWP12T U30 ( .A1(write1_in[30]), .A2(n2920), .B(n2922), .ZN(n2931) );
  INVD1BWP12T U31 ( .I(n1617), .ZN(n1443) );
  INVD1BWP12T U32 ( .I(n1615), .ZN(n1521) );
  INR2D1BWP12T U33 ( .A1(n181), .B1(n286), .ZN(n1614) );
  NR2D1BWP12T U34 ( .A1(n152), .A2(n153), .ZN(n1617) );
  INVD1BWP12T U35 ( .I(n1607), .ZN(n1475) );
  INR2D1BWP12T U36 ( .A1(n175), .B1(n299), .ZN(n1607) );
  NR2D1BWP12T U37 ( .A1(n165), .A2(n166), .ZN(n1609) );
  NR2D1BWP12T U38 ( .A1(n177), .A2(n178), .ZN(n1599) );
  INVD1BWP12T U39 ( .I(n1436), .ZN(n1597) );
  NR3D1BWP12T U40 ( .A1(n289), .A2(n291), .A3(n288), .ZN(n1510) );
  INVD1BWP12T U41 ( .I(n1508), .ZN(n1530) );
  INVD1BWP12T U42 ( .I(n1510), .ZN(n1533) );
  INVD1BWP12T U43 ( .I(n1514), .ZN(n1526) );
  ND2D1BWP12T U44 ( .A1(n285), .A2(n175), .ZN(n1527) );
  INVD1BWP12T U45 ( .I(n1591), .ZN(n1481) );
  INR2D1BWP12T U46 ( .A1(n191), .B1(n286), .ZN(n1591) );
  NR2D1BWP12T U47 ( .A1(n193), .A2(n194), .ZN(n1594) );
  ND2D1BWP12T U48 ( .A1(n191), .A2(n175), .ZN(n1478) );
  NR2D1BWP12T U49 ( .A1(n162), .A2(n163), .ZN(n1604) );
  INVD1BWP12T U50 ( .I(n1478), .ZN(n1602) );
  NR2D1BWP12T U51 ( .A1(n170), .A2(n171), .ZN(n1570) );
  INVD1BWP12T U52 ( .I(n1451), .ZN(n1567) );
  INVD1BWP12T U53 ( .I(n1555), .ZN(n1490) );
  INR2D1BWP12T U54 ( .A1(n187), .B1(n299), .ZN(n1555) );
  INVD1BWP12T U55 ( .I(n1444), .ZN(n1558) );
  NR2D1BWP12T U56 ( .A1(n185), .A2(n186), .ZN(n1564) );
  INVD1BWP12T U57 ( .I(n1445), .ZN(n1561) );
  NR2D1BWP12T U58 ( .A1(n167), .A2(n168), .ZN(n1582) );
  INVD1BWP12T U59 ( .I(n1449), .ZN(n1579) );
  AN3XD1BWP12T U60 ( .A1(n150), .A2(n902), .A3(n149), .Z(n1504) );
  INVD1BWP12T U61 ( .I(n1457), .ZN(n1573) );
  AN3XD1BWP12T U62 ( .A1(n144), .A2(n902), .A3(n143), .Z(n1511) );
  ND2D1BWP12T U63 ( .A1(n187), .A2(n285), .ZN(n1523) );
  INVD1BWP12T U64 ( .I(n1511), .ZN(n1522) );
  NR2D1BWP12T U65 ( .A1(n179), .A2(n180), .ZN(n1588) );
  INVD1BWP12T U66 ( .I(write1_in[12]), .ZN(n535) );
  INVD1BWP12T U67 ( .I(write1_in[20]), .ZN(n1423) );
  INVD1BWP12T U68 ( .I(write1_in[21]), .ZN(n1456) );
  INVD1BWP12T U69 ( .I(write1_in[28]), .ZN(n523) );
  INVD1BWP12T U70 ( .I(write1_in[29]), .ZN(n1482) );
  INVD1BWP12T U71 ( .I(write1_in[30]), .ZN(n1491) );
  BUFFD2BWP12T U72 ( .I(write1_in[31]), .Z(n1621) );
  NR2D1BWP12T U73 ( .A1(n173), .A2(n174), .ZN(n1552) );
  INVD1BWP12T U74 ( .I(n1249), .ZN(n1322) );
  INVD1BWP12T U75 ( .I(n1170), .ZN(n1321) );
  INVD1BWP12T U76 ( .I(n1304), .ZN(n1280) );
  INVD1BWP12T U77 ( .I(n1303), .ZN(n1279) );
  INVD1BWP12T U78 ( .I(n1308), .ZN(n1281) );
  INVD1BWP12T U79 ( .I(n1309), .ZN(n1282) );
  INVD1BWP12T U80 ( .I(n1301), .ZN(n1275) );
  INVD1BWP12T U81 ( .I(n1302), .ZN(n1276) );
  INVD1BWP12T U82 ( .I(n1306), .ZN(n1277) );
  INVD1BWP12T U83 ( .I(n1307), .ZN(n1278) );
  INVD1BWP12T U84 ( .I(n1287), .ZN(n1320) );
  INVD1BWP12T U85 ( .I(readC_sel[4]), .ZN(n1295) );
  INR3D0BWP12T U86 ( .A1(n457), .B1(n456), .B2(n455), .ZN(n458) );
  INR3D0BWP12T U87 ( .A1(n447), .B1(n446), .B2(n445), .ZN(n459) );
  NR2D2BWP12T U88 ( .A1(readB_sel[1]), .A2(readB_sel[2]), .ZN(n126) );
  INVD2BWP12T U89 ( .I(n2864), .ZN(n2808) );
  INVD2BWP12T U90 ( .I(n309), .ZN(n2135) );
  INVD1BWP12T U91 ( .I(n225), .ZN(n2666) );
  INVD2BWP12T U92 ( .I(n2749), .ZN(n2671) );
  INVD2BWP12T U93 ( .I(n2761), .ZN(n2679) );
  INR2D2BWP12T U94 ( .A1(n124), .B1(n125), .ZN(n2747) );
  INVD2BWP12T U95 ( .I(n210), .ZN(n2754) );
  INR2XD2BWP12T U96 ( .A1(n124), .B1(n130), .ZN(n2755) );
  INR2XD2BWP12T U97 ( .A1(n128), .B1(n130), .ZN(n2764) );
  ND2D3BWP12T U98 ( .A1(n348), .A2(n351), .ZN(n2868) );
  AN2D1BWP12T U99 ( .A1(next_cpsr_in[2]), .A2(n902), .Z(cpsrin[2]) );
  NR2D1BWP12T U100 ( .A1(n1722), .A2(n1721), .ZN(n1729) );
  AOI22D1BWP12T U101 ( .A1(r3[16]), .A2(n2810), .B1(n2809), .B2(r5[16]), .ZN(
        n355) );
  AOI22D1BWP12T U102 ( .A1(r3[19]), .A2(n2810), .B1(n2809), .B2(r5[19]), .ZN(
        n826) );
  AOI22D1BWP12T U103 ( .A1(n2814), .A2(r1[19]), .B1(n2708), .B2(r12[19]), .ZN(
        n824) );
  INR2D1BWP12T U104 ( .A1(r7[3]), .B1(n2868), .ZN(n879) );
  MAOI22D0BWP12T U105 ( .A1(n2814), .A2(r1[28]), .B1(n1791), .B2(n2851), .ZN(
        n1792) );
  OAI22D1BWP12T U106 ( .A1(n1929), .A2(n2680), .B1(n2679), .B2(n1928), .ZN(
        n1939) );
  NR4D0BWP12T U107 ( .A1(n2677), .A2(n2676), .A3(n2675), .A4(n2674), .ZN(n2699) );
  INR3D0BWP12T U108 ( .A1(n882), .B1(n881), .B2(n880), .ZN(n886) );
  ND2D1BWP12T U109 ( .A1(n654), .A2(n653), .ZN(n656) );
  AN2D1BWP12T U110 ( .A1(n878), .A2(n877), .Z(n887) );
  IND3D0BWP12T U111 ( .A1(n155), .B1(write1_sel[3]), .B2(n141), .ZN(n286) );
  NR2D0BWP12T U112 ( .A1(n298), .A2(write1_sel[4]), .ZN(n175) );
  INR3D0BWP12T U113 ( .A1(write1_sel[4]), .B1(n299), .B2(n298), .ZN(n1620) );
  INR2D0BWP12T U114 ( .A1(n193), .B1(n194), .ZN(n1507) );
  INR2D0BWP12T U115 ( .A1(n170), .B1(n171), .ZN(n1505) );
  IND2D0BWP12T U116 ( .A1(n569), .B1(n902), .ZN(n65) );
  AOI21D0BWP12T U117 ( .A1(r9[2]), .A2(n2819), .B(n1876), .ZN(n1) );
  AOI22D0BWP12T U118 ( .A1(r2[2]), .A2(n2890), .B1(r4[2]), .B2(n2791), .ZN(n2)
         );
  OAI211D0BWP12T U119 ( .A1(n2884), .A2(n1877), .B(n1), .C(n2), .ZN(n1878) );
  AO22D1BWP12T U120 ( .A1(write2_in[23]), .A2(n2916), .B1(n2920), .B2(
        write1_in[23]), .Z(n2900) );
  IND2D0BWP12T U121 ( .A1(n65), .B1(next_pc_en_BAR), .ZN(n2924) );
  IND2D0BWP12T U122 ( .A1(n286), .B1(n285), .ZN(n1532) );
  MAOI22D0BWP12T U123 ( .A1(n1469), .A2(n1468), .B1(n1469), .B2(n1468), .ZN(n3) );
  AO222D0BWP12T U124 ( .A1(pc_out[13]), .A2(n1690), .B1(n3), .B2(n2914), .C1(
        next_pc_in[13]), .C2(n1488), .Z(n2182) );
  AOI22D0BWP12T U125 ( .A1(n2809), .A2(r5[30]), .B1(n2810), .B2(r3[30]), .ZN(
        n4) );
  AOI22D0BWP12T U126 ( .A1(n2807), .A2(n[2938]), .B1(r11[30]), .B2(n2808), 
        .ZN(n5) );
  AN4XD1BWP12T U127 ( .A1(n4), .A2(n5), .A3(n818), .A4(n819), .Z(n822) );
  MAOI22D0BWP12T U128 ( .A1(n2791), .A2(r4[9]), .B1(n2789), .B2(n543), .ZN(n93) );
  INR2D0BWP12T U129 ( .A1(write2_in[28]), .B1(n2920), .ZN(n2910) );
  MOAI22D0BWP12T U130 ( .A1(n2901), .A2(n2924), .B1(next_pc_in[24]), .B2(n1488), .ZN(n2902) );
  IND2D0BWP12T U131 ( .A1(n299), .B1(n182), .ZN(n1451) );
  IND2D0BWP12T U132 ( .A1(n144), .B1(n143), .ZN(n1524) );
  MAOI22D0BWP12T U133 ( .A1(n1494), .A2(n1493), .B1(n1494), .B2(n1493), .ZN(n6) );
  AO222D0BWP12T U134 ( .A1(pc_out[14]), .A2(n1690), .B1(n6), .B2(n2914), .C1(
        next_pc_in[14]), .C2(n1488), .Z(n2183) );
  MOAI22D0BWP12T U135 ( .A1(n2868), .A2(n2010), .B1(n2811), .B2(pc_out[4]), 
        .ZN(n1860) );
  INR2D0BWP12T U136 ( .A1(write2_in[30]), .B1(n2920), .ZN(n2922) );
  MOAI22D0BWP12T U137 ( .A1(n1634), .A2(n2924), .B1(next_pc_in[25]), .B2(n1488), .ZN(n1635) );
  NR2D0BWP12T U138 ( .A1(write2_sel[2]), .A2(n290), .ZN(n7) );
  AOI211D1BWP12T U139 ( .A1(n292), .A2(n7), .B(n291), .C(reset), .ZN(n1508) );
  INR2D0BWP12T U140 ( .A1(n162), .B1(n163), .ZN(n1603) );
  INR2D0BWP12T U141 ( .A1(n185), .B1(n186), .ZN(n1520) );
  MAOI22D0BWP12T U142 ( .A1(n438), .A2(n437), .B1(n438), .B2(n437), .ZN(n8) );
  AO222D0BWP12T U143 ( .A1(pc_out[3]), .A2(n1690), .B1(n8), .B2(n2914), .C1(
        next_pc_in[3]), .C2(n1488), .Z(n2172) );
  NR2D0BWP12T U144 ( .A1(n1494), .A2(n1493), .ZN(n9) );
  MOAI22D0BWP12T U145 ( .A1(n9), .A2(n1492), .B1(n9), .B2(n1492), .ZN(n10) );
  AO222D0BWP12T U146 ( .A1(n10), .A2(n2914), .B1(next_pc_in[15]), .B2(n1488), 
        .C1(pc_out[15]), .C2(n1690), .Z(n2184) );
  MAOI22D0BWP12T U147 ( .A1(n2813), .A2(r12[2]), .B1(n2872), .B2(n1885), .ZN(
        n1886) );
  OAI22D0BWP12T U148 ( .A1(n1856), .A2(n1857), .B1(n1855), .B2(r2[4]), .ZN(n11) );
  OAI31D0BWP12T U149 ( .A1(readA_sel[1]), .A2(readA_sel[2]), .A3(r0[4]), .B(
        n1853), .ZN(n12) );
  AOI21D0BWP12T U150 ( .A1(r9[4]), .A2(n2819), .B(n1858), .ZN(n13) );
  OAI21D0BWP12T U151 ( .A1(n11), .A2(n12), .B(n13), .ZN(n1859) );
  INR3D0BWP12T U152 ( .A1(write1_sel[2]), .B1(reset), .B2(write1_sel[1]), .ZN(
        n181) );
  MAOI22D0BWP12T U153 ( .A1(n1488), .A2(next_pc_in[26]), .B1(n2924), .B2(n1707), .ZN(n1708) );
  INR2D0BWP12T U154 ( .A1(n1719), .B1(n1725), .ZN(n1721) );
  MAOI22D0BWP12T U155 ( .A1(n1368), .A2(n1367), .B1(n1368), .B2(n1367), .ZN(
        n14) );
  AO222D0BWP12T U156 ( .A1(n2914), .A2(n14), .B1(pc_out[4]), .B2(n1690), .C1(
        next_pc_in[4]), .C2(n1488), .Z(n2173) );
  MOAI22D0BWP12T U157 ( .A1(n1535), .A2(n1534), .B1(n1535), .B2(n1534), .ZN(
        n15) );
  AO222D0BWP12T U158 ( .A1(n15), .A2(n2914), .B1(next_pc_in[16]), .B2(n1488), 
        .C1(pc_out[16]), .C2(n1690), .Z(n2185) );
  MAOI22D0BWP12T U159 ( .A1(n2776), .A2(pc_out[2]), .B1(n2868), .B2(n1881), 
        .ZN(n1890) );
  MAOI22D0BWP12T U160 ( .A1(n2891), .A2(lr[11]), .B1(n2822), .B2(n1933), .ZN(
        n795) );
  MAOI22D0BWP12T U161 ( .A1(n2791), .A2(r4[1]), .B1(n2884), .B2(n849), .ZN(
        n864) );
  AN2D0BWP12T U162 ( .A1(write1_sel[2]), .A2(write1_sel[1]), .Z(n164) );
  MOAI22D0BWP12T U163 ( .A1(n2864), .A2(n1412), .B1(n2807), .B2(n[2951]), .ZN(
        n446) );
  AO22D1BWP12T U164 ( .A1(write2_in[22]), .A2(n2916), .B1(n2920), .B2(
        write1_in[22]), .Z(n1748) );
  INR2D0BWP12T U165 ( .A1(pc_out[28]), .B1(n2924), .ZN(n1737) );
  INR2D0BWP12T U166 ( .A1(n165), .B1(n166), .ZN(n1608) );
  INR3D0BWP12T U167 ( .A1(n158), .B1(n159), .B2(reset), .ZN(n1514) );
  INR2D0BWP12T U168 ( .A1(n167), .B1(n168), .ZN(n1518) );
  INR2D0BWP12T U169 ( .A1(n179), .B1(n180), .ZN(n1517) );
  OAI22D0BWP12T U170 ( .A1(write1_in[0]), .A2(n2916), .B1(n583), .B2(n2920), 
        .ZN(n16) );
  AOI22D0BWP12T U171 ( .A1(pc_out[0]), .A2(n1690), .B1(next_pc_in[0]), .B2(
        n1488), .ZN(n17) );
  OAI21D0BWP12T U172 ( .A1(n2919), .A2(n16), .B(n17), .ZN(n2169) );
  MAOI22D0BWP12T U173 ( .A1(n1415), .A2(n1414), .B1(n1415), .B2(n1414), .ZN(
        n18) );
  AO222D0BWP12T U174 ( .A1(n2914), .A2(n18), .B1(pc_out[6]), .B2(n1690), .C1(
        next_pc_in[6]), .C2(n1488), .Z(n2175) );
  MAOI22D1BWP12T U175 ( .A1(n1613), .A2(n1612), .B1(n1613), .B2(n1612), .ZN(
        n19) );
  AO222D1BWP12T U176 ( .A1(pc_out[18]), .A2(n1690), .B1(n19), .B2(n2914), .C1(
        next_pc_in[18]), .C2(n1488), .Z(n2187) );
  MAOI22D0BWP12T U177 ( .A1(n2813), .A2(r12[9]), .B1(n2884), .B2(n546), .ZN(
        n72) );
  IND2D0BWP12T U178 ( .A1(write1_sel[3]), .B1(n141), .ZN(n146) );
  MAOI22D0BWP12T U179 ( .A1(n2891), .A2(lr[2]), .B1(n2822), .B2(n1873), .ZN(
        n1880) );
  CKND0BWP12T U180 ( .I(r6[15]), .ZN(n20) );
  MOAI22D0BWP12T U181 ( .A1(n2826), .A2(n20), .B1(n2893), .B2(r10[15]), .ZN(
        n591) );
  MAOI22D0BWP12T U182 ( .A1(n2791), .A2(r4[7]), .B1(n2884), .B2(n617), .ZN(
        n626) );
  NR2D0BWP12T U183 ( .A1(write2_sel[0]), .A2(n300), .ZN(n21) );
  ND4D0BWP12T U184 ( .A1(write2_en), .A2(write2_sel[4]), .A3(write2_sel[3]), 
        .A4(n21), .ZN(n301) );
  INR2D0BWP12T U185 ( .A1(n287), .B1(reset), .ZN(n285) );
  IND2D0BWP12T U186 ( .A1(n1636), .B1(n1749), .ZN(n1638) );
  CKND0BWP12T U187 ( .I(pc_out[29]), .ZN(n22) );
  MOAI22D0BWP12T U188 ( .A1(n2924), .A2(n22), .B1(n1488), .B2(next_pc_in[29]), 
        .ZN(n1682) );
  IOA21D0BWP12T U189 ( .A1(n1663), .A2(n1664), .B(n2912), .ZN(n1667) );
  IND2D0BWP12T U190 ( .A1(n153), .B1(n152), .ZN(n1615) );
  MAOI22D0BWP12T U191 ( .A1(n434), .A2(n570), .B1(n434), .B2(n570), .ZN(n23)
         );
  AO222D0BWP12T U192 ( .A1(n23), .A2(n2914), .B1(n1690), .B2(pc_out[2]), .C1(
        next_pc_in[2]), .C2(n1488), .Z(n2171) );
  MAOI22D0BWP12T U193 ( .A1(n1409), .A2(n1410), .B1(n1409), .B2(n1410), .ZN(
        n24) );
  AO222D0BWP12T U194 ( .A1(n1690), .A2(pc_out[5]), .B1(n1488), .B2(
        next_pc_in[5]), .C1(n2914), .C2(n24), .Z(n2174) );
  MAOI22D0BWP12T U195 ( .A1(n1427), .A2(n1425), .B1(n1427), .B2(n1425), .ZN(
        n25) );
  AO222D0BWP12T U196 ( .A1(n2914), .A2(n25), .B1(pc_out[8]), .B2(n1690), .C1(
        next_pc_in[8]), .C2(n1488), .Z(n2177) );
  MAOI22D0BWP12T U197 ( .A1(n1467), .A2(n1465), .B1(n1467), .B2(n1465), .ZN(
        n26) );
  AO222D0BWP12T U198 ( .A1(pc_out[11]), .A2(n1690), .B1(n26), .B2(n2914), .C1(
        next_pc_in[11]), .C2(n1488), .Z(n2180) );
  NR2D0BWP12T U199 ( .A1(n1541), .A2(n1540), .ZN(n27) );
  MUX2ND0BWP12T U200 ( .I0(write2_in[20]), .I1(write1_in[20]), .S(n2920), .ZN(
        n28) );
  MAOI22D0BWP12T U201 ( .A1(n27), .A2(n28), .B1(n27), .B2(n28), .ZN(n29) );
  AOI22D0BWP12T U202 ( .A1(pc_out[20]), .A2(n1690), .B1(n1488), .B2(
        next_pc_in[20]), .ZN(n30) );
  OAI21D0BWP12T U203 ( .A1(n2919), .A2(n29), .B(n30), .ZN(n2189) );
  AOI22D0BWP12T U204 ( .A1(r9[30]), .A2(n1321), .B1(r10[30]), .B2(n1322), .ZN(
        n31) );
  AOI22D0BWP12T U205 ( .A1(n[2938]), .A2(n1168), .B1(lr[30]), .B2(n1319), .ZN(
        n32) );
  AOI22D0BWP12T U206 ( .A1(r4[30]), .A2(n1275), .B1(r7[30]), .B2(n1276), .ZN(
        n33) );
  AOI22D0BWP12T U207 ( .A1(r6[30]), .A2(n1277), .B1(r2[30]), .B2(n1278), .ZN(
        n34) );
  AOI22D0BWP12T U208 ( .A1(r1[30]), .A2(n1279), .B1(r5[30]), .B2(n1280), .ZN(
        n35) );
  AOI22D0BWP12T U209 ( .A1(r0[30]), .A2(n1282), .B1(r3[30]), .B2(n1281), .ZN(
        n36) );
  ND4D0BWP12T U210 ( .A1(n33), .A2(n34), .A3(n35), .A4(n36), .ZN(n37) );
  MOAI22D0BWP12T U211 ( .A1(n2923), .A2(n1268), .B1(r8[30]), .B2(n1323), .ZN(
        n38) );
  CKND0BWP12T U212 ( .I(r12[30]), .ZN(n39) );
  CKND0BWP12T U213 ( .I(r11[30]), .ZN(n40) );
  OAI22D0BWP12T U214 ( .A1(n1238), .A2(n39), .B1(n1287), .B2(n40), .ZN(n41) );
  AOI211D0BWP12T U215 ( .A1(n1295), .A2(n37), .B(n38), .C(n41), .ZN(n42) );
  ND3D0BWP12T U216 ( .A1(n31), .A2(n32), .A3(n42), .ZN(regC_out[30]) );
  MAOI22D0BWP12T U217 ( .A1(n2809), .A2(r5[2]), .B1(n2860), .B2(n1884), .ZN(
        n1887) );
  MAOI22D0BWP12T U218 ( .A1(n2893), .A2(r10[11]), .B1(n2826), .B2(n1934), .ZN(
        n794) );
  MOAI22D0BWP12T U219 ( .A1(n2826), .A2(n1874), .B1(n2893), .B2(r10[2]), .ZN(
        n1879) );
  OA22D0BWP12T U220 ( .A1(n2867), .A2(n2019), .B1(n2864), .B2(n1852), .Z(n1861) );
  MOAI22D0BWP12T U221 ( .A1(n2864), .A2(n839), .B1(n2807), .B2(n[2967]), .ZN(
        n847) );
  MAOI22D0BWP12T U222 ( .A1(n2891), .A2(lr[15]), .B1(n1943), .B2(n1055), .ZN(
        n592) );
  AOI33D0BWP12T U223 ( .A1(n348), .A2(n854), .A3(r1[9]), .B1(n363), .B2(n81), 
        .B3(r10[9]), .ZN(n43) );
  IOA21D0BWP12T U224 ( .A1(n2894), .A2(r6[9]), .B(n43), .ZN(n78) );
  MAOI22D0BWP12T U225 ( .A1(n2791), .A2(r4[17]), .B1(n2884), .B2(n448), .ZN(
        n457) );
  IND2D0BWP12T U226 ( .A1(n1534), .B1(n1535), .ZN(n1543) );
  CKND0BWP12T U227 ( .I(pc_out[31]), .ZN(n44) );
  MOAI22D0BWP12T U228 ( .A1(n2924), .A2(n44), .B1(next_pc_in[31]), .B2(n1488), 
        .ZN(n1669) );
  INR2D0BWP12T U229 ( .A1(n177), .B1(n178), .ZN(n1598) );
  INR2D0BWP12T U230 ( .A1(n189), .B1(n190), .ZN(n1519) );
  INR2D0BWP12T U231 ( .A1(n149), .B1(n150), .ZN(n1576) );
  INR2D0BWP12T U232 ( .A1(n173), .B1(n174), .ZN(n1506) );
  NR2D0BWP12T U233 ( .A1(n1427), .A2(n1425), .ZN(n45) );
  MOAI22D0BWP12T U234 ( .A1(n45), .A2(n1426), .B1(n45), .B2(n1426), .ZN(n46)
         );
  AO222D0BWP12T U235 ( .A1(n46), .A2(n2914), .B1(next_pc_in[9]), .B2(n1488), 
        .C1(pc_out[9]), .C2(n1690), .Z(n2178) );
  NR2D0BWP12T U236 ( .A1(n1467), .A2(n1465), .ZN(n47) );
  MOAI22D0BWP12T U237 ( .A1(n47), .A2(n1466), .B1(n47), .B2(n1466), .ZN(n48)
         );
  AO222D0BWP12T U238 ( .A1(n48), .A2(n2914), .B1(pc_out[12]), .B2(n1690), .C1(
        next_pc_in[12]), .C2(n1488), .Z(n2181) );
  MAOI22D0BWP12T U239 ( .A1(n1656), .A2(n1630), .B1(n1656), .B2(n1630), .ZN(
        n49) );
  AOI22D0BWP12T U240 ( .A1(pc_out[21]), .A2(n1690), .B1(n1488), .B2(
        next_pc_in[21]), .ZN(n50) );
  OAI21D0BWP12T U241 ( .A1(n49), .A2(n2919), .B(n50), .ZN(n2190) );
  AOI22D0BWP12T U242 ( .A1(r8[7]), .A2(n1382), .B1(r4[7]), .B2(n1381), .ZN(n51) );
  AOI22D0BWP12T U243 ( .A1(r10[7]), .A2(n1383), .B1(n[2961]), .B2(n1384), .ZN(
        n52) );
  AOI22D0BWP12T U244 ( .A1(r3[7]), .A2(n1399), .B1(r2[7]), .B2(n1398), .ZN(n53) );
  AOI22D0BWP12T U245 ( .A1(pc_out[7]), .A2(n1400), .B1(r0[7]), .B2(n1401), 
        .ZN(n54) );
  OAI211D0BWP12T U246 ( .A1(n768), .A2(n1404), .B(n53), .C(n54), .ZN(n55) );
  AOI22D0BWP12T U247 ( .A1(r9[7]), .A2(n1389), .B1(lr[7]), .B2(n1390), .ZN(n56) );
  AOI22D0BWP12T U248 ( .A1(r7[7]), .A2(n1388), .B1(r5[7]), .B2(n1387), .ZN(n57) );
  AOI22D0BWP12T U249 ( .A1(r6[7]), .A2(n1392), .B1(r11[7]), .B2(n1391), .ZN(
        n58) );
  ND3D0BWP12T U250 ( .A1(n56), .A2(n57), .A3(n58), .ZN(n59) );
  AOI211D0BWP12T U251 ( .A1(r12[7]), .A2(n1393), .B(n55), .C(n59), .ZN(n60) );
  CKND0BWP12T U252 ( .I(n1405), .ZN(n61) );
  AOI31D0BWP12T U253 ( .A1(n51), .A2(n52), .A3(n60), .B(n61), .ZN(regD_out[7])
         );
  TPNR2D1BWP12T U254 ( .A1(n1739), .A2(n2919), .ZN(n1718) );
  CKND2D2BWP12T U255 ( .A1(n1705), .A2(n1704), .ZN(n1739) );
  TPND2D2BWP12T U256 ( .A1(n1663), .A2(n1664), .ZN(n2911) );
  CKND2D2BWP12T U257 ( .A1(n98), .A2(n97), .ZN(regA_out[9]) );
  TPNR3D1BWP12T U258 ( .A1(n79), .A2(n78), .A3(n77), .ZN(n98) );
  TPAOI21D1BWP12T U259 ( .A1(write1_in[11]), .A2(n2920), .B(n1434), .ZN(n1465)
         );
  TPND2D1BWP12T U260 ( .A1(n1703), .A2(n1702), .ZN(n1720) );
  ND4D1BWP12T U261 ( .A1(n888), .A2(n887), .A3(n886), .A4(n885), .ZN(
        regA_out[3]) );
  TPOAI22D1BWP12T U262 ( .A1(n2693), .A2(n1140), .B1(n2691), .B2(n858), .ZN(
        n135) );
  OAI21D1BWP12T U263 ( .A1(write1_in[30]), .A2(n2916), .B(n1644), .ZN(n1658)
         );
  INVD4BWP12T U264 ( .I(n118), .ZN(n2680) );
  NR3XD3BWP12T U265 ( .A1(n1494), .A2(n1493), .A3(n1492), .ZN(n1535) );
  ND3XD4BWP12T U266 ( .A1(n120), .A2(n100), .A3(readB_sel[3]), .ZN(n125) );
  INVD3BWP12T U267 ( .I(readB_sel[0]), .ZN(n100) );
  NR2XD3BWP12T U268 ( .A1(n1631), .A2(n1630), .ZN(n1749) );
  NR3XD3BWP12T U269 ( .A1(n1541), .A2(n1540), .A3(n1539), .ZN(n1656) );
  ND2XD4BWP12T U270 ( .A1(n1535), .A2(n1545), .ZN(n1540) );
  INVD6BWP12T U271 ( .I(n2684), .ZN(n2763) );
  ND2D3BWP12T U272 ( .A1(n124), .A2(n123), .ZN(n2684) );
  NR2D2BWP12T U273 ( .A1(n122), .A2(n121), .ZN(n123) );
  CKND2D2BWP12T U274 ( .A1(n2003), .A2(n2002), .ZN(regA_out[18]) );
  TPND2D1BWP12T U275 ( .A1(n901), .A2(n900), .ZN(regB_out[19]) );
  ND2D3BWP12T U276 ( .A1(n413), .A2(n412), .ZN(regA_out[14]) );
  INR2XD2BWP12T U277 ( .A1(n126), .B1(n130), .ZN(n105) );
  ND4D2BWP12T U278 ( .A1(n496), .A2(n495), .A3(n494), .A4(n493), .ZN(
        regB_out[31]) );
  ND4D3BWP12T U279 ( .A1(n823), .A2(n822), .A3(n821), .A4(n820), .ZN(
        regA_out[30]) );
  ND4D2BWP12T U280 ( .A1(n380), .A2(n379), .A3(n378), .A4(n377), .ZN(
        regB_out[29]) );
  INVD1BWP12T U281 ( .I(n2919), .ZN(n2914) );
  ND2D1BWP12T U282 ( .A1(n569), .A2(n902), .ZN(n2919) );
  INR2XD2BWP12T U283 ( .A1(n126), .B1(n117), .ZN(n118) );
  ND2D4BWP12T U284 ( .A1(n735), .A2(n734), .ZN(regA_out[13]) );
  INVD2BWP12T U285 ( .I(readB_sel[3]), .ZN(n119) );
  OR2XD1BWP12T U286 ( .A1(n2880), .A2(n867), .Z(n62) );
  CKND0BWP12T U287 ( .I(readB_sel[0]), .ZN(n121) );
  INR2D1BWP12T U288 ( .A1(write2_en), .B1(write2_sel[4]), .ZN(n142) );
  AN2XD1BWP12T U289 ( .A1(write2_sel[0]), .A2(n142), .Z(n148) );
  ND2D1BWP12T U290 ( .A1(n148), .A2(write2_sel[3]), .ZN(n289) );
  ND2D1BWP12T U291 ( .A1(write2_sel[2]), .A2(write2_sel[1]), .ZN(n300) );
  INR2D1BWP12T U292 ( .A1(write1_en), .B1(write1_sel[4]), .ZN(n141) );
  INVD1BWP12T U293 ( .I(write1_sel[0]), .ZN(n155) );
  INR2D1BWP12T U294 ( .A1(n164), .B1(n286), .ZN(n63) );
  INVD2BWP12T U295 ( .I(n63), .ZN(n2916) );
  OAI21D1BWP12T U296 ( .A1(n289), .A2(n300), .B(n2916), .ZN(n569) );
  INVD2BWP12T U297 ( .I(reset), .ZN(n902) );
  INVD3BWP12T U298 ( .I(n2916), .ZN(n2920) );
  CKAN2D1BWP12T U299 ( .A1(write2_in[2]), .A2(n2916), .Z(n433) );
  AN2XD0BWP12T U300 ( .A1(write2_in[1]), .A2(n2916), .Z(n64) );
  TPAOI21D1BWP12T U301 ( .A1(write1_in[1]), .A2(n2920), .B(n64), .ZN(n570) );
  NR2D1BWP12T U302 ( .A1(next_pc_en_BAR), .A2(n65), .ZN(n1488) );
  DCCKND4BWP12T U303 ( .I(readA_sel[3]), .ZN(n66) );
  TPNR3D3BWP12T U304 ( .A1(n66), .A2(readA_sel[0]), .A3(readA_sel[4]), .ZN(n81) );
  INVD3BWP12T U305 ( .I(n81), .ZN(n856) );
  INR2D4BWP12T U306 ( .A1(readA_sel[2]), .B1(readA_sel[1]), .ZN(n86) );
  DCCKND4BWP12T U307 ( .I(n86), .ZN(n396) );
  OR2D4BWP12T U308 ( .A1(n856), .A2(n396), .Z(n2875) );
  CKND4BWP12T U309 ( .I(n2875), .ZN(n2813) );
  TPNR3D8BWP12T U310 ( .A1(readA_sel[3]), .A2(readA_sel[0]), .A3(readA_sel[4]), 
        .ZN(n1853) );
  TPNR2D4BWP12T U311 ( .A1(readA_sel[2]), .A2(readA_sel[1]), .ZN(n854) );
  ND2D4BWP12T U312 ( .A1(n1853), .A2(n854), .ZN(n2884) );
  INVD1BWP12T U313 ( .I(r0[9]), .ZN(n546) );
  INVD3BWP12T U314 ( .I(readA_sel[4]), .ZN(n67) );
  ND3D4BWP12T U315 ( .A1(n67), .A2(readA_sel[3]), .A3(readA_sel[0]), .ZN(n350)
         );
  INR2D2BWP12T U316 ( .A1(n86), .B1(n350), .ZN(n68) );
  CKND3BWP12T U317 ( .I(n68), .ZN(n2867) );
  INVD6BWP12T U318 ( .I(n2867), .ZN(n2807) );
  ND2D1BWP12T U319 ( .A1(n2807), .A2(n[2959]), .ZN(n71) );
  INR2D2BWP12T U320 ( .A1(n854), .B1(n350), .ZN(n69) );
  INVD3BWP12T U321 ( .I(n69), .ZN(n2883) );
  INVD4BWP12T U322 ( .I(n2883), .ZN(n2819) );
  ND2D1BWP12T U323 ( .A1(n2819), .A2(r9[9]), .ZN(n70) );
  ND3D1BWP12T U324 ( .A1(n72), .A2(n71), .A3(n70), .ZN(n79) );
  INR2D4BWP12T U325 ( .A1(readA_sel[1]), .B1(n1856), .ZN(n351) );
  ND2D4BWP12T U326 ( .A1(n1853), .A2(n351), .ZN(n2826) );
  INVD2BWP12T U327 ( .I(n2826), .ZN(n2894) );
  INR2D4BWP12T U328 ( .A1(readA_sel[1]), .B1(readA_sel[2]), .ZN(n363) );
  DCCKND4BWP12T U329 ( .I(readA_sel[0]), .ZN(n73) );
  TPNR3D4BWP12T U330 ( .A1(n73), .A2(readA_sel[3]), .A3(readA_sel[4]), .ZN(
        n348) );
  INR3D2BWP12T U331 ( .A1(readA_sel[4]), .B1(readA_sel[0]), .B2(n1856), .ZN(
        n75) );
  INVD1BWP12T U332 ( .I(readA_sel[1]), .ZN(n1855) );
  INR2D2BWP12T U333 ( .A1(readA_sel[3]), .B1(n1855), .ZN(n74) );
  ND2D4BWP12T U334 ( .A1(n75), .A2(n74), .ZN(n2880) );
  INVD1BWP12T U335 ( .I(tmp1[9]), .ZN(n209) );
  INVD1P75BWP12T U336 ( .I(n350), .ZN(n80) );
  ND3XD0BWP12T U337 ( .A1(n80), .A2(pc_out[9]), .A3(n351), .ZN(n76) );
  OAI21D1BWP12T U338 ( .A1(n2880), .A2(n209), .B(n76), .ZN(n77) );
  ND2XD4BWP12T U339 ( .A1(n80), .A2(n363), .ZN(n2864) );
  INVD1BWP12T U340 ( .I(r11[9]), .ZN(n432) );
  NR2D1BWP12T U341 ( .A1(n2864), .A2(n432), .ZN(n84) );
  TPND2D2BWP12T U342 ( .A1(n81), .A2(n854), .ZN(n82) );
  INVD2BWP12T U343 ( .I(n82), .ZN(n584) );
  INVD4BWP12T U344 ( .I(n584), .ZN(n2822) );
  INVD1BWP12T U345 ( .I(r8[9]), .ZN(n1034) );
  NR2D1BWP12T U346 ( .A1(n2822), .A2(n1034), .ZN(n83) );
  NR2D1BWP12T U347 ( .A1(n84), .A2(n83), .ZN(n96) );
  INVD1BWP12T U348 ( .I(r7[9]), .ZN(n542) );
  INVD1P75BWP12T U349 ( .I(n348), .ZN(n85) );
  INR2D2BWP12T U350 ( .A1(n86), .B1(n85), .ZN(n87) );
  INVD4BWP12T U351 ( .I(n87), .ZN(n2863) );
  INVD6BWP12T U352 ( .I(n2863), .ZN(n2809) );
  ND2D1BWP12T U353 ( .A1(n2809), .A2(r5[9]), .ZN(n88) );
  OAI21D1BWP12T U354 ( .A1(n2868), .A2(n542), .B(n88), .ZN(n95) );
  INR2D8BWP12T U355 ( .A1(n1853), .B1(n396), .ZN(n2791) );
  TPND2D4BWP12T U356 ( .A1(n363), .A2(n1853), .ZN(n2789) );
  INVD1BWP12T U357 ( .I(r2[9]), .ZN(n543) );
  INVD1P75BWP12T U358 ( .I(n351), .ZN(n89) );
  TPNR2D4BWP12T U359 ( .A1(n856), .A2(n89), .ZN(n2891) );
  TPND2D2BWP12T U360 ( .A1(n348), .A2(n363), .ZN(n90) );
  INVD2BWP12T U361 ( .I(n90), .ZN(n349) );
  CKND1BWP12T U362 ( .I(n349), .ZN(n593) );
  INVD1BWP12T U363 ( .I(r3[9]), .ZN(n431) );
  NR2D1BWP12T U364 ( .A1(n593), .A2(n431), .ZN(n91) );
  RCAOI21D0BWP12T U365 ( .A1(n2891), .A2(lr[9]), .B(n91), .ZN(n92) );
  ND2D1BWP12T U366 ( .A1(n93), .A2(n92), .ZN(n94) );
  INR3D0BWP12T U367 ( .A1(n96), .B1(n95), .B2(n94), .ZN(n97) );
  INVD1BWP12T U368 ( .I(r5[1]), .ZN(n577) );
  INR2D2BWP12T U369 ( .A1(readB_sel[2]), .B1(readB_sel[1]), .ZN(n128) );
  INVD3BWP12T U370 ( .I(readB_sel[4]), .ZN(n120) );
  AN3XD2BWP12T U371 ( .A1(n119), .A2(n120), .A3(readB_sel[0]), .Z(n99) );
  INVD2BWP12T U372 ( .I(n99), .ZN(n117) );
  INR2XD2BWP12T U373 ( .A1(n128), .B1(n117), .ZN(n2748) );
  INVD3BWP12T U374 ( .I(n2748), .ZN(n2664) );
  INR2D4BWP12T U375 ( .A1(readB_sel[1]), .B1(readB_sel[2]), .ZN(n124) );
  INVD3BWP12T U376 ( .I(n2747), .ZN(n2663) );
  INVD1BWP12T U377 ( .I(r10[1]), .ZN(n573) );
  OAI22D1BWP12T U378 ( .A1(n577), .A2(n2664), .B1(n2663), .B2(n573), .ZN(n116)
         );
  INVD1BWP12T U379 ( .I(tmp1[1]), .ZN(n850) );
  INVD1P75BWP12T U380 ( .I(readB_sel[1]), .ZN(n101) );
  INR2D4BWP12T U381 ( .A1(readB_sel[2]), .B1(n101), .ZN(n131) );
  INR2D1BWP12T U382 ( .A1(readB_sel[4]), .B1(n119), .ZN(n102) );
  ND2D1BWP12T U383 ( .A1(n131), .A2(n102), .ZN(n103) );
  INR2D1BWP12T U384 ( .A1(n121), .B1(n103), .ZN(n225) );
  INR2D1BWP12T U385 ( .A1(readB_sel[0]), .B1(n103), .ZN(n104) );
  INVD4BWP12T U386 ( .I(n309), .ZN(n2730) );
  MOAI22D0BWP12T U387 ( .A1(n850), .A2(n2666), .B1(n2730), .B2(
        immediate2_in[1]), .ZN(n115) );
  ND3D4BWP12T U388 ( .A1(n120), .A2(readB_sel[3]), .A3(readB_sel[0]), .ZN(n130) );
  NR2D1BWP12T U389 ( .A1(readB_sel[3]), .A2(readB_sel[0]), .ZN(n106) );
  CKND2D2BWP12T U390 ( .A1(n106), .A2(n120), .ZN(n133) );
  INVD1BWP12T U391 ( .I(n128), .ZN(n107) );
  TPNR2D1BWP12T U392 ( .A1(n133), .A2(n107), .ZN(n108) );
  BUFFD6BWP12T U393 ( .I(n108), .Z(n2753) );
  INR2D2BWP12T U394 ( .A1(n126), .B1(n133), .ZN(n109) );
  INVD3BWP12T U395 ( .I(n109), .ZN(n210) );
  INVD4BWP12T U396 ( .I(n210), .ZN(n2650) );
  AOI22D1BWP12T U397 ( .A1(r11[1]), .A2(n2755), .B1(n2650), .B2(r0[1]), .ZN(
        n110) );
  ND2D1BWP12T U398 ( .A1(n111), .A2(n110), .ZN(n114) );
  INR2XD2BWP12T U399 ( .A1(n131), .B1(n117), .ZN(n2750) );
  INVD3BWP12T U400 ( .I(n2750), .ZN(n2673) );
  INVD1BWP12T U401 ( .I(r7[1]), .ZN(n837) );
  INVD1BWP12T U402 ( .I(n124), .ZN(n112) );
  TPNR2D3BWP12T U403 ( .A1(n133), .A2(n112), .ZN(n2749) );
  INVD1BWP12T U404 ( .I(r2[1]), .ZN(n574) );
  OAI22D1BWP12T U405 ( .A1(n2673), .A2(n837), .B1(n2671), .B2(n574), .ZN(n113)
         );
  NR4D0BWP12T U406 ( .A1(n116), .A2(n115), .A3(n114), .A4(n113), .ZN(n140) );
  INVD1BWP12T U407 ( .I(r1[1]), .ZN(n842) );
  INR2XD2BWP12T U408 ( .A1(n128), .B1(n125), .ZN(n2761) );
  INVD1BWP12T U409 ( .I(r12[1]), .ZN(n1139) );
  INVD1BWP12T U410 ( .I(r3[1]), .ZN(n840) );
  CKND2D1BWP12T U411 ( .A1(n120), .A2(n119), .ZN(n122) );
  INR2D4BWP12T U412 ( .A1(n131), .B1(n125), .ZN(n2762) );
  INVD3BWP12T U413 ( .I(n2762), .ZN(n2683) );
  INVD1BWP12T U414 ( .I(lr[1]), .ZN(n1138) );
  OAI22D1BWP12T U415 ( .A1(n840), .A2(n2684), .B1(n2683), .B2(n1138), .ZN(n137) );
  INR2D1BWP12T U416 ( .A1(n126), .B1(n125), .ZN(n127) );
  BUFFD3BWP12T U417 ( .I(n127), .Z(n2765) );
  INVD2BWP12T U418 ( .I(n2765), .ZN(n2689) );
  INVD1BWP12T U419 ( .I(r8[1]), .ZN(n1137) );
  INVD3BWP12T U420 ( .I(n2764), .ZN(n2687) );
  INVD1BWP12T U421 ( .I(n[2967]), .ZN(n129) );
  OAI22D1BWP12T U422 ( .A1(n2689), .A2(n1137), .B1(n2687), .B2(n129), .ZN(n136) );
  INR2D4BWP12T U423 ( .A1(n131), .B1(n130), .ZN(n2767) );
  INVD3BWP12T U424 ( .I(n2767), .ZN(n2693) );
  INVD1BWP12T U425 ( .I(pc_out[1]), .ZN(n1140) );
  INVD1BWP12T U426 ( .I(n131), .ZN(n132) );
  TPNR2D1BWP12T U427 ( .A1(n133), .A2(n132), .ZN(n134) );
  BUFFXD4BWP12T U428 ( .I(n134), .Z(n2766) );
  INVD4BWP12T U429 ( .I(n2766), .ZN(n2691) );
  INVD1BWP12T U430 ( .I(r6[1]), .ZN(n858) );
  NR4D0BWP12T U431 ( .A1(n138), .A2(n137), .A3(n136), .A4(n135), .ZN(n139) );
  TPND2D1BWP12T U432 ( .A1(n140), .A2(n139), .ZN(regB_out[1]) );
  INR2D1BWP12T U433 ( .A1(n155), .B1(n146), .ZN(n187) );
  INR2D1BWP12T U434 ( .A1(write1_sel[1]), .B1(write1_sel[2]), .ZN(n287) );
  INR2D1BWP12T U435 ( .A1(n142), .B1(write2_sel[0]), .ZN(n156) );
  INVD1BWP12T U436 ( .I(write2_sel[3]), .ZN(n147) );
  ND2D1BWP12T U437 ( .A1(n156), .A2(n147), .ZN(n188) );
  INVD1BWP12T U438 ( .I(n188), .ZN(n172) );
  INVD1BWP12T U439 ( .I(write2_sel[1]), .ZN(n290) );
  NR3D1BWP12T U440 ( .A1(n290), .A2(reset), .A3(write2_sel[2]), .ZN(n157) );
  CKND2D1BWP12T U441 ( .A1(n172), .A2(n157), .ZN(n144) );
  TPND2D0BWP12T U442 ( .A1(n187), .A2(n287), .ZN(n143) );
  INVD1BWP12T U443 ( .I(n1524), .ZN(n1513) );
  AOI22D0BWP12T U444 ( .A1(write2_in[30]), .A2(n1513), .B1(n1511), .B2(r2[30]), 
        .ZN(n145) );
  TPOAI21D0BWP12T U445 ( .A1(n1491), .A2(n1523), .B(n145), .ZN(n2583) );
  INR2D1BWP12T U446 ( .A1(write1_sel[0]), .B1(n146), .ZN(n182) );
  CKND2D1BWP12T U447 ( .A1(n182), .A2(n285), .ZN(n1457) );
  AN2XD1BWP12T U448 ( .A1(n148), .A2(n147), .Z(n184) );
  CKND2D1BWP12T U449 ( .A1(n184), .A2(n157), .ZN(n150) );
  TPND2D0BWP12T U450 ( .A1(n182), .A2(n287), .ZN(n149) );
  AOI22D0BWP12T U451 ( .A1(write2_in[29]), .A2(n1576), .B1(r3[29]), .B2(n1504), 
        .ZN(n151) );
  TPOAI21D0BWP12T U452 ( .A1(n1482), .A2(n1457), .B(n151), .ZN(n2550) );
  INVD1BWP12T U453 ( .I(n1614), .ZN(n1442) );
  INVD1BWP12T U454 ( .I(n289), .ZN(n292) );
  INR2D1BWP12T U455 ( .A1(write2_sel[2]), .B1(write2_sel[1]), .ZN(n183) );
  CKND2D1BWP12T U456 ( .A1(n292), .A2(n183), .ZN(n152) );
  ND2D1BWP12T U457 ( .A1(n1442), .A2(n902), .ZN(n153) );
  AOI22D0BWP12T U458 ( .A1(write2_in[29]), .A2(n1617), .B1(n[2939]), .B2(n1521), .ZN(n154) );
  TPOAI21D0BWP12T U459 ( .A1(n1482), .A2(n1442), .B(n154), .ZN(spin[29]) );
  ND3D1BWP12T U460 ( .A1(write1_sel[3]), .A2(write1_en), .A3(n155), .ZN(n298)
         );
  ND2D1BWP12T U461 ( .A1(n156), .A2(write2_sel[3]), .ZN(n161) );
  INVD1BWP12T U462 ( .I(n157), .ZN(n288) );
  NR2D1BWP12T U463 ( .A1(n161), .A2(n288), .ZN(n159) );
  TPND2D0BWP12T U464 ( .A1(n287), .A2(n175), .ZN(n158) );
  ND2D1BWP12T U465 ( .A1(n159), .A2(n158), .ZN(n1528) );
  INVD1BWP12T U466 ( .I(n1528), .ZN(n1516) );
  AOI22D0BWP12T U467 ( .A1(write2_in[30]), .A2(n1516), .B1(n1514), .B2(r10[30]), .ZN(n160) );
  TPOAI21D0BWP12T U468 ( .A1(n1491), .A2(n1527), .B(n160), .ZN(n2327) );
  INVD1BWP12T U469 ( .I(n161), .ZN(n176) );
  NR2D1BWP12T U470 ( .A1(write2_sel[2]), .A2(write2_sel[1]), .ZN(n192) );
  CKND2D1BWP12T U471 ( .A1(n176), .A2(n192), .ZN(n162) );
  ND2D1BWP12T U472 ( .A1(n1478), .A2(n902), .ZN(n163) );
  INVD1BWP12T U473 ( .I(n1604), .ZN(n1441) );
  INVD1BWP12T U474 ( .I(write2_in[20]), .ZN(n1537) );
  INVD1BWP12T U475 ( .I(n1603), .ZN(n1440) );
  INVD1BWP12T U476 ( .I(r8[20]), .ZN(n2072) );
  OAI222D0BWP12T U477 ( .A1(n1423), .A2(n1478), .B1(n1441), .B2(n1537), .C1(
        n1440), .C2(n2072), .ZN(n2381) );
  INVD1BWP12T U478 ( .I(n1576), .ZN(n1458) );
  INVD1BWP12T U479 ( .I(n1504), .ZN(n1574) );
  INVD1BWP12T U480 ( .I(r3[20]), .ZN(n2070) );
  OAI222D0BWP12T U481 ( .A1(n1423), .A2(n1457), .B1(n1458), .B2(n1537), .C1(
        n1574), .C2(n2070), .ZN(n2541) );
  ND2D1BWP12T U482 ( .A1(n164), .A2(n902), .ZN(n299) );
  INVD1BWP12T U483 ( .I(n300), .ZN(n169) );
  ND2D1BWP12T U484 ( .A1(n176), .A2(n169), .ZN(n165) );
  ND2D1BWP12T U485 ( .A1(n1475), .A2(n902), .ZN(n166) );
  INVD1BWP12T U486 ( .I(n1609), .ZN(n1439) );
  INVD1BWP12T U487 ( .I(n1608), .ZN(n1438) );
  INVD1BWP12T U488 ( .I(lr[20]), .ZN(n2069) );
  OAI222D0BWP12T U489 ( .A1(n1423), .A2(n1475), .B1(n1439), .B2(n1537), .C1(
        n1438), .C2(n2069), .ZN(n2221) );
  CKND2D1BWP12T U490 ( .A1(n187), .A2(n181), .ZN(n1449) );
  CKND2D1BWP12T U491 ( .A1(n172), .A2(n183), .ZN(n167) );
  ND2D1BWP12T U492 ( .A1(n1449), .A2(n902), .ZN(n168) );
  INVD1BWP12T U493 ( .I(n1582), .ZN(n1450) );
  INVD1BWP12T U494 ( .I(n1518), .ZN(n1580) );
  INVD1BWP12T U495 ( .I(r4[20]), .ZN(n1979) );
  OAI222D0BWP12T U496 ( .A1(n1423), .A2(n1449), .B1(n1450), .B2(n1537), .C1(
        n1580), .C2(n1979), .ZN(n2509) );
  ND2D1BWP12T U497 ( .A1(n184), .A2(n169), .ZN(n170) );
  ND2D1BWP12T U498 ( .A1(n1451), .A2(n902), .ZN(n171) );
  INVD1BWP12T U499 ( .I(n1570), .ZN(n1452) );
  INVD1BWP12T U500 ( .I(n1505), .ZN(n1568) );
  INVD1BWP12T U501 ( .I(r7[20]), .ZN(n2062) );
  OAI222D0BWP12T U502 ( .A1(n1423), .A2(n1451), .B1(n1452), .B2(n1537), .C1(
        n1568), .C2(n2062), .ZN(n2413) );
  ND2D1BWP12T U503 ( .A1(n187), .A2(n191), .ZN(n1454) );
  CKND2D1BWP12T U504 ( .A1(n172), .A2(n192), .ZN(n173) );
  ND2D1BWP12T U505 ( .A1(n1454), .A2(n902), .ZN(n174) );
  INVD1BWP12T U506 ( .I(n1552), .ZN(n1455) );
  INVD1BWP12T U507 ( .I(n1506), .ZN(n1550) );
  INVD1BWP12T U508 ( .I(r0[20]), .ZN(n1978) );
  OAI222D0BWP12T U509 ( .A1(n1423), .A2(n1454), .B1(n1455), .B2(n1537), .C1(
        n1550), .C2(n1978), .ZN(n2637) );
  ND2D1BWP12T U510 ( .A1(n181), .A2(n175), .ZN(n1436) );
  ND2D1BWP12T U511 ( .A1(n176), .A2(n183), .ZN(n177) );
  ND2D1BWP12T U512 ( .A1(n1436), .A2(n902), .ZN(n178) );
  INVD1BWP12T U513 ( .I(n1599), .ZN(n1437) );
  INVD1BWP12T U514 ( .I(n1598), .ZN(n1435) );
  INVD1BWP12T U515 ( .I(r12[20]), .ZN(n2067) );
  OAI222D0BWP12T U516 ( .A1(n1423), .A2(n1436), .B1(n1437), .B2(n1537), .C1(
        n1435), .C2(n2067), .ZN(n2253) );
  ND2D1BWP12T U517 ( .A1(n182), .A2(n191), .ZN(n1447) );
  CKND2D1BWP12T U518 ( .A1(n184), .A2(n192), .ZN(n179) );
  ND2D1BWP12T U519 ( .A1(n1447), .A2(n902), .ZN(n180) );
  INVD1BWP12T U520 ( .I(n1588), .ZN(n1448) );
  INVD1BWP12T U521 ( .I(n1517), .ZN(n1586) );
  INVD1BWP12T U522 ( .I(r1[20]), .ZN(n2068) );
  OAI222D0BWP12T U523 ( .A1(n1423), .A2(n1447), .B1(n1448), .B2(n1537), .C1(
        n1586), .C2(n2068), .ZN(n2605) );
  CKND2D1BWP12T U524 ( .A1(n182), .A2(n181), .ZN(n1445) );
  CKND2D1BWP12T U525 ( .A1(n184), .A2(n183), .ZN(n185) );
  ND2D1BWP12T U526 ( .A1(n1445), .A2(n902), .ZN(n186) );
  INVD1BWP12T U527 ( .I(n1564), .ZN(n1446) );
  INVD1BWP12T U528 ( .I(n1520), .ZN(n1562) );
  INVD1BWP12T U529 ( .I(r5[20]), .ZN(n2057) );
  OAI222D0BWP12T U530 ( .A1(n1423), .A2(n1445), .B1(n1446), .B2(n1537), .C1(
        n1562), .C2(n2057), .ZN(n2477) );
  NR2D1BWP12T U531 ( .A1(n188), .A2(n300), .ZN(n190) );
  NR2D1BWP12T U532 ( .A1(n1555), .A2(reset), .ZN(n189) );
  ND2D1BWP12T U533 ( .A1(n190), .A2(n189), .ZN(n1444) );
  INVD1BWP12T U534 ( .I(n1519), .ZN(n1556) );
  INVD1BWP12T U535 ( .I(r6[20]), .ZN(n2073) );
  OAI222D0BWP12T U536 ( .A1(n1423), .A2(n1490), .B1(n1444), .B2(n1537), .C1(
        n1556), .C2(n2073), .ZN(n2445) );
  CKND2D1BWP12T U537 ( .A1(n292), .A2(n192), .ZN(n193) );
  ND2D1BWP12T U538 ( .A1(n1481), .A2(n902), .ZN(n194) );
  INVD1BWP12T U539 ( .I(n1594), .ZN(n1453) );
  INVD1BWP12T U540 ( .I(n1507), .ZN(n1592) );
  INVD1BWP12T U541 ( .I(r9[20]), .ZN(n1977) );
  OAI222D0BWP12T U542 ( .A1(n1423), .A2(n1481), .B1(n1453), .B2(n1537), .C1(
        n1592), .C2(n1977), .ZN(n2349) );
  INVD1BWP12T U543 ( .I(write2_in[17]), .ZN(n1418) );
  INVD3BWP12T U544 ( .I(write1_in[17]), .ZN(n1498) );
  INVD1BWP12T U545 ( .I(r5[17]), .ZN(n2665) );
  OAI222D0BWP12T U546 ( .A1(n1446), .A2(n1418), .B1(n1445), .B2(n1498), .C1(
        n1562), .C2(n2665), .ZN(n2474) );
  INVD1BWP12T U547 ( .I(r8[17]), .ZN(n2688) );
  OAI222D0BWP12T U548 ( .A1(n1441), .A2(n1418), .B1(n1478), .B2(n1498), .C1(
        n1440), .C2(n2688), .ZN(n2378) );
  INVD1BWP12T U549 ( .I(r0[17]), .ZN(n448) );
  OAI222D0BWP12T U550 ( .A1(n1455), .A2(n1418), .B1(n1454), .B2(n1498), .C1(
        n1550), .C2(n448), .ZN(n2634) );
  INVD1BWP12T U551 ( .I(r12[17]), .ZN(n2678) );
  OAI222D0BWP12T U552 ( .A1(n1437), .A2(n1418), .B1(n1436), .B2(n1498), .C1(
        n1435), .C2(n2678), .ZN(n2250) );
  INVD1BWP12T U553 ( .I(r7[17]), .ZN(n2672) );
  OAI222D0BWP12T U554 ( .A1(n1452), .A2(n1418), .B1(n1451), .B2(n1498), .C1(
        n1568), .C2(n2672), .ZN(n2410) );
  INVD1BWP12T U555 ( .I(r1[17]), .ZN(n2681) );
  OAI222D0BWP12T U556 ( .A1(n1448), .A2(n1418), .B1(n1447), .B2(n1498), .C1(
        n1586), .C2(n2681), .ZN(n2602) );
  CKND0BWP12T U557 ( .I(r4[17]), .ZN(n195) );
  OAI222D0BWP12T U558 ( .A1(n1450), .A2(n1418), .B1(n1449), .B2(n1498), .C1(
        n1580), .C2(n195), .ZN(n2506) );
  AO222D0BWP12T U559 ( .A1(n1614), .A2(write1_in[15]), .B1(n1521), .B2(n[2953]), .C1(write2_in[15]), .C2(n1617), .Z(spin[15]) );
  INVD1BWP12T U560 ( .I(r5[12]), .ZN(n536) );
  INVD1BWP12T U561 ( .I(r10[12]), .ZN(n429) );
  OAI22D1BWP12T U562 ( .A1(n536), .A2(n2664), .B1(n2663), .B2(n429), .ZN(n201)
         );
  INVD1BWP12T U563 ( .I(tmp1[12]), .ZN(n1947) );
  MOAI22D0BWP12T U564 ( .A1(n1947), .A2(n2666), .B1(n2730), .B2(
        immediate2_in[12]), .ZN(n200) );
  AOI22D1BWP12T U565 ( .A1(r9[12]), .A2(n105), .B1(n2753), .B2(r4[12]), .ZN(
        n197) );
  AOI22D1BWP12T U566 ( .A1(r11[12]), .A2(n2755), .B1(n2754), .B2(r0[12]), .ZN(
        n196) );
  ND2D1BWP12T U567 ( .A1(n197), .A2(n196), .ZN(n199) );
  INVD1BWP12T U568 ( .I(r7[12]), .ZN(n1957) );
  INVD1BWP12T U569 ( .I(r2[12]), .ZN(n428) );
  OAI22D1BWP12T U570 ( .A1(n2673), .A2(n1957), .B1(n2671), .B2(n428), .ZN(n198) );
  NR4D0BWP12T U571 ( .A1(n201), .A2(n200), .A3(n199), .A4(n198), .ZN(n208) );
  INVD1BWP12T U572 ( .I(r1[12]), .ZN(n1963) );
  INVD1BWP12T U573 ( .I(r12[12]), .ZN(n1125) );
  OAI22D1BWP12T U574 ( .A1(n1963), .A2(n2680), .B1(n2679), .B2(n1125), .ZN(
        n206) );
  INVD1BWP12T U575 ( .I(r3[12]), .ZN(n1961) );
  INVD1BWP12T U576 ( .I(lr[12]), .ZN(n530) );
  OAI22D1BWP12T U577 ( .A1(n1961), .A2(n2684), .B1(n2683), .B2(n530), .ZN(n205) );
  INVD1BWP12T U578 ( .I(r8[12]), .ZN(n1942) );
  INVD1BWP12T U579 ( .I(n[2956]), .ZN(n202) );
  OAI22D1BWP12T U580 ( .A1(n2689), .A2(n1942), .B1(n2687), .B2(n202), .ZN(n204) );
  INVD1BWP12T U581 ( .I(pc_out[12]), .ZN(n1126) );
  INVD1BWP12T U582 ( .I(r6[12]), .ZN(n1946) );
  OAI22D1BWP12T U583 ( .A1(n2693), .A2(n1126), .B1(n2691), .B2(n1946), .ZN(
        n203) );
  NR4D0BWP12T U584 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(n207) );
  CKND2D1BWP12T U585 ( .A1(n208), .A2(n207), .ZN(regB_out[12]) );
  CKND1BWP12T U586 ( .I(r5[9]), .ZN(n548) );
  INVD1BWP12T U587 ( .I(r10[9]), .ZN(n545) );
  OAI22D1BWP12T U588 ( .A1(n548), .A2(n2664), .B1(n2663), .B2(n545), .ZN(n216)
         );
  MOAI22D0BWP12T U589 ( .A1(n209), .A2(n2666), .B1(n2730), .B2(
        immediate2_in[9]), .ZN(n215) );
  AOI22D1BWP12T U590 ( .A1(r9[9]), .A2(n105), .B1(n2753), .B2(r4[9]), .ZN(n212) );
  INVD4BWP12T U591 ( .I(n210), .ZN(n2733) );
  AOI22D1BWP12T U592 ( .A1(r11[9]), .A2(n2755), .B1(n2733), .B2(r0[9]), .ZN(
        n211) );
  ND2D1BWP12T U593 ( .A1(n212), .A2(n211), .ZN(n214) );
  OAI22D1BWP12T U594 ( .A1(n2673), .A2(n542), .B1(n2671), .B2(n543), .ZN(n213)
         );
  NR4D0BWP12T U595 ( .A1(n216), .A2(n215), .A3(n214), .A4(n213), .ZN(n224) );
  INVD1BWP12T U596 ( .I(r1[9]), .ZN(n540) );
  INVD1BWP12T U597 ( .I(r12[9]), .ZN(n541) );
  OAI22D1BWP12T U598 ( .A1(n540), .A2(n2680), .B1(n2679), .B2(n541), .ZN(n222)
         );
  INVD1BWP12T U599 ( .I(lr[9]), .ZN(n539) );
  OAI22D1BWP12T U600 ( .A1(n431), .A2(n2684), .B1(n2683), .B2(n539), .ZN(n221)
         );
  INVD1BWP12T U601 ( .I(n[2959]), .ZN(n217) );
  OAI22D1BWP12T U602 ( .A1(n2689), .A2(n1034), .B1(n2687), .B2(n217), .ZN(n220) );
  INVD0BWP12T U603 ( .I(pc_out[9]), .ZN(n218) );
  INVD1BWP12T U604 ( .I(r6[9]), .ZN(n430) );
  OAI22D1BWP12T U605 ( .A1(n2693), .A2(n218), .B1(n2691), .B2(n430), .ZN(n219)
         );
  NR4D0BWP12T U606 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(n223) );
  CKND2D1BWP12T U607 ( .A1(n224), .A2(n223), .ZN(regB_out[9]) );
  BUFFD2BWP12T U608 ( .I(n225), .Z(n2746) );
  AOI22D1BWP12T U609 ( .A1(tmp1[0]), .A2(n2746), .B1(n2135), .B2(
        immediate2_in[0]), .ZN(n232) );
  AOI22D1BWP12T U610 ( .A1(r5[0]), .A2(n2748), .B1(n2747), .B2(r10[0]), .ZN(
        n227) );
  AOI22D1BWP12T U611 ( .A1(r7[0]), .A2(n2750), .B1(n2749), .B2(r2[0]), .ZN(
        n226) );
  ND2D1BWP12T U612 ( .A1(n227), .A2(n226), .ZN(n231) );
  AOI22D1BWP12T U613 ( .A1(r9[0]), .A2(n105), .B1(n2753), .B2(r4[0]), .ZN(n229) );
  AOI22D1BWP12T U614 ( .A1(r11[0]), .A2(n2755), .B1(n2754), .B2(r0[0]), .ZN(
        n228) );
  ND2D1BWP12T U615 ( .A1(n229), .A2(n228), .ZN(n230) );
  INR3XD0BWP12T U616 ( .A1(n232), .B1(n231), .B2(n230), .ZN(n238) );
  AOI22D1BWP12T U617 ( .A1(r1[0]), .A2(n118), .B1(n2761), .B2(r12[0]), .ZN(
        n236) );
  AOI22D1BWP12T U618 ( .A1(r3[0]), .A2(n2763), .B1(n2762), .B2(lr[0]), .ZN(
        n235) );
  AOI22D1BWP12T U619 ( .A1(r8[0]), .A2(n2765), .B1(n2764), .B2(n[2968]), .ZN(
        n234) );
  AOI22D1BWP12T U620 ( .A1(pc_out[0]), .A2(n2767), .B1(n2766), .B2(r6[0]), 
        .ZN(n233) );
  AN4XD1BWP12T U621 ( .A1(n236), .A2(n235), .A3(n234), .A4(n233), .Z(n237) );
  ND2D1BWP12T U622 ( .A1(n238), .A2(n237), .ZN(regB_out[0]) );
  NR2D1BWP12T U623 ( .A1(readD_sel[1]), .A2(readD_sel[0]), .ZN(n252) );
  INVD1BWP12T U624 ( .I(n252), .ZN(n243) );
  IND2D1BWP12T U625 ( .A1(readD_sel[2]), .B1(readD_sel[3]), .ZN(n242) );
  NR2D1BWP12T U626 ( .A1(n243), .A2(n242), .ZN(n1382) );
  IND2D1BWP12T U627 ( .A1(readD_sel[3]), .B1(readD_sel[2]), .ZN(n241) );
  NR2D1BWP12T U628 ( .A1(n243), .A2(n241), .ZN(n1381) );
  AOI22D0BWP12T U629 ( .A1(r8[2]), .A2(n1382), .B1(n1381), .B2(r4[2]), .ZN(
        n240) );
  ND2D1BWP12T U630 ( .A1(readD_sel[3]), .A2(readD_sel[2]), .ZN(n254) );
  IND2D1BWP12T U631 ( .A1(readD_sel[1]), .B1(readD_sel[0]), .ZN(n248) );
  NR2D1BWP12T U632 ( .A1(n254), .A2(n248), .ZN(n1384) );
  IND2D1BWP12T U633 ( .A1(readD_sel[0]), .B1(readD_sel[1]), .ZN(n250) );
  NR2D1BWP12T U634 ( .A1(n242), .A2(n250), .ZN(n1383) );
  AOI22D0BWP12T U635 ( .A1(n[2966]), .A2(n1384), .B1(n1383), .B2(r10[2]), .ZN(
        n239) );
  CKND2D1BWP12T U636 ( .A1(n240), .A2(n239), .ZN(n259) );
  ND2D1BWP12T U637 ( .A1(readD_sel[1]), .A2(readD_sel[0]), .ZN(n253) );
  NR2D1BWP12T U638 ( .A1(n253), .A2(n241), .ZN(n1388) );
  NR2D1BWP12T U639 ( .A1(n248), .A2(n241), .ZN(n1387) );
  AOI22D0BWP12T U640 ( .A1(r7[2]), .A2(n1388), .B1(n1387), .B2(r5[2]), .ZN(
        n247) );
  NR2D1BWP12T U641 ( .A1(n254), .A2(n250), .ZN(n1390) );
  NR2D1BWP12T U642 ( .A1(n242), .A2(n248), .ZN(n1389) );
  AOI22D0BWP12T U643 ( .A1(lr[2]), .A2(n1390), .B1(n1389), .B2(r9[2]), .ZN(
        n246) );
  NR2D1BWP12T U644 ( .A1(n250), .A2(n241), .ZN(n1392) );
  NR2D1BWP12T U645 ( .A1(n242), .A2(n253), .ZN(n1391) );
  AOI22D0BWP12T U646 ( .A1(r6[2]), .A2(n1392), .B1(n1391), .B2(r11[2]), .ZN(
        n245) );
  NR2D1BWP12T U647 ( .A1(n254), .A2(n243), .ZN(n1393) );
  CKND2D0BWP12T U648 ( .A1(n1393), .A2(r12[2]), .ZN(n244) );
  ND4D1BWP12T U649 ( .A1(n247), .A2(n246), .A3(n245), .A4(n244), .ZN(n258) );
  INVD1BWP12T U650 ( .I(r1[2]), .ZN(n1885) );
  NR2D1BWP12T U651 ( .A1(readD_sel[3]), .A2(readD_sel[2]), .ZN(n251) );
  INVD1BWP12T U652 ( .I(n251), .ZN(n249) );
  OR2XD1BWP12T U653 ( .A1(n248), .A2(n249), .Z(n1404) );
  NR2D1BWP12T U654 ( .A1(n253), .A2(n249), .ZN(n1399) );
  NR2D1BWP12T U655 ( .A1(n250), .A2(n249), .ZN(n1398) );
  AOI22D0BWP12T U656 ( .A1(r3[2]), .A2(n1399), .B1(n1398), .B2(r2[2]), .ZN(
        n256) );
  AN2XD1BWP12T U657 ( .A1(n252), .A2(n251), .Z(n1401) );
  NR2D1BWP12T U658 ( .A1(n254), .A2(n253), .ZN(n1400) );
  AOI22D0BWP12T U659 ( .A1(n1401), .A2(r0[2]), .B1(pc_out[2]), .B2(n1400), 
        .ZN(n255) );
  OAI211D0BWP12T U660 ( .A1(n1885), .A2(n1404), .B(n256), .C(n255), .ZN(n257)
         );
  INVD1BWP12T U661 ( .I(readD_sel[4]), .ZN(n1405) );
  OA31D1BWP12T U662 ( .A1(n259), .A2(n258), .A3(n257), .B(n1405), .Z(
        regD_out[2]) );
  AOI22D0BWP12T U663 ( .A1(r8[5]), .A2(n1382), .B1(n1381), .B2(r4[5]), .ZN(
        n261) );
  AOI22D0BWP12T U664 ( .A1(n[2963]), .A2(n1384), .B1(n1383), .B2(r10[5]), .ZN(
        n260) );
  CKND2D1BWP12T U665 ( .A1(n261), .A2(n260), .ZN(n270) );
  AOI22D0BWP12T U666 ( .A1(r7[5]), .A2(n1388), .B1(n1387), .B2(r5[5]), .ZN(
        n265) );
  AOI22D0BWP12T U667 ( .A1(lr[5]), .A2(n1390), .B1(n1389), .B2(r9[5]), .ZN(
        n264) );
  AOI22D0BWP12T U668 ( .A1(r6[5]), .A2(n1392), .B1(n1391), .B2(r11[5]), .ZN(
        n263) );
  CKND2D0BWP12T U669 ( .A1(n1393), .A2(r12[5]), .ZN(n262) );
  ND4D1BWP12T U670 ( .A1(n265), .A2(n264), .A3(n263), .A4(n262), .ZN(n269) );
  INVD1BWP12T U671 ( .I(r1[5]), .ZN(n2114) );
  AOI22D0BWP12T U672 ( .A1(r3[5]), .A2(n1399), .B1(n1398), .B2(r2[5]), .ZN(
        n267) );
  AOI22D0BWP12T U673 ( .A1(n1401), .A2(r0[5]), .B1(pc_out[5]), .B2(n1400), 
        .ZN(n266) );
  OAI211D0BWP12T U674 ( .A1(n2114), .A2(n1404), .B(n267), .C(n266), .ZN(n268)
         );
  OA31D1BWP12T U675 ( .A1(n270), .A2(n269), .A3(n268), .B(n1405), .Z(
        regD_out[5]) );
  AOI22D0BWP12T U676 ( .A1(r8[4]), .A2(n1382), .B1(n1381), .B2(r4[4]), .ZN(
        n272) );
  AOI22D0BWP12T U677 ( .A1(n[2964]), .A2(n1384), .B1(n1383), .B2(r10[4]), .ZN(
        n271) );
  CKND2D1BWP12T U678 ( .A1(n272), .A2(n271), .ZN(n281) );
  AOI22D0BWP12T U679 ( .A1(r7[4]), .A2(n1388), .B1(n1387), .B2(r5[4]), .ZN(
        n276) );
  AOI22D0BWP12T U680 ( .A1(lr[4]), .A2(n1390), .B1(n1389), .B2(r9[4]), .ZN(
        n275) );
  AOI22D0BWP12T U681 ( .A1(r6[4]), .A2(n1392), .B1(n1391), .B2(r11[4]), .ZN(
        n274) );
  CKND2D0BWP12T U682 ( .A1(n1393), .A2(r12[4]), .ZN(n273) );
  ND4D1BWP12T U683 ( .A1(n276), .A2(n275), .A3(n274), .A4(n273), .ZN(n280) );
  INVD1BWP12T U684 ( .I(r1[4]), .ZN(n2016) );
  AOI22D0BWP12T U685 ( .A1(r3[4]), .A2(n1399), .B1(n1398), .B2(r2[4]), .ZN(
        n278) );
  AOI22D0BWP12T U686 ( .A1(n1401), .A2(r0[4]), .B1(pc_out[4]), .B2(n1400), 
        .ZN(n277) );
  OAI211D0BWP12T U687 ( .A1(n2016), .A2(n1404), .B(n278), .C(n277), .ZN(n279)
         );
  OA31D1BWP12T U688 ( .A1(n281), .A2(n280), .A3(n279), .B(n1405), .Z(
        regD_out[4]) );
  AOI22D0BWP12T U689 ( .A1(write2_in[30]), .A2(n1588), .B1(n1517), .B2(r1[30]), 
        .ZN(n282) );
  TPOAI21D0BWP12T U690 ( .A1(n1491), .A2(n1447), .B(n282), .ZN(n2615) );
  AOI22D0BWP12T U691 ( .A1(write2_in[29]), .A2(n1588), .B1(r1[29]), .B2(n1517), 
        .ZN(n283) );
  TPOAI21D0BWP12T U692 ( .A1(n1482), .A2(n1447), .B(n283), .ZN(n2614) );
  AOI22D0BWP12T U693 ( .A1(write2_in[29]), .A2(n1552), .B1(r0[29]), .B2(n1506), 
        .ZN(n284) );
  TPOAI21D0BWP12T U694 ( .A1(n1482), .A2(n1454), .B(n284), .ZN(n2646) );
  INR2D1BWP12T U695 ( .A1(n287), .B1(n286), .ZN(n291) );
  AOI22D0BWP12T U696 ( .A1(write2_in[30]), .A2(n1510), .B1(n1508), .B2(r11[30]), .ZN(n293) );
  TPOAI21D0BWP12T U697 ( .A1(n1491), .A2(n1532), .B(n293), .ZN(n2295) );
  AOI22D0BWP12T U698 ( .A1(write2_in[29]), .A2(n1570), .B1(r7[29]), .B2(n1505), 
        .ZN(n294) );
  TPOAI21D0BWP12T U699 ( .A1(n1482), .A2(n1451), .B(n294), .ZN(n2422) );
  AOI22D0BWP12T U700 ( .A1(write2_in[30]), .A2(n1609), .B1(n1608), .B2(lr[30]), 
        .ZN(n295) );
  TPOAI21D0BWP12T U701 ( .A1(n1491), .A2(n1475), .B(n295), .ZN(n2231) );
  AOI22D0BWP12T U702 ( .A1(write2_in[30]), .A2(n1594), .B1(n1507), .B2(r9[30]), 
        .ZN(n296) );
  TPOAI21D0BWP12T U703 ( .A1(n1491), .A2(n1481), .B(n296), .ZN(n2359) );
  AOI22D0BWP12T U704 ( .A1(write2_in[30]), .A2(n1576), .B1(n1504), .B2(r3[30]), 
        .ZN(n297) );
  TPOAI21D0BWP12T U705 ( .A1(n1491), .A2(n1457), .B(n297), .ZN(n2551) );
  INVD1BWP12T U706 ( .I(n1620), .ZN(n427) );
  ND2D1BWP12T U707 ( .A1(n427), .A2(n902), .ZN(n303) );
  INVD1BWP12T U708 ( .I(n301), .ZN(n302) );
  AOI22D0BWP12T U709 ( .A1(write2_in[30]), .A2(n1625), .B1(n1622), .B2(
        tmp1[30]), .ZN(n304) );
  TPOAI21D0BWP12T U710 ( .A1(n1491), .A2(n427), .B(n304), .ZN(n2167) );
  AOI22D0BWP12T U711 ( .A1(write2_in[30]), .A2(n1570), .B1(n1505), .B2(r7[30]), 
        .ZN(n305) );
  TPOAI21D0BWP12T U712 ( .A1(n1491), .A2(n1451), .B(n305), .ZN(n2423) );
  AOI22D0BWP12T U713 ( .A1(write2_in[29]), .A2(n1582), .B1(r4[29]), .B2(n1518), 
        .ZN(n306) );
  TPOAI21D0BWP12T U714 ( .A1(n1482), .A2(n1449), .B(n306), .ZN(n2518) );
  AOI22D0BWP12T U715 ( .A1(write2_in[30]), .A2(n1552), .B1(n1506), .B2(r0[30]), 
        .ZN(n307) );
  TPOAI21D0BWP12T U716 ( .A1(n1491), .A2(n1454), .B(n307), .ZN(n2647) );
  AOI22D0BWP12T U717 ( .A1(write2_in[29]), .A2(n1564), .B1(r5[29]), .B2(n1520), 
        .ZN(n308) );
  TPOAI21D0BWP12T U718 ( .A1(n1482), .A2(n1445), .B(n308), .ZN(n2486) );
  INVD1BWP12T U719 ( .I(n[2948]), .ZN(n2071) );
  OAI222D0BWP12T U720 ( .A1(n1423), .A2(n1442), .B1(n1443), .B2(n1537), .C1(
        n1615), .C2(n2071), .ZN(spin[20]) );
  INVD1BWP12T U721 ( .I(n[2951]), .ZN(n2686) );
  OAI222D0BWP12T U722 ( .A1(n1443), .A2(n1418), .B1(n1442), .B2(n1498), .C1(
        n1615), .C2(n2686), .ZN(spin[17]) );
  INVD1BWP12T U723 ( .I(write2_in[12]), .ZN(n1363) );
  OAI222D0BWP12T U724 ( .A1(n1363), .A2(n1458), .B1(n535), .B2(n1457), .C1(
        n1574), .C2(n1961), .ZN(n2533) );
  INVD1BWP12T U725 ( .I(r5[5]), .ZN(n2109) );
  INVD1BWP12T U726 ( .I(r10[5]), .ZN(n2127) );
  OAI22D1BWP12T U727 ( .A1(n2109), .A2(n2664), .B1(n2663), .B2(n2127), .ZN(
        n315) );
  INVD1BWP12T U728 ( .I(tmp1[5]), .ZN(n2120) );
  INVD4BWP12T U729 ( .I(n309), .ZN(n2745) );
  MOAI22D0BWP12T U730 ( .A1(n2120), .A2(n2666), .B1(n2745), .B2(
        immediate2_in[5]), .ZN(n314) );
  AOI22D1BWP12T U731 ( .A1(r9[5]), .A2(n105), .B1(n2753), .B2(r4[5]), .ZN(n311) );
  AOI22D1BWP12T U732 ( .A1(r11[5]), .A2(n2755), .B1(n2650), .B2(r0[5]), .ZN(
        n310) );
  ND2D1BWP12T U733 ( .A1(n311), .A2(n310), .ZN(n313) );
  INVD1BWP12T U734 ( .I(r7[5]), .ZN(n2112) );
  INVD1BWP12T U735 ( .I(r2[5]), .ZN(n553) );
  OAI22D1BWP12T U736 ( .A1(n2673), .A2(n2112), .B1(n2671), .B2(n553), .ZN(n312) );
  NR4D0BWP12T U737 ( .A1(n315), .A2(n314), .A3(n313), .A4(n312), .ZN(n321) );
  INVD1BWP12T U738 ( .I(r12[5]), .ZN(n2115) );
  OAI22D1BWP12T U739 ( .A1(n2114), .A2(n2680), .B1(n2679), .B2(n2115), .ZN(
        n319) );
  INVD1BWP12T U740 ( .I(r3[5]), .ZN(n2108) );
  INVD1BWP12T U741 ( .I(lr[5]), .ZN(n2129) );
  OAI22D1BWP12T U742 ( .A1(n2108), .A2(n2684), .B1(n2683), .B2(n2129), .ZN(
        n318) );
  INVD1BWP12T U743 ( .I(r8[5]), .ZN(n2128) );
  INVD1BWP12T U744 ( .I(n[2963]), .ZN(n2111) );
  OAI22D1BWP12T U745 ( .A1(n2689), .A2(n2128), .B1(n2687), .B2(n2111), .ZN(
        n317) );
  INVD1BWP12T U746 ( .I(pc_out[5]), .ZN(n2113) );
  INVD1BWP12T U747 ( .I(r6[5]), .ZN(n2126) );
  OAI22D1BWP12T U748 ( .A1(n2693), .A2(n2113), .B1(n2691), .B2(n2126), .ZN(
        n316) );
  NR4D0BWP12T U749 ( .A1(n319), .A2(n318), .A3(n317), .A4(n316), .ZN(n320) );
  CKND2D1BWP12T U750 ( .A1(n321), .A2(n320), .ZN(regB_out[5]) );
  INVD1BWP12T U751 ( .I(r5[6]), .ZN(n2082) );
  INVD1BWP12T U752 ( .I(r10[6]), .ZN(n2100) );
  OAI22D1BWP12T U753 ( .A1(n2082), .A2(n2664), .B1(n2663), .B2(n2100), .ZN(
        n327) );
  INVD1BWP12T U754 ( .I(tmp1[6]), .ZN(n2093) );
  MOAI22D0BWP12T U755 ( .A1(n2093), .A2(n2666), .B1(n2135), .B2(
        immediate2_in[6]), .ZN(n326) );
  AOI22D1BWP12T U756 ( .A1(r9[6]), .A2(n105), .B1(n2753), .B2(r4[6]), .ZN(n323) );
  AOI22D1BWP12T U757 ( .A1(r11[6]), .A2(n2755), .B1(n2754), .B2(r0[6]), .ZN(
        n322) );
  ND2D1BWP12T U758 ( .A1(n323), .A2(n322), .ZN(n325) );
  INVD1BWP12T U759 ( .I(r7[6]), .ZN(n2085) );
  INVD1BWP12T U760 ( .I(r2[6]), .ZN(n557) );
  OAI22D1BWP12T U761 ( .A1(n2673), .A2(n2085), .B1(n2671), .B2(n557), .ZN(n324) );
  NR4D0BWP12T U762 ( .A1(n327), .A2(n326), .A3(n325), .A4(n324), .ZN(n333) );
  INVD1BWP12T U763 ( .I(r1[6]), .ZN(n2087) );
  INVD1BWP12T U764 ( .I(r12[6]), .ZN(n2088) );
  OAI22D1BWP12T U765 ( .A1(n2087), .A2(n2680), .B1(n2679), .B2(n2088), .ZN(
        n331) );
  INVD1BWP12T U766 ( .I(r3[6]), .ZN(n2081) );
  INVD1BWP12T U767 ( .I(lr[6]), .ZN(n2102) );
  OAI22D1BWP12T U768 ( .A1(n2081), .A2(n2684), .B1(n2683), .B2(n2102), .ZN(
        n330) );
  INVD1BWP12T U769 ( .I(r8[6]), .ZN(n2101) );
  INVD1BWP12T U770 ( .I(n[2962]), .ZN(n2084) );
  OAI22D1BWP12T U771 ( .A1(n2689), .A2(n2101), .B1(n2687), .B2(n2084), .ZN(
        n329) );
  INVD1BWP12T U772 ( .I(pc_out[6]), .ZN(n2086) );
  INVD1BWP12T U773 ( .I(r6[6]), .ZN(n2099) );
  OAI22D1BWP12T U774 ( .A1(n2693), .A2(n2086), .B1(n2691), .B2(n2099), .ZN(
        n328) );
  NR4D0BWP12T U775 ( .A1(n331), .A2(n330), .A3(n329), .A4(n328), .ZN(n332) );
  CKND2D1BWP12T U776 ( .A1(n333), .A2(n332), .ZN(regB_out[6]) );
  INVD1BWP12T U777 ( .I(r5[8]), .ZN(n564) );
  INVD1BWP12T U778 ( .I(r10[8]), .ZN(n558) );
  OAI22D1BWP12T U779 ( .A1(n564), .A2(n2664), .B1(n2663), .B2(n558), .ZN(n339)
         );
  INVD1BWP12T U780 ( .I(tmp1[8]), .ZN(n2716) );
  MOAI22D0BWP12T U781 ( .A1(n2716), .A2(n2666), .B1(n2135), .B2(
        immediate2_in[8]), .ZN(n338) );
  AOI22D1BWP12T U782 ( .A1(r9[8]), .A2(n105), .B1(n2753), .B2(r4[8]), .ZN(n335) );
  AOI22D1BWP12T U783 ( .A1(r11[8]), .A2(n2755), .B1(n2733), .B2(r0[8]), .ZN(
        n334) );
  ND2D1BWP12T U784 ( .A1(n335), .A2(n334), .ZN(n337) );
  INVD1BWP12T U785 ( .I(r7[8]), .ZN(n2700) );
  INVD1BWP12T U786 ( .I(r2[8]), .ZN(n439) );
  OAI22D1BWP12T U787 ( .A1(n2673), .A2(n2700), .B1(n2671), .B2(n439), .ZN(n336) );
  NR4D0BWP12T U788 ( .A1(n339), .A2(n338), .A3(n337), .A4(n336), .ZN(n347) );
  INVD1BWP12T U789 ( .I(r1[8]), .ZN(n2706) );
  INVD1BWP12T U790 ( .I(r12[8]), .ZN(n1067) );
  OAI22D1BWP12T U791 ( .A1(n2706), .A2(n2680), .B1(n2679), .B2(n1067), .ZN(
        n345) );
  INVD1BWP12T U792 ( .I(r3[8]), .ZN(n2704) );
  INVD1BWP12T U793 ( .I(lr[8]), .ZN(n562) );
  OAI22D1BWP12T U794 ( .A1(n2704), .A2(n2684), .B1(n2683), .B2(n562), .ZN(n344) );
  INVD1BWP12T U795 ( .I(r8[8]), .ZN(n2719) );
  INVD0BWP12T U796 ( .I(n[2960]), .ZN(n340) );
  OAI22D1BWP12T U797 ( .A1(n2689), .A2(n2719), .B1(n2687), .B2(n340), .ZN(n343) );
  INVD1BWP12T U798 ( .I(pc_out[8]), .ZN(n341) );
  INVD1BWP12T U799 ( .I(r6[8]), .ZN(n2721) );
  OAI22D1BWP12T U800 ( .A1(n2693), .A2(n341), .B1(n2691), .B2(n2721), .ZN(n342) );
  NR4D0BWP12T U801 ( .A1(n345), .A2(n344), .A3(n343), .A4(n342), .ZN(n346) );
  CKND2D1BWP12T U802 ( .A1(n347), .A2(n346), .ZN(regB_out[8]) );
  TPND2D3BWP12T U803 ( .A1(n348), .A2(n854), .ZN(n2872) );
  INVD3BWP12T U804 ( .I(n2872), .ZN(n2814) );
  AOI22D1BWP12T U805 ( .A1(n2814), .A2(r1[16]), .B1(n2813), .B2(r12[16]), .ZN(
        n356) );
  CKND4BWP12T U806 ( .I(n349), .ZN(n2860) );
  INVD4BWP12T U807 ( .I(n2860), .ZN(n2810) );
  INVD2BWP12T U808 ( .I(n2868), .ZN(n2812) );
  INR2D2BWP12T U809 ( .A1(n351), .B1(n350), .ZN(n394) );
  INVD2BWP12T U810 ( .I(n394), .ZN(n352) );
  INVD2BWP12T U811 ( .I(n352), .ZN(n2811) );
  AOI22D1BWP12T U812 ( .A1(n2812), .A2(r7[16]), .B1(n2811), .B2(pc_out[16]), 
        .ZN(n354) );
  AOI22D1BWP12T U813 ( .A1(n2808), .A2(r11[16]), .B1(n2807), .B2(n[2952]), 
        .ZN(n353) );
  AN4XD1BWP12T U814 ( .A1(n356), .A2(n355), .A3(n354), .A4(n353), .Z(n369) );
  INVD3BWP12T U815 ( .I(n2789), .ZN(n2890) );
  INVD1BWP12T U816 ( .I(r9[16]), .ZN(n358) );
  INVD1BWP12T U817 ( .I(tmp1[16]), .ZN(n357) );
  OAI22D1BWP12T U818 ( .A1(n2883), .A2(n358), .B1(n357), .B2(n2880), .ZN(n362)
         );
  INVD3BWP12T U819 ( .I(n2791), .ZN(n2887) );
  INVD1BWP12T U820 ( .I(r4[16]), .ZN(n360) );
  INVD1BWP12T U821 ( .I(r0[16]), .ZN(n359) );
  OAI22D1BWP12T U822 ( .A1(n2887), .A2(n360), .B1(n359), .B2(n2884), .ZN(n361)
         );
  RCAOI211D0BWP12T U823 ( .A1(r2[16]), .A2(n2890), .B(n362), .C(n361), .ZN(
        n368) );
  INVD2BWP12T U824 ( .I(n2822), .ZN(n2892) );
  AOI22D1BWP12T U825 ( .A1(n2892), .A2(r8[16]), .B1(n2891), .B2(lr[16]), .ZN(
        n366) );
  INVD1P75BWP12T U826 ( .I(n363), .ZN(n364) );
  TPNR2D4BWP12T U827 ( .A1(n856), .A2(n364), .ZN(n2893) );
  AOI22D1BWP12T U828 ( .A1(r6[16]), .A2(n2894), .B1(n2893), .B2(r10[16]), .ZN(
        n365) );
  AN2XD1BWP12T U829 ( .A1(n366), .A2(n365), .Z(n367) );
  AOI22D1BWP12T U830 ( .A1(r1[29]), .A2(n118), .B1(n2761), .B2(r12[29]), .ZN(
        n373) );
  AOI22D1BWP12T U831 ( .A1(r3[29]), .A2(n2763), .B1(n2762), .B2(lr[29]), .ZN(
        n372) );
  RCAOI22D0BWP12T U832 ( .A1(r8[29]), .A2(n2765), .B1(n2764), .B2(n[2939]), 
        .ZN(n371) );
  AOI22D1BWP12T U833 ( .A1(pc_out[29]), .A2(n2767), .B1(n2766), .B2(r6[29]), 
        .ZN(n370) );
  AN4XD1BWP12T U834 ( .A1(n373), .A2(n372), .A3(n371), .A4(n370), .Z(n380) );
  AOI22D1BWP12T U835 ( .A1(tmp1[29]), .A2(n2746), .B1(n2745), .B2(
        immediate2_in[29]), .ZN(n376) );
  AOI22D1BWP12T U836 ( .A1(r9[29]), .A2(n105), .B1(n2753), .B2(r4[29]), .ZN(
        n375) );
  AOI22D1BWP12T U837 ( .A1(r11[29]), .A2(n2755), .B1(n2754), .B2(r0[29]), .ZN(
        n374) );
  AOI22D1BWP12T U838 ( .A1(r5[29]), .A2(n2748), .B1(n2747), .B2(r10[29]), .ZN(
        n378) );
  AOI22D1BWP12T U839 ( .A1(r7[29]), .A2(n2750), .B1(n2749), .B2(r2[29]), .ZN(
        n377) );
  AOI22D1BWP12T U840 ( .A1(r1[25]), .A2(n118), .B1(n2761), .B2(r12[25]), .ZN(
        n384) );
  AOI22D1BWP12T U841 ( .A1(r3[25]), .A2(n2763), .B1(n2762), .B2(lr[25]), .ZN(
        n383) );
  AOI22D1BWP12T U842 ( .A1(r8[25]), .A2(n2765), .B1(n2764), .B2(n[2943]), .ZN(
        n382) );
  AOI22D1BWP12T U843 ( .A1(pc_out[25]), .A2(n2767), .B1(n2766), .B2(r6[25]), 
        .ZN(n381) );
  AN4XD1BWP12T U844 ( .A1(n384), .A2(n383), .A3(n382), .A4(n381), .Z(n391) );
  AOI22D1BWP12T U845 ( .A1(tmp1[25]), .A2(n2746), .B1(n2745), .B2(
        immediate2_in[25]), .ZN(n387) );
  AOI22D1BWP12T U846 ( .A1(r9[25]), .A2(n105), .B1(n2753), .B2(r4[25]), .ZN(
        n386) );
  AOI22D1BWP12T U847 ( .A1(r11[25]), .A2(n2755), .B1(n2650), .B2(r0[25]), .ZN(
        n385) );
  AN3XD1BWP12T U848 ( .A1(n387), .A2(n386), .A3(n385), .Z(n390) );
  AOI22D1BWP12T U849 ( .A1(r5[25]), .A2(n2748), .B1(n2747), .B2(r10[25]), .ZN(
        n389) );
  AOI22D1BWP12T U850 ( .A1(r7[25]), .A2(n2750), .B1(n2749), .B2(r2[25]), .ZN(
        n388) );
  INVD1BWP12T U851 ( .I(r5[14]), .ZN(n668) );
  INVD1BWP12T U852 ( .I(r3[14]), .ZN(n392) );
  OAI22D1BWP12T U853 ( .A1(n2863), .A2(n668), .B1(n392), .B2(n2860), .ZN(n402)
         );
  INVD1BWP12T U854 ( .I(n[2954]), .ZN(n1253) );
  INVD1BWP12T U855 ( .I(r11[14]), .ZN(n393) );
  OAI22D0BWP12T U856 ( .A1(n2867), .A2(n1253), .B1(n393), .B2(n2864), .ZN(n401) );
  INVD3BWP12T U857 ( .I(n394), .ZN(n2871) );
  INVD0BWP12T U858 ( .I(pc_out[14]), .ZN(n395) );
  INVD1BWP12T U859 ( .I(r7[14]), .ZN(n673) );
  OAI22D1BWP12T U860 ( .A1(n2871), .A2(n395), .B1(n673), .B2(n2868), .ZN(n400)
         );
  OR2D2BWP12T U861 ( .A1(n856), .A2(n396), .Z(n2851) );
  INVD1BWP12T U862 ( .I(r12[14]), .ZN(n398) );
  INVD1BWP12T U863 ( .I(r1[14]), .ZN(n397) );
  OAI22D1BWP12T U864 ( .A1(n2851), .A2(n398), .B1(n397), .B2(n2872), .ZN(n399)
         );
  NR4D0BWP12T U865 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .ZN(n413) );
  INVD1BWP12T U866 ( .I(tmp1[14]), .ZN(n669) );
  NR2D1BWP12T U867 ( .A1(n2880), .A2(n669), .ZN(n404) );
  INVD1BWP12T U868 ( .I(r2[14]), .ZN(n672) );
  TPNR2D0BWP12T U869 ( .A1(n2789), .A2(n672), .ZN(n403) );
  AO211D1BWP12T U870 ( .A1(n2819), .A2(r9[14]), .B(n404), .C(n403), .Z(n411)
         );
  INVD3BWP12T U871 ( .I(n2891), .ZN(n2825) );
  INVD1BWP12T U872 ( .I(lr[14]), .ZN(n1252) );
  INVD1BWP12T U873 ( .I(r8[14]), .ZN(n1251) );
  OAI22D1BWP12T U874 ( .A1(n2825), .A2(n1252), .B1(n1251), .B2(n2822), .ZN(
        n410) );
  INVD3BWP12T U875 ( .I(n2893), .ZN(n2829) );
  INVD1BWP12T U876 ( .I(r10[14]), .ZN(n1250) );
  INVD1BWP12T U877 ( .I(r6[14]), .ZN(n405) );
  OAI22D1BWP12T U878 ( .A1(n2829), .A2(n1250), .B1(n405), .B2(n2826), .ZN(n409) );
  INVD1BWP12T U879 ( .I(r4[14]), .ZN(n407) );
  INVD1BWP12T U880 ( .I(r0[14]), .ZN(n406) );
  OAI22D1BWP12T U881 ( .A1(n2887), .A2(n407), .B1(n406), .B2(n2884), .ZN(n408)
         );
  NR4D1BWP12T U882 ( .A1(n411), .A2(n410), .A3(n409), .A4(n408), .ZN(n412) );
  AOI22D0BWP12T U883 ( .A1(r8[6]), .A2(n1382), .B1(n1381), .B2(r4[6]), .ZN(
        n415) );
  AOI22D0BWP12T U884 ( .A1(n[2962]), .A2(n1384), .B1(n1383), .B2(r10[6]), .ZN(
        n414) );
  CKND2D1BWP12T U885 ( .A1(n415), .A2(n414), .ZN(n424) );
  AOI22D0BWP12T U886 ( .A1(r7[6]), .A2(n1388), .B1(n1387), .B2(r5[6]), .ZN(
        n419) );
  AOI22D0BWP12T U887 ( .A1(lr[6]), .A2(n1390), .B1(n1389), .B2(r9[6]), .ZN(
        n418) );
  AOI22D0BWP12T U888 ( .A1(r6[6]), .A2(n1392), .B1(n1391), .B2(r11[6]), .ZN(
        n417) );
  CKND2D0BWP12T U889 ( .A1(n1393), .A2(r12[6]), .ZN(n416) );
  ND4D1BWP12T U890 ( .A1(n419), .A2(n418), .A3(n417), .A4(n416), .ZN(n423) );
  AOI22D0BWP12T U891 ( .A1(r3[6]), .A2(n1399), .B1(n1398), .B2(r2[6]), .ZN(
        n421) );
  AOI22D0BWP12T U892 ( .A1(n1401), .A2(r0[6]), .B1(pc_out[6]), .B2(n1400), 
        .ZN(n420) );
  OAI211D0BWP12T U893 ( .A1(n2087), .A2(n1404), .B(n421), .C(n420), .ZN(n422)
         );
  OA31D1BWP12T U894 ( .A1(n424), .A2(n423), .A3(n422), .B(n1405), .Z(
        regD_out[6]) );
  AOI22D0BWP12T U895 ( .A1(write2_in[29]), .A2(n1625), .B1(tmp1[29]), .B2(
        n1622), .ZN(n425) );
  TPOAI21D0BWP12T U896 ( .A1(n1482), .A2(n427), .B(n425), .ZN(n2166) );
  AOI22D0BWP12T U897 ( .A1(write2_in[28]), .A2(n1625), .B1(n1622), .B2(
        tmp1[28]), .ZN(n426) );
  TPOAI21D0BWP12T U898 ( .A1(n523), .A2(n427), .B(n426), .ZN(n2165) );
  INVD1BWP12T U899 ( .I(write2_in[11]), .ZN(n1366) );
  INVD1BWP12T U900 ( .I(write1_in[11]), .ZN(n537) );
  INVD1BWP12T U901 ( .I(r3[11]), .ZN(n1931) );
  OAI222D0BWP12T U902 ( .A1(n1366), .A2(n1458), .B1(n537), .B2(n1457), .C1(
        n1574), .C2(n1931), .ZN(n2532) );
  INVD1BWP12T U903 ( .I(r2[11]), .ZN(n1922) );
  OAI222D0BWP12T U904 ( .A1(n1366), .A2(n1524), .B1(n537), .B2(n1523), .C1(
        n1522), .C2(n1922), .ZN(n2564) );
  OAI222D0BWP12T U905 ( .A1(n1363), .A2(n1524), .B1(n535), .B2(n1523), .C1(
        n1522), .C2(n428), .ZN(n2565) );
  OAI222D0BWP12T U906 ( .A1(n1363), .A2(n1528), .B1(n535), .B2(n1527), .C1(
        n1526), .C2(n429), .ZN(n2309) );
  INVD1BWP12T U907 ( .I(r10[11]), .ZN(n1917) );
  OAI222D0BWP12T U908 ( .A1(n1366), .A2(n1528), .B1(n537), .B2(n1527), .C1(
        n1526), .C2(n1917), .ZN(n2308) );
  OAI222D0BWP12T U909 ( .A1(n1946), .A2(n1556), .B1(n535), .B2(n1490), .C1(
        n1363), .C2(n1444), .ZN(n2437) );
  INVD1BWP12T U910 ( .I(r11[12]), .ZN(n1960) );
  OAI222D0BWP12T U911 ( .A1(n1363), .A2(n1533), .B1(n535), .B2(n1532), .C1(
        n1530), .C2(n1960), .ZN(n2277) );
  INVD1BWP12T U912 ( .I(r6[11]), .ZN(n1934) );
  OAI222D0BWP12T U913 ( .A1(n1934), .A2(n1556), .B1(n537), .B2(n1490), .C1(
        n1366), .C2(n1444), .ZN(n2436) );
  INVD1BWP12T U914 ( .I(r11[11]), .ZN(n797) );
  OAI222D0BWP12T U915 ( .A1(n1366), .A2(n1533), .B1(n537), .B2(n1532), .C1(
        n1530), .C2(n797), .ZN(n2276) );
  INVD1BWP12T U916 ( .I(write1_in[9]), .ZN(n549) );
  INVD1BWP12T U917 ( .I(write2_in[9]), .ZN(n1338) );
  OAI222D0BWP12T U918 ( .A1(n430), .A2(n1556), .B1(n549), .B2(n1490), .C1(
        n1338), .C2(n1444), .ZN(n2434) );
  OAI222D0BWP12T U919 ( .A1(n1338), .A2(n1458), .B1(n549), .B2(n1457), .C1(
        n1574), .C2(n431), .ZN(n2530) );
  OAI222D0BWP12T U920 ( .A1(n1338), .A2(n1533), .B1(n549), .B2(n1532), .C1(
        n1530), .C2(n432), .ZN(n2274) );
  INVD1BWP12T U921 ( .I(write2_in[10]), .ZN(n1335) );
  INVD1BWP12T U922 ( .I(write1_in[10]), .ZN(n547) );
  INVD1BWP12T U923 ( .I(r11[10]), .ZN(n2778) );
  OAI222D0BWP12T U924 ( .A1(n1335), .A2(n1533), .B1(n547), .B2(n1532), .C1(
        n1530), .C2(n2778), .ZN(n2275) );
  INVD1BWP12T U925 ( .I(r6[10]), .ZN(n2798) );
  OAI222D0BWP12T U926 ( .A1(n2798), .A2(n1556), .B1(n547), .B2(n1490), .C1(
        n1335), .C2(n1444), .ZN(n2435) );
  INVD1BWP12T U927 ( .I(r3[10]), .ZN(n2779) );
  OAI222D0BWP12T U928 ( .A1(n1335), .A2(n1458), .B1(n547), .B2(n1457), .C1(
        n1574), .C2(n2779), .ZN(n2531) );
  TPNR2D2BWP12T U929 ( .A1(n434), .A2(n570), .ZN(n438) );
  CKND2D0BWP12T U930 ( .A1(write2_in[3]), .A2(n2916), .ZN(n435) );
  IOA21D2BWP12T U931 ( .A1(write1_in[3]), .A2(n2920), .B(n435), .ZN(n437) );
  TPND2D1BWP12T U932 ( .A1(n438), .A2(n437), .ZN(n1368) );
  AN2XD0BWP12T U933 ( .A1(write2_in[4]), .A2(n2916), .Z(n436) );
  TPAOI21D1BWP12T U934 ( .A1(write1_in[4]), .A2(n2920), .B(n436), .ZN(n1367)
         );
  INVD1BWP12T U935 ( .I(write2_in[5]), .ZN(n1028) );
  INVD1BWP12T U936 ( .I(write1_in[5]), .ZN(n555) );
  OAI222D0BWP12T U937 ( .A1(n1028), .A2(n1458), .B1(n555), .B2(n1457), .C1(
        n1574), .C2(n2108), .ZN(n2526) );
  INVD1BWP12T U938 ( .I(write2_in[7]), .ZN(n1203) );
  INVD1BWP12T U939 ( .I(write1_in[7]), .ZN(n565) );
  INVD1BWP12T U940 ( .I(r3[7]), .ZN(n694) );
  OAI222D0BWP12T U941 ( .A1(n1203), .A2(n1458), .B1(n565), .B2(n1457), .C1(
        n1574), .C2(n694), .ZN(n2528) );
  INVD1BWP12T U942 ( .I(write2_in[8]), .ZN(n1332) );
  INVD1BWP12T U943 ( .I(write1_in[8]), .ZN(n566) );
  OAI222D0BWP12T U944 ( .A1(n1332), .A2(n1458), .B1(n566), .B2(n1457), .C1(
        n1574), .C2(n2704), .ZN(n2529) );
  INVD1BWP12T U945 ( .I(write2_in[4]), .ZN(n1262) );
  INVD1BWP12T U946 ( .I(write1_in[4]), .ZN(n554) );
  INVD1BWP12T U947 ( .I(r3[4]), .ZN(n2018) );
  OAI222D0BWP12T U948 ( .A1(n1262), .A2(n1458), .B1(n554), .B2(n1457), .C1(
        n1574), .C2(n2018), .ZN(n2525) );
  INVD1BWP12T U949 ( .I(r11[5]), .ZN(n2110) );
  OAI222D0BWP12T U950 ( .A1(n1028), .A2(n1533), .B1(n555), .B2(n1532), .C1(
        n1530), .C2(n2110), .ZN(n2270) );
  INVD1BWP12T U951 ( .I(r11[4]), .ZN(n1852) );
  OAI222D0BWP12T U952 ( .A1(n1262), .A2(n1533), .B1(n554), .B2(n1532), .C1(
        n1530), .C2(n1852), .ZN(n2269) );
  OAI222D0BWP12T U953 ( .A1(n2721), .A2(n1556), .B1(n566), .B2(n1490), .C1(
        n1332), .C2(n1444), .ZN(n2433) );
  INVD1BWP12T U954 ( .I(r11[8]), .ZN(n2703) );
  OAI222D0BWP12T U955 ( .A1(n1332), .A2(n1533), .B1(n566), .B2(n1532), .C1(
        n1530), .C2(n2703), .ZN(n2273) );
  OAI222D0BWP12T U956 ( .A1(n1332), .A2(n1524), .B1(n566), .B2(n1523), .C1(
        n1522), .C2(n439), .ZN(n2561) );
  INVD1BWP12T U957 ( .I(write2_in[6]), .ZN(n1149) );
  INVD1BWP12T U958 ( .I(write1_in[6]), .ZN(n568) );
  INVD1BWP12T U959 ( .I(r11[6]), .ZN(n2083) );
  OAI222D0BWP12T U960 ( .A1(n1149), .A2(n1533), .B1(n568), .B2(n1532), .C1(
        n1530), .C2(n2083), .ZN(n2271) );
  OAI222D0BWP12T U961 ( .A1(n1149), .A2(n1458), .B1(n568), .B2(n1457), .C1(
        n1574), .C2(n2081), .ZN(n2527) );
  INVD3BWP12T U962 ( .I(n2871), .ZN(n2776) );
  NR2D1BWP12T U963 ( .A1(n2868), .A2(n2672), .ZN(n440) );
  AOI21D1BWP12T U964 ( .A1(n2776), .A2(pc_out[17]), .B(n440), .ZN(n447) );
  INVD1BWP12T U965 ( .I(r11[17]), .ZN(n1412) );
  INVD1BWP12T U966 ( .I(r3[17]), .ZN(n2685) );
  NR2D1BWP12T U967 ( .A1(n2860), .A2(n2685), .ZN(n441) );
  AOI21D1BWP12T U968 ( .A1(n2809), .A2(r5[17]), .B(n441), .ZN(n444) );
  INVD4BWP12T U969 ( .I(n2875), .ZN(n2708) );
  NR2D1BWP12T U970 ( .A1(n2872), .A2(n2681), .ZN(n442) );
  AOI21D1BWP12T U971 ( .A1(n2708), .A2(r12[17]), .B(n442), .ZN(n443) );
  ND2D1BWP12T U972 ( .A1(n444), .A2(n443), .ZN(n445) );
  INVD1BWP12T U973 ( .I(tmp1[17]), .ZN(n2667) );
  NR2D1BWP12T U974 ( .A1(n2880), .A2(n2667), .ZN(n449) );
  AOI21D1BWP12T U975 ( .A1(n2819), .A2(r9[17]), .B(n449), .ZN(n450) );
  IOA21D1BWP12T U976 ( .A1(n2890), .A2(r2[17]), .B(n450), .ZN(n456) );
  NR2D1BWP12T U977 ( .A1(n2822), .A2(n2688), .ZN(n451) );
  AOI21D1BWP12T U978 ( .A1(n2891), .A2(lr[17]), .B(n451), .ZN(n454) );
  INVD1BWP12T U979 ( .I(r6[17]), .ZN(n2690) );
  NR2D1BWP12T U980 ( .A1(n2826), .A2(n2690), .ZN(n452) );
  TPAOI21D0BWP12T U981 ( .A1(n2893), .A2(r10[17]), .B(n452), .ZN(n453) );
  ND2D1BWP12T U982 ( .A1(n454), .A2(n453), .ZN(n455) );
  CKND2D2BWP12T U983 ( .A1(n459), .A2(n458), .ZN(regA_out[17]) );
  INVD1BWP12T U984 ( .I(r5[2]), .ZN(n905) );
  INVD1BWP12T U985 ( .I(r10[2]), .ZN(n578) );
  OAI22D1BWP12T U986 ( .A1(n905), .A2(n2664), .B1(n2663), .B2(n578), .ZN(n465)
         );
  INVD1BWP12T U987 ( .I(tmp1[2]), .ZN(n1875) );
  AOI22D1BWP12T U988 ( .A1(r9[2]), .A2(n105), .B1(n2753), .B2(r4[2]), .ZN(n461) );
  AOI22D1BWP12T U989 ( .A1(r11[2]), .A2(n2755), .B1(n2650), .B2(r0[2]), .ZN(
        n460) );
  AO22D1BWP12T U990 ( .A1(n2750), .A2(r7[2]), .B1(n2749), .B2(r2[2]), .Z(n462)
         );
  NR4D1BWP12T U991 ( .A1(n465), .A2(n464), .A3(n463), .A4(n462), .ZN(n472) );
  INVD1BWP12T U992 ( .I(r12[2]), .ZN(n579) );
  OAI22D1BWP12T U993 ( .A1(n1885), .A2(n2680), .B1(n2679), .B2(n579), .ZN(n470) );
  INVD1BWP12T U994 ( .I(r3[2]), .ZN(n1884) );
  INVD1BWP12T U995 ( .I(lr[2]), .ZN(n580) );
  OAI22D1BWP12T U996 ( .A1(n1884), .A2(n2684), .B1(n2683), .B2(n580), .ZN(n469) );
  INVD1BWP12T U997 ( .I(r8[2]), .ZN(n1873) );
  INVD1BWP12T U998 ( .I(n[2966]), .ZN(n466) );
  OAI22D1BWP12T U999 ( .A1(n2689), .A2(n1873), .B1(n2687), .B2(n466), .ZN(n468) );
  INVD1BWP12T U1000 ( .I(pc_out[2]), .ZN(n913) );
  INVD1BWP12T U1001 ( .I(r6[2]), .ZN(n1874) );
  OAI22D1BWP12T U1002 ( .A1(n2693), .A2(n913), .B1(n2691), .B2(n1874), .ZN(
        n467) );
  NR4D0BWP12T U1003 ( .A1(n470), .A2(n469), .A3(n468), .A4(n467), .ZN(n471) );
  ND2D1BWP12T U1004 ( .A1(n472), .A2(n471), .ZN(regB_out[2]) );
  INVD1BWP12T U1005 ( .I(r5[24]), .ZN(n2845) );
  INVD1BWP12T U1006 ( .I(r10[24]), .ZN(n1193) );
  OAI22D1BWP12T U1007 ( .A1(n2845), .A2(n2664), .B1(n2663), .B2(n1193), .ZN(
        n479) );
  INVD1BWP12T U1008 ( .I(tmp1[24]), .ZN(n2838) );
  MOAI22D0BWP12T U1009 ( .A1(n2838), .A2(n2666), .B1(n2135), .B2(
        immediate2_in[24]), .ZN(n478) );
  AOI22D1BWP12T U1010 ( .A1(r9[24]), .A2(n105), .B1(n2753), .B2(r4[24]), .ZN(
        n474) );
  AOI22D1BWP12T U1011 ( .A1(r11[24]), .A2(n2755), .B1(n2650), .B2(r0[24]), 
        .ZN(n473) );
  ND2D1BWP12T U1012 ( .A1(n474), .A2(n473), .ZN(n477) );
  INVD1BWP12T U1013 ( .I(r7[24]), .ZN(n2848) );
  INVD1BWP12T U1014 ( .I(r2[24]), .ZN(n475) );
  OAI22D1BWP12T U1015 ( .A1(n2673), .A2(n2848), .B1(n2671), .B2(n475), .ZN(
        n476) );
  NR4D0BWP12T U1016 ( .A1(n479), .A2(n478), .A3(n477), .A4(n476), .ZN(n485) );
  AOI22D1BWP12T U1017 ( .A1(r1[24]), .A2(n118), .B1(n2761), .B2(r12[24]), .ZN(
        n483) );
  AOI22D1BWP12T U1018 ( .A1(r3[24]), .A2(n2763), .B1(n2762), .B2(lr[24]), .ZN(
        n482) );
  AOI22D1BWP12T U1019 ( .A1(r8[24]), .A2(n2765), .B1(n2764), .B2(n[2944]), 
        .ZN(n481) );
  AOI22D1BWP12T U1020 ( .A1(pc_out[24]), .A2(n2767), .B1(n2766), .B2(r6[24]), 
        .ZN(n480) );
  AN4XD1BWP12T U1021 ( .A1(n483), .A2(n482), .A3(n481), .A4(n480), .Z(n484) );
  ND2D1BWP12T U1022 ( .A1(n485), .A2(n484), .ZN(regB_out[24]) );
  AOI22D1BWP12T U1023 ( .A1(r1[31]), .A2(n118), .B1(n2761), .B2(r12[31]), .ZN(
        n489) );
  AOI22D1BWP12T U1024 ( .A1(r3[31]), .A2(n2763), .B1(n2762), .B2(lr[31]), .ZN(
        n488) );
  RCAOI22D0BWP12T U1025 ( .A1(r8[31]), .A2(n2765), .B1(n2764), .B2(n[2937]), 
        .ZN(n487) );
  AOI22D1BWP12T U1026 ( .A1(pc_out[31]), .A2(n2767), .B1(n2766), .B2(r6[31]), 
        .ZN(n486) );
  AN4XD1BWP12T U1027 ( .A1(n489), .A2(n488), .A3(n487), .A4(n486), .Z(n496) );
  AOI22D1BWP12T U1028 ( .A1(tmp1[31]), .A2(n2746), .B1(n2745), .B2(
        immediate2_in[31]), .ZN(n492) );
  AOI22D1BWP12T U1029 ( .A1(r9[31]), .A2(n105), .B1(n2753), .B2(r4[31]), .ZN(
        n491) );
  AOI22D1BWP12T U1030 ( .A1(r11[31]), .A2(n2755), .B1(n2733), .B2(r0[31]), 
        .ZN(n490) );
  AN3XD1BWP12T U1031 ( .A1(n492), .A2(n491), .A3(n490), .Z(n495) );
  AOI22D1BWP12T U1032 ( .A1(r5[31]), .A2(n2748), .B1(n2747), .B2(r10[31]), 
        .ZN(n494) );
  AOI22D1BWP12T U1033 ( .A1(r7[31]), .A2(n2750), .B1(n2749), .B2(r2[31]), .ZN(
        n493) );
  AOI22D0BWP12T U1034 ( .A1(r8[9]), .A2(n1382), .B1(n1381), .B2(r4[9]), .ZN(
        n498) );
  AOI22D0BWP12T U1035 ( .A1(n[2959]), .A2(n1384), .B1(n1383), .B2(r10[9]), 
        .ZN(n497) );
  CKND2D1BWP12T U1036 ( .A1(n498), .A2(n497), .ZN(n507) );
  AOI22D0BWP12T U1037 ( .A1(r7[9]), .A2(n1388), .B1(n1387), .B2(r5[9]), .ZN(
        n502) );
  AOI22D0BWP12T U1038 ( .A1(lr[9]), .A2(n1390), .B1(n1389), .B2(r9[9]), .ZN(
        n501) );
  AOI22D0BWP12T U1039 ( .A1(r6[9]), .A2(n1392), .B1(n1391), .B2(r11[9]), .ZN(
        n500) );
  CKND2D0BWP12T U1040 ( .A1(n1393), .A2(r12[9]), .ZN(n499) );
  ND4D1BWP12T U1041 ( .A1(n502), .A2(n501), .A3(n500), .A4(n499), .ZN(n506) );
  AOI22D0BWP12T U1042 ( .A1(r3[9]), .A2(n1399), .B1(n1398), .B2(r2[9]), .ZN(
        n504) );
  AOI22D0BWP12T U1043 ( .A1(n1401), .A2(r0[9]), .B1(pc_out[9]), .B2(n1400), 
        .ZN(n503) );
  OAI211D0BWP12T U1044 ( .A1(n540), .A2(n1404), .B(n504), .C(n503), .ZN(n505)
         );
  OA31D1BWP12T U1045 ( .A1(n507), .A2(n506), .A3(n505), .B(n1405), .Z(
        regD_out[9]) );
  AOI22D0BWP12T U1046 ( .A1(write2_in[28]), .A2(n1513), .B1(n1511), .B2(r2[28]), .ZN(n508) );
  TPOAI21D0BWP12T U1047 ( .A1(n523), .A2(n1523), .B(n508), .ZN(n2581) );
  AOI22D0BWP12T U1048 ( .A1(write2_in[28]), .A2(n1594), .B1(n1507), .B2(r9[28]), .ZN(n509) );
  TPOAI21D0BWP12T U1049 ( .A1(n523), .A2(n1481), .B(n509), .ZN(n2357) );
  AOI22D0BWP12T U1050 ( .A1(write2_in[28]), .A2(n1558), .B1(n1519), .B2(r6[28]), .ZN(n510) );
  TPOAI21D0BWP12T U1051 ( .A1(n523), .A2(n1490), .B(n510), .ZN(n2453) );
  AOI22D0BWP12T U1052 ( .A1(write2_in[28]), .A2(n1570), .B1(n1505), .B2(r7[28]), .ZN(n511) );
  TPOAI21D0BWP12T U1053 ( .A1(n523), .A2(n1451), .B(n511), .ZN(n2421) );
  AOI22D0BWP12T U1054 ( .A1(write2_in[28]), .A2(n1510), .B1(n1508), .B2(
        r11[28]), .ZN(n512) );
  TPOAI21D0BWP12T U1055 ( .A1(n523), .A2(n1532), .B(n512), .ZN(n2293) );
  AOI22D0BWP12T U1056 ( .A1(write2_in[28]), .A2(n1604), .B1(n1603), .B2(r8[28]), .ZN(n513) );
  TPOAI21D0BWP12T U1057 ( .A1(n523), .A2(n1478), .B(n513), .ZN(n2389) );
  AOI22D0BWP12T U1058 ( .A1(write2_in[28]), .A2(n1564), .B1(n1520), .B2(r5[28]), .ZN(n514) );
  TPOAI21D0BWP12T U1059 ( .A1(n523), .A2(n1445), .B(n514), .ZN(n2485) );
  AOI22D0BWP12T U1060 ( .A1(write2_in[28]), .A2(n1552), .B1(n1506), .B2(r0[28]), .ZN(n515) );
  TPOAI21D0BWP12T U1061 ( .A1(n523), .A2(n1454), .B(n515), .ZN(n2645) );
  AOI22D0BWP12T U1062 ( .A1(write2_in[28]), .A2(n1609), .B1(n1608), .B2(lr[28]), .ZN(n516) );
  TPOAI21D0BWP12T U1063 ( .A1(n523), .A2(n1475), .B(n516), .ZN(n2229) );
  AOI22D0BWP12T U1064 ( .A1(write2_in[28]), .A2(n1617), .B1(n1521), .B2(
        n[2940]), .ZN(n517) );
  TPOAI21D0BWP12T U1065 ( .A1(n523), .A2(n1442), .B(n517), .ZN(spin[28]) );
  AOI22D0BWP12T U1066 ( .A1(write2_in[28]), .A2(n1516), .B1(n1514), .B2(
        r10[28]), .ZN(n518) );
  TPOAI21D0BWP12T U1067 ( .A1(n523), .A2(n1527), .B(n518), .ZN(n2325) );
  AOI22D0BWP12T U1068 ( .A1(write2_in[28]), .A2(n1599), .B1(n1598), .B2(
        r12[28]), .ZN(n519) );
  TPOAI21D0BWP12T U1069 ( .A1(n523), .A2(n1436), .B(n519), .ZN(n2261) );
  AOI22D0BWP12T U1070 ( .A1(write2_in[28]), .A2(n1588), .B1(n1517), .B2(r1[28]), .ZN(n520) );
  TPOAI21D0BWP12T U1071 ( .A1(n523), .A2(n1447), .B(n520), .ZN(n2613) );
  AOI22D0BWP12T U1072 ( .A1(write2_in[28]), .A2(n1576), .B1(n1504), .B2(r3[28]), .ZN(n521) );
  TPOAI21D0BWP12T U1073 ( .A1(n523), .A2(n1457), .B(n521), .ZN(n2549) );
  AOI22D0BWP12T U1074 ( .A1(write2_in[28]), .A2(n1582), .B1(n1518), .B2(r4[28]), .ZN(n522) );
  TPOAI21D0BWP12T U1075 ( .A1(n523), .A2(n1449), .B(n522), .ZN(n2517) );
  AOI22D0BWP12T U1076 ( .A1(write2_in[30]), .A2(n1617), .B1(n1521), .B2(
        n[2938]), .ZN(n524) );
  TPOAI21D0BWP12T U1077 ( .A1(n1491), .A2(n1442), .B(n524), .ZN(spin[30]) );
  AOI22D0BWP12T U1078 ( .A1(write2_in[30]), .A2(n1604), .B1(n1603), .B2(r8[30]), .ZN(n525) );
  TPOAI21D0BWP12T U1079 ( .A1(n1491), .A2(n1478), .B(n525), .ZN(n2391) );
  AOI22D0BWP12T U1080 ( .A1(write2_in[30]), .A2(n1582), .B1(n1518), .B2(r4[30]), .ZN(n526) );
  TPOAI21D0BWP12T U1081 ( .A1(n1491), .A2(n1449), .B(n526), .ZN(n2519) );
  AOI22D0BWP12T U1082 ( .A1(write2_in[30]), .A2(n1564), .B1(n1520), .B2(r5[30]), .ZN(n527) );
  TPOAI21D0BWP12T U1083 ( .A1(n1491), .A2(n1445), .B(n527), .ZN(n2487) );
  AOI22D0BWP12T U1084 ( .A1(write2_in[29]), .A2(n1599), .B1(r12[29]), .B2(
        n1598), .ZN(n528) );
  TPOAI21D0BWP12T U1085 ( .A1(n1482), .A2(n1436), .B(n528), .ZN(n2262) );
  AOI22D0BWP12T U1086 ( .A1(write2_in[30]), .A2(n1599), .B1(n1598), .B2(
        r12[30]), .ZN(n529) );
  TPOAI21D0BWP12T U1087 ( .A1(n1491), .A2(n1436), .B(n529), .ZN(n2263) );
  INVD1BWP12T U1088 ( .I(n1527), .ZN(n1515) );
  BUFFD6BWP12T U1089 ( .I(write1_in[14]), .Z(n1471) );
  AO222D1BWP12T U1090 ( .A1(n1515), .A2(n1471), .B1(n1516), .B2(write2_in[14]), 
        .C1(n1514), .C2(r10[14]), .Z(n2311) );
  AO222D1BWP12T U1091 ( .A1(n1567), .A2(n1471), .B1(n1505), .B2(r7[14]), .C1(
        write2_in[14]), .C2(n1570), .Z(n2407) );
  AO222D1BWP12T U1092 ( .A1(n1573), .A2(n1471), .B1(n1576), .B2(write2_in[14]), 
        .C1(n1504), .C2(r3[14]), .Z(n2535) );
  AO222D1BWP12T U1093 ( .A1(n1561), .A2(n1471), .B1(n1520), .B2(r5[14]), .C1(
        write2_in[14]), .C2(n1564), .Z(n2471) );
  INVD1BWP12T U1094 ( .I(n1523), .ZN(n1512) );
  AO222D1BWP12T U1095 ( .A1(n1512), .A2(n1471), .B1(n1513), .B2(write2_in[14]), 
        .C1(n1511), .C2(r2[14]), .Z(n2567) );
  AO222D1BWP12T U1096 ( .A1(n1602), .A2(n1471), .B1(n1603), .B2(r8[14]), .C1(
        write2_in[14]), .C2(n1604), .Z(n2375) );
  AO222D1BWP12T U1097 ( .A1(n1579), .A2(n1471), .B1(n1518), .B2(r4[14]), .C1(
        write2_in[14]), .C2(n1582), .Z(n2503) );
  INVD1BWP12T U1098 ( .I(n1447), .ZN(n1585) );
  AO222D1BWP12T U1099 ( .A1(n1585), .A2(n1471), .B1(n1517), .B2(r1[14]), .C1(
        write2_in[14]), .C2(n1588), .Z(n2599) );
  AO222D1BWP12T U1100 ( .A1(n1597), .A2(n1471), .B1(n1598), .B2(r12[14]), .C1(
        write2_in[14]), .C2(n1599), .Z(n2247) );
  INVD1BWP12T U1101 ( .I(n1532), .ZN(n1509) );
  AO222D1BWP12T U1102 ( .A1(n1509), .A2(n1471), .B1(n1510), .B2(write2_in[14]), 
        .C1(n1508), .C2(r11[14]), .Z(n2279) );
  INVD1BWP12T U1103 ( .I(n1454), .ZN(n1549) );
  AO222D1BWP12T U1104 ( .A1(n1549), .A2(n1471), .B1(n1506), .B2(r0[14]), .C1(
        write2_in[14]), .C2(n1552), .Z(n2631) );
  OAI222D0BWP12T U1105 ( .A1(n530), .A2(n1438), .B1(n535), .B2(n1475), .C1(
        n1363), .C2(n1439), .ZN(n2213) );
  OAI222D0BWP12T U1106 ( .A1(n1125), .A2(n1435), .B1(n535), .B2(n1436), .C1(
        n1363), .C2(n1437), .ZN(n2245) );
  INVD1BWP12T U1107 ( .I(lr[11]), .ZN(n1930) );
  OAI222D0BWP12T U1108 ( .A1(n1930), .A2(n1438), .B1(n537), .B2(n1475), .C1(
        n1366), .C2(n1439), .ZN(n2212) );
  CKND0BWP12T U1109 ( .I(r9[11]), .ZN(n531) );
  OAI222D0BWP12T U1110 ( .A1(n531), .A2(n1592), .B1(n537), .B2(n1481), .C1(
        n1366), .C2(n1453), .ZN(n2340) );
  CKND0BWP12T U1111 ( .I(r4[12]), .ZN(n532) );
  OAI222D0BWP12T U1112 ( .A1(n532), .A2(n1580), .B1(n535), .B2(n1449), .C1(
        n1363), .C2(n1450), .ZN(n2501) );
  CKND0BWP12T U1113 ( .I(r9[12]), .ZN(n533) );
  OAI222D0BWP12T U1114 ( .A1(n533), .A2(n1592), .B1(n535), .B2(n1481), .C1(
        n1363), .C2(n1453), .ZN(n2341) );
  CKND0BWP12T U1115 ( .I(r4[11]), .ZN(n534) );
  OAI222D0BWP12T U1116 ( .A1(n534), .A2(n1580), .B1(n537), .B2(n1449), .C1(
        n1366), .C2(n1450), .ZN(n2500) );
  INVD1BWP12T U1117 ( .I(r12[11]), .ZN(n1928) );
  OAI222D0BWP12T U1118 ( .A1(n1928), .A2(n1435), .B1(n537), .B2(n1436), .C1(
        n1366), .C2(n1437), .ZN(n2244) );
  INVD1BWP12T U1119 ( .I(r1[11]), .ZN(n1929) );
  OAI222D0BWP12T U1120 ( .A1(n1929), .A2(n1586), .B1(n537), .B2(n1447), .C1(
        n1366), .C2(n1448), .ZN(n2596) );
  INVD1BWP12T U1121 ( .I(r8[11]), .ZN(n1933) );
  OAI222D0BWP12T U1122 ( .A1(n1933), .A2(n1440), .B1(n537), .B2(n1478), .C1(
        n1366), .C2(n1441), .ZN(n2372) );
  OAI222D0BWP12T U1123 ( .A1(n1963), .A2(n1586), .B1(n535), .B2(n1447), .C1(
        n1363), .C2(n1448), .ZN(n2597) );
  OAI222D0BWP12T U1124 ( .A1(n1957), .A2(n1568), .B1(n535), .B2(n1451), .C1(
        n1363), .C2(n1452), .ZN(n2405) );
  INVD1BWP12T U1125 ( .I(r7[11]), .ZN(n1923) );
  OAI222D0BWP12T U1126 ( .A1(n1923), .A2(n1568), .B1(n537), .B2(n1451), .C1(
        n1366), .C2(n1452), .ZN(n2404) );
  INVD1BWP12T U1127 ( .I(r0[12]), .ZN(n1949) );
  OAI222D0BWP12T U1128 ( .A1(n1949), .A2(n1550), .B1(n535), .B2(n1454), .C1(
        n1363), .C2(n1455), .ZN(n2629) );
  INVD1BWP12T U1129 ( .I(r5[11]), .ZN(n1918) );
  OAI222D0BWP12T U1130 ( .A1(n1918), .A2(n1562), .B1(n537), .B2(n1445), .C1(
        n1366), .C2(n1446), .ZN(n2468) );
  OAI222D0BWP12T U1131 ( .A1(n1942), .A2(n1440), .B1(n535), .B2(n1478), .C1(
        n1363), .C2(n1441), .ZN(n2373) );
  OAI222D0BWP12T U1132 ( .A1(n536), .A2(n1562), .B1(n535), .B2(n1445), .C1(
        n1363), .C2(n1446), .ZN(n2469) );
  CKND0BWP12T U1133 ( .I(r0[11]), .ZN(n538) );
  OAI222D0BWP12T U1134 ( .A1(n538), .A2(n1550), .B1(n537), .B2(n1454), .C1(
        n1366), .C2(n1455), .ZN(n2628) );
  AO222D1BWP12T U1135 ( .A1(n1509), .A2(write1_in[13]), .B1(n1510), .B2(
        write2_in[13]), .C1(n1508), .C2(r11[13]), .Z(n2278) );
  AO222D1BWP12T U1136 ( .A1(n1561), .A2(write1_in[13]), .B1(n1520), .B2(r5[13]), .C1(write2_in[13]), .C2(n1564), .Z(n2470) );
  AO222D1BWP12T U1137 ( .A1(n1573), .A2(write1_in[13]), .B1(n1576), .B2(
        write2_in[13]), .C1(n1504), .C2(r3[13]), .Z(n2534) );
  AO222D0BWP12T U1138 ( .A1(n1620), .A2(write1_in[11]), .B1(n1625), .B2(
        write2_in[11]), .C1(n1622), .C2(tmp1[11]), .Z(n2148) );
  AO222D0BWP12T U1139 ( .A1(n1620), .A2(write1_in[12]), .B1(n1625), .B2(
        write2_in[12]), .C1(n1622), .C2(tmp1[12]), .Z(n2149) );
  AO222D1BWP12T U1140 ( .A1(n1512), .A2(write1_in[13]), .B1(n1513), .B2(
        write2_in[13]), .C1(n1511), .C2(r2[13]), .Z(n2566) );
  AO222D1BWP12T U1141 ( .A1(n1515), .A2(write1_in[13]), .B1(n1516), .B2(
        write2_in[13]), .C1(n1514), .C2(r10[13]), .Z(n2310) );
  OAI222D0BWP12T U1142 ( .A1(n539), .A2(n1438), .B1(n549), .B2(n1475), .C1(
        n1338), .C2(n1439), .ZN(n2210) );
  INVD1BWP12T U1143 ( .I(r2[10]), .ZN(n2788) );
  OAI222D0BWP12T U1144 ( .A1(n1335), .A2(n1524), .B1(n547), .B2(n1523), .C1(
        n1522), .C2(n2788), .ZN(n2563) );
  INVD1BWP12T U1145 ( .I(lr[10]), .ZN(n712) );
  OAI222D0BWP12T U1146 ( .A1(n712), .A2(n1438), .B1(n547), .B2(n1475), .C1(
        n1335), .C2(n1439), .ZN(n2211) );
  CKND0BWP12T U1147 ( .I(r9[9]), .ZN(n1033) );
  OAI222D0BWP12T U1148 ( .A1(n1033), .A2(n1592), .B1(n549), .B2(n1481), .C1(
        n1338), .C2(n1453), .ZN(n2338) );
  OAI222D0BWP12T U1149 ( .A1(n540), .A2(n1586), .B1(n549), .B2(n1447), .C1(
        n1338), .C2(n1448), .ZN(n2594) );
  INVD1BWP12T U1150 ( .I(r7[10]), .ZN(n2774) );
  OAI222D0BWP12T U1151 ( .A1(n2774), .A2(n1568), .B1(n547), .B2(n1451), .C1(
        n1335), .C2(n1452), .ZN(n2403) );
  OAI222D0BWP12T U1152 ( .A1(n541), .A2(n1435), .B1(n549), .B2(n1436), .C1(
        n1338), .C2(n1437), .ZN(n2242) );
  INVD1BWP12T U1153 ( .I(r12[10]), .ZN(n711) );
  OAI222D0BWP12T U1154 ( .A1(n711), .A2(n1435), .B1(n547), .B2(n1436), .C1(
        n1335), .C2(n1437), .ZN(n2243) );
  OAI222D0BWP12T U1155 ( .A1(n542), .A2(n1568), .B1(n549), .B2(n1451), .C1(
        n1338), .C2(n1452), .ZN(n2402) );
  INVD1BWP12T U1156 ( .I(r1[10]), .ZN(n2781) );
  OAI222D0BWP12T U1157 ( .A1(n2781), .A2(n1586), .B1(n547), .B2(n1447), .C1(
        n1335), .C2(n1448), .ZN(n2595) );
  OAI222D0BWP12T U1158 ( .A1(n1338), .A2(n1524), .B1(n549), .B2(n1523), .C1(
        n1522), .C2(n543), .ZN(n2562) );
  CKND0BWP12T U1159 ( .I(r9[10]), .ZN(n544) );
  OAI222D0BWP12T U1160 ( .A1(n544), .A2(n1592), .B1(n547), .B2(n1481), .C1(
        n1335), .C2(n1453), .ZN(n2339) );
  INVD1BWP12T U1161 ( .I(r10[10]), .ZN(n704) );
  OAI222D0BWP12T U1162 ( .A1(n1335), .A2(n1528), .B1(n547), .B2(n1527), .C1(
        n1526), .C2(n704), .ZN(n2307) );
  OAI222D0BWP12T U1163 ( .A1(n1338), .A2(n1528), .B1(n549), .B2(n1527), .C1(
        n1526), .C2(n545), .ZN(n2306) );
  CKND0BWP12T U1164 ( .I(r4[10]), .ZN(n1300) );
  OAI222D0BWP12T U1165 ( .A1(n1300), .A2(n1580), .B1(n547), .B2(n1449), .C1(
        n1335), .C2(n1450), .ZN(n2499) );
  OAI222D0BWP12T U1166 ( .A1(n546), .A2(n1550), .B1(n549), .B2(n1454), .C1(
        n1338), .C2(n1455), .ZN(n2626) );
  INVD1BWP12T U1167 ( .I(r8[10]), .ZN(n2796) );
  OAI222D0BWP12T U1168 ( .A1(n2796), .A2(n1440), .B1(n547), .B2(n1478), .C1(
        n1335), .C2(n1441), .ZN(n2371) );
  INVD1BWP12T U1169 ( .I(r5[10]), .ZN(n1305) );
  OAI222D0BWP12T U1170 ( .A1(n1305), .A2(n1562), .B1(n547), .B2(n1445), .C1(
        n1335), .C2(n1446), .ZN(n2467) );
  CKND0BWP12T U1171 ( .I(r0[10]), .ZN(n1310) );
  OAI222D0BWP12T U1172 ( .A1(n1310), .A2(n1550), .B1(n547), .B2(n1454), .C1(
        n1335), .C2(n1455), .ZN(n2627) );
  OAI222D0BWP12T U1173 ( .A1(n1034), .A2(n1440), .B1(n549), .B2(n1478), .C1(
        n1338), .C2(n1441), .ZN(n2370) );
  OAI222D0BWP12T U1174 ( .A1(n548), .A2(n1562), .B1(n549), .B2(n1445), .C1(
        n1338), .C2(n1446), .ZN(n2466) );
  CKND0BWP12T U1175 ( .I(r4[9]), .ZN(n550) );
  OAI222D0BWP12T U1176 ( .A1(n550), .A2(n1580), .B1(n549), .B2(n1449), .C1(
        n1338), .C2(n1450), .ZN(n2498) );
  INVD1BWP12T U1177 ( .I(r8[4]), .ZN(n2020) );
  OAI222D0BWP12T U1178 ( .A1(n2020), .A2(n1440), .B1(n554), .B2(n1478), .C1(
        n1262), .C2(n1441), .ZN(n2365) );
  INVD1BWP12T U1179 ( .I(r5[4]), .ZN(n2005) );
  OAI222D0BWP12T U1180 ( .A1(n2005), .A2(n1562), .B1(n554), .B2(n1445), .C1(
        n1262), .C2(n1446), .ZN(n2461) );
  INVD1BWP12T U1181 ( .I(r4[5]), .ZN(n2123) );
  OAI222D0BWP12T U1182 ( .A1(n2123), .A2(n1580), .B1(n555), .B2(n1449), .C1(
        n1028), .C2(n1450), .ZN(n2494) );
  INVD1BWP12T U1183 ( .I(r7[4]), .ZN(n2010) );
  OAI222D0BWP12T U1184 ( .A1(n2010), .A2(n1568), .B1(n554), .B2(n1451), .C1(
        n1262), .C2(n1452), .ZN(n2397) );
  OAI222D0BWP12T U1185 ( .A1(n2112), .A2(n1568), .B1(n555), .B2(n1451), .C1(
        n1028), .C2(n1452), .ZN(n2398) );
  CKND0BWP12T U1186 ( .I(r9[4]), .ZN(n551) );
  OAI222D0BWP12T U1187 ( .A1(n551), .A2(n1592), .B1(n554), .B2(n1481), .C1(
        n1262), .C2(n1453), .ZN(n2333) );
  CKND0BWP12T U1188 ( .I(r0[4]), .ZN(n552) );
  OAI222D0BWP12T U1189 ( .A1(n552), .A2(n1550), .B1(n554), .B2(n1454), .C1(
        n1262), .C2(n1455), .ZN(n2621) );
  AO222D0BWP12T U1190 ( .A1(n1620), .A2(write1_in[9]), .B1(n1625), .B2(
        write2_in[9]), .C1(n1622), .C2(tmp1[9]), .Z(n2146) );
  CKND1BWP12T U1191 ( .I(r4[4]), .ZN(n1854) );
  OAI222D0BWP12T U1192 ( .A1(n1854), .A2(n1580), .B1(n554), .B2(n1449), .C1(
        n1262), .C2(n1450), .ZN(n2493) );
  INVD1BWP12T U1193 ( .I(r9[5]), .ZN(n2121) );
  OAI222D0BWP12T U1194 ( .A1(n2121), .A2(n1592), .B1(n555), .B2(n1481), .C1(
        n1028), .C2(n1453), .ZN(n2334) );
  OAI222D0BWP12T U1195 ( .A1(n2128), .A2(n1440), .B1(n555), .B2(n1478), .C1(
        n1028), .C2(n1441), .ZN(n2366) );
  AO222D0BWP12T U1196 ( .A1(n1620), .A2(write1_in[10]), .B1(n1625), .B2(
        write2_in[10]), .C1(n1622), .C2(tmp1[10]), .Z(n2147) );
  INVD1BWP12T U1197 ( .I(r10[4]), .ZN(n2004) );
  OAI222D0BWP12T U1198 ( .A1(n1262), .A2(n1528), .B1(n554), .B2(n1527), .C1(
        n1526), .C2(n2004), .ZN(n2301) );
  INVD1BWP12T U1199 ( .I(r0[5]), .ZN(n2122) );
  OAI222D0BWP12T U1200 ( .A1(n2122), .A2(n1550), .B1(n555), .B2(n1454), .C1(
        n1028), .C2(n1455), .ZN(n2622) );
  INVD1BWP12T U1201 ( .I(r6[4]), .ZN(n2021) );
  OAI222D0BWP12T U1202 ( .A1(n2021), .A2(n1556), .B1(n554), .B2(n1490), .C1(
        n1262), .C2(n1444), .ZN(n2429) );
  INVD1BWP12T U1203 ( .I(r12[4]), .ZN(n2015) );
  OAI222D0BWP12T U1204 ( .A1(n2015), .A2(n1435), .B1(n554), .B2(n1436), .C1(
        n1262), .C2(n1437), .ZN(n2237) );
  OAI222D0BWP12T U1205 ( .A1(n1028), .A2(n1528), .B1(n555), .B2(n1527), .C1(
        n1526), .C2(n2127), .ZN(n2302) );
  OAI222D0BWP12T U1206 ( .A1(n2115), .A2(n1435), .B1(n555), .B2(n1436), .C1(
        n1028), .C2(n1437), .ZN(n2238) );
  INVD1BWP12T U1207 ( .I(r2[4]), .ZN(n2009) );
  OAI222D0BWP12T U1208 ( .A1(n1262), .A2(n1524), .B1(n554), .B2(n1523), .C1(
        n1522), .C2(n2009), .ZN(n2557) );
  OAI222D0BWP12T U1209 ( .A1(n2016), .A2(n1586), .B1(n554), .B2(n1447), .C1(
        n1262), .C2(n1448), .ZN(n2589) );
  OAI222D0BWP12T U1210 ( .A1(n1028), .A2(n1524), .B1(n555), .B2(n1523), .C1(
        n1522), .C2(n553), .ZN(n2558) );
  OAI222D0BWP12T U1211 ( .A1(n2129), .A2(n1438), .B1(n555), .B2(n1475), .C1(
        n1028), .C2(n1439), .ZN(n2206) );
  OAI222D0BWP12T U1212 ( .A1(n2126), .A2(n1556), .B1(n555), .B2(n1490), .C1(
        n1028), .C2(n1444), .ZN(n2430) );
  OAI222D0BWP12T U1213 ( .A1(n2109), .A2(n1562), .B1(n555), .B2(n1445), .C1(
        n1028), .C2(n1446), .ZN(n2462) );
  INVD1BWP12T U1214 ( .I(lr[4]), .ZN(n2017) );
  OAI222D0BWP12T U1215 ( .A1(n2017), .A2(n1438), .B1(n554), .B2(n1475), .C1(
        n1262), .C2(n1439), .ZN(n2205) );
  OAI222D0BWP12T U1216 ( .A1(n2114), .A2(n1586), .B1(n555), .B2(n1447), .C1(
        n1028), .C2(n1448), .ZN(n2590) );
  INVD1BWP12T U1217 ( .I(r2[7]), .ZN(n688) );
  OAI222D0BWP12T U1218 ( .A1(n1203), .A2(n1524), .B1(n565), .B2(n1523), .C1(
        n1522), .C2(n688), .ZN(n2560) );
  INVD1BWP12T U1219 ( .I(write2_in[3]), .ZN(n1163) );
  INVD1BWP12T U1220 ( .I(write1_in[3]), .ZN(n567) );
  INVD1BWP12T U1221 ( .I(r10[3]), .ZN(n871) );
  OAI222D0BWP12T U1222 ( .A1(n1163), .A2(n1528), .B1(n567), .B2(n1527), .C1(
        n1526), .C2(n871), .ZN(n2300) );
  INVD1BWP12T U1223 ( .I(r6[7]), .ZN(n696) );
  OAI222D0BWP12T U1224 ( .A1(n696), .A2(n1556), .B1(n565), .B2(n1490), .C1(
        n1203), .C2(n1444), .ZN(n2432) );
  INVD1BWP12T U1225 ( .I(r8[3]), .ZN(n870) );
  OAI222D0BWP12T U1226 ( .A1(n870), .A2(n1440), .B1(n567), .B2(n1478), .C1(
        n1163), .C2(n1441), .ZN(n2364) );
  OAI222D0BWP12T U1227 ( .A1(n1149), .A2(n1528), .B1(n568), .B2(n1527), .C1(
        n1526), .C2(n2100), .ZN(n2303) );
  CKND0BWP12T U1228 ( .I(r9[8]), .ZN(n556) );
  OAI222D0BWP12T U1229 ( .A1(n556), .A2(n1592), .B1(n566), .B2(n1481), .C1(
        n1332), .C2(n1453), .ZN(n2337) );
  OAI222D0BWP12T U1230 ( .A1(n1149), .A2(n1524), .B1(n568), .B2(n1523), .C1(
        n1522), .C2(n557), .ZN(n2559) );
  OAI222D0BWP12T U1231 ( .A1(n1332), .A2(n1528), .B1(n566), .B2(n1527), .C1(
        n1526), .C2(n558), .ZN(n2305) );
  INVD1BWP12T U1232 ( .I(r7[3]), .ZN(n928) );
  OAI222D0BWP12T U1233 ( .A1(n928), .A2(n1568), .B1(n567), .B2(n1451), .C1(
        n1163), .C2(n1452), .ZN(n2396) );
  OAI222D0BWP12T U1234 ( .A1(n2099), .A2(n1556), .B1(n568), .B2(n1490), .C1(
        n1149), .C2(n1444), .ZN(n2431) );
  CKND0BWP12T U1235 ( .I(r4[8]), .ZN(n559) );
  OAI222D0BWP12T U1236 ( .A1(n559), .A2(n1580), .B1(n566), .B2(n1449), .C1(
        n1332), .C2(n1450), .ZN(n2497) );
  CKND0BWP12T U1237 ( .I(r9[7]), .ZN(n560) );
  OAI222D0BWP12T U1238 ( .A1(n560), .A2(n1592), .B1(n565), .B2(n1481), .C1(
        n1203), .C2(n1453), .ZN(n2336) );
  OAI222D0BWP12T U1239 ( .A1(n2085), .A2(n1568), .B1(n568), .B2(n1451), .C1(
        n1149), .C2(n1452), .ZN(n2399) );
  INVD1BWP12T U1240 ( .I(r6[3]), .ZN(n931) );
  OAI222D0BWP12T U1241 ( .A1(n931), .A2(n1556), .B1(n567), .B2(n1490), .C1(
        n1163), .C2(n1444), .ZN(n2428) );
  INVD1BWP12T U1242 ( .I(r7[7]), .ZN(n689) );
  OAI222D0BWP12T U1243 ( .A1(n689), .A2(n1568), .B1(n565), .B2(n1451), .C1(
        n1203), .C2(n1452), .ZN(n2400) );
  CKND0BWP12T U1244 ( .I(r4[7]), .ZN(n561) );
  OAI222D0BWP12T U1245 ( .A1(n561), .A2(n1580), .B1(n565), .B2(n1449), .C1(
        n1203), .C2(n1450), .ZN(n2496) );
  INVD1BWP12T U1246 ( .I(r5[3]), .ZN(n930) );
  OAI222D0BWP12T U1247 ( .A1(n930), .A2(n1562), .B1(n567), .B2(n1445), .C1(
        n1163), .C2(n1446), .ZN(n2460) );
  OAI222D0BWP12T U1248 ( .A1(n2700), .A2(n1568), .B1(n566), .B2(n1451), .C1(
        n1332), .C2(n1452), .ZN(n2401) );
  OAI222D0BWP12T U1249 ( .A1(n1067), .A2(n1435), .B1(n566), .B2(n1436), .C1(
        n1332), .C2(n1437), .ZN(n2241) );
  INVD1BWP12T U1250 ( .I(r12[7]), .ZN(n1090) );
  OAI222D0BWP12T U1251 ( .A1(n1090), .A2(n1435), .B1(n565), .B2(n1436), .C1(
        n1203), .C2(n1437), .ZN(n2240) );
  INVD1BWP12T U1252 ( .I(r4[6]), .ZN(n2096) );
  OAI222D0BWP12T U1253 ( .A1(n2096), .A2(n1580), .B1(n568), .B2(n1449), .C1(
        n1149), .C2(n1450), .ZN(n2495) );
  INVD1BWP12T U1254 ( .I(r10[7]), .ZN(n1091) );
  OAI222D0BWP12T U1255 ( .A1(n1203), .A2(n1528), .B1(n565), .B2(n1527), .C1(
        n1526), .C2(n1091), .ZN(n2304) );
  OAI222D0BWP12T U1256 ( .A1(n2088), .A2(n1435), .B1(n568), .B2(n1436), .C1(
        n1149), .C2(n1437), .ZN(n2239) );
  INVD1BWP12T U1257 ( .I(r9[6]), .ZN(n2094) );
  OAI222D0BWP12T U1258 ( .A1(n2094), .A2(n1592), .B1(n568), .B2(n1481), .C1(
        n1149), .C2(n1453), .ZN(n2335) );
  CKND0BWP12T U1259 ( .I(r4[3]), .ZN(n927) );
  OAI222D0BWP12T U1260 ( .A1(n927), .A2(n1580), .B1(n567), .B2(n1449), .C1(
        n1163), .C2(n1450), .ZN(n2492) );
  INVD1BWP12T U1261 ( .I(r12[3]), .ZN(n659) );
  OAI222D0BWP12T U1262 ( .A1(n659), .A2(n1435), .B1(n567), .B2(n1436), .C1(
        n1163), .C2(n1437), .ZN(n2236) );
  OAI222D0BWP12T U1263 ( .A1(n562), .A2(n1438), .B1(n566), .B2(n1475), .C1(
        n1332), .C2(n1439), .ZN(n2209) );
  INVD1BWP12T U1264 ( .I(r1[3]), .ZN(n929) );
  OAI222D0BWP12T U1265 ( .A1(n929), .A2(n1586), .B1(n567), .B2(n1447), .C1(
        n1163), .C2(n1448), .ZN(n2588) );
  OAI222D0BWP12T U1266 ( .A1(n2087), .A2(n1586), .B1(n568), .B2(n1447), .C1(
        n1149), .C2(n1448), .ZN(n2591) );
  INVD1BWP12T U1267 ( .I(r0[8]), .ZN(n2714) );
  OAI222D0BWP12T U1268 ( .A1(n2714), .A2(n1550), .B1(n566), .B2(n1454), .C1(
        n1332), .C2(n1455), .ZN(n2625) );
  CKND0BWP12T U1269 ( .I(r9[3]), .ZN(n563) );
  OAI222D0BWP12T U1270 ( .A1(n563), .A2(n1592), .B1(n567), .B2(n1481), .C1(
        n1163), .C2(n1453), .ZN(n2332) );
  INVD1BWP12T U1271 ( .I(r1[7]), .ZN(n768) );
  OAI222D0BWP12T U1272 ( .A1(n768), .A2(n1586), .B1(n565), .B2(n1447), .C1(
        n1203), .C2(n1448), .ZN(n2592) );
  INVD1BWP12T U1273 ( .I(r0[7]), .ZN(n617) );
  OAI222D0BWP12T U1274 ( .A1(n617), .A2(n1550), .B1(n565), .B2(n1454), .C1(
        n1203), .C2(n1455), .ZN(n2624) );
  INVD1BWP12T U1275 ( .I(lr[7]), .ZN(n1092) );
  OAI222D0BWP12T U1276 ( .A1(n1092), .A2(n1438), .B1(n565), .B2(n1475), .C1(
        n1203), .C2(n1439), .ZN(n2208) );
  OAI222D0BWP12T U1277 ( .A1(n2706), .A2(n1586), .B1(n566), .B2(n1447), .C1(
        n1332), .C2(n1448), .ZN(n2593) );
  INVD1BWP12T U1278 ( .I(r0[6]), .ZN(n2095) );
  OAI222D0BWP12T U1279 ( .A1(n2095), .A2(n1550), .B1(n568), .B2(n1454), .C1(
        n1149), .C2(n1455), .ZN(n2623) );
  INVD1BWP12T U1280 ( .I(lr[3]), .ZN(n660) );
  OAI222D0BWP12T U1281 ( .A1(n660), .A2(n1438), .B1(n567), .B2(n1475), .C1(
        n1163), .C2(n1439), .ZN(n2204) );
  INVD1BWP12T U1282 ( .I(r0[3]), .ZN(n934) );
  OAI222D0BWP12T U1283 ( .A1(n934), .A2(n1550), .B1(n567), .B2(n1454), .C1(
        n1163), .C2(n1455), .ZN(n2620) );
  OAI222D0BWP12T U1284 ( .A1(n2102), .A2(n1438), .B1(n568), .B2(n1475), .C1(
        n1149), .C2(n1439), .ZN(n2207) );
  OAI222D0BWP12T U1285 ( .A1(n564), .A2(n1562), .B1(n566), .B2(n1445), .C1(
        n1332), .C2(n1446), .ZN(n2465) );
  INVD1BWP12T U1286 ( .I(r5[7]), .ZN(n684) );
  OAI222D0BWP12T U1287 ( .A1(n684), .A2(n1562), .B1(n565), .B2(n1445), .C1(
        n1203), .C2(n1446), .ZN(n2464) );
  OAI222D0BWP12T U1288 ( .A1(n2082), .A2(n1562), .B1(n568), .B2(n1445), .C1(
        n1149), .C2(n1446), .ZN(n2463) );
  AO222D0BWP12T U1289 ( .A1(n1620), .A2(write1_in[5]), .B1(n1625), .B2(
        write2_in[5]), .C1(n1622), .C2(tmp1[5]), .Z(n2142) );
  INVD1BWP12T U1290 ( .I(r2[3]), .ZN(n932) );
  OAI222D0BWP12T U1291 ( .A1(n1163), .A2(n1524), .B1(n567), .B2(n1523), .C1(
        n1522), .C2(n932), .ZN(n2556) );
  INVD1BWP12T U1292 ( .I(r3[3]), .ZN(n933) );
  OAI222D0BWP12T U1293 ( .A1(n1163), .A2(n1458), .B1(n567), .B2(n1457), .C1(
        n1574), .C2(n933), .ZN(n2524) );
  INVD1BWP12T U1294 ( .I(r8[7]), .ZN(n1089) );
  OAI222D0BWP12T U1295 ( .A1(n1089), .A2(n1440), .B1(n565), .B2(n1478), .C1(
        n1203), .C2(n1441), .ZN(n2368) );
  INVD1BWP12T U1296 ( .I(r11[7]), .ZN(n609) );
  OAI222D0BWP12T U1297 ( .A1(n1203), .A2(n1533), .B1(n565), .B2(n1532), .C1(
        n1530), .C2(n609), .ZN(n2272) );
  OAI222D0BWP12T U1298 ( .A1(n2719), .A2(n1440), .B1(n566), .B2(n1478), .C1(
        n1332), .C2(n1441), .ZN(n2369) );
  INVD1BWP12T U1299 ( .I(r11[3]), .ZN(n884) );
  OAI222D0BWP12T U1300 ( .A1(n1163), .A2(n1533), .B1(n567), .B2(n1532), .C1(
        n1530), .C2(n884), .ZN(n2268) );
  OAI222D0BWP12T U1301 ( .A1(n2101), .A2(n1440), .B1(n568), .B2(n1478), .C1(
        n1149), .C2(n1441), .ZN(n2367) );
  CKND2D0BWP12T U1302 ( .A1(n570), .A2(n569), .ZN(n572) );
  TPAOI21D0BWP12T U1303 ( .A1(n1488), .A2(next_pc_in[1]), .B(reset), .ZN(n571)
         );
  OAI211D0BWP12T U1304 ( .A1(n2924), .A2(n1140), .B(n572), .C(n571), .ZN(n2170) );
  AO222D0BWP12T U1305 ( .A1(n1620), .A2(write1_in[8]), .B1(n1625), .B2(
        write2_in[8]), .C1(n1622), .C2(tmp1[8]), .Z(n2145) );
  AO222D0BWP12T U1306 ( .A1(n1620), .A2(write1_in[6]), .B1(n1625), .B2(
        write2_in[6]), .C1(n1622), .C2(tmp1[6]), .Z(n2143) );
  AO222D0BWP12T U1307 ( .A1(n1620), .A2(write1_in[3]), .B1(n1625), .B2(
        write2_in[3]), .C1(n1622), .C2(tmp1[3]), .Z(n2140) );
  INVD1BWP12T U1308 ( .I(write2_in[1]), .ZN(n1022) );
  INVD1BWP12T U1309 ( .I(write1_in[1]), .ZN(n576) );
  OAI222D0BWP12T U1310 ( .A1(n1022), .A2(n1528), .B1(n576), .B2(n1527), .C1(
        n1526), .C2(n573), .ZN(n2298) );
  OAI222D0BWP12T U1311 ( .A1(n1137), .A2(n1440), .B1(n576), .B2(n1478), .C1(
        n1022), .C2(n1441), .ZN(n2362) );
  OAI222D0BWP12T U1312 ( .A1(n1022), .A2(n1524), .B1(n576), .B2(n1523), .C1(
        n1522), .C2(n574), .ZN(n2554) );
  OAI222D0BWP12T U1313 ( .A1(n1022), .A2(n1458), .B1(n576), .B2(n1457), .C1(
        n1574), .C2(n840), .ZN(n2522) );
  INVD1BWP12T U1314 ( .I(r11[1]), .ZN(n839) );
  OAI222D0BWP12T U1315 ( .A1(n1022), .A2(n1533), .B1(n576), .B2(n1532), .C1(
        n1530), .C2(n839), .ZN(n2266) );
  OAI222D0BWP12T U1316 ( .A1(n837), .A2(n1568), .B1(n576), .B2(n1451), .C1(
        n1022), .C2(n1452), .ZN(n2394) );
  INVD1BWP12T U1317 ( .I(r9[1]), .ZN(n852) );
  OAI222D0BWP12T U1318 ( .A1(n852), .A2(n1592), .B1(n576), .B2(n1481), .C1(
        n1022), .C2(n1453), .ZN(n2330) );
  CKND0BWP12T U1319 ( .I(r4[1]), .ZN(n575) );
  OAI222D0BWP12T U1320 ( .A1(n575), .A2(n1580), .B1(n576), .B2(n1449), .C1(
        n1022), .C2(n1450), .ZN(n2490) );
  OAI222D0BWP12T U1321 ( .A1(n842), .A2(n1586), .B1(n576), .B2(n1447), .C1(
        n1022), .C2(n1448), .ZN(n2586) );
  OAI222D0BWP12T U1322 ( .A1(n858), .A2(n1556), .B1(n576), .B2(n1490), .C1(
        n1022), .C2(n1444), .ZN(n2426) );
  OAI222D0BWP12T U1323 ( .A1(n1139), .A2(n1435), .B1(n576), .B2(n1436), .C1(
        n1022), .C2(n1437), .ZN(n2234) );
  OAI222D0BWP12T U1324 ( .A1(n1138), .A2(n1438), .B1(n576), .B2(n1475), .C1(
        n1022), .C2(n1439), .ZN(n2202) );
  INVD1BWP12T U1325 ( .I(r0[1]), .ZN(n849) );
  OAI222D0BWP12T U1326 ( .A1(n849), .A2(n1550), .B1(n576), .B2(n1454), .C1(
        n1022), .C2(n1455), .ZN(n2618) );
  OAI222D0BWP12T U1327 ( .A1(n577), .A2(n1562), .B1(n576), .B2(n1445), .C1(
        n1022), .C2(n1446), .ZN(n2458) );
  INVD1BWP12T U1328 ( .I(write2_in[2]), .ZN(n1025) );
  INVD1BWP12T U1329 ( .I(write1_in[2]), .ZN(n582) );
  OAI222D0BWP12T U1330 ( .A1(n1025), .A2(n1528), .B1(n582), .B2(n1527), .C1(
        n1526), .C2(n578), .ZN(n2299) );
  CKND0BWP12T U1331 ( .I(r4[2]), .ZN(n903) );
  OAI222D0BWP12T U1332 ( .A1(n903), .A2(n1580), .B1(n582), .B2(n1449), .C1(
        n1025), .C2(n1450), .ZN(n2491) );
  OAI222D0BWP12T U1333 ( .A1(n579), .A2(n1435), .B1(n582), .B2(n1436), .C1(
        n1025), .C2(n1437), .ZN(n2235) );
  INVD1BWP12T U1334 ( .I(r7[2]), .ZN(n1881) );
  OAI222D0BWP12T U1335 ( .A1(n1881), .A2(n1568), .B1(n582), .B2(n1451), .C1(
        n1025), .C2(n1452), .ZN(n2395) );
  OAI222D0BWP12T U1336 ( .A1(n1885), .A2(n1586), .B1(n582), .B2(n1447), .C1(
        n1025), .C2(n1448), .ZN(n2587) );
  OAI222D0BWP12T U1337 ( .A1(n580), .A2(n1438), .B1(n582), .B2(n1475), .C1(
        n1025), .C2(n1439), .ZN(n2203) );
  OAI222D0BWP12T U1338 ( .A1(n905), .A2(n1562), .B1(n582), .B2(n1445), .C1(
        n1025), .C2(n1446), .ZN(n2459) );
  OAI222D0BWP12T U1339 ( .A1(n1874), .A2(n1556), .B1(n582), .B2(n1490), .C1(
        n1025), .C2(n1444), .ZN(n2427) );
  INVD1BWP12T U1340 ( .I(r0[2]), .ZN(n1877) );
  OAI222D0BWP12T U1341 ( .A1(n1877), .A2(n1550), .B1(n582), .B2(n1454), .C1(
        n1025), .C2(n1455), .ZN(n2619) );
  CKND0BWP12T U1342 ( .I(r9[2]), .ZN(n581) );
  OAI222D0BWP12T U1343 ( .A1(n581), .A2(n1592), .B1(n582), .B2(n1481), .C1(
        n1025), .C2(n1453), .ZN(n2331) );
  OAI222D0BWP12T U1344 ( .A1(n1025), .A2(n1458), .B1(n582), .B2(n1457), .C1(
        n1574), .C2(n1884), .ZN(n2523) );
  AO222D0BWP12T U1345 ( .A1(n1620), .A2(write1_in[1]), .B1(n1625), .B2(
        write2_in[1]), .C1(n1622), .C2(tmp1[1]), .Z(n2138) );
  INVD1BWP12T U1346 ( .I(r11[2]), .ZN(n1883) );
  OAI222D0BWP12T U1347 ( .A1(n1025), .A2(n1533), .B1(n582), .B2(n1532), .C1(
        n1530), .C2(n1883), .ZN(n2267) );
  CKND0BWP12T U1348 ( .I(r2[2]), .ZN(n907) );
  OAI222D0BWP12T U1349 ( .A1(n1025), .A2(n1524), .B1(n582), .B2(n1523), .C1(
        n1522), .C2(n907), .ZN(n2555) );
  OAI222D0BWP12T U1350 ( .A1(n1873), .A2(n1440), .B1(n582), .B2(n1478), .C1(
        n1025), .C2(n1441), .ZN(n2363) );
  BUFFD1BWP12T U1351 ( .I(write2_in[0]), .Z(n583) );
  AO222D0BWP12T U1352 ( .A1(n1620), .A2(write1_in[2]), .B1(n1625), .B2(
        write2_in[2]), .C1(n1622), .C2(tmp1[2]), .Z(n2139) );
  AO222D0BWP12T U1353 ( .A1(n1579), .A2(write1_in[0]), .B1(n1518), .B2(r4[0]), 
        .C1(n583), .C2(n1582), .Z(n2489) );
  AO222D0BWP12T U1354 ( .A1(n1602), .A2(write1_in[0]), .B1(n1603), .B2(r8[0]), 
        .C1(n583), .C2(n1604), .Z(n2361) );
  AO222D0BWP12T U1355 ( .A1(n1515), .A2(write1_in[0]), .B1(n1516), .B2(n583), 
        .C1(n1514), .C2(r10[0]), .Z(n2297) );
  AO222D0BWP12T U1356 ( .A1(n1585), .A2(write1_in[0]), .B1(n1517), .B2(r1[0]), 
        .C1(n583), .C2(n1588), .Z(n2585) );
  AO222D0BWP12T U1357 ( .A1(n1597), .A2(write1_in[0]), .B1(n1598), .B2(r12[0]), 
        .C1(n583), .C2(n1599), .Z(n2233) );
  AO222D0BWP12T U1358 ( .A1(n1607), .A2(write1_in[0]), .B1(n1608), .B2(lr[0]), 
        .C1(n583), .C2(n1609), .Z(n2201) );
  AO222D0BWP12T U1359 ( .A1(n1567), .A2(write1_in[0]), .B1(n1505), .B2(r7[0]), 
        .C1(n583), .C2(n1570), .Z(n2393) );
  AO222D0BWP12T U1360 ( .A1(n1614), .A2(write1_in[0]), .B1(n1521), .B2(n[2968]), .C1(n583), .C2(n1617), .Z(spin[0]) );
  AO222D0BWP12T U1361 ( .A1(n1573), .A2(write1_in[0]), .B1(n1576), .B2(n583), 
        .C1(n1504), .C2(r3[0]), .Z(n2521) );
  AO222D0BWP12T U1362 ( .A1(n1620), .A2(write1_in[0]), .B1(n1625), .B2(n583), 
        .C1(n1622), .C2(tmp1[0]), .Z(n2136) );
  AO222D0BWP12T U1363 ( .A1(n1591), .A2(write1_in[0]), .B1(n1507), .B2(r9[0]), 
        .C1(n583), .C2(n1594), .Z(n2329) );
  AO222D0BWP12T U1364 ( .A1(n1509), .A2(write1_in[0]), .B1(n1510), .B2(n583), 
        .C1(n1508), .C2(r11[0]), .Z(n2265) );
  AO222D0BWP12T U1365 ( .A1(n1561), .A2(write1_in[0]), .B1(n1520), .B2(r5[0]), 
        .C1(n583), .C2(n1564), .Z(n2457) );
  AO222D0BWP12T U1366 ( .A1(n1555), .A2(write1_in[0]), .B1(n1519), .B2(r6[0]), 
        .C1(n583), .C2(n1558), .Z(n2425) );
  AO222D0BWP12T U1367 ( .A1(n1549), .A2(write1_in[0]), .B1(n1506), .B2(r0[0]), 
        .C1(n583), .C2(n1552), .Z(n2617) );
  AO222D0BWP12T U1368 ( .A1(n1512), .A2(write1_in[0]), .B1(n1513), .B2(n583), 
        .C1(n1511), .C2(r2[0]), .Z(n2553) );
  CKND1BWP12T U1369 ( .I(n584), .ZN(n1943) );
  INVD1BWP12T U1370 ( .I(r8[15]), .ZN(n1055) );
  INR2D1BWP12T U1371 ( .A1(tmp1[15]), .B1(n2880), .ZN(n585) );
  AOI21D1BWP12T U1372 ( .A1(n2819), .A2(r9[15]), .B(n585), .ZN(n589) );
  INR2D1BWP12T U1373 ( .A1(r2[15]), .B1(n2789), .ZN(n586) );
  AOI21D1BWP12T U1374 ( .A1(n2791), .A2(r4[15]), .B(n586), .ZN(n588) );
  INVD1P75BWP12T U1375 ( .I(n2884), .ZN(n2795) );
  ND2D1BWP12T U1376 ( .A1(n2795), .A2(r0[15]), .ZN(n587) );
  INR3D2BWP12T U1377 ( .A1(n592), .B1(n591), .B2(n590), .ZN(n606) );
  INR2D1BWP12T U1378 ( .A1(r3[15]), .B1(n593), .ZN(n594) );
  AOI21D1BWP12T U1379 ( .A1(n2809), .A2(r5[15]), .B(n594), .ZN(n597) );
  INR2D1BWP12T U1380 ( .A1(r1[15]), .B1(n2872), .ZN(n595) );
  AOI21D1BWP12T U1381 ( .A1(n2708), .A2(r12[15]), .B(n595), .ZN(n596) );
  ND2D1BWP12T U1382 ( .A1(n597), .A2(n596), .ZN(n604) );
  INVD1BWP12T U1383 ( .I(r11[15]), .ZN(n599) );
  ND2D1BWP12T U1384 ( .A1(n2807), .A2(n[2953]), .ZN(n598) );
  OAI21D1BWP12T U1385 ( .A1(n2864), .A2(n599), .B(n598), .ZN(n603) );
  INVD1BWP12T U1386 ( .I(r7[15]), .ZN(n601) );
  ND2D1BWP12T U1387 ( .A1(n2811), .A2(pc_out[15]), .ZN(n600) );
  OAI21D1BWP12T U1388 ( .A1(n2868), .A2(n601), .B(n600), .ZN(n602) );
  TPNR3D1BWP12T U1389 ( .A1(n604), .A2(n603), .A3(n602), .ZN(n605) );
  ND2D2BWP12T U1390 ( .A1(n606), .A2(n605), .ZN(regA_out[15]) );
  NR2D1BWP12T U1391 ( .A1(n2868), .A2(n689), .ZN(n607) );
  AOI21D1BWP12T U1392 ( .A1(n2776), .A2(pc_out[7]), .B(n607), .ZN(n616) );
  ND2D1BWP12T U1393 ( .A1(n2807), .A2(n[2961]), .ZN(n608) );
  OAI21D1BWP12T U1394 ( .A1(n2864), .A2(n609), .B(n608), .ZN(n615) );
  NR2D1BWP12T U1395 ( .A1(n2860), .A2(n694), .ZN(n610) );
  AOI21D1BWP12T U1396 ( .A1(n2809), .A2(r5[7]), .B(n610), .ZN(n613) );
  NR2D1BWP12T U1397 ( .A1(n2872), .A2(n768), .ZN(n611) );
  AOI21D1BWP12T U1398 ( .A1(n2813), .A2(r12[7]), .B(n611), .ZN(n612) );
  ND2D1BWP12T U1399 ( .A1(n613), .A2(n612), .ZN(n614) );
  INR3D2BWP12T U1400 ( .A1(n616), .B1(n615), .B2(n614), .ZN(n628) );
  INVD1BWP12T U1401 ( .I(tmp1[7]), .ZN(n685) );
  IOA21D1BWP12T U1402 ( .A1(n2890), .A2(r2[7]), .B(n619), .ZN(n625) );
  NR2D1BWP12T U1403 ( .A1(n2822), .A2(n1089), .ZN(n620) );
  AOI21D1BWP12T U1404 ( .A1(n2891), .A2(lr[7]), .B(n620), .ZN(n623) );
  NR2D1BWP12T U1405 ( .A1(n2826), .A2(n696), .ZN(n621) );
  AOI21D1BWP12T U1406 ( .A1(n2893), .A2(r10[7]), .B(n621), .ZN(n622) );
  ND2D1BWP12T U1407 ( .A1(n623), .A2(n622), .ZN(n624) );
  INR3D0BWP12T U1408 ( .A1(n626), .B1(n625), .B2(n624), .ZN(n627) );
  CKND2D2BWP12T U1409 ( .A1(n628), .A2(n627), .ZN(regA_out[7]) );
  INVD1BWP12T U1410 ( .I(r5[23]), .ZN(n2862) );
  INVD1BWP12T U1411 ( .I(r10[23]), .ZN(n1430) );
  OAI22D1BWP12T U1412 ( .A1(n2862), .A2(n2664), .B1(n2663), .B2(n1430), .ZN(
        n634) );
  INVD1BWP12T U1413 ( .I(tmp1[23]), .ZN(n2881) );
  MOAI22D0BWP12T U1414 ( .A1(n2881), .A2(n2666), .B1(n2745), .B2(
        immediate2_in[23]), .ZN(n633) );
  AOI22D1BWP12T U1415 ( .A1(r9[23]), .A2(n105), .B1(n2753), .B2(r4[23]), .ZN(
        n630) );
  AOI22D1BWP12T U1416 ( .A1(r11[23]), .A2(n2755), .B1(n2754), .B2(r0[23]), 
        .ZN(n629) );
  ND2D1BWP12T U1417 ( .A1(n630), .A2(n629), .ZN(n632) );
  INVD1BWP12T U1418 ( .I(r7[23]), .ZN(n2869) );
  INVD1BWP12T U1419 ( .I(r2[23]), .ZN(n1429) );
  OAI22D1BWP12T U1420 ( .A1(n2673), .A2(n2869), .B1(n2671), .B2(n1429), .ZN(
        n631) );
  NR4D0BWP12T U1421 ( .A1(n634), .A2(n633), .A3(n632), .A4(n631), .ZN(n640) );
  AOI22D1BWP12T U1422 ( .A1(r1[23]), .A2(n118), .B1(n2761), .B2(r12[23]), .ZN(
        n638) );
  AOI22D1BWP12T U1423 ( .A1(r3[23]), .A2(n2763), .B1(n2762), .B2(lr[23]), .ZN(
        n637) );
  AOI22D1BWP12T U1424 ( .A1(r8[23]), .A2(n2765), .B1(n2764), .B2(n[2945]), 
        .ZN(n636) );
  AOI22D1BWP12T U1425 ( .A1(pc_out[23]), .A2(n2767), .B1(n2766), .B2(r6[23]), 
        .ZN(n635) );
  AN4XD1BWP12T U1426 ( .A1(n638), .A2(n637), .A3(n636), .A4(n635), .Z(n639) );
  CKND2D1BWP12T U1427 ( .A1(n640), .A2(n639), .ZN(regB_out[23]) );
  INVD1BWP12T U1428 ( .I(r5[22]), .ZN(n737) );
  INVD1BWP12T U1429 ( .I(r10[22]), .ZN(n1460) );
  OAI22D1BWP12T U1430 ( .A1(n737), .A2(n2664), .B1(n2663), .B2(n1460), .ZN(
        n646) );
  INVD1BWP12T U1431 ( .I(tmp1[22]), .ZN(n745) );
  MOAI22D0BWP12T U1432 ( .A1(n745), .A2(n2666), .B1(n2730), .B2(
        immediate2_in[22]), .ZN(n645) );
  AOI22D1BWP12T U1433 ( .A1(r9[22]), .A2(n105), .B1(n2753), .B2(r4[22]), .ZN(
        n642) );
  AOI22D1BWP12T U1434 ( .A1(r11[22]), .A2(n2755), .B1(n2650), .B2(r0[22]), 
        .ZN(n641) );
  ND2D1BWP12T U1435 ( .A1(n642), .A2(n641), .ZN(n644) );
  INVD1BWP12T U1436 ( .I(r7[22]), .ZN(n738) );
  INVD1BWP12T U1437 ( .I(r2[22]), .ZN(n1462) );
  OAI22D1BWP12T U1438 ( .A1(n2673), .A2(n738), .B1(n2671), .B2(n1462), .ZN(
        n643) );
  NR4D0BWP12T U1439 ( .A1(n646), .A2(n645), .A3(n644), .A4(n643), .ZN(n652) );
  AOI22D1BWP12T U1440 ( .A1(r1[22]), .A2(n118), .B1(n2761), .B2(r12[22]), .ZN(
        n650) );
  AOI22D1BWP12T U1441 ( .A1(r3[22]), .A2(n2763), .B1(n2762), .B2(lr[22]), .ZN(
        n649) );
  AOI22D1BWP12T U1442 ( .A1(r8[22]), .A2(n2765), .B1(n2764), .B2(n[2946]), 
        .ZN(n648) );
  AOI22D1BWP12T U1443 ( .A1(pc_out[22]), .A2(n2767), .B1(n2766), .B2(r6[22]), 
        .ZN(n647) );
  AN4XD1BWP12T U1444 ( .A1(n650), .A2(n649), .A3(n648), .A4(n647), .Z(n651) );
  CKND2D1BWP12T U1445 ( .A1(n652), .A2(n651), .ZN(regB_out[22]) );
  OAI22D1BWP12T U1446 ( .A1(n930), .A2(n2664), .B1(n2663), .B2(n871), .ZN(n658) );
  INVD1BWP12T U1447 ( .I(tmp1[3]), .ZN(n867) );
  MOAI22D0BWP12T U1448 ( .A1(n867), .A2(n2666), .B1(n2745), .B2(
        immediate2_in[3]), .ZN(n657) );
  AOI22D1BWP12T U1449 ( .A1(r9[3]), .A2(n105), .B1(n2753), .B2(r4[3]), .ZN(
        n654) );
  AOI22D1BWP12T U1450 ( .A1(r11[3]), .A2(n2755), .B1(n2733), .B2(r0[3]), .ZN(
        n653) );
  OAI22D1BWP12T U1451 ( .A1(n2673), .A2(n928), .B1(n2671), .B2(n932), .ZN(n655) );
  NR4D0BWP12T U1452 ( .A1(n658), .A2(n657), .A3(n656), .A4(n655), .ZN(n667) );
  OAI22D1BWP12T U1453 ( .A1(n659), .A2(n2679), .B1(n2680), .B2(n929), .ZN(n665) );
  OAI22D1BWP12T U1454 ( .A1(n933), .A2(n2684), .B1(n2683), .B2(n660), .ZN(n664) );
  INVD1BWP12T U1455 ( .I(n[2965]), .ZN(n661) );
  OAI22D1BWP12T U1456 ( .A1(n2689), .A2(n870), .B1(n2687), .B2(n661), .ZN(n663) );
  INVD1BWP12T U1457 ( .I(pc_out[3]), .ZN(n939) );
  OAI22D1BWP12T U1458 ( .A1(n2693), .A2(n939), .B1(n2691), .B2(n931), .ZN(n662) );
  NR4D0BWP12T U1459 ( .A1(n665), .A2(n664), .A3(n663), .A4(n662), .ZN(n666) );
  ND2D1BWP12T U1460 ( .A1(n667), .A2(n666), .ZN(regB_out[3]) );
  OAI22D1BWP12T U1461 ( .A1(n668), .A2(n2664), .B1(n2663), .B2(n1250), .ZN(
        n677) );
  MOAI22D0BWP12T U1462 ( .A1(n669), .A2(n2666), .B1(n2730), .B2(
        immediate2_in[14]), .ZN(n676) );
  AOI22D1BWP12T U1463 ( .A1(r9[14]), .A2(n105), .B1(n2753), .B2(r4[14]), .ZN(
        n671) );
  AOI22D1BWP12T U1464 ( .A1(r11[14]), .A2(n2755), .B1(n2650), .B2(r0[14]), 
        .ZN(n670) );
  ND2D1BWP12T U1465 ( .A1(n671), .A2(n670), .ZN(n675) );
  OAI22D1BWP12T U1466 ( .A1(n2673), .A2(n673), .B1(n2671), .B2(n672), .ZN(n674) );
  NR4D0BWP12T U1467 ( .A1(n677), .A2(n676), .A3(n675), .A4(n674), .ZN(n683) );
  AOI22D1BWP12T U1468 ( .A1(r1[14]), .A2(n118), .B1(n2761), .B2(r12[14]), .ZN(
        n681) );
  AOI22D1BWP12T U1469 ( .A1(r3[14]), .A2(n2763), .B1(n2762), .B2(lr[14]), .ZN(
        n680) );
  AOI22D1BWP12T U1470 ( .A1(r8[14]), .A2(n2765), .B1(n2764), .B2(n[2954]), 
        .ZN(n679) );
  AOI22D1BWP12T U1471 ( .A1(pc_out[14]), .A2(n2767), .B1(n2766), .B2(r6[14]), 
        .ZN(n678) );
  AN4XD1BWP12T U1472 ( .A1(n681), .A2(n680), .A3(n679), .A4(n678), .Z(n682) );
  CKND2D1BWP12T U1473 ( .A1(n683), .A2(n682), .ZN(regB_out[14]) );
  OAI22D1BWP12T U1474 ( .A1(n684), .A2(n2664), .B1(n2663), .B2(n1091), .ZN(
        n693) );
  MOAI22D0BWP12T U1475 ( .A1(n685), .A2(n2666), .B1(n2730), .B2(
        immediate2_in[7]), .ZN(n692) );
  AOI22D1BWP12T U1476 ( .A1(r9[7]), .A2(n105), .B1(n2753), .B2(r4[7]), .ZN(
        n687) );
  AOI22D1BWP12T U1477 ( .A1(r11[7]), .A2(n2755), .B1(n2733), .B2(r0[7]), .ZN(
        n686) );
  ND2D1BWP12T U1478 ( .A1(n687), .A2(n686), .ZN(n691) );
  OAI22D1BWP12T U1479 ( .A1(n2673), .A2(n689), .B1(n2671), .B2(n688), .ZN(n690) );
  NR4D0BWP12T U1480 ( .A1(n693), .A2(n692), .A3(n691), .A4(n690), .ZN(n703) );
  OAI22D1BWP12T U1481 ( .A1(n768), .A2(n2680), .B1(n2679), .B2(n1090), .ZN(
        n701) );
  OAI22D1BWP12T U1482 ( .A1(n694), .A2(n2684), .B1(n2683), .B2(n1092), .ZN(
        n700) );
  INVD0BWP12T U1483 ( .I(n[2961]), .ZN(n695) );
  OAI22D1BWP12T U1484 ( .A1(n2689), .A2(n1089), .B1(n2687), .B2(n695), .ZN(
        n699) );
  INVD0BWP12T U1485 ( .I(pc_out[7]), .ZN(n697) );
  OAI22D1BWP12T U1486 ( .A1(n2693), .A2(n697), .B1(n2691), .B2(n696), .ZN(n698) );
  NR4D0BWP12T U1487 ( .A1(n701), .A2(n700), .A3(n699), .A4(n698), .ZN(n702) );
  CKND2D1BWP12T U1488 ( .A1(n703), .A2(n702), .ZN(regB_out[7]) );
  OAI22D1BWP12T U1489 ( .A1(n1305), .A2(n2664), .B1(n2663), .B2(n704), .ZN(
        n710) );
  INVD1BWP12T U1490 ( .I(tmp1[10]), .ZN(n2792) );
  MOAI22D0BWP12T U1491 ( .A1(n2792), .A2(n2666), .B1(n2135), .B2(
        immediate2_in[10]), .ZN(n709) );
  AOI22D1BWP12T U1492 ( .A1(r9[10]), .A2(n105), .B1(n2753), .B2(r4[10]), .ZN(
        n706) );
  AOI22D1BWP12T U1493 ( .A1(r11[10]), .A2(n2755), .B1(n2754), .B2(r0[10]), 
        .ZN(n705) );
  ND2D1BWP12T U1494 ( .A1(n706), .A2(n705), .ZN(n708) );
  OAI22D1BWP12T U1495 ( .A1(n2673), .A2(n2774), .B1(n2671), .B2(n2788), .ZN(
        n707) );
  NR4D0BWP12T U1496 ( .A1(n710), .A2(n709), .A3(n708), .A4(n707), .ZN(n719) );
  OAI22D1BWP12T U1497 ( .A1(n2781), .A2(n2680), .B1(n2679), .B2(n711), .ZN(
        n717) );
  OAI22D1BWP12T U1498 ( .A1(n2779), .A2(n2684), .B1(n2683), .B2(n712), .ZN(
        n716) );
  INVD1BWP12T U1499 ( .I(n[2958]), .ZN(n1315) );
  OAI22D1BWP12T U1500 ( .A1(n2689), .A2(n2796), .B1(n2687), .B2(n1315), .ZN(
        n715) );
  INVD1BWP12T U1501 ( .I(pc_out[10]), .ZN(n713) );
  OAI22D1BWP12T U1502 ( .A1(n2693), .A2(n713), .B1(n2691), .B2(n2798), .ZN(
        n714) );
  NR4D0BWP12T U1503 ( .A1(n717), .A2(n716), .A3(n715), .A4(n714), .ZN(n718) );
  CKND2D1BWP12T U1504 ( .A1(n719), .A2(n718), .ZN(regB_out[10]) );
  AOI22D1BWP12T U1505 ( .A1(n2808), .A2(r11[13]), .B1(n2807), .B2(n[2955]), 
        .ZN(n723) );
  AOI22D1BWP12T U1506 ( .A1(r3[13]), .A2(n2810), .B1(n2809), .B2(r5[13]), .ZN(
        n722) );
  AOI22D1BWP12T U1507 ( .A1(n2812), .A2(r7[13]), .B1(n2811), .B2(pc_out[13]), 
        .ZN(n721) );
  AN4D2BWP12T U1508 ( .A1(n723), .A2(n722), .A3(n721), .A4(n720), .Z(n735) );
  INVD2BWP12T U1509 ( .I(n2880), .ZN(n2820) );
  AOI22D1BWP12T U1510 ( .A1(tmp1[13]), .A2(n2820), .B1(n2819), .B2(r9[13]), 
        .ZN(n724) );
  IOA21D1BWP12T U1511 ( .A1(r2[13]), .A2(n2890), .B(n724), .ZN(n733) );
  INVD1BWP12T U1512 ( .I(lr[13]), .ZN(n1004) );
  INVD1BWP12T U1513 ( .I(r8[13]), .ZN(n725) );
  OAI22D1BWP12T U1514 ( .A1(n2825), .A2(n1004), .B1(n725), .B2(n2822), .ZN(
        n732) );
  INVD1BWP12T U1515 ( .I(r10[13]), .ZN(n727) );
  INVD1BWP12T U1516 ( .I(r6[13]), .ZN(n726) );
  OAI22D1BWP12T U1517 ( .A1(n2829), .A2(n727), .B1(n726), .B2(n2826), .ZN(n731) );
  INVD1BWP12T U1518 ( .I(r4[13]), .ZN(n729) );
  INVD1BWP12T U1519 ( .I(r0[13]), .ZN(n728) );
  OAI22D1BWP12T U1520 ( .A1(n2887), .A2(n729), .B1(n728), .B2(n2884), .ZN(n730) );
  NR4D2BWP12T U1521 ( .A1(n733), .A2(n732), .A3(n731), .A4(n730), .ZN(n734) );
  INVD1BWP12T U1522 ( .I(r3[22]), .ZN(n736) );
  OAI22D1BWP12T U1523 ( .A1(n2863), .A2(n737), .B1(n736), .B2(n2860), .ZN(n744) );
  INVD1BWP12T U1524 ( .I(n[2946]), .ZN(n1292) );
  INVD1BWP12T U1525 ( .I(r11[22]), .ZN(n1461) );
  OAI22D0BWP12T U1526 ( .A1(n2867), .A2(n1292), .B1(n1461), .B2(n2864), .ZN(
        n743) );
  INVD1BWP12T U1527 ( .I(pc_out[22]), .ZN(n1750) );
  OAI22D1BWP12T U1528 ( .A1(n2871), .A2(n1750), .B1(n738), .B2(n2868), .ZN(
        n742) );
  INVD1BWP12T U1529 ( .I(r12[22]), .ZN(n740) );
  INVD1BWP12T U1530 ( .I(r1[22]), .ZN(n739) );
  OAI22D1BWP12T U1531 ( .A1(n2875), .A2(n740), .B1(n739), .B2(n2872), .ZN(n741) );
  NR4D0BWP12T U1532 ( .A1(n744), .A2(n743), .A3(n742), .A4(n741), .ZN(n756) );
  NR2D1BWP12T U1533 ( .A1(n2880), .A2(n745), .ZN(n747) );
  NR2D1BWP12T U1534 ( .A1(n2789), .A2(n1462), .ZN(n746) );
  AO211D1BWP12T U1535 ( .A1(n2819), .A2(r9[22]), .B(n747), .C(n746), .Z(n754)
         );
  INVD1BWP12T U1536 ( .I(lr[22]), .ZN(n1288) );
  INVD1BWP12T U1537 ( .I(r8[22]), .ZN(n1290) );
  OAI22D1BWP12T U1538 ( .A1(n2825), .A2(n1288), .B1(n1290), .B2(n2822), .ZN(
        n753) );
  INVD1BWP12T U1539 ( .I(r6[22]), .ZN(n748) );
  OAI22D1BWP12T U1540 ( .A1(n2829), .A2(n1460), .B1(n748), .B2(n2826), .ZN(
        n752) );
  INVD1BWP12T U1541 ( .I(r4[22]), .ZN(n750) );
  INVD1BWP12T U1542 ( .I(r0[22]), .ZN(n749) );
  OAI22D1BWP12T U1543 ( .A1(n2887), .A2(n750), .B1(n749), .B2(n2884), .ZN(n751) );
  NR4D0BWP12T U1544 ( .A1(n754), .A2(n753), .A3(n752), .A4(n751), .ZN(n755) );
  CKND2D1BWP12T U1545 ( .A1(n756), .A2(n755), .ZN(regA_out[22]) );
  AOI22D1BWP12T U1546 ( .A1(r1[28]), .A2(n118), .B1(n2761), .B2(r12[28]), .ZN(
        n760) );
  AOI22D1BWP12T U1547 ( .A1(r3[28]), .A2(n2763), .B1(n2762), .B2(lr[28]), .ZN(
        n759) );
  AOI22D1BWP12T U1548 ( .A1(r8[28]), .A2(n2765), .B1(n2764), .B2(n[2940]), 
        .ZN(n758) );
  AOI22D1BWP12T U1549 ( .A1(pc_out[28]), .A2(n2767), .B1(n2766), .B2(r6[28]), 
        .ZN(n757) );
  AN4XD1BWP12T U1550 ( .A1(n760), .A2(n759), .A3(n758), .A4(n757), .Z(n767) );
  AOI22D1BWP12T U1551 ( .A1(tmp1[28]), .A2(n2746), .B1(n2135), .B2(
        immediate2_in[28]), .ZN(n763) );
  AOI22D1BWP12T U1552 ( .A1(r9[28]), .A2(n105), .B1(n2753), .B2(r4[28]), .ZN(
        n762) );
  AOI22D1BWP12T U1553 ( .A1(r11[28]), .A2(n2755), .B1(n2754), .B2(r0[28]), 
        .ZN(n761) );
  AN3XD1BWP12T U1554 ( .A1(n763), .A2(n762), .A3(n761), .Z(n766) );
  AOI22D1BWP12T U1555 ( .A1(r5[28]), .A2(n2748), .B1(n2747), .B2(r10[28]), 
        .ZN(n765) );
  AOI22D1BWP12T U1556 ( .A1(r7[28]), .A2(n2750), .B1(n2749), .B2(r2[28]), .ZN(
        n764) );
  ND4D1BWP12T U1557 ( .A1(n767), .A2(n766), .A3(n765), .A4(n764), .ZN(
        regB_out[28]) );
  AOI22D0BWP12T U1558 ( .A1(r8[3]), .A2(n1382), .B1(n1381), .B2(r4[3]), .ZN(
        n770) );
  AOI22D0BWP12T U1559 ( .A1(n[2965]), .A2(n1384), .B1(n1383), .B2(r10[3]), 
        .ZN(n769) );
  CKND2D1BWP12T U1560 ( .A1(n770), .A2(n769), .ZN(n779) );
  AOI22D0BWP12T U1561 ( .A1(r7[3]), .A2(n1388), .B1(n1387), .B2(r5[3]), .ZN(
        n774) );
  AOI22D0BWP12T U1562 ( .A1(lr[3]), .A2(n1390), .B1(n1389), .B2(r9[3]), .ZN(
        n773) );
  AOI22D0BWP12T U1563 ( .A1(r6[3]), .A2(n1392), .B1(n1391), .B2(r11[3]), .ZN(
        n772) );
  CKND2D0BWP12T U1564 ( .A1(n1393), .A2(r12[3]), .ZN(n771) );
  ND4D1BWP12T U1565 ( .A1(n774), .A2(n773), .A3(n772), .A4(n771), .ZN(n778) );
  AOI22D0BWP12T U1566 ( .A1(r3[3]), .A2(n1399), .B1(n1398), .B2(r2[3]), .ZN(
        n776) );
  AOI22D0BWP12T U1567 ( .A1(n1401), .A2(r0[3]), .B1(pc_out[3]), .B2(n1400), 
        .ZN(n775) );
  OAI211D0BWP12T U1568 ( .A1(n929), .A2(n1404), .B(n776), .C(n775), .ZN(n777)
         );
  OA31D0BWP12T U1569 ( .A1(n779), .A2(n778), .A3(n777), .B(n1405), .Z(
        regD_out[3]) );
  AO222D0BWP12T U1570 ( .A1(write1_in[23]), .A2(n1620), .B1(write2_in[23]), 
        .B2(n1625), .C1(n1622), .C2(tmp1[23]), .Z(n2160) );
  AO222D0BWP12T U1571 ( .A1(write1_in[23]), .A2(n1614), .B1(write2_in[23]), 
        .B2(n1617), .C1(n1521), .C2(n[2945]), .Z(spin[23]) );
  AO222D0BWP12T U1572 ( .A1(write1_in[23]), .A2(n1555), .B1(write2_in[23]), 
        .B2(n1558), .C1(n1519), .C2(r6[23]), .Z(n2448) );
  AO222D0BWP12T U1573 ( .A1(write1_in[23]), .A2(n1607), .B1(write2_in[23]), 
        .B2(n1609), .C1(n1608), .C2(lr[23]), .Z(n2224) );
  AO222D0BWP12T U1574 ( .A1(write1_in[23]), .A2(n1597), .B1(write2_in[23]), 
        .B2(n1599), .C1(n1598), .C2(r12[23]), .Z(n2256) );
  AO222D0BWP12T U1575 ( .A1(write1_in[23]), .A2(n1567), .B1(write2_in[23]), 
        .B2(n1570), .C1(n1505), .C2(r7[23]), .Z(n2416) );
  AO222D0BWP12T U1576 ( .A1(write1_in[23]), .A2(n1549), .B1(write2_in[23]), 
        .B2(n1552), .C1(n1506), .C2(r0[23]), .Z(n2640) );
  AO222D0BWP12T U1577 ( .A1(n1591), .A2(n1471), .B1(n1507), .B2(r9[14]), .C1(
        write2_in[14]), .C2(n1594), .Z(n2343) );
  AO222D0BWP12T U1578 ( .A1(n1607), .A2(n1471), .B1(n1608), .B2(lr[14]), .C1(
        write2_in[14]), .C2(n1609), .Z(n2215) );
  AO222D0BWP12T U1579 ( .A1(n1555), .A2(n1471), .B1(n1519), .B2(r6[14]), .C1(
        write2_in[14]), .C2(n1558), .Z(n2439) );
  AO222D0BWP12T U1580 ( .A1(n1614), .A2(n1471), .B1(n1521), .B2(n[2954]), .C1(
        write2_in[14]), .C2(n1617), .Z(spin[14]) );
  AO222D0BWP12T U1581 ( .A1(n1620), .A2(n1471), .B1(n1625), .B2(write2_in[14]), 
        .C1(n1622), .C2(tmp1[14]), .Z(n2151) );
  AOI22D1BWP12T U1582 ( .A1(n2808), .A2(r11[27]), .B1(n2807), .B2(n[2941]), 
        .ZN(n783) );
  AOI22D1BWP12T U1583 ( .A1(r3[27]), .A2(n2810), .B1(n2809), .B2(r5[27]), .ZN(
        n782) );
  AOI22D1BWP12T U1584 ( .A1(n2812), .A2(r7[27]), .B1(n2776), .B2(pc_out[27]), 
        .ZN(n781) );
  AOI22D1BWP12T U1585 ( .A1(n2814), .A2(r1[27]), .B1(n2708), .B2(r12[27]), 
        .ZN(n780) );
  AN4XD1BWP12T U1586 ( .A1(n783), .A2(n782), .A3(n781), .A4(n780), .Z(n790) );
  INVD1BWP12T U1587 ( .I(r2[27]), .ZN(n1483) );
  AOI22D1BWP12T U1588 ( .A1(r4[27]), .A2(n2791), .B1(n2795), .B2(r0[27]), .ZN(
        n785) );
  AOI22D1BWP12T U1589 ( .A1(tmp1[27]), .A2(n2820), .B1(n2819), .B2(r9[27]), 
        .ZN(n784) );
  OA211D1BWP12T U1590 ( .A1(n1483), .A2(n2789), .B(n785), .C(n784), .Z(n789)
         );
  AOI22D1BWP12T U1591 ( .A1(n2892), .A2(r8[27]), .B1(n2891), .B2(lr[27]), .ZN(
        n787) );
  AOI22D1BWP12T U1592 ( .A1(r6[27]), .A2(n2894), .B1(n2893), .B2(r10[27]), 
        .ZN(n786) );
  AN2XD1BWP12T U1593 ( .A1(n787), .A2(n786), .Z(n788) );
  AO222D0BWP12T U1594 ( .A1(n1620), .A2(write1_in[7]), .B1(n1625), .B2(
        write2_in[7]), .C1(n1622), .C2(tmp1[7]), .Z(n2144) );
  AO222D0BWP12T U1595 ( .A1(n1620), .A2(write1_in[4]), .B1(n1625), .B2(
        write2_in[4]), .C1(n1622), .C2(tmp1[4]), .Z(n2141) );
  ND2D1BWP12T U1596 ( .A1(n2708), .A2(r12[11]), .ZN(n793) );
  ND2D1BWP12T U1597 ( .A1(n2819), .A2(r9[11]), .ZN(n792) );
  OR2D0BWP12T U1598 ( .A1(n2872), .A2(n1929), .Z(n791) );
  AN3XD1BWP12T U1599 ( .A1(n793), .A2(n792), .A3(n791), .Z(n813) );
  ND2D1BWP12T U1600 ( .A1(n795), .A2(n794), .ZN(n803) );
  NR2D1BWP12T U1601 ( .A1(n2860), .A2(n1931), .ZN(n796) );
  AOI21D1BWP12T U1602 ( .A1(n2809), .A2(r5[11]), .B(n796), .ZN(n801) );
  OAI22D1BWP12T U1603 ( .A1(n2789), .A2(n1922), .B1(n797), .B2(n2864), .ZN(
        n799) );
  INVD1BWP12T U1604 ( .I(tmp1[11]), .ZN(n1919) );
  NR2D1BWP12T U1605 ( .A1(n2880), .A2(n1919), .ZN(n798) );
  NR2D1BWP12T U1606 ( .A1(n799), .A2(n798), .ZN(n800) );
  ND2D1BWP12T U1607 ( .A1(n801), .A2(n800), .ZN(n802) );
  NR2XD0BWP12T U1608 ( .A1(n803), .A2(n802), .ZN(n812) );
  INR2D1BWP12T U1609 ( .A1(r0[11]), .B1(n2884), .ZN(n804) );
  INVD1BWP12T U1610 ( .I(n804), .ZN(n810) );
  AN2D1BWP12T U1611 ( .A1(n2791), .A2(r4[11]), .Z(n809) );
  NR2D1BWP12T U1612 ( .A1(n2868), .A2(n1923), .ZN(n805) );
  AOI21D1BWP12T U1613 ( .A1(n2776), .A2(pc_out[11]), .B(n805), .ZN(n807) );
  CKND2D1BWP12T U1614 ( .A1(n2807), .A2(n[2957]), .ZN(n806) );
  ND2D1BWP12T U1615 ( .A1(n807), .A2(n806), .ZN(n808) );
  INR3D2BWP12T U1616 ( .A1(n810), .B1(n809), .B2(n808), .ZN(n811) );
  ND3D2BWP12T U1617 ( .A1(n813), .A2(n812), .A3(n811), .ZN(regA_out[11]) );
  AO222D0BWP12T U1618 ( .A1(n1620), .A2(write1_in[13]), .B1(n1625), .B2(
        write2_in[13]), .C1(n1622), .C2(tmp1[13]), .Z(n2150) );
  AO222D0BWP12T U1619 ( .A1(n1614), .A2(write1_in[13]), .B1(n1521), .B2(
        n[2955]), .C1(write2_in[13]), .C2(n1617), .Z(spin[13]) );
  AO222D0BWP12T U1620 ( .A1(n1585), .A2(write1_in[13]), .B1(n1517), .B2(r1[13]), .C1(write2_in[13]), .C2(n1588), .Z(n2598) );
  AO222D0BWP12T U1621 ( .A1(n1555), .A2(write1_in[13]), .B1(n1519), .B2(r6[13]), .C1(write2_in[13]), .C2(n1558), .Z(n2438) );
  AO222D0BWP12T U1622 ( .A1(n1591), .A2(write1_in[13]), .B1(n1507), .B2(r9[13]), .C1(write2_in[13]), .C2(n1594), .Z(n2342) );
  AO222D0BWP12T U1623 ( .A1(n1579), .A2(write1_in[13]), .B1(n1518), .B2(r4[13]), .C1(write2_in[13]), .C2(n1582), .Z(n2502) );
  AO222D0BWP12T U1624 ( .A1(n1602), .A2(write1_in[13]), .B1(n1603), .B2(r8[13]), .C1(write2_in[13]), .C2(n1604), .Z(n2374) );
  AO222D0BWP12T U1625 ( .A1(n1597), .A2(write1_in[13]), .B1(n1598), .B2(
        r12[13]), .C1(write2_in[13]), .C2(n1599), .Z(n2246) );
  AO222D0BWP12T U1626 ( .A1(n1549), .A2(write1_in[13]), .B1(n1506), .B2(r0[13]), .C1(write2_in[13]), .C2(n1552), .Z(n2630) );
  AO222D0BWP12T U1627 ( .A1(n1607), .A2(write1_in[13]), .B1(n1608), .B2(lr[13]), .C1(write2_in[13]), .C2(n1609), .Z(n2214) );
  AO222D0BWP12T U1628 ( .A1(n1567), .A2(write1_in[13]), .B1(n1505), .B2(r7[13]), .C1(write2_in[13]), .C2(n1570), .Z(n2406) );
  INVD1BWP12T U1629 ( .I(r2[30]), .ZN(n817) );
  CKND0BWP12T U1630 ( .I(n2887), .ZN(n814) );
  AOI22D1BWP12T U1631 ( .A1(n814), .A2(r4[30]), .B1(n2795), .B2(r0[30]), .ZN(
        n816) );
  AOI22D1BWP12T U1632 ( .A1(tmp1[30]), .A2(n2820), .B1(n2819), .B2(r9[30]), 
        .ZN(n815) );
  OA211D1BWP12T U1633 ( .A1(n817), .A2(n2789), .B(n816), .C(n815), .Z(n823) );
  AOI22D1BWP12T U1634 ( .A1(r7[30]), .A2(n2812), .B1(n2776), .B2(pc_out[30]), 
        .ZN(n819) );
  AOI22D1BWP12T U1635 ( .A1(n2814), .A2(r1[30]), .B1(r12[30]), .B2(n2813), 
        .ZN(n818) );
  AOI22D1BWP12T U1636 ( .A1(n2892), .A2(r8[30]), .B1(n2891), .B2(lr[30]), .ZN(
        n821) );
  AOI22D1BWP12T U1637 ( .A1(n2894), .A2(r6[30]), .B1(n2893), .B2(r10[30]), 
        .ZN(n820) );
  AOI22D1BWP12T U1638 ( .A1(n2808), .A2(r11[19]), .B1(n2807), .B2(n[2949]), 
        .ZN(n827) );
  AOI22D1BWP12T U1639 ( .A1(n2812), .A2(r7[19]), .B1(n2811), .B2(pc_out[19]), 
        .ZN(n825) );
  AN4XD1BWP12T U1640 ( .A1(n827), .A2(n826), .A3(n825), .A4(n824), .Z(n836) );
  INVD1BWP12T U1641 ( .I(r9[19]), .ZN(n961) );
  INVD1BWP12T U1642 ( .I(tmp1[19]), .ZN(n828) );
  OAI22D1BWP12T U1643 ( .A1(n2883), .A2(n961), .B1(n828), .B2(n2880), .ZN(n832) );
  INVD1BWP12T U1644 ( .I(r4[19]), .ZN(n830) );
  INVD1BWP12T U1645 ( .I(r0[19]), .ZN(n829) );
  OAI22D1BWP12T U1646 ( .A1(n2887), .A2(n830), .B1(n829), .B2(n2884), .ZN(n831) );
  RCAOI211D0BWP12T U1647 ( .A1(r2[19]), .A2(n2890), .B(n832), .C(n831), .ZN(
        n835) );
  AOI22D1BWP12T U1648 ( .A1(n2892), .A2(r8[19]), .B1(n2891), .B2(lr[19]), .ZN(
        n834) );
  AOI22D1BWP12T U1649 ( .A1(r6[19]), .A2(n2894), .B1(n2893), .B2(r10[19]), 
        .ZN(n833) );
  NR2D1BWP12T U1650 ( .A1(n2868), .A2(n837), .ZN(n838) );
  AOI21D1BWP12T U1651 ( .A1(n2776), .A2(pc_out[1]), .B(n838), .ZN(n848) );
  AOI21D1BWP12T U1652 ( .A1(n2809), .A2(r5[1]), .B(n841), .ZN(n845) );
  NR2D1BWP12T U1653 ( .A1(n2872), .A2(n842), .ZN(n843) );
  AOI21D1BWP12T U1654 ( .A1(n2708), .A2(r12[1]), .B(n843), .ZN(n844) );
  ND2D1BWP12T U1655 ( .A1(n845), .A2(n844), .ZN(n846) );
  INR3D0BWP12T U1656 ( .A1(n848), .B1(n847), .B2(n846), .ZN(n866) );
  NR2D1BWP12T U1657 ( .A1(n2880), .A2(n850), .ZN(n851) );
  RCIAO21D0BWP12T U1658 ( .A1(n2883), .A2(n852), .B(n851), .ZN(n853) );
  IOA21D1BWP12T U1659 ( .A1(n2890), .A2(r2[1]), .B(n853), .ZN(n863) );
  TPND2D0BWP12T U1660 ( .A1(n854), .A2(r8[1]), .ZN(n855) );
  NR2D1BWP12T U1661 ( .A1(n856), .A2(n855), .ZN(n857) );
  AOI21D1BWP12T U1662 ( .A1(n2891), .A2(lr[1]), .B(n857), .ZN(n861) );
  NR2D1BWP12T U1663 ( .A1(n2826), .A2(n858), .ZN(n859) );
  AOI21D1BWP12T U1664 ( .A1(n2893), .A2(r10[1]), .B(n859), .ZN(n860) );
  ND2D1BWP12T U1665 ( .A1(n861), .A2(n860), .ZN(n862) );
  INR3D0BWP12T U1666 ( .A1(n864), .B1(n863), .B2(n862), .ZN(n865) );
  TPND2D1BWP12T U1667 ( .A1(n866), .A2(n865), .ZN(regA_out[1]) );
  CKND2D1BWP12T U1668 ( .A1(n2819), .A2(r9[3]), .ZN(n869) );
  CKND2D1BWP12T U1669 ( .A1(n2791), .A2(r4[3]), .ZN(n868) );
  ND3D1BWP12T U1670 ( .A1(n62), .A2(n869), .A3(n868), .ZN(n874) );
  NR2D1BWP12T U1671 ( .A1(n2822), .A2(n870), .ZN(n873) );
  OAI22D1BWP12T U1672 ( .A1(n2829), .A2(n871), .B1(n2871), .B2(n939), .ZN(n872) );
  NR3D1BWP12T U1673 ( .A1(n874), .A2(n873), .A3(n872), .ZN(n888) );
  NR2D1BWP12T U1674 ( .A1(n2860), .A2(n933), .ZN(n875) );
  AOI21D1BWP12T U1675 ( .A1(n2809), .A2(r5[3]), .B(n875), .ZN(n878) );
  NR2D1BWP12T U1676 ( .A1(n2872), .A2(n929), .ZN(n876) );
  AOI21D1BWP12T U1677 ( .A1(n2813), .A2(r12[3]), .B(n876), .ZN(n877) );
  AOI21D1BWP12T U1678 ( .A1(lr[3]), .A2(n2891), .B(n879), .ZN(n882) );
  OAI22D1BWP12T U1679 ( .A1(n2884), .A2(n934), .B1(n2789), .B2(n932), .ZN(n881) );
  NR2D1BWP12T U1680 ( .A1(n2826), .A2(n931), .ZN(n880) );
  ND2D1BWP12T U1681 ( .A1(n2807), .A2(n[2965]), .ZN(n883) );
  OA21D1BWP12T U1682 ( .A1(n2864), .A2(n884), .B(n883), .Z(n885) );
  AO222D0BWP12T U1683 ( .A1(write1_in[17]), .A2(n1620), .B1(write2_in[17]), 
        .B2(n1625), .C1(n1622), .C2(tmp1[17]), .Z(n2154) );
  AOI22D1BWP12T U1684 ( .A1(tmp1[19]), .A2(n2746), .B1(n2730), .B2(
        immediate2_in[19]), .ZN(n895) );
  AOI22D1BWP12T U1685 ( .A1(r5[19]), .A2(n2748), .B1(n2747), .B2(r10[19]), 
        .ZN(n890) );
  AOI22D1BWP12T U1686 ( .A1(r7[19]), .A2(n2750), .B1(n2749), .B2(r2[19]), .ZN(
        n889) );
  ND2D1BWP12T U1687 ( .A1(n890), .A2(n889), .ZN(n894) );
  AOI22D1BWP12T U1688 ( .A1(r9[19]), .A2(n105), .B1(n2753), .B2(r4[19]), .ZN(
        n892) );
  AOI22D1BWP12T U1689 ( .A1(r11[19]), .A2(n2755), .B1(n2733), .B2(r0[19]), 
        .ZN(n891) );
  ND2D1BWP12T U1690 ( .A1(n892), .A2(n891), .ZN(n893) );
  INR3XD0BWP12T U1691 ( .A1(n895), .B1(n894), .B2(n893), .ZN(n901) );
  AOI22D1BWP12T U1692 ( .A1(r1[19]), .A2(n118), .B1(n2761), .B2(r12[19]), .ZN(
        n899) );
  AOI22D1BWP12T U1693 ( .A1(r3[19]), .A2(n2763), .B1(n2762), .B2(lr[19]), .ZN(
        n898) );
  AOI22D1BWP12T U1694 ( .A1(r8[19]), .A2(n2765), .B1(n2764), .B2(n[2949]), 
        .ZN(n897) );
  AOI22D1BWP12T U1695 ( .A1(pc_out[19]), .A2(n2767), .B1(n2766), .B2(r6[19]), 
        .ZN(n896) );
  AN4XD1BWP12T U1696 ( .A1(n899), .A2(n898), .A3(n897), .A4(n896), .Z(n900) );
  AO222D1BWP12T U1697 ( .A1(write1_in[27]), .A2(n1591), .B1(write2_in[27]), 
        .B2(n1594), .C1(n1507), .C2(r9[27]), .Z(n2356) );
  AN2XD2BWP12T U1698 ( .A1(next_cpsr_in[3]), .A2(n902), .Z(cpsrin[3]) );
  AN2XD2BWP12T U1699 ( .A1(next_cpsr_in[1]), .A2(n902), .Z(cpsrin[1]) );
  AN2XD2BWP12T U1700 ( .A1(next_cpsr_in[0]), .A2(n902), .Z(cpsrin[0]) );
  IND2D1BWP12T U1701 ( .A1(readC_sel[0]), .B1(readC_sel[1]), .ZN(n919) );
  ND3D1BWP12T U1702 ( .A1(readC_sel[2]), .A2(readC_sel[3]), .A3(n1295), .ZN(
        n921) );
  NR2D1BWP12T U1703 ( .A1(n919), .A2(n921), .ZN(n1319) );
  CKND0BWP12T U1704 ( .I(readC_sel[3]), .ZN(n904) );
  TPND2D0BWP12T U1705 ( .A1(readC_sel[2]), .A2(n904), .ZN(n906) );
  ND2D1BWP12T U1706 ( .A1(readC_sel[1]), .A2(readC_sel[0]), .ZN(n917) );
  OR2XD1BWP12T U1707 ( .A1(n906), .A2(n917), .Z(n1302) );
  OR2XD1BWP12T U1708 ( .A1(readC_sel[0]), .A2(readC_sel[1]), .Z(n920) );
  OR2XD1BWP12T U1709 ( .A1(n906), .A2(n920), .Z(n1301) );
  OAI22D0BWP12T U1710 ( .A1(n1881), .A2(n1302), .B1(n1301), .B2(n903), .ZN(
        n912) );
  IND2D1BWP12T U1711 ( .A1(readC_sel[1]), .B1(readC_sel[0]), .ZN(n922) );
  OR2XD1BWP12T U1712 ( .A1(n922), .A2(n906), .Z(n1304) );
  INVD1BWP12T U1713 ( .I(readC_sel[2]), .ZN(n916) );
  CKND2D1BWP12T U1714 ( .A1(n916), .A2(n904), .ZN(n908) );
  OR2XD1BWP12T U1715 ( .A1(n922), .A2(n908), .Z(n1303) );
  OAI22D0BWP12T U1716 ( .A1(n905), .A2(n1304), .B1(n1303), .B2(n1885), .ZN(
        n911) );
  OR2XD1BWP12T U1717 ( .A1(n919), .A2(n908), .Z(n1307) );
  OR2XD1BWP12T U1718 ( .A1(n906), .A2(n919), .Z(n1306) );
  OAI22D0BWP12T U1719 ( .A1(n1307), .A2(n907), .B1(n1306), .B2(n1874), .ZN(
        n910) );
  OR2XD1BWP12T U1720 ( .A1(n908), .A2(n920), .Z(n1309) );
  OR2XD1BWP12T U1721 ( .A1(n908), .A2(n917), .Z(n1308) );
  OAI22D0BWP12T U1722 ( .A1(n1877), .A2(n1309), .B1(n1308), .B2(n1884), .ZN(
        n909) );
  NR4D0BWP12T U1723 ( .A1(n912), .A2(n911), .A3(n910), .A4(n909), .ZN(n914) );
  OR2XD1BWP12T U1724 ( .A1(n917), .A2(n921), .Z(n1268) );
  OAI22D0BWP12T U1725 ( .A1(n914), .A2(readC_sel[4]), .B1(n1268), .B2(n913), 
        .ZN(n915) );
  AOI21D0BWP12T U1726 ( .A1(lr[2]), .A2(n1319), .B(n915), .ZN(n926) );
  ND3D1BWP12T U1727 ( .A1(readC_sel[3]), .A2(n1295), .A3(n916), .ZN(n918) );
  OR2XD1BWP12T U1728 ( .A1(n922), .A2(n918), .Z(n1170) );
  OR2XD1BWP12T U1729 ( .A1(n917), .A2(n918), .Z(n1287) );
  AOI22D0BWP12T U1730 ( .A1(r9[2]), .A2(n1321), .B1(n1320), .B2(r11[2]), .ZN(
        n925) );
  NR2D1BWP12T U1731 ( .A1(n920), .A2(n918), .ZN(n1323) );
  OR2XD1BWP12T U1732 ( .A1(n919), .A2(n918), .Z(n1249) );
  AOI22D0BWP12T U1733 ( .A1(r8[2]), .A2(n1323), .B1(n1322), .B2(r10[2]), .ZN(
        n924) );
  NR2D1BWP12T U1734 ( .A1(n920), .A2(n921), .ZN(n1325) );
  NR2D1BWP12T U1735 ( .A1(n922), .A2(n921), .ZN(n1168) );
  AOI22D0BWP12T U1736 ( .A1(r12[2]), .A2(n1325), .B1(n1168), .B2(n[2966]), 
        .ZN(n923) );
  ND4D1BWP12T U1737 ( .A1(n926), .A2(n925), .A3(n924), .A4(n923), .ZN(
        regC_out[2]) );
  OAI22D0BWP12T U1738 ( .A1(n928), .A2(n1302), .B1(n1301), .B2(n927), .ZN(n938) );
  OAI22D0BWP12T U1739 ( .A1(n930), .A2(n1304), .B1(n1303), .B2(n929), .ZN(n937) );
  OAI22D0BWP12T U1740 ( .A1(n1307), .A2(n932), .B1(n1306), .B2(n931), .ZN(n936) );
  OAI22D0BWP12T U1741 ( .A1(n934), .A2(n1309), .B1(n1308), .B2(n933), .ZN(n935) );
  NR4D0BWP12T U1742 ( .A1(n938), .A2(n937), .A3(n936), .A4(n935), .ZN(n940) );
  OAI22D0BWP12T U1743 ( .A1(n940), .A2(readC_sel[4]), .B1(n1268), .B2(n939), 
        .ZN(n941) );
  AOI21D0BWP12T U1744 ( .A1(lr[3]), .A2(n1319), .B(n941), .ZN(n945) );
  AOI22D0BWP12T U1745 ( .A1(r9[3]), .A2(n1321), .B1(n1320), .B2(r11[3]), .ZN(
        n944) );
  AOI22D0BWP12T U1746 ( .A1(r8[3]), .A2(n1323), .B1(n1322), .B2(r10[3]), .ZN(
        n943) );
  AOI22D0BWP12T U1747 ( .A1(r12[3]), .A2(n1325), .B1(n1168), .B2(n[2965]), 
        .ZN(n942) );
  ND4D1BWP12T U1748 ( .A1(n945), .A2(n944), .A3(n943), .A4(n942), .ZN(
        regC_out[3]) );
  INVD1BWP12T U1749 ( .I(n1268), .ZN(n1324) );
  AOI22D0BWP12T U1750 ( .A1(r12[31]), .A2(n1325), .B1(n1324), .B2(pc_out[31]), 
        .ZN(n956) );
  AOI22D0BWP12T U1751 ( .A1(lr[31]), .A2(n1319), .B1(n1168), .B2(n[2937]), 
        .ZN(n955) );
  AOI22D0BWP12T U1752 ( .A1(r8[31]), .A2(n1323), .B1(n1320), .B2(r11[31]), 
        .ZN(n954) );
  AOI22D0BWP12T U1753 ( .A1(r7[31]), .A2(n1276), .B1(n1275), .B2(r4[31]), .ZN(
        n949) );
  AOI22D0BWP12T U1754 ( .A1(r2[31]), .A2(n1278), .B1(n1277), .B2(r6[31]), .ZN(
        n948) );
  AOI22D0BWP12T U1755 ( .A1(r5[31]), .A2(n1280), .B1(n1279), .B2(r1[31]), .ZN(
        n947) );
  AOI22D0BWP12T U1756 ( .A1(r0[31]), .A2(n1282), .B1(n1281), .B2(r3[31]), .ZN(
        n946) );
  ND4D1BWP12T U1757 ( .A1(n949), .A2(n948), .A3(n947), .A4(n946), .ZN(n952) );
  CKND0BWP12T U1758 ( .I(r9[31]), .ZN(n950) );
  CKND0BWP12T U1759 ( .I(r10[31]), .ZN(n1525) );
  OAI22D0BWP12T U1760 ( .A1(n1170), .A2(n950), .B1(n1525), .B2(n1249), .ZN(
        n951) );
  AOI21D0BWP12T U1761 ( .A1(n952), .A2(n1295), .B(n951), .ZN(n953) );
  ND4D1BWP12T U1762 ( .A1(n956), .A2(n955), .A3(n954), .A4(n953), .ZN(
        regC_out[31]) );
  AOI22D0BWP12T U1763 ( .A1(pc_out[19]), .A2(n1324), .B1(n1323), .B2(r8[19]), 
        .ZN(n968) );
  AOI22D0BWP12T U1764 ( .A1(n[2949]), .A2(n1168), .B1(n1325), .B2(r12[19]), 
        .ZN(n967) );
  AOI22D0BWP12T U1765 ( .A1(r10[19]), .A2(n1322), .B1(n1320), .B2(r11[19]), 
        .ZN(n966) );
  AOI22D0BWP12T U1766 ( .A1(r7[19]), .A2(n1276), .B1(n1275), .B2(r4[19]), .ZN(
        n960) );
  AOI22D0BWP12T U1767 ( .A1(r2[19]), .A2(n1278), .B1(n1277), .B2(r6[19]), .ZN(
        n959) );
  AOI22D0BWP12T U1768 ( .A1(r5[19]), .A2(n1280), .B1(n1279), .B2(r1[19]), .ZN(
        n958) );
  AOI22D0BWP12T U1769 ( .A1(r0[19]), .A2(n1282), .B1(n1281), .B2(r3[19]), .ZN(
        n957) );
  ND4D1BWP12T U1770 ( .A1(n960), .A2(n959), .A3(n958), .A4(n957), .ZN(n964) );
  INVD1BWP12T U1771 ( .I(n1319), .ZN(n1289) );
  CKND0BWP12T U1772 ( .I(lr[19]), .ZN(n962) );
  OAI22D0BWP12T U1773 ( .A1(n1289), .A2(n962), .B1(n961), .B2(n1170), .ZN(n963) );
  AOI21D0BWP12T U1774 ( .A1(n964), .A2(n1295), .B(n963), .ZN(n965) );
  ND4D1BWP12T U1775 ( .A1(n968), .A2(n967), .A3(n966), .A4(n965), .ZN(
        regC_out[19]) );
  AOI22D0BWP12T U1776 ( .A1(pc_out[0]), .A2(n1324), .B1(n1323), .B2(r8[0]), 
        .ZN(n978) );
  AOI22D0BWP12T U1777 ( .A1(n[2968]), .A2(n1168), .B1(n1325), .B2(r12[0]), 
        .ZN(n977) );
  AOI22D0BWP12T U1778 ( .A1(r9[0]), .A2(n1321), .B1(n1320), .B2(r11[0]), .ZN(
        n976) );
  AOI22D0BWP12T U1779 ( .A1(r7[0]), .A2(n1276), .B1(n1275), .B2(r4[0]), .ZN(
        n972) );
  AOI22D0BWP12T U1780 ( .A1(r2[0]), .A2(n1278), .B1(n1277), .B2(r6[0]), .ZN(
        n971) );
  AOI22D0BWP12T U1781 ( .A1(r5[0]), .A2(n1280), .B1(n1279), .B2(r1[0]), .ZN(
        n970) );
  AOI22D0BWP12T U1782 ( .A1(r0[0]), .A2(n1282), .B1(n1281), .B2(r3[0]), .ZN(
        n969) );
  ND4D1BWP12T U1783 ( .A1(n972), .A2(n971), .A3(n970), .A4(n969), .ZN(n974) );
  INVD1BWP12T U1784 ( .I(lr[0]), .ZN(n1828) );
  INVD1BWP12T U1785 ( .I(r10[0]), .ZN(n1830) );
  OAI22D0BWP12T U1786 ( .A1(n1289), .A2(n1828), .B1(n1830), .B2(n1249), .ZN(
        n973) );
  AOI21D0BWP12T U1787 ( .A1(n974), .A2(n1295), .B(n973), .ZN(n975) );
  ND4D1BWP12T U1788 ( .A1(n978), .A2(n977), .A3(n976), .A4(n975), .ZN(
        regC_out[0]) );
  AOI22D0BWP12T U1789 ( .A1(pc_out[5]), .A2(n1324), .B1(n1323), .B2(r8[5]), 
        .ZN(n988) );
  AOI22D0BWP12T U1790 ( .A1(r12[5]), .A2(n1325), .B1(n1168), .B2(n[2963]), 
        .ZN(n987) );
  AOI22D0BWP12T U1791 ( .A1(r10[5]), .A2(n1322), .B1(n1320), .B2(r11[5]), .ZN(
        n986) );
  AOI22D0BWP12T U1792 ( .A1(r7[5]), .A2(n1276), .B1(n1275), .B2(r4[5]), .ZN(
        n982) );
  AOI22D0BWP12T U1793 ( .A1(r2[5]), .A2(n1278), .B1(n1277), .B2(r6[5]), .ZN(
        n981) );
  AOI22D0BWP12T U1794 ( .A1(r5[5]), .A2(n1280), .B1(n1279), .B2(r1[5]), .ZN(
        n980) );
  AOI22D0BWP12T U1795 ( .A1(r0[5]), .A2(n1282), .B1(n1281), .B2(r3[5]), .ZN(
        n979) );
  ND4D1BWP12T U1796 ( .A1(n982), .A2(n981), .A3(n980), .A4(n979), .ZN(n984) );
  OAI22D0BWP12T U1797 ( .A1(n1289), .A2(n2129), .B1(n2121), .B2(n1170), .ZN(
        n983) );
  AOI21D0BWP12T U1798 ( .A1(n984), .A2(n1295), .B(n983), .ZN(n985) );
  ND4D1BWP12T U1799 ( .A1(n988), .A2(n987), .A3(n986), .A4(n985), .ZN(
        regC_out[5]) );
  AOI22D0BWP12T U1800 ( .A1(r8[4]), .A2(n1323), .B1(n1322), .B2(r10[4]), .ZN(
        n998) );
  AOI22D0BWP12T U1801 ( .A1(r12[4]), .A2(n1325), .B1(n1168), .B2(n[2964]), 
        .ZN(n997) );
  AOI22D0BWP12T U1802 ( .A1(r9[4]), .A2(n1321), .B1(n1320), .B2(r11[4]), .ZN(
        n996) );
  AOI22D0BWP12T U1803 ( .A1(r7[4]), .A2(n1276), .B1(n1275), .B2(r4[4]), .ZN(
        n992) );
  AOI22D0BWP12T U1804 ( .A1(r2[4]), .A2(n1278), .B1(n1277), .B2(r6[4]), .ZN(
        n991) );
  AOI22D0BWP12T U1805 ( .A1(r5[4]), .A2(n1280), .B1(n1279), .B2(r1[4]), .ZN(
        n990) );
  AOI22D0BWP12T U1806 ( .A1(r0[4]), .A2(n1282), .B1(n1281), .B2(r3[4]), .ZN(
        n989) );
  ND4D1BWP12T U1807 ( .A1(n992), .A2(n991), .A3(n990), .A4(n989), .ZN(n994) );
  INVD1BWP12T U1808 ( .I(pc_out[4]), .ZN(n2022) );
  OAI22D0BWP12T U1809 ( .A1(n2022), .A2(n1268), .B1(n1289), .B2(n2017), .ZN(
        n993) );
  AOI21D0BWP12T U1810 ( .A1(n994), .A2(n1295), .B(n993), .ZN(n995) );
  ND4D1BWP12T U1811 ( .A1(n998), .A2(n997), .A3(n996), .A4(n995), .ZN(
        regC_out[4]) );
  AOI22D0BWP12T U1812 ( .A1(r7[13]), .A2(n1276), .B1(n1275), .B2(r4[13]), .ZN(
        n1002) );
  AOI22D0BWP12T U1813 ( .A1(r2[13]), .A2(n1278), .B1(n1277), .B2(r6[13]), .ZN(
        n1001) );
  AOI22D0BWP12T U1814 ( .A1(r5[13]), .A2(n1280), .B1(n1279), .B2(r1[13]), .ZN(
        n1000) );
  AOI22D0BWP12T U1815 ( .A1(r0[13]), .A2(n1282), .B1(n1281), .B2(r3[13]), .ZN(
        n999) );
  ND4D1BWP12T U1816 ( .A1(n1002), .A2(n1001), .A3(n1000), .A4(n999), .ZN(n1003) );
  MOAI22D0BWP12T U1817 ( .A1(n1289), .A2(n1004), .B1(n1003), .B2(n1295), .ZN(
        n1005) );
  AOI21D0BWP12T U1818 ( .A1(n[2955]), .A2(n1168), .B(n1005), .ZN(n1009) );
  AOI22D0BWP12T U1819 ( .A1(r10[13]), .A2(n1322), .B1(n1320), .B2(r11[13]), 
        .ZN(n1008) );
  AOI22D0BWP12T U1820 ( .A1(r8[13]), .A2(n1323), .B1(n1321), .B2(r9[13]), .ZN(
        n1007) );
  AOI22D0BWP12T U1821 ( .A1(r12[13]), .A2(n1325), .B1(n1324), .B2(pc_out[13]), 
        .ZN(n1006) );
  ND4D1BWP12T U1822 ( .A1(n1009), .A2(n1008), .A3(n1007), .A4(n1006), .ZN(
        regC_out[13]) );
  AOI22D0BWP12T U1823 ( .A1(r7[21]), .A2(n1276), .B1(n1275), .B2(r4[21]), .ZN(
        n1013) );
  AOI22D0BWP12T U1824 ( .A1(r2[21]), .A2(n1278), .B1(n1277), .B2(r6[21]), .ZN(
        n1012) );
  AOI22D0BWP12T U1825 ( .A1(r5[21]), .A2(n1280), .B1(n1279), .B2(r1[21]), .ZN(
        n1011) );
  AOI22D0BWP12T U1826 ( .A1(r0[21]), .A2(n1282), .B1(n1281), .B2(r3[21]), .ZN(
        n1010) );
  ND4D1BWP12T U1827 ( .A1(n1013), .A2(n1012), .A3(n1011), .A4(n1010), .ZN(
        n1019) );
  AOI22D0BWP12T U1828 ( .A1(r8[21]), .A2(n1323), .B1(n1321), .B2(r9[21]), .ZN(
        n1017) );
  AOI22D0BWP12T U1829 ( .A1(lr[21]), .A2(n1319), .B1(n1168), .B2(n[2947]), 
        .ZN(n1016) );
  AOI22D0BWP12T U1830 ( .A1(r12[21]), .A2(n1325), .B1(n1324), .B2(pc_out[21]), 
        .ZN(n1015) );
  AOI22D0BWP12T U1831 ( .A1(r10[21]), .A2(n1322), .B1(n1320), .B2(r11[21]), 
        .ZN(n1014) );
  ND4D1BWP12T U1832 ( .A1(n1017), .A2(n1016), .A3(n1015), .A4(n1014), .ZN(
        n1018) );
  AO21D1BWP12T U1833 ( .A1(n1295), .A2(n1019), .B(n1018), .Z(regC_out[21]) );
  CKND2D0BWP12T U1834 ( .A1(write1_in[1]), .A2(n1614), .ZN(n1021) );
  AOI21D0BWP12T U1835 ( .A1(n1521), .A2(n[2967]), .B(reset), .ZN(n1020) );
  OAI211D1BWP12T U1836 ( .A1(n1022), .A2(n1443), .B(n1021), .C(n1020), .ZN(
        spin[1]) );
  CKND2D0BWP12T U1837 ( .A1(write1_in[2]), .A2(n1614), .ZN(n1024) );
  AOI21D0BWP12T U1838 ( .A1(n1521), .A2(n[2966]), .B(reset), .ZN(n1023) );
  OAI211D1BWP12T U1839 ( .A1(n1025), .A2(n1443), .B(n1024), .C(n1023), .ZN(
        spin[2]) );
  CKND2D0BWP12T U1840 ( .A1(write1_in[5]), .A2(n1614), .ZN(n1027) );
  AOI21D0BWP12T U1841 ( .A1(n1521), .A2(n[2963]), .B(reset), .ZN(n1026) );
  OAI211D1BWP12T U1842 ( .A1(n1028), .A2(n1443), .B(n1027), .C(n1026), .ZN(
        spin[5]) );
  AOI22D0BWP12T U1843 ( .A1(r12[9]), .A2(n1325), .B1(n1324), .B2(pc_out[9]), 
        .ZN(n1040) );
  AOI22D0BWP12T U1844 ( .A1(lr[9]), .A2(n1319), .B1(n1168), .B2(n[2959]), .ZN(
        n1039) );
  AOI22D0BWP12T U1845 ( .A1(r10[9]), .A2(n1322), .B1(n1320), .B2(r11[9]), .ZN(
        n1038) );
  AOI22D0BWP12T U1846 ( .A1(r7[9]), .A2(n1276), .B1(n1275), .B2(r4[9]), .ZN(
        n1032) );
  AOI22D0BWP12T U1847 ( .A1(r2[9]), .A2(n1278), .B1(n1277), .B2(r6[9]), .ZN(
        n1031) );
  AOI22D0BWP12T U1848 ( .A1(r5[9]), .A2(n1280), .B1(n1279), .B2(r1[9]), .ZN(
        n1030) );
  AOI22D0BWP12T U1849 ( .A1(r0[9]), .A2(n1282), .B1(n1281), .B2(r3[9]), .ZN(
        n1029) );
  ND4D1BWP12T U1850 ( .A1(n1032), .A2(n1031), .A3(n1030), .A4(n1029), .ZN(
        n1036) );
  INVD1BWP12T U1851 ( .I(n1323), .ZN(n1291) );
  OAI22D0BWP12T U1852 ( .A1(n1291), .A2(n1034), .B1(n1033), .B2(n1170), .ZN(
        n1035) );
  AOI21D0BWP12T U1853 ( .A1(n1036), .A2(n1295), .B(n1035), .ZN(n1037) );
  ND4D1BWP12T U1854 ( .A1(n1040), .A2(n1039), .A3(n1038), .A4(n1037), .ZN(
        regC_out[9]) );
  INVD0BWP12T U1855 ( .I(pc_out[30]), .ZN(n2923) );
  INVD1BWP12T U1856 ( .I(n1325), .ZN(n1238) );
  AOI22D0BWP12T U1857 ( .A1(r12[25]), .A2(n1325), .B1(n1321), .B2(r9[25]), 
        .ZN(n1050) );
  AOI22D0BWP12T U1858 ( .A1(lr[25]), .A2(n1319), .B1(n1168), .B2(n[2943]), 
        .ZN(n1049) );
  AOI22D0BWP12T U1859 ( .A1(r10[25]), .A2(n1322), .B1(n1320), .B2(r11[25]), 
        .ZN(n1048) );
  AOI22D0BWP12T U1860 ( .A1(r7[25]), .A2(n1276), .B1(n1275), .B2(r4[25]), .ZN(
        n1044) );
  AOI22D0BWP12T U1861 ( .A1(r2[25]), .A2(n1278), .B1(n1277), .B2(r6[25]), .ZN(
        n1043) );
  AOI22D0BWP12T U1862 ( .A1(r5[25]), .A2(n1280), .B1(n1279), .B2(r1[25]), .ZN(
        n1042) );
  AOI22D0BWP12T U1863 ( .A1(r0[25]), .A2(n1282), .B1(n1281), .B2(r3[25]), .ZN(
        n1041) );
  ND4D1BWP12T U1864 ( .A1(n1044), .A2(n1043), .A3(n1042), .A4(n1041), .ZN(
        n1046) );
  CKND0BWP12T U1865 ( .I(pc_out[25]), .ZN(n1634) );
  INVD1BWP12T U1866 ( .I(r8[25]), .ZN(n2823) );
  OAI22D0BWP12T U1867 ( .A1(n1634), .A2(n1268), .B1(n1291), .B2(n2823), .ZN(
        n1045) );
  AOI21D0BWP12T U1868 ( .A1(n1046), .A2(n1295), .B(n1045), .ZN(n1047) );
  ND4D1BWP12T U1869 ( .A1(n1050), .A2(n1049), .A3(n1048), .A4(n1047), .ZN(
        regC_out[25]) );
  AOI22D0BWP12T U1870 ( .A1(pc_out[15]), .A2(n1324), .B1(n1322), .B2(r10[15]), 
        .ZN(n1062) );
  AOI22D0BWP12T U1871 ( .A1(n[2953]), .A2(n1168), .B1(n1325), .B2(r12[15]), 
        .ZN(n1061) );
  AOI22D0BWP12T U1872 ( .A1(r9[15]), .A2(n1321), .B1(n1320), .B2(r11[15]), 
        .ZN(n1060) );
  AOI22D0BWP12T U1873 ( .A1(r7[15]), .A2(n1276), .B1(n1275), .B2(r4[15]), .ZN(
        n1054) );
  AOI22D0BWP12T U1874 ( .A1(r2[15]), .A2(n1278), .B1(n1277), .B2(r6[15]), .ZN(
        n1053) );
  AOI22D0BWP12T U1875 ( .A1(r5[15]), .A2(n1280), .B1(n1279), .B2(r1[15]), .ZN(
        n1052) );
  AOI22D0BWP12T U1876 ( .A1(r0[15]), .A2(n1282), .B1(n1281), .B2(r3[15]), .ZN(
        n1051) );
  ND4D1BWP12T U1877 ( .A1(n1054), .A2(n1053), .A3(n1052), .A4(n1051), .ZN(
        n1058) );
  CKND0BWP12T U1878 ( .I(lr[15]), .ZN(n1056) );
  OAI22D0BWP12T U1879 ( .A1(n1289), .A2(n1056), .B1(n1055), .B2(n1291), .ZN(
        n1057) );
  AOI21D0BWP12T U1880 ( .A1(n1058), .A2(n1295), .B(n1057), .ZN(n1059) );
  ND4D1BWP12T U1881 ( .A1(n1062), .A2(n1061), .A3(n1060), .A4(n1059), .ZN(
        regC_out[15]) );
  AOI22D0BWP12T U1882 ( .A1(pc_out[8]), .A2(n1324), .B1(n1321), .B2(r9[8]), 
        .ZN(n1073) );
  AOI22D0BWP12T U1883 ( .A1(lr[8]), .A2(n1319), .B1(n1168), .B2(n[2960]), .ZN(
        n1072) );
  AOI22D0BWP12T U1884 ( .A1(r10[8]), .A2(n1322), .B1(n1320), .B2(r11[8]), .ZN(
        n1071) );
  AOI22D0BWP12T U1885 ( .A1(r7[8]), .A2(n1276), .B1(n1275), .B2(r4[8]), .ZN(
        n1066) );
  AOI22D0BWP12T U1886 ( .A1(r2[8]), .A2(n1278), .B1(n1277), .B2(r6[8]), .ZN(
        n1065) );
  AOI22D0BWP12T U1887 ( .A1(r5[8]), .A2(n1280), .B1(n1279), .B2(r1[8]), .ZN(
        n1064) );
  AOI22D0BWP12T U1888 ( .A1(r0[8]), .A2(n1282), .B1(n1281), .B2(r3[8]), .ZN(
        n1063) );
  ND4D1BWP12T U1889 ( .A1(n1066), .A2(n1065), .A3(n1064), .A4(n1063), .ZN(
        n1069) );
  OAI22D0BWP12T U1890 ( .A1(n1238), .A2(n1067), .B1(n2719), .B2(n1291), .ZN(
        n1068) );
  AOI21D0BWP12T U1891 ( .A1(n1069), .A2(n1295), .B(n1068), .ZN(n1070) );
  ND4D1BWP12T U1892 ( .A1(n1073), .A2(n1072), .A3(n1071), .A4(n1070), .ZN(
        regC_out[8]) );
  AOI22D0BWP12T U1893 ( .A1(pc_out[18]), .A2(n1324), .B1(n1321), .B2(r9[18]), 
        .ZN(n1084) );
  AOI22D0BWP12T U1894 ( .A1(lr[18]), .A2(n1319), .B1(n1168), .B2(n[2950]), 
        .ZN(n1083) );
  AOI22D0BWP12T U1895 ( .A1(r10[18]), .A2(n1322), .B1(n1320), .B2(r11[18]), 
        .ZN(n1082) );
  AOI22D0BWP12T U1896 ( .A1(r7[18]), .A2(n1276), .B1(n1275), .B2(r4[18]), .ZN(
        n1077) );
  AOI22D0BWP12T U1897 ( .A1(r2[18]), .A2(n1278), .B1(n1277), .B2(r6[18]), .ZN(
        n1076) );
  AOI22D0BWP12T U1898 ( .A1(r5[18]), .A2(n1280), .B1(n1279), .B2(r1[18]), .ZN(
        n1075) );
  AOI22D0BWP12T U1899 ( .A1(r0[18]), .A2(n1282), .B1(n1281), .B2(r3[18]), .ZN(
        n1074) );
  ND4D1BWP12T U1900 ( .A1(n1077), .A2(n1076), .A3(n1075), .A4(n1074), .ZN(
        n1080) );
  CKND0BWP12T U1901 ( .I(r12[18]), .ZN(n1078) );
  INVD1BWP12T U1902 ( .I(r8[18]), .ZN(n1992) );
  OAI22D0BWP12T U1903 ( .A1(n1238), .A2(n1078), .B1(n1992), .B2(n1291), .ZN(
        n1079) );
  AOI21D0BWP12T U1904 ( .A1(n1080), .A2(n1295), .B(n1079), .ZN(n1081) );
  ND4D1BWP12T U1905 ( .A1(n1084), .A2(n1083), .A3(n1082), .A4(n1081), .ZN(
        regC_out[18]) );
  AOI22D0BWP12T U1906 ( .A1(n[2961]), .A2(n1168), .B1(n1324), .B2(pc_out[7]), 
        .ZN(n1098) );
  AOI22D0BWP12T U1907 ( .A1(r9[7]), .A2(n1321), .B1(n1320), .B2(r11[7]), .ZN(
        n1097) );
  AOI22D0BWP12T U1908 ( .A1(r7[7]), .A2(n1276), .B1(n1275), .B2(r4[7]), .ZN(
        n1088) );
  AOI22D0BWP12T U1909 ( .A1(r2[7]), .A2(n1278), .B1(n1277), .B2(r6[7]), .ZN(
        n1087) );
  AOI22D0BWP12T U1910 ( .A1(r5[7]), .A2(n1280), .B1(n1279), .B2(r1[7]), .ZN(
        n1086) );
  AOI22D0BWP12T U1911 ( .A1(r0[7]), .A2(n1282), .B1(n1281), .B2(r3[7]), .ZN(
        n1085) );
  ND4D1BWP12T U1912 ( .A1(n1088), .A2(n1087), .A3(n1086), .A4(n1085), .ZN(
        n1095) );
  OAI22D0BWP12T U1913 ( .A1(n1238), .A2(n1090), .B1(n1089), .B2(n1291), .ZN(
        n1094) );
  OAI22D0BWP12T U1914 ( .A1(n1289), .A2(n1092), .B1(n1091), .B2(n1249), .ZN(
        n1093) );
  AOI211D0BWP12T U1915 ( .A1(n1095), .A2(n1295), .B(n1094), .C(n1093), .ZN(
        n1096) );
  ND3D1BWP12T U1916 ( .A1(n1098), .A2(n1097), .A3(n1096), .ZN(regC_out[7]) );
  AOI22D0BWP12T U1917 ( .A1(r8[28]), .A2(n1323), .B1(n1322), .B2(r10[28]), 
        .ZN(n1109) );
  AOI22D0BWP12T U1918 ( .A1(n[2940]), .A2(n1168), .B1(n1324), .B2(pc_out[28]), 
        .ZN(n1108) );
  AOI22D0BWP12T U1919 ( .A1(r9[28]), .A2(n1321), .B1(n1320), .B2(r11[28]), 
        .ZN(n1107) );
  AOI22D0BWP12T U1920 ( .A1(r7[28]), .A2(n1276), .B1(n1275), .B2(r4[28]), .ZN(
        n1102) );
  AOI22D0BWP12T U1921 ( .A1(r2[28]), .A2(n1278), .B1(n1277), .B2(r6[28]), .ZN(
        n1101) );
  AOI22D0BWP12T U1922 ( .A1(r5[28]), .A2(n1280), .B1(n1279), .B2(r1[28]), .ZN(
        n1100) );
  AOI22D0BWP12T U1923 ( .A1(r0[28]), .A2(n1282), .B1(n1281), .B2(r3[28]), .ZN(
        n1099) );
  ND4D1BWP12T U1924 ( .A1(n1102), .A2(n1101), .A3(n1100), .A4(n1099), .ZN(
        n1105) );
  CKND0BWP12T U1925 ( .I(lr[28]), .ZN(n1103) );
  TPOAI22D0BWP12T U1926 ( .A1(n1289), .A2(n1103), .B1(n1791), .B2(n1238), .ZN(
        n1104) );
  AOI21D0BWP12T U1927 ( .A1(n1105), .A2(n1295), .B(n1104), .ZN(n1106) );
  ND4D1BWP12T U1928 ( .A1(n1109), .A2(n1108), .A3(n1107), .A4(n1106), .ZN(
        regC_out[28]) );
  CKND0BWP12T U1929 ( .I(r8[23]), .ZN(n1115) );
  AOI22D0BWP12T U1930 ( .A1(r7[23]), .A2(n1276), .B1(n1275), .B2(r4[23]), .ZN(
        n1113) );
  AOI22D0BWP12T U1931 ( .A1(r2[23]), .A2(n1278), .B1(n1277), .B2(r6[23]), .ZN(
        n1112) );
  AOI22D0BWP12T U1932 ( .A1(r5[23]), .A2(n1280), .B1(n1279), .B2(r1[23]), .ZN(
        n1111) );
  AOI22D0BWP12T U1933 ( .A1(r0[23]), .A2(n1282), .B1(n1281), .B2(r3[23]), .ZN(
        n1110) );
  ND4D1BWP12T U1934 ( .A1(n1113), .A2(n1112), .A3(n1111), .A4(n1110), .ZN(
        n1114) );
  MOAI22D0BWP12T U1935 ( .A1(n1291), .A2(n1115), .B1(n1114), .B2(n1295), .ZN(
        n1116) );
  AOI21D0BWP12T U1936 ( .A1(lr[23]), .A2(n1319), .B(n1116), .ZN(n1120) );
  AOI22D0BWP12T U1937 ( .A1(r9[23]), .A2(n1321), .B1(n1320), .B2(r11[23]), 
        .ZN(n1119) );
  AOI22D0BWP12T U1938 ( .A1(pc_out[23]), .A2(n1324), .B1(n1322), .B2(r10[23]), 
        .ZN(n1118) );
  AOI22D0BWP12T U1939 ( .A1(n[2945]), .A2(n1168), .B1(n1325), .B2(r12[23]), 
        .ZN(n1117) );
  ND4D1BWP12T U1940 ( .A1(n1120), .A2(n1119), .A3(n1118), .A4(n1117), .ZN(
        regC_out[23]) );
  AOI22D0BWP12T U1941 ( .A1(r8[12]), .A2(n1323), .B1(n1321), .B2(r9[12]), .ZN(
        n1132) );
  AOI22D0BWP12T U1942 ( .A1(lr[12]), .A2(n1319), .B1(n1168), .B2(n[2956]), 
        .ZN(n1131) );
  AOI22D0BWP12T U1943 ( .A1(r10[12]), .A2(n1322), .B1(n1320), .B2(r11[12]), 
        .ZN(n1130) );
  AOI22D0BWP12T U1944 ( .A1(r7[12]), .A2(n1276), .B1(n1275), .B2(r4[12]), .ZN(
        n1124) );
  AOI22D0BWP12T U1945 ( .A1(r2[12]), .A2(n1278), .B1(n1277), .B2(r6[12]), .ZN(
        n1123) );
  AOI22D0BWP12T U1946 ( .A1(r5[12]), .A2(n1280), .B1(n1279), .B2(r1[12]), .ZN(
        n1122) );
  AOI22D0BWP12T U1947 ( .A1(r0[12]), .A2(n1282), .B1(n1281), .B2(r3[12]), .ZN(
        n1121) );
  ND4D1BWP12T U1948 ( .A1(n1124), .A2(n1123), .A3(n1122), .A4(n1121), .ZN(
        n1128) );
  OAI22D0BWP12T U1949 ( .A1(n1126), .A2(n1268), .B1(n1238), .B2(n1125), .ZN(
        n1127) );
  AOI21D0BWP12T U1950 ( .A1(n1128), .A2(n1295), .B(n1127), .ZN(n1129) );
  ND4D1BWP12T U1951 ( .A1(n1132), .A2(n1131), .A3(n1130), .A4(n1129), .ZN(
        regC_out[12]) );
  AOI22D0BWP12T U1952 ( .A1(n[2967]), .A2(n1168), .B1(n1322), .B2(r10[1]), 
        .ZN(n1146) );
  AOI22D0BWP12T U1953 ( .A1(r9[1]), .A2(n1321), .B1(n1320), .B2(r11[1]), .ZN(
        n1145) );
  AOI22D0BWP12T U1954 ( .A1(r7[1]), .A2(n1276), .B1(n1275), .B2(r4[1]), .ZN(
        n1136) );
  AOI22D0BWP12T U1955 ( .A1(r2[1]), .A2(n1278), .B1(n1277), .B2(r6[1]), .ZN(
        n1135) );
  AOI22D0BWP12T U1956 ( .A1(r5[1]), .A2(n1280), .B1(n1279), .B2(r1[1]), .ZN(
        n1134) );
  AOI22D0BWP12T U1957 ( .A1(r0[1]), .A2(n1282), .B1(n1281), .B2(r3[1]), .ZN(
        n1133) );
  ND4D1BWP12T U1958 ( .A1(n1136), .A2(n1135), .A3(n1134), .A4(n1133), .ZN(
        n1143) );
  OAI22D0BWP12T U1959 ( .A1(n1289), .A2(n1138), .B1(n1137), .B2(n1291), .ZN(
        n1142) );
  OAI22D0BWP12T U1960 ( .A1(n1140), .A2(n1268), .B1(n1238), .B2(n1139), .ZN(
        n1141) );
  AOI211D0BWP12T U1961 ( .A1(n1143), .A2(n1295), .B(n1142), .C(n1141), .ZN(
        n1144) );
  ND3D1BWP12T U1962 ( .A1(n1146), .A2(n1145), .A3(n1144), .ZN(regC_out[1]) );
  CKND2D0BWP12T U1963 ( .A1(write1_in[6]), .A2(n1614), .ZN(n1148) );
  TPAOI21D0BWP12T U1964 ( .A1(n1521), .A2(n[2962]), .B(reset), .ZN(n1147) );
  OAI211D1BWP12T U1965 ( .A1(n1149), .A2(n1443), .B(n1148), .C(n1147), .ZN(
        spin[6]) );
  CKND0BWP12T U1966 ( .I(r12[16]), .ZN(n1155) );
  AOI22D0BWP12T U1967 ( .A1(r7[16]), .A2(n1276), .B1(n1275), .B2(r4[16]), .ZN(
        n1153) );
  AOI22D0BWP12T U1968 ( .A1(r2[16]), .A2(n1278), .B1(n1277), .B2(r6[16]), .ZN(
        n1152) );
  AOI22D0BWP12T U1969 ( .A1(r5[16]), .A2(n1280), .B1(n1279), .B2(r1[16]), .ZN(
        n1151) );
  AOI22D0BWP12T U1970 ( .A1(r0[16]), .A2(n1282), .B1(n1281), .B2(r3[16]), .ZN(
        n1150) );
  ND4D1BWP12T U1971 ( .A1(n1153), .A2(n1152), .A3(n1151), .A4(n1150), .ZN(
        n1154) );
  MOAI22D0BWP12T U1972 ( .A1(n1238), .A2(n1155), .B1(n1154), .B2(n1295), .ZN(
        n1156) );
  AOI21D0BWP12T U1973 ( .A1(lr[16]), .A2(n1319), .B(n1156), .ZN(n1160) );
  AOI22D0BWP12T U1974 ( .A1(r9[16]), .A2(n1321), .B1(n1320), .B2(r11[16]), 
        .ZN(n1159) );
  AOI22D0BWP12T U1975 ( .A1(r8[16]), .A2(n1323), .B1(n1322), .B2(r10[16]), 
        .ZN(n1158) );
  AOI22D0BWP12T U1976 ( .A1(n[2952]), .A2(n1168), .B1(n1324), .B2(pc_out[16]), 
        .ZN(n1157) );
  ND4D1BWP12T U1977 ( .A1(n1160), .A2(n1159), .A3(n1158), .A4(n1157), .ZN(
        regC_out[16]) );
  CKND2D0BWP12T U1978 ( .A1(write1_in[3]), .A2(n1614), .ZN(n1162) );
  AOI21D0BWP12T U1979 ( .A1(n1521), .A2(n[2965]), .B(reset), .ZN(n1161) );
  OAI211D1BWP12T U1980 ( .A1(n1163), .A2(n1443), .B(n1162), .C(n1161), .ZN(
        spin[3]) );
  AOI22D0BWP12T U1981 ( .A1(pc_out[29]), .A2(n1324), .B1(n1323), .B2(r8[29]), 
        .ZN(n1177) );
  AOI22D0BWP12T U1982 ( .A1(lr[29]), .A2(n1319), .B1(n1325), .B2(r12[29]), 
        .ZN(n1176) );
  AOI22D0BWP12T U1983 ( .A1(r10[29]), .A2(n1322), .B1(n1320), .B2(r11[29]), 
        .ZN(n1175) );
  AOI22D0BWP12T U1984 ( .A1(r7[29]), .A2(n1276), .B1(n1275), .B2(r4[29]), .ZN(
        n1167) );
  AOI22D0BWP12T U1985 ( .A1(r2[29]), .A2(n1278), .B1(n1277), .B2(r6[29]), .ZN(
        n1166) );
  AOI22D0BWP12T U1986 ( .A1(r5[29]), .A2(n1280), .B1(n1279), .B2(r1[29]), .ZN(
        n1165) );
  AOI22D0BWP12T U1987 ( .A1(r0[29]), .A2(n1282), .B1(n1281), .B2(r3[29]), .ZN(
        n1164) );
  ND4D1BWP12T U1988 ( .A1(n1167), .A2(n1166), .A3(n1165), .A4(n1164), .ZN(
        n1173) );
  CKND0BWP12T U1989 ( .I(n[2939]), .ZN(n1171) );
  INVD1BWP12T U1990 ( .I(n1168), .ZN(n1316) );
  CKND0BWP12T U1991 ( .I(r9[29]), .ZN(n1169) );
  OAI22D0BWP12T U1992 ( .A1(n1171), .A2(n1316), .B1(n1170), .B2(n1169), .ZN(
        n1172) );
  AOI21D0BWP12T U1993 ( .A1(n1173), .A2(n1295), .B(n1172), .ZN(n1174) );
  ND4D1BWP12T U1994 ( .A1(n1177), .A2(n1176), .A3(n1175), .A4(n1174), .ZN(
        regC_out[29]) );
  AOI22D0BWP12T U1995 ( .A1(pc_out[27]), .A2(n1324), .B1(n1323), .B2(r8[27]), 
        .ZN(n1188) );
  AOI22D0BWP12T U1996 ( .A1(lr[27]), .A2(n1319), .B1(n1325), .B2(r12[27]), 
        .ZN(n1187) );
  AOI22D0BWP12T U1997 ( .A1(r9[27]), .A2(n1321), .B1(n1322), .B2(r10[27]), 
        .ZN(n1186) );
  AOI22D0BWP12T U1998 ( .A1(r7[27]), .A2(n1276), .B1(n1275), .B2(r4[27]), .ZN(
        n1181) );
  AOI22D0BWP12T U1999 ( .A1(r2[27]), .A2(n1278), .B1(n1277), .B2(r6[27]), .ZN(
        n1180) );
  AOI22D0BWP12T U2000 ( .A1(r5[27]), .A2(n1280), .B1(n1279), .B2(r1[27]), .ZN(
        n1179) );
  AOI22D0BWP12T U2001 ( .A1(r0[27]), .A2(n1282), .B1(n1281), .B2(r3[27]), .ZN(
        n1178) );
  ND4D1BWP12T U2002 ( .A1(n1181), .A2(n1180), .A3(n1179), .A4(n1178), .ZN(
        n1184) );
  CKND0BWP12T U2003 ( .I(n[2941]), .ZN(n1182) );
  CKND0BWP12T U2004 ( .I(r11[27]), .ZN(n1485) );
  OAI22D0BWP12T U2005 ( .A1(n1182), .A2(n1316), .B1(n1287), .B2(n1485), .ZN(
        n1183) );
  AOI21D0BWP12T U2006 ( .A1(n1184), .A2(n1295), .B(n1183), .ZN(n1185) );
  ND4D1BWP12T U2007 ( .A1(n1188), .A2(n1187), .A3(n1186), .A4(n1185), .ZN(
        regC_out[27]) );
  AOI22D0BWP12T U2008 ( .A1(pc_out[24]), .A2(n1324), .B1(n1323), .B2(r8[24]), 
        .ZN(n1200) );
  AOI22D0BWP12T U2009 ( .A1(r9[24]), .A2(n1321), .B1(n1320), .B2(r11[24]), 
        .ZN(n1199) );
  AOI22D0BWP12T U2010 ( .A1(r7[24]), .A2(n1276), .B1(n1275), .B2(r4[24]), .ZN(
        n1192) );
  AOI22D0BWP12T U2011 ( .A1(r2[24]), .A2(n1278), .B1(n1277), .B2(r6[24]), .ZN(
        n1191) );
  AOI22D0BWP12T U2012 ( .A1(r5[24]), .A2(n1280), .B1(n1279), .B2(r1[24]), .ZN(
        n1190) );
  AOI22D0BWP12T U2013 ( .A1(r0[24]), .A2(n1282), .B1(n1281), .B2(r3[24]), .ZN(
        n1189) );
  ND4D1BWP12T U2014 ( .A1(n1192), .A2(n1191), .A3(n1190), .A4(n1189), .ZN(
        n1197) );
  INVD1BWP12T U2015 ( .I(r12[24]), .ZN(n2850) );
  OAI22D0BWP12T U2016 ( .A1(n1238), .A2(n2850), .B1(n1193), .B2(n1249), .ZN(
        n1196) );
  INVD1BWP12T U2017 ( .I(n[2944]), .ZN(n2847) );
  CKND0BWP12T U2018 ( .I(lr[24]), .ZN(n1194) );
  OAI22D0BWP12T U2019 ( .A1(n2847), .A2(n1316), .B1(n1289), .B2(n1194), .ZN(
        n1195) );
  AOI211D0BWP12T U2020 ( .A1(n1197), .A2(n1295), .B(n1196), .C(n1195), .ZN(
        n1198) );
  ND3D1BWP12T U2021 ( .A1(n1200), .A2(n1199), .A3(n1198), .ZN(regC_out[24]) );
  CKND2D0BWP12T U2022 ( .A1(write1_in[7]), .A2(n1614), .ZN(n1202) );
  AOI21D0BWP12T U2023 ( .A1(n1521), .A2(n[2961]), .B(reset), .ZN(n1201) );
  OAI211D1BWP12T U2024 ( .A1(n1203), .A2(n1443), .B(n1202), .C(n1201), .ZN(
        spin[7]) );
  AOI22D0BWP12T U2025 ( .A1(r8[17]), .A2(n1323), .B1(n1322), .B2(r10[17]), 
        .ZN(n1213) );
  AOI22D0BWP12T U2026 ( .A1(r12[17]), .A2(n1325), .B1(n1324), .B2(pc_out[17]), 
        .ZN(n1212) );
  AOI22D0BWP12T U2027 ( .A1(r9[17]), .A2(n1321), .B1(n1320), .B2(r11[17]), 
        .ZN(n1211) );
  AOI22D0BWP12T U2028 ( .A1(r7[17]), .A2(n1276), .B1(n1275), .B2(r4[17]), .ZN(
        n1207) );
  AOI22D0BWP12T U2029 ( .A1(r2[17]), .A2(n1278), .B1(n1277), .B2(r6[17]), .ZN(
        n1206) );
  AOI22D0BWP12T U2030 ( .A1(r5[17]), .A2(n1280), .B1(n1279), .B2(r1[17]), .ZN(
        n1205) );
  AOI22D0BWP12T U2031 ( .A1(r0[17]), .A2(n1282), .B1(n1281), .B2(r3[17]), .ZN(
        n1204) );
  ND4D1BWP12T U2032 ( .A1(n1207), .A2(n1206), .A3(n1205), .A4(n1204), .ZN(
        n1209) );
  INVD1BWP12T U2033 ( .I(lr[17]), .ZN(n2682) );
  OAI22D0BWP12T U2034 ( .A1(n2686), .A2(n1316), .B1(n1289), .B2(n2682), .ZN(
        n1208) );
  AOI21D0BWP12T U2035 ( .A1(n1209), .A2(n1295), .B(n1208), .ZN(n1210) );
  ND4D1BWP12T U2036 ( .A1(n1213), .A2(n1212), .A3(n1211), .A4(n1210), .ZN(
        regC_out[17]) );
  AOI22D0BWP12T U2037 ( .A1(pc_out[20]), .A2(n1324), .B1(n1323), .B2(r8[20]), 
        .ZN(n1223) );
  AOI22D0BWP12T U2038 ( .A1(lr[20]), .A2(n1319), .B1(n1325), .B2(r12[20]), 
        .ZN(n1222) );
  AOI22D0BWP12T U2039 ( .A1(r9[20]), .A2(n1321), .B1(n1322), .B2(r10[20]), 
        .ZN(n1221) );
  AOI22D0BWP12T U2040 ( .A1(r7[20]), .A2(n1276), .B1(n1275), .B2(r4[20]), .ZN(
        n1217) );
  AOI22D0BWP12T U2041 ( .A1(r2[20]), .A2(n1278), .B1(n1277), .B2(r6[20]), .ZN(
        n1216) );
  AOI22D0BWP12T U2042 ( .A1(r5[20]), .A2(n1280), .B1(n1279), .B2(r1[20]), .ZN(
        n1215) );
  AOI22D0BWP12T U2043 ( .A1(r0[20]), .A2(n1282), .B1(n1281), .B2(r3[20]), .ZN(
        n1214) );
  ND4D1BWP12T U2044 ( .A1(n1217), .A2(n1216), .A3(n1215), .A4(n1214), .ZN(
        n1219) );
  INVD1BWP12T U2045 ( .I(r11[20]), .ZN(n1972) );
  OAI22D0BWP12T U2046 ( .A1(n2071), .A2(n1316), .B1(n1287), .B2(n1972), .ZN(
        n1218) );
  AOI21D0BWP12T U2047 ( .A1(n1219), .A2(n1295), .B(n1218), .ZN(n1220) );
  ND4D1BWP12T U2048 ( .A1(n1223), .A2(n1222), .A3(n1221), .A4(n1220), .ZN(
        regC_out[20]) );
  AOI22D0BWP12T U2049 ( .A1(r8[11]), .A2(n1323), .B1(n1321), .B2(r9[11]), .ZN(
        n1233) );
  AOI22D0BWP12T U2050 ( .A1(lr[11]), .A2(n1319), .B1(n1324), .B2(pc_out[11]), 
        .ZN(n1232) );
  AOI22D0BWP12T U2051 ( .A1(r10[11]), .A2(n1322), .B1(n1320), .B2(r11[11]), 
        .ZN(n1231) );
  AOI22D0BWP12T U2052 ( .A1(r7[11]), .A2(n1276), .B1(n1275), .B2(r4[11]), .ZN(
        n1227) );
  AOI22D0BWP12T U2053 ( .A1(r2[11]), .A2(n1278), .B1(n1277), .B2(r6[11]), .ZN(
        n1226) );
  AOI22D0BWP12T U2054 ( .A1(r5[11]), .A2(n1280), .B1(n1279), .B2(r1[11]), .ZN(
        n1225) );
  AOI22D0BWP12T U2055 ( .A1(r0[11]), .A2(n1282), .B1(n1281), .B2(r3[11]), .ZN(
        n1224) );
  ND4D1BWP12T U2056 ( .A1(n1227), .A2(n1226), .A3(n1225), .A4(n1224), .ZN(
        n1229) );
  INVD1BWP12T U2057 ( .I(n[2957]), .ZN(n1932) );
  OAI22D0BWP12T U2058 ( .A1(n1932), .A2(n1316), .B1(n1238), .B2(n1928), .ZN(
        n1228) );
  AOI21D0BWP12T U2059 ( .A1(n1229), .A2(n1295), .B(n1228), .ZN(n1230) );
  ND4D1BWP12T U2060 ( .A1(n1233), .A2(n1232), .A3(n1231), .A4(n1230), .ZN(
        regC_out[11]) );
  AOI22D0BWP12T U2061 ( .A1(r8[6]), .A2(n1323), .B1(n1321), .B2(r9[6]), .ZN(
        n1244) );
  AOI22D0BWP12T U2062 ( .A1(lr[6]), .A2(n1319), .B1(n1324), .B2(pc_out[6]), 
        .ZN(n1243) );
  AOI22D0BWP12T U2063 ( .A1(r10[6]), .A2(n1322), .B1(n1320), .B2(r11[6]), .ZN(
        n1242) );
  AOI22D0BWP12T U2064 ( .A1(r7[6]), .A2(n1276), .B1(n1275), .B2(r4[6]), .ZN(
        n1237) );
  AOI22D0BWP12T U2065 ( .A1(r2[6]), .A2(n1278), .B1(n1277), .B2(r6[6]), .ZN(
        n1236) );
  AOI22D0BWP12T U2066 ( .A1(r5[6]), .A2(n1280), .B1(n1279), .B2(r1[6]), .ZN(
        n1235) );
  AOI22D0BWP12T U2067 ( .A1(r0[6]), .A2(n1282), .B1(n1281), .B2(r3[6]), .ZN(
        n1234) );
  ND4D1BWP12T U2068 ( .A1(n1237), .A2(n1236), .A3(n1235), .A4(n1234), .ZN(
        n1240) );
  OAI22D0BWP12T U2069 ( .A1(n2084), .A2(n1316), .B1(n1238), .B2(n2088), .ZN(
        n1239) );
  AOI21D0BWP12T U2070 ( .A1(n1240), .A2(n1295), .B(n1239), .ZN(n1241) );
  ND4D1BWP12T U2071 ( .A1(n1244), .A2(n1243), .A3(n1242), .A4(n1241), .ZN(
        regC_out[6]) );
  AOI22D0BWP12T U2072 ( .A1(r12[14]), .A2(n1325), .B1(n1324), .B2(pc_out[14]), 
        .ZN(n1259) );
  AOI22D0BWP12T U2073 ( .A1(r9[14]), .A2(n1321), .B1(n1320), .B2(r11[14]), 
        .ZN(n1258) );
  AOI22D0BWP12T U2074 ( .A1(r7[14]), .A2(n1276), .B1(n1275), .B2(r4[14]), .ZN(
        n1248) );
  AOI22D0BWP12T U2075 ( .A1(r2[14]), .A2(n1278), .B1(n1277), .B2(r6[14]), .ZN(
        n1247) );
  AOI22D0BWP12T U2076 ( .A1(r5[14]), .A2(n1280), .B1(n1279), .B2(r1[14]), .ZN(
        n1246) );
  AOI22D0BWP12T U2077 ( .A1(r0[14]), .A2(n1282), .B1(n1281), .B2(r3[14]), .ZN(
        n1245) );
  ND4D1BWP12T U2078 ( .A1(n1248), .A2(n1247), .A3(n1246), .A4(n1245), .ZN(
        n1256) );
  OAI22D0BWP12T U2079 ( .A1(n1291), .A2(n1251), .B1(n1250), .B2(n1249), .ZN(
        n1255) );
  OAI22D0BWP12T U2080 ( .A1(n1253), .A2(n1316), .B1(n1289), .B2(n1252), .ZN(
        n1254) );
  AOI211D0BWP12T U2081 ( .A1(n1256), .A2(n1295), .B(n1255), .C(n1254), .ZN(
        n1257) );
  ND3D1BWP12T U2082 ( .A1(n1259), .A2(n1258), .A3(n1257), .ZN(regC_out[14]) );
  CKND2D0BWP12T U2083 ( .A1(write1_in[4]), .A2(n1614), .ZN(n1261) );
  AOI21D0BWP12T U2084 ( .A1(n1521), .A2(n[2964]), .B(reset), .ZN(n1260) );
  OAI211D1BWP12T U2085 ( .A1(n1262), .A2(n1443), .B(n1261), .C(n1260), .ZN(
        spin[4]) );
  AOI22D0BWP12T U2086 ( .A1(r8[26]), .A2(n1323), .B1(n1321), .B2(r9[26]), .ZN(
        n1274) );
  AOI22D0BWP12T U2087 ( .A1(lr[26]), .A2(n1319), .B1(n1325), .B2(r12[26]), 
        .ZN(n1273) );
  AOI22D0BWP12T U2088 ( .A1(r10[26]), .A2(n1322), .B1(n1320), .B2(r11[26]), 
        .ZN(n1272) );
  AOI22D0BWP12T U2089 ( .A1(r7[26]), .A2(n1276), .B1(n1275), .B2(r4[26]), .ZN(
        n1266) );
  AOI22D0BWP12T U2090 ( .A1(r2[26]), .A2(n1278), .B1(n1277), .B2(r6[26]), .ZN(
        n1265) );
  AOI22D0BWP12T U2091 ( .A1(r5[26]), .A2(n1280), .B1(n1279), .B2(r1[26]), .ZN(
        n1264) );
  AOI22D0BWP12T U2092 ( .A1(r0[26]), .A2(n1282), .B1(n1281), .B2(r3[26]), .ZN(
        n1263) );
  ND4D1BWP12T U2093 ( .A1(n1266), .A2(n1265), .A3(n1264), .A4(n1263), .ZN(
        n1270) );
  CKND0BWP12T U2094 ( .I(pc_out[26]), .ZN(n1707) );
  CKND0BWP12T U2095 ( .I(n[2942]), .ZN(n1267) );
  OAI22D0BWP12T U2096 ( .A1(n1707), .A2(n1268), .B1(n1267), .B2(n1316), .ZN(
        n1269) );
  AOI21D0BWP12T U2097 ( .A1(n1270), .A2(n1295), .B(n1269), .ZN(n1271) );
  ND4D1BWP12T U2098 ( .A1(n1274), .A2(n1273), .A3(n1272), .A4(n1271), .ZN(
        regC_out[26]) );
  AOI22D0BWP12T U2099 ( .A1(r12[22]), .A2(n1325), .B1(n1324), .B2(pc_out[22]), 
        .ZN(n1299) );
  AOI22D0BWP12T U2100 ( .A1(r9[22]), .A2(n1321), .B1(n1322), .B2(r10[22]), 
        .ZN(n1298) );
  AOI22D0BWP12T U2101 ( .A1(r7[22]), .A2(n1276), .B1(n1275), .B2(r4[22]), .ZN(
        n1286) );
  AOI22D0BWP12T U2102 ( .A1(r2[22]), .A2(n1278), .B1(n1277), .B2(r6[22]), .ZN(
        n1285) );
  AOI22D0BWP12T U2103 ( .A1(r5[22]), .A2(n1280), .B1(n1279), .B2(r1[22]), .ZN(
        n1284) );
  AOI22D0BWP12T U2104 ( .A1(r0[22]), .A2(n1282), .B1(n1281), .B2(r3[22]), .ZN(
        n1283) );
  ND4D1BWP12T U2105 ( .A1(n1286), .A2(n1285), .A3(n1284), .A4(n1283), .ZN(
        n1296) );
  OAI22D0BWP12T U2106 ( .A1(n1289), .A2(n1288), .B1(n1461), .B2(n1287), .ZN(
        n1294) );
  OAI22D0BWP12T U2107 ( .A1(n1292), .A2(n1316), .B1(n1291), .B2(n1290), .ZN(
        n1293) );
  AOI211D0BWP12T U2108 ( .A1(n1296), .A2(n1295), .B(n1294), .C(n1293), .ZN(
        n1297) );
  ND3D1BWP12T U2109 ( .A1(n1299), .A2(n1298), .A3(n1297), .ZN(regC_out[22]) );
  OAI22D0BWP12T U2110 ( .A1(n2774), .A2(n1302), .B1(n1301), .B2(n1300), .ZN(
        n1314) );
  OAI22D0BWP12T U2111 ( .A1(n1305), .A2(n1304), .B1(n1303), .B2(n2781), .ZN(
        n1313) );
  OAI22D0BWP12T U2112 ( .A1(n1307), .A2(n2788), .B1(n1306), .B2(n2798), .ZN(
        n1312) );
  OAI22D0BWP12T U2113 ( .A1(n1310), .A2(n1309), .B1(n1308), .B2(n2779), .ZN(
        n1311) );
  NR4D0BWP12T U2114 ( .A1(n1314), .A2(n1313), .A3(n1312), .A4(n1311), .ZN(
        n1317) );
  OAI22D0BWP12T U2115 ( .A1(n1317), .A2(readC_sel[4]), .B1(n1316), .B2(n1315), 
        .ZN(n1318) );
  AOI21D0BWP12T U2116 ( .A1(lr[10]), .A2(n1319), .B(n1318), .ZN(n1329) );
  AOI22D0BWP12T U2117 ( .A1(r9[10]), .A2(n1321), .B1(n1320), .B2(r11[10]), 
        .ZN(n1328) );
  AOI22D0BWP12T U2118 ( .A1(r8[10]), .A2(n1323), .B1(n1322), .B2(r10[10]), 
        .ZN(n1327) );
  AOI22D0BWP12T U2119 ( .A1(r12[10]), .A2(n1325), .B1(n1324), .B2(pc_out[10]), 
        .ZN(n1326) );
  ND4D1BWP12T U2120 ( .A1(n1329), .A2(n1328), .A3(n1327), .A4(n1326), .ZN(
        regC_out[10]) );
  CKND2D0BWP12T U2121 ( .A1(write1_in[8]), .A2(n1614), .ZN(n1331) );
  AOI21D0BWP12T U2122 ( .A1(n1521), .A2(n[2960]), .B(reset), .ZN(n1330) );
  OAI211D1BWP12T U2123 ( .A1(n1332), .A2(n1443), .B(n1331), .C(n1330), .ZN(
        spin[8]) );
  CKND2D0BWP12T U2124 ( .A1(write1_in[10]), .A2(n1614), .ZN(n1334) );
  AOI21D0BWP12T U2125 ( .A1(n1521), .A2(n[2958]), .B(reset), .ZN(n1333) );
  OAI211D1BWP12T U2126 ( .A1(n1335), .A2(n1443), .B(n1334), .C(n1333), .ZN(
        spin[10]) );
  CKND2D0BWP12T U2127 ( .A1(write1_in[9]), .A2(n1614), .ZN(n1337) );
  AOI21D0BWP12T U2128 ( .A1(n1521), .A2(n[2959]), .B(reset), .ZN(n1336) );
  OAI211D1BWP12T U2129 ( .A1(n1338), .A2(n1443), .B(n1337), .C(n1336), .ZN(
        spin[9]) );
  AOI22D0BWP12T U2130 ( .A1(r8[8]), .A2(n1382), .B1(n1381), .B2(r4[8]), .ZN(
        n1340) );
  AOI22D0BWP12T U2131 ( .A1(n[2960]), .A2(n1384), .B1(n1383), .B2(r10[8]), 
        .ZN(n1339) );
  CKND2D1BWP12T U2132 ( .A1(n1340), .A2(n1339), .ZN(n1349) );
  AOI22D0BWP12T U2133 ( .A1(r7[8]), .A2(n1388), .B1(n1387), .B2(r5[8]), .ZN(
        n1344) );
  AOI22D0BWP12T U2134 ( .A1(lr[8]), .A2(n1390), .B1(n1389), .B2(r9[8]), .ZN(
        n1343) );
  AOI22D0BWP12T U2135 ( .A1(r6[8]), .A2(n1392), .B1(n1391), .B2(r11[8]), .ZN(
        n1342) );
  CKND2D0BWP12T U2136 ( .A1(n1393), .A2(r12[8]), .ZN(n1341) );
  ND4D1BWP12T U2137 ( .A1(n1344), .A2(n1343), .A3(n1342), .A4(n1341), .ZN(
        n1348) );
  AOI22D0BWP12T U2138 ( .A1(r3[8]), .A2(n1399), .B1(n1398), .B2(r2[8]), .ZN(
        n1346) );
  AOI22D0BWP12T U2139 ( .A1(n1401), .A2(r0[8]), .B1(pc_out[8]), .B2(n1400), 
        .ZN(n1345) );
  OAI211D0BWP12T U2140 ( .A1(n2706), .A2(n1404), .B(n1346), .C(n1345), .ZN(
        n1347) );
  OA31D1BWP12T U2141 ( .A1(n1349), .A2(n1348), .A3(n1347), .B(n1405), .Z(
        regD_out[8]) );
  AOI22D0BWP12T U2142 ( .A1(r8[10]), .A2(n1382), .B1(n1381), .B2(r4[10]), .ZN(
        n1351) );
  AOI22D0BWP12T U2143 ( .A1(n[2958]), .A2(n1384), .B1(n1383), .B2(r10[10]), 
        .ZN(n1350) );
  CKND2D1BWP12T U2144 ( .A1(n1351), .A2(n1350), .ZN(n1360) );
  AOI22D0BWP12T U2145 ( .A1(r7[10]), .A2(n1388), .B1(n1387), .B2(r5[10]), .ZN(
        n1355) );
  AOI22D0BWP12T U2146 ( .A1(lr[10]), .A2(n1390), .B1(n1389), .B2(r9[10]), .ZN(
        n1354) );
  AOI22D0BWP12T U2147 ( .A1(r6[10]), .A2(n1392), .B1(n1391), .B2(r11[10]), 
        .ZN(n1353) );
  CKND2D0BWP12T U2148 ( .A1(n1393), .A2(r12[10]), .ZN(n1352) );
  ND4D1BWP12T U2149 ( .A1(n1355), .A2(n1354), .A3(n1353), .A4(n1352), .ZN(
        n1359) );
  AOI22D0BWP12T U2150 ( .A1(r3[10]), .A2(n1399), .B1(n1398), .B2(r2[10]), .ZN(
        n1357) );
  AOI22D0BWP12T U2151 ( .A1(n1401), .A2(r0[10]), .B1(pc_out[10]), .B2(n1400), 
        .ZN(n1356) );
  OAI211D0BWP12T U2152 ( .A1(n2781), .A2(n1404), .B(n1357), .C(n1356), .ZN(
        n1358) );
  OA31D1BWP12T U2153 ( .A1(n1360), .A2(n1359), .A3(n1358), .B(n1405), .Z(
        regD_out[10]) );
  CKND2D0BWP12T U2154 ( .A1(write1_in[12]), .A2(n1614), .ZN(n1362) );
  TPAOI21D0BWP12T U2155 ( .A1(n1521), .A2(n[2956]), .B(reset), .ZN(n1361) );
  OAI211D1BWP12T U2156 ( .A1(n1363), .A2(n1443), .B(n1362), .C(n1361), .ZN(
        spin[12]) );
  CKND2D0BWP12T U2157 ( .A1(write1_in[11]), .A2(n1614), .ZN(n1365) );
  TPAOI21D0BWP12T U2158 ( .A1(n1521), .A2(n[2957]), .B(reset), .ZN(n1364) );
  OAI211D1BWP12T U2159 ( .A1(n1366), .A2(n1443), .B(n1365), .C(n1364), .ZN(
        spin[11]) );
  TPNR2D2BWP12T U2160 ( .A1(n1368), .A2(n1367), .ZN(n1409) );
  CKND2D0BWP12T U2161 ( .A1(write2_in[5]), .A2(n2916), .ZN(n1369) );
  IOA21D1BWP12T U2162 ( .A1(write1_in[5]), .A2(n2920), .B(n1369), .ZN(n1410)
         );
  AOI22D0BWP12T U2163 ( .A1(r8[12]), .A2(n1382), .B1(n1381), .B2(r4[12]), .ZN(
        n1371) );
  AOI22D0BWP12T U2164 ( .A1(n[2956]), .A2(n1384), .B1(n1383), .B2(r10[12]), 
        .ZN(n1370) );
  CKND2D1BWP12T U2165 ( .A1(n1371), .A2(n1370), .ZN(n1380) );
  AOI22D0BWP12T U2166 ( .A1(r7[12]), .A2(n1388), .B1(n1387), .B2(r5[12]), .ZN(
        n1375) );
  AOI22D0BWP12T U2167 ( .A1(lr[12]), .A2(n1390), .B1(n1389), .B2(r9[12]), .ZN(
        n1374) );
  AOI22D0BWP12T U2168 ( .A1(r6[12]), .A2(n1392), .B1(n1391), .B2(r11[12]), 
        .ZN(n1373) );
  CKND2D0BWP12T U2169 ( .A1(n1393), .A2(r12[12]), .ZN(n1372) );
  ND4D1BWP12T U2170 ( .A1(n1375), .A2(n1374), .A3(n1373), .A4(n1372), .ZN(
        n1379) );
  AOI22D0BWP12T U2171 ( .A1(r3[12]), .A2(n1399), .B1(n1398), .B2(r2[12]), .ZN(
        n1377) );
  AOI22D0BWP12T U2172 ( .A1(n1401), .A2(r0[12]), .B1(pc_out[12]), .B2(n1400), 
        .ZN(n1376) );
  OAI211D0BWP12T U2173 ( .A1(n1963), .A2(n1404), .B(n1377), .C(n1376), .ZN(
        n1378) );
  OA31D1BWP12T U2174 ( .A1(n1380), .A2(n1379), .A3(n1378), .B(n1405), .Z(
        regD_out[12]) );
  AOI22D0BWP12T U2175 ( .A1(r8[11]), .A2(n1382), .B1(n1381), .B2(r4[11]), .ZN(
        n1386) );
  AOI22D0BWP12T U2176 ( .A1(n[2957]), .A2(n1384), .B1(n1383), .B2(r10[11]), 
        .ZN(n1385) );
  CKND2D1BWP12T U2177 ( .A1(n1386), .A2(n1385), .ZN(n1408) );
  AOI22D0BWP12T U2178 ( .A1(r7[11]), .A2(n1388), .B1(n1387), .B2(r5[11]), .ZN(
        n1397) );
  AOI22D0BWP12T U2179 ( .A1(lr[11]), .A2(n1390), .B1(n1389), .B2(r9[11]), .ZN(
        n1396) );
  AOI22D0BWP12T U2180 ( .A1(r6[11]), .A2(n1392), .B1(n1391), .B2(r11[11]), 
        .ZN(n1395) );
  CKND2D0BWP12T U2181 ( .A1(n1393), .A2(r12[11]), .ZN(n1394) );
  ND4D1BWP12T U2182 ( .A1(n1397), .A2(n1396), .A3(n1395), .A4(n1394), .ZN(
        n1407) );
  AOI22D0BWP12T U2183 ( .A1(r3[11]), .A2(n1399), .B1(n1398), .B2(r2[11]), .ZN(
        n1403) );
  AOI22D0BWP12T U2184 ( .A1(n1401), .A2(r0[11]), .B1(pc_out[11]), .B2(n1400), 
        .ZN(n1402) );
  OAI211D0BWP12T U2185 ( .A1(n1929), .A2(n1404), .B(n1403), .C(n1402), .ZN(
        n1406) );
  OA31D1BWP12T U2186 ( .A1(n1408), .A2(n1407), .A3(n1406), .B(n1405), .Z(
        regD_out[11]) );
  TPND2D1BWP12T U2187 ( .A1(n1410), .A2(n1409), .ZN(n1415) );
  AN2XD0BWP12T U2188 ( .A1(write2_in[6]), .A2(n2916), .Z(n1411) );
  AOI21D1BWP12T U2189 ( .A1(write1_in[6]), .A2(n2920), .B(n1411), .ZN(n1414)
         );
  AO222D1BWP12T U2190 ( .A1(n1512), .A2(write1_in[15]), .B1(n1513), .B2(
        write2_in[15]), .C1(n1511), .C2(r2[15]), .Z(n2568) );
  AO222D1BWP12T U2191 ( .A1(n1515), .A2(write1_in[15]), .B1(n1516), .B2(
        write2_in[15]), .C1(n1514), .C2(r10[15]), .Z(n2312) );
  AO222D1BWP12T U2192 ( .A1(n1509), .A2(write1_in[15]), .B1(n1510), .B2(
        write2_in[15]), .C1(n1508), .C2(r11[15]), .Z(n2280) );
  AO222D1BWP12T U2193 ( .A1(n1607), .A2(write1_in[15]), .B1(n1608), .B2(lr[15]), .C1(write2_in[15]), .C2(n1609), .Z(n2216) );
  AO222D1BWP12T U2194 ( .A1(n1602), .A2(write1_in[15]), .B1(n1603), .B2(r8[15]), .C1(write2_in[15]), .C2(n1604), .Z(n2376) );
  AO222D1BWP12T U2195 ( .A1(n1597), .A2(write1_in[15]), .B1(n1598), .B2(
        r12[15]), .C1(write2_in[15]), .C2(n1599), .Z(n2248) );
  AO222D1BWP12T U2196 ( .A1(n1573), .A2(write1_in[15]), .B1(n1576), .B2(
        write2_in[15]), .C1(n1504), .C2(r3[15]), .Z(n2536) );
  AO222D1BWP12T U2197 ( .A1(n1555), .A2(write1_in[15]), .B1(n1519), .B2(r6[15]), .C1(write2_in[15]), .C2(n1558), .Z(n2440) );
  AO222D1BWP12T U2198 ( .A1(n1561), .A2(write1_in[15]), .B1(n1520), .B2(r5[15]), .C1(write2_in[15]), .C2(n1564), .Z(n2472) );
  AO222D1BWP12T U2199 ( .A1(n1567), .A2(write1_in[15]), .B1(n1505), .B2(r7[15]), .C1(write2_in[15]), .C2(n1570), .Z(n2408) );
  AO222D1BWP12T U2200 ( .A1(n1585), .A2(write1_in[15]), .B1(n1517), .B2(r1[15]), .C1(write2_in[15]), .C2(n1588), .Z(n2600) );
  AO222D1BWP12T U2201 ( .A1(n1579), .A2(write1_in[15]), .B1(n1518), .B2(r4[15]), .C1(write2_in[15]), .C2(n1582), .Z(n2504) );
  AO222D1BWP12T U2202 ( .A1(n1591), .A2(write1_in[15]), .B1(n1507), .B2(r9[15]), .C1(write2_in[15]), .C2(n1594), .Z(n2344) );
  AO222D1BWP12T U2203 ( .A1(n1549), .A2(write1_in[15]), .B1(n1506), .B2(r0[15]), .C1(write2_in[15]), .C2(n1552), .Z(n2632) );
  AO222D1BWP12T U2204 ( .A1(n1620), .A2(write1_in[15]), .B1(n1625), .B2(
        write2_in[15]), .C1(n1622), .C2(tmp1[15]), .Z(n2152) );
  INVD1BWP12T U2205 ( .I(r2[17]), .ZN(n2670) );
  OAI222D1BWP12T U2206 ( .A1(n1524), .A2(n1418), .B1(n1523), .B2(n1498), .C1(
        n1522), .C2(n2670), .ZN(n2570) );
  OAI222D1BWP12T U2207 ( .A1(n1439), .A2(n1418), .B1(n1475), .B2(n1498), .C1(
        n1438), .C2(n2682), .ZN(n2218) );
  OAI222D1BWP12T U2208 ( .A1(n1533), .A2(n1418), .B1(n1532), .B2(n1498), .C1(
        n1530), .C2(n1412), .ZN(n2282) );
  INVD1BWP12T U2209 ( .I(r10[17]), .ZN(n2662) );
  OAI222D1BWP12T U2210 ( .A1(n1528), .A2(n1418), .B1(n1527), .B2(n1498), .C1(
        n1526), .C2(n2662), .ZN(n2314) );
  BUFFD3BWP12T U2211 ( .I(write1_in[16]), .Z(n1496) );
  AO222D1BWP12T U2212 ( .A1(n1597), .A2(n1496), .B1(n1598), .B2(r12[16]), .C1(
        write2_in[16]), .C2(n1599), .Z(n2249) );
  AO222D1BWP12T U2213 ( .A1(n1607), .A2(n1496), .B1(n1608), .B2(lr[16]), .C1(
        write2_in[16]), .C2(n1609), .Z(n2217) );
  AO222D1BWP12T U2214 ( .A1(n1602), .A2(n1496), .B1(n1603), .B2(r8[16]), .C1(
        write2_in[16]), .C2(n1604), .Z(n2377) );
  AO222D1BWP12T U2215 ( .A1(n1555), .A2(n1496), .B1(n1519), .B2(r6[16]), .C1(
        write2_in[16]), .C2(n1558), .Z(n2441) );
  AO222D1BWP12T U2216 ( .A1(n1561), .A2(n1496), .B1(n1520), .B2(r5[16]), .C1(
        write2_in[16]), .C2(n1564), .Z(n2473) );
  AO222D1BWP12T U2217 ( .A1(n1579), .A2(n1496), .B1(n1518), .B2(r4[16]), .C1(
        write2_in[16]), .C2(n1582), .Z(n2505) );
  AO222D1BWP12T U2218 ( .A1(n1585), .A2(n1496), .B1(n1517), .B2(r1[16]), .C1(
        write2_in[16]), .C2(n1588), .Z(n2601) );
  AO222D1BWP12T U2219 ( .A1(n1567), .A2(n1496), .B1(n1505), .B2(r7[16]), .C1(
        write2_in[16]), .C2(n1570), .Z(n2409) );
  AO222D1BWP12T U2220 ( .A1(n1549), .A2(n1496), .B1(n1506), .B2(r0[16]), .C1(
        write2_in[16]), .C2(n1552), .Z(n2633) );
  AO222D1BWP12T U2221 ( .A1(n1591), .A2(n1496), .B1(n1507), .B2(r9[16]), .C1(
        write2_in[16]), .C2(n1594), .Z(n2345) );
  AO222D1BWP12T U2222 ( .A1(n1515), .A2(n1496), .B1(n1516), .B2(write2_in[16]), 
        .C1(n1514), .C2(r10[16]), .Z(n2313) );
  AO222D1BWP12T U2223 ( .A1(n1509), .A2(n1496), .B1(n1510), .B2(write2_in[16]), 
        .C1(n1508), .C2(r11[16]), .Z(n2281) );
  AO222D1BWP12T U2224 ( .A1(n1512), .A2(n1496), .B1(n1513), .B2(write2_in[16]), 
        .C1(n1511), .C2(r2[16]), .Z(n2569) );
  AO222D1BWP12T U2225 ( .A1(n1573), .A2(n1496), .B1(n1576), .B2(write2_in[16]), 
        .C1(n1504), .C2(r3[16]), .Z(n2537) );
  AO222D1BWP12T U2226 ( .A1(n1614), .A2(n1496), .B1(n1521), .B2(n[2952]), .C1(
        write2_in[16]), .C2(n1617), .Z(spin[16]) );
  CKND2D0BWP12T U2227 ( .A1(write2_in[7]), .A2(n2916), .ZN(n1413) );
  IOA21D1BWP12T U2228 ( .A1(write1_in[7]), .A2(n2920), .B(n1413), .ZN(n1421)
         );
  TPNR2D1BWP12T U2229 ( .A1(n1415), .A2(n1414), .ZN(n1420) );
  XOR2XD1BWP12T U2230 ( .A1(n1421), .A2(n1420), .Z(n1416) );
  AO222D1BWP12T U2231 ( .A1(n1416), .A2(n2914), .B1(n1488), .B2(next_pc_in[7]), 
        .C1(n1690), .C2(pc_out[7]), .Z(n2176) );
  OAI222D1BWP12T U2232 ( .A1(n1444), .A2(n1418), .B1(n1490), .B2(n1498), .C1(
        n1556), .C2(n2690), .ZN(n2442) );
  AO222D1BWP12T U2233 ( .A1(n1620), .A2(n1496), .B1(n1625), .B2(write2_in[16]), 
        .C1(n1622), .C2(tmp1[16]), .Z(n2153) );
  OAI222D1BWP12T U2234 ( .A1(n1458), .A2(n1418), .B1(n1457), .B2(n1498), .C1(
        n1574), .C2(n2685), .ZN(n2538) );
  CKND0BWP12T U2235 ( .I(r9[17]), .ZN(n1417) );
  OAI222D1BWP12T U2236 ( .A1(n1453), .A2(n1418), .B1(n1481), .B2(n1498), .C1(
        n1592), .C2(n1417), .ZN(n2346) );
  AO222D1BWP12T U2237 ( .A1(write2_in[18]), .A2(n1617), .B1(n1614), .B2(
        write1_in[18]), .C1(n1521), .C2(n[2950]), .Z(spin[18]) );
  AO222D1BWP12T U2238 ( .A1(write2_in[18]), .A2(n1552), .B1(n1549), .B2(
        write1_in[18]), .C1(n1506), .C2(r0[18]), .Z(n2635) );
  AO222D1BWP12T U2239 ( .A1(write2_in[18]), .A2(n1609), .B1(n1607), .B2(
        write1_in[18]), .C1(n1608), .C2(lr[18]), .Z(n2219) );
  AO222D1BWP12T U2240 ( .A1(write2_in[18]), .A2(n1588), .B1(n1585), .B2(
        write1_in[18]), .C1(n1517), .C2(r1[18]), .Z(n2603) );
  AO222D1BWP12T U2241 ( .A1(write2_in[18]), .A2(n1513), .B1(n1512), .B2(
        write1_in[18]), .C1(n1511), .C2(r2[18]), .Z(n2571) );
  AO222D1BWP12T U2242 ( .A1(write2_in[18]), .A2(n1510), .B1(n1509), .B2(
        write1_in[18]), .C1(n1508), .C2(r11[18]), .Z(n2283) );
  AO222D1BWP12T U2243 ( .A1(write2_in[18]), .A2(n1594), .B1(n1591), .B2(
        write1_in[18]), .C1(n1507), .C2(r9[18]), .Z(n2347) );
  AO222D1BWP12T U2244 ( .A1(write2_in[18]), .A2(n1516), .B1(n1515), .B2(
        write1_in[18]), .C1(n1514), .C2(r10[18]), .Z(n2315) );
  AO222D1BWP12T U2245 ( .A1(write2_in[18]), .A2(n1570), .B1(n1567), .B2(
        write1_in[18]), .C1(n1505), .C2(r7[18]), .Z(n2411) );
  AO222D1BWP12T U2246 ( .A1(write2_in[18]), .A2(n1582), .B1(n1579), .B2(
        write1_in[18]), .C1(n1518), .C2(r4[18]), .Z(n2507) );
  AO222D1BWP12T U2247 ( .A1(write2_in[18]), .A2(n1599), .B1(n1597), .B2(
        write1_in[18]), .C1(n1598), .C2(r12[18]), .Z(n2251) );
  AO222D1BWP12T U2248 ( .A1(write2_in[18]), .A2(n1604), .B1(n1602), .B2(
        write1_in[18]), .C1(n1603), .C2(r8[18]), .Z(n2379) );
  AO222D1BWP12T U2249 ( .A1(write2_in[18]), .A2(n1558), .B1(n1555), .B2(
        write1_in[18]), .C1(n1519), .C2(r6[18]), .Z(n2443) );
  AO222D1BWP12T U2250 ( .A1(write2_in[18]), .A2(n1564), .B1(n1561), .B2(
        write1_in[18]), .C1(n1520), .C2(r5[18]), .Z(n2475) );
  AO222D1BWP12T U2251 ( .A1(write2_in[18]), .A2(n1576), .B1(n1573), .B2(
        write1_in[18]), .C1(n1504), .C2(r3[18]), .Z(n2539) );
  AO222D1BWP12T U2252 ( .A1(write2_in[18]), .A2(n1625), .B1(n1620), .B2(
        write1_in[18]), .C1(n1622), .C2(tmp1[18]), .Z(n2155) );
  AN2XD0BWP12T U2253 ( .A1(write2_in[8]), .A2(n2916), .Z(n1419) );
  AOI21D1BWP12T U2254 ( .A1(write1_in[8]), .A2(n2920), .B(n1419), .ZN(n1427)
         );
  ND2D2BWP12T U2255 ( .A1(n1421), .A2(n1420), .ZN(n1425) );
  AN2XD0BWP12T U2256 ( .A1(write2_in[9]), .A2(n2916), .Z(n1422) );
  AOI21D1BWP12T U2257 ( .A1(write1_in[9]), .A2(n2920), .B(n1422), .ZN(n1426)
         );
  OAI222D1BWP12T U2258 ( .A1(n1423), .A2(n1532), .B1(n1533), .B2(n1537), .C1(
        n1530), .C2(n1972), .ZN(n2285) );
  INVD1BWP12T U2259 ( .I(r10[20]), .ZN(n2056) );
  OAI222D1BWP12T U2260 ( .A1(n1423), .A2(n1527), .B1(n1528), .B2(n1537), .C1(
        n1526), .C2(n2056), .ZN(n2317) );
  INVD1BWP12T U2261 ( .I(r2[20]), .ZN(n2061) );
  OAI222D1BWP12T U2262 ( .A1(n1423), .A2(n1523), .B1(n1524), .B2(n1537), .C1(
        n1522), .C2(n2061), .ZN(n2573) );
  AO222D1BWP12T U2263 ( .A1(write1_in[21]), .A2(n1620), .B1(write2_in[21]), 
        .B2(n1625), .C1(n1622), .C2(tmp1[21]), .Z(n2158) );
  AO222D1BWP12T U2264 ( .A1(write2_in[20]), .A2(n1625), .B1(n1620), .B2(
        write1_in[20]), .C1(n1622), .C2(tmp1[20]), .Z(n2157) );
  AO222D1BWP12T U2265 ( .A1(write2_in[19]), .A2(n1510), .B1(n1509), .B2(
        write1_in[19]), .C1(n1508), .C2(r11[19]), .Z(n2284) );
  AO222D1BWP12T U2266 ( .A1(write2_in[19]), .A2(n1558), .B1(n1555), .B2(
        write1_in[19]), .C1(n1519), .C2(r6[19]), .Z(n2444) );
  AO222D1BWP12T U2267 ( .A1(write2_in[19]), .A2(n1513), .B1(n1512), .B2(
        write1_in[19]), .C1(n1511), .C2(r2[19]), .Z(n2572) );
  AO222D1BWP12T U2268 ( .A1(write2_in[19]), .A2(n1516), .B1(n1515), .B2(
        write1_in[19]), .C1(n1514), .C2(r10[19]), .Z(n2316) );
  AO222D1BWP12T U2269 ( .A1(write2_in[19]), .A2(n1609), .B1(n1607), .B2(
        write1_in[19]), .C1(n1608), .C2(lr[19]), .Z(n2220) );
  AO222D1BWP12T U2270 ( .A1(write2_in[19]), .A2(n1576), .B1(n1573), .B2(
        write1_in[19]), .C1(n1504), .C2(r3[19]), .Z(n2540) );
  AO222D1BWP12T U2271 ( .A1(write2_in[19]), .A2(n1604), .B1(n1602), .B2(
        write1_in[19]), .C1(n1603), .C2(r8[19]), .Z(n2380) );
  AO222D1BWP12T U2272 ( .A1(write2_in[19]), .A2(n1617), .B1(n1614), .B2(
        write1_in[19]), .C1(n1521), .C2(n[2949]), .Z(spin[19]) );
  AO222D1BWP12T U2273 ( .A1(write2_in[19]), .A2(n1564), .B1(n1561), .B2(
        write1_in[19]), .C1(n1520), .C2(r5[19]), .Z(n2476) );
  AO222D1BWP12T U2274 ( .A1(write2_in[19]), .A2(n1594), .B1(n1591), .B2(
        write1_in[19]), .C1(n1507), .C2(r9[19]), .Z(n2348) );
  AO222D1BWP12T U2275 ( .A1(write2_in[19]), .A2(n1552), .B1(n1549), .B2(
        write1_in[19]), .C1(n1506), .C2(r0[19]), .Z(n2636) );
  AO222D1BWP12T U2276 ( .A1(write2_in[19]), .A2(n1582), .B1(n1579), .B2(
        write1_in[19]), .C1(n1518), .C2(r4[19]), .Z(n2508) );
  AO222D1BWP12T U2277 ( .A1(write2_in[19]), .A2(n1570), .B1(n1567), .B2(
        write1_in[19]), .C1(n1505), .C2(r7[19]), .Z(n2412) );
  AO222D1BWP12T U2278 ( .A1(write2_in[19]), .A2(n1588), .B1(n1585), .B2(
        write1_in[19]), .C1(n1517), .C2(r1[19]), .Z(n2604) );
  AO222D1BWP12T U2279 ( .A1(write2_in[19]), .A2(n1599), .B1(n1597), .B2(
        write1_in[19]), .C1(n1598), .C2(r12[19]), .Z(n2252) );
  AO222D1BWP12T U2280 ( .A1(write2_in[19]), .A2(n1625), .B1(n1620), .B2(
        write1_in[19]), .C1(n1622), .C2(tmp1[19]), .Z(n2156) );
  CKND2D0BWP12T U2281 ( .A1(write2_in[10]), .A2(n2916), .ZN(n1424) );
  IOA21D1BWP12T U2282 ( .A1(write1_in[10]), .A2(n2920), .B(n1424), .ZN(n1432)
         );
  TPNR3D2BWP12T U2283 ( .A1(n1427), .A2(n1426), .A3(n1425), .ZN(n1433) );
  XOR2XD1BWP12T U2284 ( .A1(n1432), .A2(n1433), .Z(n1428) );
  AO222D1BWP12T U2285 ( .A1(n1428), .A2(n2914), .B1(n1488), .B2(next_pc_in[10]), .C1(n1690), .C2(pc_out[10]), .Z(n2179) );
  INVD1BWP12T U2286 ( .I(write2_in[23]), .ZN(n1649) );
  CKND1BWP12T U2287 ( .I(write1_in[23]), .ZN(n1431) );
  OAI222D1BWP12T U2288 ( .A1(n1524), .A2(n1649), .B1(n1523), .B2(n1431), .C1(
        n1522), .C2(n1429), .ZN(n2576) );
  INVD1BWP12T U2289 ( .I(r11[23]), .ZN(n2865) );
  OAI222D1BWP12T U2290 ( .A1(n1533), .A2(n1649), .B1(n1532), .B2(n1431), .C1(
        n1530), .C2(n2865), .ZN(n2288) );
  OAI222D1BWP12T U2291 ( .A1(n1528), .A2(n1649), .B1(n1527), .B2(n1431), .C1(
        n1526), .C2(n1430), .ZN(n2320) );
  TPND2D2BWP12T U2292 ( .A1(n1433), .A2(n1432), .ZN(n1467) );
  AN2XD0BWP12T U2293 ( .A1(write2_in[11]), .A2(n2916), .Z(n1434) );
  BUFFD6BWP12T U2294 ( .I(write1_in[24]), .Z(n1674) );
  AO222D1BWP12T U2295 ( .A1(n1674), .A2(n1573), .B1(write2_in[24]), .B2(n1576), 
        .C1(n1504), .C2(r3[24]), .Z(n2545) );
  AO222D1BWP12T U2296 ( .A1(n1674), .A2(n1515), .B1(write2_in[24]), .B2(n1516), 
        .C1(n1514), .C2(r10[24]), .Z(n2321) );
  AO222D1BWP12T U2297 ( .A1(n1674), .A2(n1512), .B1(write2_in[24]), .B2(n1513), 
        .C1(n1511), .C2(r2[24]), .Z(n2577) );
  AO222D1BWP12T U2298 ( .A1(n1674), .A2(n1509), .B1(write2_in[24]), .B2(n1510), 
        .C1(n1508), .C2(r11[24]), .Z(n2289) );
  AO222D1BWP12T U2299 ( .A1(n1674), .A2(n1602), .B1(write2_in[24]), .B2(n1604), 
        .C1(n1603), .C2(r8[24]), .Z(n2385) );
  AO222D1BWP12T U2300 ( .A1(n1674), .A2(n1561), .B1(write2_in[24]), .B2(n1564), 
        .C1(n1520), .C2(r5[24]), .Z(n2481) );
  AO222D1BWP12T U2301 ( .A1(n1674), .A2(n1591), .B1(write2_in[24]), .B2(n1594), 
        .C1(n1507), .C2(r9[24]), .Z(n2353) );
  AO222D1BWP12T U2302 ( .A1(n1674), .A2(n1549), .B1(write2_in[24]), .B2(n1552), 
        .C1(n1506), .C2(r0[24]), .Z(n2641) );
  AO222D1BWP12T U2303 ( .A1(n1674), .A2(n1585), .B1(write2_in[24]), .B2(n1588), 
        .C1(n1517), .C2(r1[24]), .Z(n2609) );
  AO222D1BWP12T U2304 ( .A1(n1674), .A2(n1567), .B1(write2_in[24]), .B2(n1570), 
        .C1(n1505), .C2(r7[24]), .Z(n2417) );
  AO222D1BWP12T U2305 ( .A1(n1674), .A2(n1579), .B1(write2_in[24]), .B2(n1582), 
        .C1(n1518), .C2(r4[24]), .Z(n2513) );
  AO222D1BWP12T U2306 ( .A1(n1674), .A2(n1597), .B1(write2_in[24]), .B2(n1599), 
        .C1(n1598), .C2(r12[24]), .Z(n2257) );
  AO222D1BWP12T U2307 ( .A1(n1674), .A2(n1607), .B1(write2_in[24]), .B2(n1609), 
        .C1(n1608), .C2(lr[24]), .Z(n2225) );
  AO222D1BWP12T U2308 ( .A1(n1674), .A2(n1555), .B1(write2_in[24]), .B2(n1558), 
        .C1(n1519), .C2(r6[24]), .Z(n2449) );
  AO222D1BWP12T U2309 ( .A1(n1674), .A2(n1614), .B1(write2_in[24]), .B2(n1617), 
        .C1(n1521), .C2(n[2944]), .Z(spin[24]) );
  AO222D1BWP12T U2310 ( .A1(n1674), .A2(n1620), .B1(write2_in[24]), .B2(n1625), 
        .C1(n1622), .C2(tmp1[24]), .Z(n2161) );
  INVD1BWP12T U2311 ( .I(write2_in[21]), .ZN(n1651) );
  INVD1BWP12T U2312 ( .I(r12[21]), .ZN(n2036) );
  OAI222D1BWP12T U2313 ( .A1(n1437), .A2(n1651), .B1(n1436), .B2(n1456), .C1(
        n1435), .C2(n2036), .ZN(n2254) );
  INVD1BWP12T U2314 ( .I(lr[21]), .ZN(n2050) );
  OAI222D1BWP12T U2315 ( .A1(n1439), .A2(n1651), .B1(n1475), .B2(n1456), .C1(
        n1438), .C2(n2050), .ZN(n2222) );
  INVD1BWP12T U2316 ( .I(r8[21]), .ZN(n2049) );
  OAI222D1BWP12T U2317 ( .A1(n1441), .A2(n1651), .B1(n1478), .B2(n1456), .C1(
        n1440), .C2(n2049), .ZN(n2382) );
  INVD1BWP12T U2318 ( .I(r10[21]), .ZN(n2048) );
  OAI222D1BWP12T U2319 ( .A1(n1528), .A2(n1651), .B1(n1527), .B2(n1456), .C1(
        n1526), .C2(n2048), .ZN(n2318) );
  INVD1BWP12T U2320 ( .I(r2[21]), .ZN(n1841) );
  OAI222D1BWP12T U2321 ( .A1(n1524), .A2(n1651), .B1(n1523), .B2(n1456), .C1(
        n1522), .C2(n1841), .ZN(n2574) );
  INVD1BWP12T U2322 ( .I(r11[21]), .ZN(n2031) );
  OAI222D1BWP12T U2323 ( .A1(n1533), .A2(n1651), .B1(n1532), .B2(n1456), .C1(
        n1530), .C2(n2031), .ZN(n2286) );
  AO222D1BWP12T U2324 ( .A1(write1_in[23]), .A2(n1602), .B1(write2_in[23]), 
        .B2(n1604), .C1(n1603), .C2(r8[23]), .Z(n2384) );
  AO222D1BWP12T U2325 ( .A1(write1_in[23]), .A2(n1573), .B1(write2_in[23]), 
        .B2(n1576), .C1(n1504), .C2(r3[23]), .Z(n2544) );
  AO222D1BWP12T U2326 ( .A1(write1_in[23]), .A2(n1561), .B1(write2_in[23]), 
        .B2(n1564), .C1(n1520), .C2(r5[23]), .Z(n2480) );
  AO222D1BWP12T U2327 ( .A1(write1_in[23]), .A2(n1579), .B1(write2_in[23]), 
        .B2(n1582), .C1(n1518), .C2(r4[23]), .Z(n2512) );
  AO222D1BWP12T U2328 ( .A1(write1_in[23]), .A2(n1585), .B1(write2_in[23]), 
        .B2(n1588), .C1(n1517), .C2(r1[23]), .Z(n2608) );
  AO222D1BWP12T U2329 ( .A1(write1_in[23]), .A2(n1591), .B1(write2_in[23]), 
        .B2(n1594), .C1(n1507), .C2(r9[23]), .Z(n2352) );
  INVD1BWP12T U2330 ( .I(n[2947]), .ZN(n2032) );
  OAI222D1BWP12T U2331 ( .A1(n1443), .A2(n1651), .B1(n1442), .B2(n1456), .C1(
        n1615), .C2(n2032), .ZN(spin[21]) );
  INVD1BWP12T U2332 ( .I(r6[21]), .ZN(n2047) );
  OAI222D1BWP12T U2333 ( .A1(n1444), .A2(n1651), .B1(n1490), .B2(n1456), .C1(
        n1556), .C2(n2047), .ZN(n2446) );
  INVD1BWP12T U2334 ( .I(r5[21]), .ZN(n2030) );
  OAI222D1BWP12T U2335 ( .A1(n1446), .A2(n1651), .B1(n1445), .B2(n1456), .C1(
        n1562), .C2(n2030), .ZN(n2478) );
  INVD1BWP12T U2336 ( .I(r1[21]), .ZN(n2035) );
  OAI222D1BWP12T U2337 ( .A1(n1448), .A2(n1651), .B1(n1447), .B2(n1456), .C1(
        n1586), .C2(n2035), .ZN(n2606) );
  INVD1BWP12T U2338 ( .I(r4[21]), .ZN(n2044) );
  OAI222D1BWP12T U2339 ( .A1(n1450), .A2(n1651), .B1(n1449), .B2(n1456), .C1(
        n1580), .C2(n2044), .ZN(n2510) );
  INVD1BWP12T U2340 ( .I(r7[21]), .ZN(n2033) );
  OAI222D1BWP12T U2341 ( .A1(n1452), .A2(n1651), .B1(n1451), .B2(n1456), .C1(
        n1568), .C2(n2033), .ZN(n2414) );
  INVD1BWP12T U2342 ( .I(r9[21]), .ZN(n2042) );
  OAI222D1BWP12T U2343 ( .A1(n1453), .A2(n1651), .B1(n1481), .B2(n1456), .C1(
        n1592), .C2(n2042), .ZN(n2350) );
  INVD1BWP12T U2344 ( .I(r0[21]), .ZN(n2043) );
  OAI222D1BWP12T U2345 ( .A1(n1455), .A2(n1651), .B1(n1454), .B2(n1456), .C1(
        n1550), .C2(n2043), .ZN(n2638) );
  INVD1BWP12T U2346 ( .I(r3[21]), .ZN(n2029) );
  OAI222D1BWP12T U2347 ( .A1(n1458), .A2(n1651), .B1(n1457), .B2(n1456), .C1(
        n1574), .C2(n2029), .ZN(n2542) );
  AO222D1BWP12T U2348 ( .A1(write1_in[22]), .A2(n1602), .B1(write2_in[22]), 
        .B2(n1604), .C1(n1603), .C2(r8[22]), .Z(n2383) );
  AO222D1BWP12T U2349 ( .A1(write1_in[22]), .A2(n1573), .B1(write2_in[22]), 
        .B2(n1576), .C1(n1504), .C2(r3[22]), .Z(n2543) );
  AO222D1BWP12T U2350 ( .A1(write1_in[22]), .A2(n1561), .B1(write2_in[22]), 
        .B2(n1564), .C1(n1520), .C2(r5[22]), .Z(n2479) );
  AO222D1BWP12T U2351 ( .A1(write1_in[22]), .A2(n1549), .B1(write2_in[22]), 
        .B2(n1552), .C1(n1506), .C2(r0[22]), .Z(n2639) );
  AO222D1BWP12T U2352 ( .A1(write1_in[22]), .A2(n1591), .B1(write2_in[22]), 
        .B2(n1594), .C1(n1507), .C2(r9[22]), .Z(n2351) );
  AO222D1BWP12T U2353 ( .A1(write1_in[22]), .A2(n1585), .B1(write2_in[22]), 
        .B2(n1588), .C1(n1517), .C2(r1[22]), .Z(n2607) );
  AO222D1BWP12T U2354 ( .A1(write1_in[22]), .A2(n1567), .B1(write2_in[22]), 
        .B2(n1570), .C1(n1505), .C2(r7[22]), .Z(n2415) );
  AO222D1BWP12T U2355 ( .A1(write1_in[22]), .A2(n1579), .B1(write2_in[22]), 
        .B2(n1582), .C1(n1518), .C2(r4[22]), .Z(n2511) );
  AO222D1BWP12T U2356 ( .A1(write1_in[22]), .A2(n1597), .B1(write2_in[22]), 
        .B2(n1599), .C1(n1598), .C2(r12[22]), .Z(n2255) );
  AO222D1BWP12T U2357 ( .A1(write1_in[22]), .A2(n1607), .B1(write2_in[22]), 
        .B2(n1609), .C1(n1608), .C2(lr[22]), .Z(n2223) );
  AO222D1BWP12T U2358 ( .A1(write1_in[22]), .A2(n1555), .B1(write2_in[22]), 
        .B2(n1558), .C1(n1519), .C2(r6[22]), .Z(n2447) );
  AO222D1BWP12T U2359 ( .A1(write1_in[22]), .A2(n1614), .B1(write2_in[22]), 
        .B2(n1617), .C1(n1521), .C2(n[2946]), .Z(spin[22]) );
  AO222D1BWP12T U2360 ( .A1(write1_in[22]), .A2(n1620), .B1(write2_in[22]), 
        .B2(n1625), .C1(n1622), .C2(tmp1[22]), .Z(n2159) );
  AN2XD0BWP12T U2361 ( .A1(write2_in[12]), .A2(n2916), .Z(n1459) );
  AOI21D2BWP12T U2362 ( .A1(write1_in[12]), .A2(n2920), .B(n1459), .ZN(n1466)
         );
  INVD1BWP12T U2363 ( .I(write2_in[22]), .ZN(n1652) );
  INVD1BWP12T U2364 ( .I(write1_in[22]), .ZN(n1463) );
  OAI222D1BWP12T U2365 ( .A1(n1528), .A2(n1652), .B1(n1527), .B2(n1463), .C1(
        n1526), .C2(n1460), .ZN(n2319) );
  OAI222D1BWP12T U2366 ( .A1(n1533), .A2(n1652), .B1(n1532), .B2(n1463), .C1(
        n1530), .C2(n1461), .ZN(n2287) );
  OAI222D1BWP12T U2367 ( .A1(n1524), .A2(n1652), .B1(n1523), .B2(n1463), .C1(
        n1522), .C2(n1462), .ZN(n2575) );
  CKND2D0BWP12T U2368 ( .A1(write2_in[13]), .A2(n2916), .ZN(n1464) );
  IOA21D2BWP12T U2369 ( .A1(write1_in[13]), .A2(n2920), .B(n1464), .ZN(n1469)
         );
  TPNR3D4BWP12T U2370 ( .A1(n1467), .A2(n1466), .A3(n1465), .ZN(n1468) );
  AO222D1BWP12T U2371 ( .A1(write1_in[26]), .A2(n1515), .B1(write2_in[26]), 
        .B2(n1516), .C1(n1514), .C2(r10[26]), .Z(n2323) );
  AO222D1BWP12T U2372 ( .A1(write1_in[26]), .A2(n1602), .B1(write2_in[26]), 
        .B2(n1604), .C1(n1603), .C2(r8[26]), .Z(n2387) );
  AO222D1BWP12T U2373 ( .A1(write1_in[26]), .A2(n1512), .B1(write2_in[26]), 
        .B2(n1513), .C1(n1511), .C2(r2[26]), .Z(n2579) );
  AO222D1BWP12T U2374 ( .A1(write1_in[26]), .A2(n1509), .B1(write2_in[26]), 
        .B2(n1510), .C1(n1508), .C2(r11[26]), .Z(n2291) );
  AO222D1BWP12T U2375 ( .A1(write1_in[26]), .A2(n1573), .B1(write2_in[26]), 
        .B2(n1576), .C1(n1504), .C2(r3[26]), .Z(n2547) );
  AO222D1BWP12T U2376 ( .A1(write1_in[26]), .A2(n1549), .B1(write2_in[26]), 
        .B2(n1552), .C1(n1506), .C2(r0[26]), .Z(n2643) );
  AO222D1BWP12T U2377 ( .A1(write1_in[26]), .A2(n1561), .B1(write2_in[26]), 
        .B2(n1564), .C1(n1520), .C2(r5[26]), .Z(n2483) );
  AO222D1BWP12T U2378 ( .A1(write1_in[26]), .A2(n1591), .B1(write2_in[26]), 
        .B2(n1594), .C1(n1507), .C2(r9[26]), .Z(n2355) );
  AO222D1BWP12T U2379 ( .A1(write1_in[26]), .A2(n1579), .B1(write2_in[26]), 
        .B2(n1582), .C1(n1518), .C2(r4[26]), .Z(n2515) );
  AO222D1BWP12T U2380 ( .A1(write1_in[26]), .A2(n1585), .B1(write2_in[26]), 
        .B2(n1588), .C1(n1517), .C2(r1[26]), .Z(n2611) );
  AO222D1BWP12T U2381 ( .A1(write1_in[26]), .A2(n1567), .B1(write2_in[26]), 
        .B2(n1570), .C1(n1505), .C2(r7[26]), .Z(n2419) );
  AO222D1BWP12T U2382 ( .A1(write1_in[26]), .A2(n1597), .B1(write2_in[26]), 
        .B2(n1599), .C1(n1598), .C2(r12[26]), .Z(n2259) );
  AO222D1BWP12T U2383 ( .A1(write1_in[26]), .A2(n1607), .B1(write2_in[26]), 
        .B2(n1609), .C1(n1608), .C2(lr[26]), .Z(n2227) );
  AO222D1BWP12T U2384 ( .A1(write1_in[26]), .A2(n1555), .B1(write2_in[26]), 
        .B2(n1558), .C1(n1519), .C2(r6[26]), .Z(n2451) );
  AO222D1BWP12T U2385 ( .A1(write1_in[26]), .A2(n1614), .B1(write2_in[26]), 
        .B2(n1617), .C1(n1521), .C2(n[2942]), .Z(spin[26]) );
  AO222D1BWP12T U2386 ( .A1(write1_in[26]), .A2(n1620), .B1(write2_in[26]), 
        .B2(n1625), .C1(n1622), .C2(tmp1[26]), .Z(n2163) );
  TPND2D3BWP12T U2387 ( .A1(n1469), .A2(n1468), .ZN(n1494) );
  CKAN2D1BWP12T U2388 ( .A1(write2_in[14]), .A2(n2916), .Z(n1470) );
  TPAOI21D4BWP12T U2389 ( .A1(n1471), .A2(n2920), .B(n1470), .ZN(n1493) );
  AOI22D0BWP12T U2390 ( .A1(write2_in[29]), .A2(n1510), .B1(r11[29]), .B2(
        n1508), .ZN(n1472) );
  OAI21D1BWP12T U2391 ( .A1(n1482), .A2(n1532), .B(n1472), .ZN(n2294) );
  AOI22D0BWP12T U2392 ( .A1(write2_in[29]), .A2(n1558), .B1(r6[29]), .B2(n1519), .ZN(n1473) );
  OAI21D1BWP12T U2393 ( .A1(n1482), .A2(n1490), .B(n1473), .ZN(n2454) );
  AOI22D0BWP12T U2394 ( .A1(write2_in[29]), .A2(n1609), .B1(lr[29]), .B2(n1608), .ZN(n1474) );
  OAI21D1BWP12T U2395 ( .A1(n1482), .A2(n1475), .B(n1474), .ZN(n2230) );
  AOI22D0BWP12T U2396 ( .A1(write2_in[29]), .A2(n1513), .B1(r2[29]), .B2(n1511), .ZN(n1476) );
  OAI21D1BWP12T U2397 ( .A1(n1482), .A2(n1523), .B(n1476), .ZN(n2582) );
  AOI22D0BWP12T U2398 ( .A1(write2_in[29]), .A2(n1604), .B1(r8[29]), .B2(n1603), .ZN(n1477) );
  OAI21D1BWP12T U2399 ( .A1(n1482), .A2(n1478), .B(n1477), .ZN(n2390) );
  AOI22D0BWP12T U2400 ( .A1(write2_in[29]), .A2(n1516), .B1(r10[29]), .B2(
        n1514), .ZN(n1479) );
  OAI21D1BWP12T U2401 ( .A1(n1482), .A2(n1527), .B(n1479), .ZN(n2326) );
  AOI22D0BWP12T U2402 ( .A1(write2_in[29]), .A2(n1594), .B1(r9[29]), .B2(n1507), .ZN(n1480) );
  OAI21D1BWP12T U2403 ( .A1(n1482), .A2(n1481), .B(n1480), .ZN(n2358) );
  INVD1BWP12T U2404 ( .I(write2_in[27]), .ZN(n1731) );
  INVD1BWP12T U2405 ( .I(write1_in[27]), .ZN(n1486) );
  OAI222D1BWP12T U2406 ( .A1(n1524), .A2(n1731), .B1(n1523), .B2(n1486), .C1(
        n1522), .C2(n1483), .ZN(n2580) );
  CKND0BWP12T U2407 ( .I(r10[27]), .ZN(n1484) );
  OAI222D1BWP12T U2408 ( .A1(n1528), .A2(n1731), .B1(n1527), .B2(n1486), .C1(
        n1526), .C2(n1484), .ZN(n2324) );
  OAI222D1BWP12T U2409 ( .A1(n1533), .A2(n1731), .B1(n1532), .B2(n1486), .C1(
        n1530), .C2(n1485), .ZN(n2292) );
  CKAN2D1BWP12T U2410 ( .A1(write2_in[15]), .A2(n2916), .Z(n1487) );
  AOI21D2BWP12T U2411 ( .A1(write1_in[15]), .A2(n2920), .B(n1487), .ZN(n1492)
         );
  AOI22D0BWP12T U2412 ( .A1(write2_in[30]), .A2(n1558), .B1(n1519), .B2(r6[30]), .ZN(n1489) );
  OAI21D1BWP12T U2413 ( .A1(n1491), .A2(n1490), .B(n1489), .ZN(n2455) );
  AO222D1BWP12T U2414 ( .A1(write1_in[27]), .A2(n1602), .B1(write2_in[27]), 
        .B2(n1604), .C1(n1603), .C2(r8[27]), .Z(n2388) );
  AO222D1BWP12T U2415 ( .A1(write1_in[27]), .A2(n1573), .B1(write2_in[27]), 
        .B2(n1576), .C1(n1504), .C2(r3[27]), .Z(n2548) );
  AO222D1BWP12T U2416 ( .A1(write1_in[27]), .A2(n1561), .B1(write2_in[27]), 
        .B2(n1564), .C1(n1520), .C2(r5[27]), .Z(n2484) );
  AO222D1BWP12T U2417 ( .A1(write1_in[27]), .A2(n1549), .B1(write2_in[27]), 
        .B2(n1552), .C1(n1506), .C2(r0[27]), .Z(n2644) );
  AO222D1BWP12T U2418 ( .A1(write1_in[27]), .A2(n1567), .B1(write2_in[27]), 
        .B2(n1570), .C1(n1505), .C2(r7[27]), .Z(n2420) );
  AO222D1BWP12T U2419 ( .A1(write1_in[27]), .A2(n1579), .B1(write2_in[27]), 
        .B2(n1582), .C1(n1518), .C2(r4[27]), .Z(n2516) );
  AO222D1BWP12T U2420 ( .A1(write1_in[27]), .A2(n1585), .B1(write2_in[27]), 
        .B2(n1588), .C1(n1517), .C2(r1[27]), .Z(n2612) );
  AO222D1BWP12T U2421 ( .A1(write1_in[27]), .A2(n1597), .B1(write2_in[27]), 
        .B2(n1599), .C1(n1598), .C2(r12[27]), .Z(n2260) );
  AO222D1BWP12T U2422 ( .A1(write1_in[27]), .A2(n1607), .B1(write2_in[27]), 
        .B2(n1609), .C1(n1608), .C2(lr[27]), .Z(n2228) );
  AO222D1BWP12T U2423 ( .A1(write1_in[27]), .A2(n1555), .B1(write2_in[27]), 
        .B2(n1558), .C1(n1519), .C2(r6[27]), .Z(n2452) );
  AO222D1BWP12T U2424 ( .A1(write1_in[27]), .A2(n1614), .B1(write2_in[27]), 
        .B2(n1617), .C1(n1521), .C2(n[2941]), .Z(spin[27]) );
  AO222D1BWP12T U2425 ( .A1(write1_in[27]), .A2(n1620), .B1(write2_in[27]), 
        .B2(n1625), .C1(n1622), .C2(tmp1[27]), .Z(n2164) );
  CKAN2D1BWP12T U2426 ( .A1(write2_in[16]), .A2(n2916), .Z(n1495) );
  AOI21D2BWP12T U2427 ( .A1(n1496), .A2(n2920), .B(n1495), .ZN(n1534) );
  AOI21D0BWP12T U2428 ( .A1(write2_in[18]), .A2(write2_in[17]), .B(n2920), 
        .ZN(n1497) );
  AOI21D1BWP12T U2429 ( .A1(n1498), .A2(n2920), .B(n1497), .ZN(n1501) );
  NR2D1BWP12T U2430 ( .A1(write1_in[18]), .A2(n2916), .ZN(n1499) );
  TPNR2D1BWP12T U2431 ( .A1(n1499), .A2(n1534), .ZN(n1500) );
  CKND2D2BWP12T U2432 ( .A1(n1501), .A2(n1500), .ZN(n1541) );
  CKND2D2BWP12T U2433 ( .A1(write1_in[19]), .A2(n2920), .ZN(n1503) );
  CKND2D0BWP12T U2434 ( .A1(write2_in[19]), .A2(n2916), .ZN(n1502) );
  ND2D2BWP12T U2435 ( .A1(n1503), .A2(n1502), .ZN(n1545) );
  AO222D1BWP12T U2436 ( .A1(write2_in[25]), .A2(n1576), .B1(n1573), .B2(
        write1_in[25]), .C1(n1504), .C2(r3[25]), .Z(n2546) );
  AO222D1BWP12T U2437 ( .A1(write2_in[25]), .A2(n1599), .B1(n1597), .B2(
        write1_in[25]), .C1(n1598), .C2(r12[25]), .Z(n2258) );
  AO222D1BWP12T U2438 ( .A1(write2_in[25]), .A2(n1570), .B1(n1567), .B2(
        write1_in[25]), .C1(n1505), .C2(r7[25]), .Z(n2418) );
  AO222D1BWP12T U2439 ( .A1(write2_in[25]), .A2(n1552), .B1(n1549), .B2(
        write1_in[25]), .C1(n1506), .C2(r0[25]), .Z(n2642) );
  AO222D1BWP12T U2440 ( .A1(write2_in[25]), .A2(n1594), .B1(n1591), .B2(
        write1_in[25]), .C1(n1507), .C2(r9[25]), .Z(n2354) );
  AO222D1BWP12T U2441 ( .A1(write2_in[25]), .A2(n1510), .B1(n1509), .B2(
        write1_in[25]), .C1(n1508), .C2(r11[25]), .Z(n2290) );
  AO222D1BWP12T U2442 ( .A1(write2_in[25]), .A2(n1513), .B1(n1512), .B2(
        write1_in[25]), .C1(n1511), .C2(r2[25]), .Z(n2578) );
  AO222D1BWP12T U2443 ( .A1(write2_in[25]), .A2(n1516), .B1(n1515), .B2(
        write1_in[25]), .C1(n1514), .C2(r10[25]), .Z(n2322) );
  AO222D1BWP12T U2444 ( .A1(write2_in[25]), .A2(n1609), .B1(n1607), .B2(
        write1_in[25]), .C1(n1608), .C2(lr[25]), .Z(n2226) );
  AO222D1BWP12T U2445 ( .A1(write2_in[25]), .A2(n1588), .B1(n1585), .B2(
        write1_in[25]), .C1(n1517), .C2(r1[25]), .Z(n2610) );
  AO222D1BWP12T U2446 ( .A1(write2_in[25]), .A2(n1604), .B1(n1602), .B2(
        write1_in[25]), .C1(n1603), .C2(r8[25]), .Z(n2386) );
  AO222D1BWP12T U2447 ( .A1(write2_in[25]), .A2(n1582), .B1(n1579), .B2(
        write1_in[25]), .C1(n1518), .C2(r4[25]), .Z(n2514) );
  AO222D1BWP12T U2448 ( .A1(write2_in[25]), .A2(n1625), .B1(n1620), .B2(
        write1_in[25]), .C1(n1622), .C2(tmp1[25]), .Z(n2162) );
  AO222D1BWP12T U2449 ( .A1(write2_in[25]), .A2(n1558), .B1(n1555), .B2(
        write1_in[25]), .C1(n1519), .C2(r6[25]), .Z(n2450) );
  AO222D1BWP12T U2450 ( .A1(write2_in[25]), .A2(n1564), .B1(n1561), .B2(
        write1_in[25]), .C1(n1520), .C2(r5[25]), .Z(n2482) );
  AO222D1BWP12T U2451 ( .A1(write2_in[25]), .A2(n1617), .B1(n1614), .B2(
        write1_in[25]), .C1(n1521), .C2(n[2943]), .Z(spin[25]) );
  INVD1BWP12T U2452 ( .I(write2_in[31]), .ZN(n1665) );
  INVD1BWP12T U2453 ( .I(write1_in[31]), .ZN(n1531) );
  INVD1BWP12T U2454 ( .I(r2[31]), .ZN(n1756) );
  OAI222D1BWP12T U2455 ( .A1(n1524), .A2(n1665), .B1(n1523), .B2(n1531), .C1(
        n1522), .C2(n1756), .ZN(n2584) );
  OAI222D1BWP12T U2456 ( .A1(n1528), .A2(n1665), .B1(n1527), .B2(n1531), .C1(
        n1526), .C2(n1525), .ZN(n2328) );
  CKND0BWP12T U2457 ( .I(r11[31]), .ZN(n1529) );
  OAI222D1BWP12T U2458 ( .A1(n1533), .A2(n1665), .B1(n1532), .B2(n1531), .C1(
        n1530), .C2(n1529), .ZN(n2296) );
  MUX2NXD0BWP12T U2459 ( .I0(write1_in[17]), .I1(write2_in[17]), .S(n2916), 
        .ZN(n1544) );
  XOR2XD1BWP12T U2460 ( .A1(n1544), .A2(n1543), .Z(n1536) );
  AO222D1BWP12T U2461 ( .A1(n1536), .A2(n2914), .B1(n1488), .B2(next_pc_in[17]), .C1(n1690), .C2(pc_out[17]), .Z(n2186) );
  CKND2D0BWP12T U2462 ( .A1(n1537), .A2(n2916), .ZN(n1538) );
  OAI21D1BWP12T U2463 ( .A1(write1_in[20]), .A2(n2916), .B(n1538), .ZN(n1539)
         );
  AN2XD0BWP12T U2464 ( .A1(write2_in[21]), .A2(n2916), .Z(n1542) );
  AOI21D1BWP12T U2465 ( .A1(write1_in[21]), .A2(n2920), .B(n1542), .ZN(n1630)
         );
  TPNR2D1BWP12T U2466 ( .A1(n1544), .A2(n1543), .ZN(n1613) );
  MUX2D1BWP12T U2467 ( .I0(write2_in[18]), .I1(write1_in[18]), .S(n2920), .Z(
        n1612) );
  CKND2D1BWP12T U2468 ( .A1(n1613), .A2(n1612), .ZN(n1546) );
  XOR2XD1BWP12T U2469 ( .A1(n1546), .A2(n1545), .Z(n1548) );
  AOI22D1BWP12T U2470 ( .A1(next_pc_in[19]), .A2(n1488), .B1(n1690), .B2(
        pc_out[19]), .ZN(n1547) );
  OAI21D1BWP12T U2471 ( .A1(n1548), .A2(n2919), .B(n1547), .ZN(n2188) );
  CKND2D1BWP12T U2472 ( .A1(n1621), .A2(n1549), .ZN(n1554) );
  INR2D0BWP12T U2473 ( .A1(r0[31]), .B1(n1550), .ZN(n1551) );
  AOI21D0BWP12T U2474 ( .A1(write2_in[31]), .A2(n1552), .B(n1551), .ZN(n1553)
         );
  ND2D1BWP12T U2475 ( .A1(n1554), .A2(n1553), .ZN(n2648) );
  CKND2D1BWP12T U2476 ( .A1(n1621), .A2(n1555), .ZN(n1560) );
  INR2D0BWP12T U2477 ( .A1(r6[31]), .B1(n1556), .ZN(n1557) );
  TPAOI21D0BWP12T U2478 ( .A1(write2_in[31]), .A2(n1558), .B(n1557), .ZN(n1559) );
  ND2D1BWP12T U2479 ( .A1(n1560), .A2(n1559), .ZN(n2456) );
  CKND2D1BWP12T U2480 ( .A1(n1621), .A2(n1561), .ZN(n1566) );
  INR2D0BWP12T U2481 ( .A1(r5[31]), .B1(n1562), .ZN(n1563) );
  AOI21D0BWP12T U2482 ( .A1(write2_in[31]), .A2(n1564), .B(n1563), .ZN(n1565)
         );
  ND2D1BWP12T U2483 ( .A1(n1566), .A2(n1565), .ZN(n2488) );
  CKND2D1BWP12T U2484 ( .A1(n1621), .A2(n1567), .ZN(n1572) );
  INR2D0BWP12T U2485 ( .A1(r7[31]), .B1(n1568), .ZN(n1569) );
  AOI21D0BWP12T U2486 ( .A1(write2_in[31]), .A2(n1570), .B(n1569), .ZN(n1571)
         );
  ND2D1BWP12T U2487 ( .A1(n1572), .A2(n1571), .ZN(n2424) );
  CKND2D1BWP12T U2488 ( .A1(n1621), .A2(n1573), .ZN(n1578) );
  INR2D0BWP12T U2489 ( .A1(r3[31]), .B1(n1574), .ZN(n1575) );
  AOI21D0BWP12T U2490 ( .A1(write2_in[31]), .A2(n1576), .B(n1575), .ZN(n1577)
         );
  ND2D1BWP12T U2491 ( .A1(n1578), .A2(n1577), .ZN(n2552) );
  CKND2D1BWP12T U2492 ( .A1(n1621), .A2(n1579), .ZN(n1584) );
  INR2D0BWP12T U2493 ( .A1(r4[31]), .B1(n1580), .ZN(n1581) );
  AOI21D0BWP12T U2494 ( .A1(write2_in[31]), .A2(n1582), .B(n1581), .ZN(n1583)
         );
  ND2D1BWP12T U2495 ( .A1(n1584), .A2(n1583), .ZN(n2520) );
  CKND2D1BWP12T U2496 ( .A1(n1621), .A2(n1585), .ZN(n1590) );
  INR2D0BWP12T U2497 ( .A1(r1[31]), .B1(n1586), .ZN(n1587) );
  AOI21D0BWP12T U2498 ( .A1(write2_in[31]), .A2(n1588), .B(n1587), .ZN(n1589)
         );
  ND2D1BWP12T U2499 ( .A1(n1590), .A2(n1589), .ZN(n2616) );
  CKND2D1BWP12T U2500 ( .A1(n1621), .A2(n1591), .ZN(n1596) );
  INR2D0BWP12T U2501 ( .A1(r9[31]), .B1(n1592), .ZN(n1593) );
  AOI21D0BWP12T U2502 ( .A1(write2_in[31]), .A2(n1594), .B(n1593), .ZN(n1595)
         );
  ND2D1BWP12T U2503 ( .A1(n1596), .A2(n1595), .ZN(n2360) );
  CKND2D1BWP12T U2504 ( .A1(n1621), .A2(n1597), .ZN(n1601) );
  AOI22D0BWP12T U2505 ( .A1(write2_in[31]), .A2(n1599), .B1(r12[31]), .B2(
        n1598), .ZN(n1600) );
  ND2D1BWP12T U2506 ( .A1(n1601), .A2(n1600), .ZN(n2264) );
  CKND2D1BWP12T U2507 ( .A1(n1621), .A2(n1602), .ZN(n1606) );
  AOI22D0BWP12T U2508 ( .A1(write2_in[31]), .A2(n1604), .B1(n1603), .B2(r8[31]), .ZN(n1605) );
  ND2D1BWP12T U2509 ( .A1(n1606), .A2(n1605), .ZN(n2392) );
  CKND2D1BWP12T U2510 ( .A1(n1621), .A2(n1607), .ZN(n1611) );
  AOI22D0BWP12T U2511 ( .A1(write2_in[31]), .A2(n1609), .B1(n1608), .B2(lr[31]), .ZN(n1610) );
  ND2D1BWP12T U2512 ( .A1(n1611), .A2(n1610), .ZN(n2232) );
  CKND2D1BWP12T U2513 ( .A1(n1621), .A2(n1614), .ZN(n1619) );
  INR2D0BWP12T U2514 ( .A1(n[2937]), .B1(n1615), .ZN(n1616) );
  AOI21D0BWP12T U2515 ( .A1(write2_in[31]), .A2(n1617), .B(n1616), .ZN(n1618)
         );
  ND2D1BWP12T U2516 ( .A1(n1619), .A2(n1618), .ZN(spin[31]) );
  CKND2D1BWP12T U2517 ( .A1(n1621), .A2(n1620), .ZN(n1627) );
  CKND0BWP12T U2518 ( .I(n1622), .ZN(n1623) );
  INR2XD0BWP12T U2519 ( .A1(tmp1[31]), .B1(n1623), .ZN(n1624) );
  AOI21D0BWP12T U2520 ( .A1(write2_in[31]), .A2(n1625), .B(n1624), .ZN(n1626)
         );
  ND2D1BWP12T U2521 ( .A1(n1627), .A2(n1626), .ZN(n2168) );
  CKND2D1BWP12T U2522 ( .A1(n1748), .A2(n2900), .ZN(n1636) );
  CKND0BWP12T U2523 ( .I(write2_in[24]), .ZN(n1628) );
  TPNR2D0BWP12T U2524 ( .A1(n1628), .A2(n2920), .ZN(n1629) );
  AOI21D1BWP12T U2525 ( .A1(n1674), .A2(n2920), .B(n1629), .ZN(n2906) );
  TPNR3D0BWP12T U2526 ( .A1(n1636), .A2(n2906), .A3(n2919), .ZN(n1632) );
  INVD2BWP12T U2527 ( .I(n1656), .ZN(n1631) );
  ND2XD0BWP12T U2528 ( .A1(write2_in[25]), .A2(n2916), .ZN(n1699) );
  INVD1BWP12T U2529 ( .I(n1699), .ZN(n1701) );
  AOI21D1BWP12T U2530 ( .A1(write1_in[25]), .A2(n2920), .B(n1701), .ZN(n1633)
         );
  TPND3D0BWP12T U2531 ( .A1(n1632), .A2(n1749), .A3(n1633), .ZN(n1641) );
  NR2D1BWP12T U2532 ( .A1(n1633), .A2(n2919), .ZN(n1637) );
  TPAOI21D0BWP12T U2533 ( .A1(n1637), .A2(n2906), .B(n1635), .ZN(n1640) );
  CKND2D1BWP12T U2534 ( .A1(n1638), .A2(n1637), .ZN(n1639) );
  ND3D1BWP12T U2535 ( .A1(n1641), .A2(n1640), .A3(n1639), .ZN(n2194) );
  AOI21D0BWP12T U2536 ( .A1(n2916), .A2(write2_in[31]), .B(n2919), .ZN(n1642)
         );
  OAI21D0BWP12T U2537 ( .A1(write2_in[30]), .A2(n2920), .B(n1642), .ZN(n1643)
         );
  RCAOI21D1BWP12T U2538 ( .A1(n2920), .A2(write1_in[31]), .B(n1643), .ZN(n1644) );
  INVD1P25BWP12T U2539 ( .I(n1674), .ZN(n1646) );
  TPNR2D1BWP12T U2540 ( .A1(n1646), .A2(n1645), .ZN(n1647) );
  ND3D1BWP12T U2541 ( .A1(n1647), .A2(write1_in[26]), .A3(write1_in[27]), .ZN(
        n1663) );
  CKND2D0BWP12T U2542 ( .A1(write2_in[24]), .A2(write2_in[26]), .ZN(n1648) );
  NR2D0BWP12T U2543 ( .A1(n1649), .A2(n1648), .ZN(n1650) );
  NR2D1BWP12T U2544 ( .A1(n1731), .A2(n2920), .ZN(n1713) );
  ND2XD0BWP12T U2545 ( .A1(n1650), .A2(n1713), .ZN(n1664) );
  INR2XD1BWP12T U2546 ( .A1(write1_in[21]), .B1(n2916), .ZN(n1654) );
  NR3D0BWP12T U2547 ( .A1(n1652), .A2(n1651), .A3(n1699), .ZN(n1653) );
  AOI31D1BWP12T U2548 ( .A1(write1_in[25]), .A2(n1654), .A3(write1_in[22]), 
        .B(n1653), .ZN(n1655) );
  INR2D4BWP12T U2549 ( .A1(n1656), .B1(n1655), .ZN(n2912) );
  CKND2D1BWP12T U2550 ( .A1(n2911), .A2(n2912), .ZN(n1657) );
  TPNR2D1BWP12T U2551 ( .A1(n1658), .A2(n1657), .ZN(n1661) );
  ND3D0BWP12T U2552 ( .A1(write1_in[28]), .A2(write1_in[29]), .A3(n2920), .ZN(
        n1660) );
  CKND2D0BWP12T U2553 ( .A1(write2_in[29]), .A2(n2916), .ZN(n2915) );
  CKND0BWP12T U2554 ( .I(n2915), .ZN(n2918) );
  CKND2D0BWP12T U2555 ( .A1(n2918), .A2(write2_in[28]), .ZN(n1659) );
  ND2D1BWP12T U2556 ( .A1(n1660), .A2(n1659), .ZN(n1662) );
  TPND2D1BWP12T U2557 ( .A1(n1661), .A2(n1662), .ZN(n1673) );
  INVD1BWP12T U2558 ( .I(n1662), .ZN(n1668) );
  AOI21D0BWP12T U2559 ( .A1(n2916), .A2(n1665), .B(n2919), .ZN(n1666) );
  OA21D1BWP12T U2560 ( .A1(write1_in[31]), .A2(n2916), .B(n1666), .Z(n1670) );
  OAI21D1BWP12T U2561 ( .A1(n1668), .A2(n1667), .B(n1670), .ZN(n1672) );
  AOI21D1BWP12T U2562 ( .A1(n1670), .A2(n2931), .B(n1669), .ZN(n1671) );
  ND3D1BWP12T U2563 ( .A1(n1673), .A2(n1672), .A3(n1671), .ZN(n2200) );
  ND3D1BWP12T U2564 ( .A1(n1674), .A2(write1_in[23]), .A3(n2920), .ZN(n1676)
         );
  IND3D0BWP12T U2565 ( .A1(n2920), .B1(write2_in[23]), .B2(write2_in[24]), 
        .ZN(n1675) );
  ND2D1BWP12T U2566 ( .A1(n1676), .A2(n1675), .ZN(n1740) );
  ND3D0BWP12T U2567 ( .A1(write1_in[27]), .A2(n2920), .A3(write1_in[26]), .ZN(
        n1677) );
  IOA21D1BWP12T U2568 ( .A1(write2_in[26]), .A2(n1713), .B(n1677), .ZN(n1678)
         );
  ND3D1BWP12T U2569 ( .A1(n2912), .A2(n1740), .A3(n1678), .ZN(n1689) );
  OA21XD0BWP12T U2570 ( .A1(write2_in[28]), .A2(n2920), .B(n2914), .Z(n1680)
         );
  OAI21D0BWP12T U2571 ( .A1(write1_in[28]), .A2(n2916), .B(n1680), .ZN(n1681)
         );
  OR2D2BWP12T U2572 ( .A1(n2927), .A2(n1681), .Z(n1688) );
  AOI21D1BWP12T U2573 ( .A1(n2920), .A2(write1_in[28]), .B(n2910), .ZN(n1741)
         );
  AOI31D1BWP12T U2574 ( .A1(n2927), .A2(n2914), .A3(n1741), .B(n1682), .ZN(
        n1687) );
  INR2XD0BWP12T U2575 ( .A1(n2920), .B1(n2919), .ZN(n1684) );
  INR2D0BWP12T U2576 ( .A1(n2914), .B1(n2915), .ZN(n1683) );
  AO21D0BWP12T U2577 ( .A1(write1_in[29]), .A2(n1684), .B(n1683), .Z(n1685) );
  ND2D1BWP12T U2578 ( .A1(n1689), .A2(n1685), .ZN(n1686) );
  OAI211D1BWP12T U2579 ( .A1(n1689), .A2(n1688), .B(n1687), .C(n1686), .ZN(
        n2198) );
  CKND2D1BWP12T U2580 ( .A1(n2900), .A2(n2914), .ZN(n1694) );
  AOI22D0BWP12T U2581 ( .A1(next_pc_in[23]), .A2(n1488), .B1(n1690), .B2(
        pc_out[23]), .ZN(n1691) );
  OA21D1BWP12T U2582 ( .A1(n1694), .A2(n1749), .B(n1691), .Z(n1698) );
  CKND1BWP12T U2583 ( .I(n2900), .ZN(n1692) );
  CKND2D1BWP12T U2584 ( .A1(n1692), .A2(n2914), .ZN(n1693) );
  CKND2D2BWP12T U2585 ( .A1(n1749), .A2(n1748), .ZN(n2905) );
  NR2D1BWP12T U2586 ( .A1(n1693), .A2(n2905), .ZN(n1696) );
  NR2D1BWP12T U2587 ( .A1(n1694), .A2(n1748), .ZN(n1695) );
  NR2D1BWP12T U2588 ( .A1(n1696), .A2(n1695), .ZN(n1697) );
  ND2D1BWP12T U2589 ( .A1(n1698), .A2(n1697), .ZN(n2192) );
  IND2XD1BWP12T U2590 ( .A1(write1_in[25]), .B1(n1699), .ZN(n1703) );
  IOA21D1BWP12T U2591 ( .A1(n1701), .A2(write2_in[22]), .B(n1700), .ZN(n1702)
         );
  TPND2D3BWP12T U2592 ( .A1(write1_in[26]), .A2(n2920), .ZN(n1705) );
  CKND2D0BWP12T U2593 ( .A1(write2_in[26]), .A2(n2916), .ZN(n1704) );
  CKND2D1BWP12T U2594 ( .A1(n1739), .A2(n2914), .ZN(n1709) );
  INVD1BWP12T U2595 ( .I(n1709), .ZN(n1706) );
  OAI21D1BWP12T U2596 ( .A1(n1735), .A2(n1720), .B(n1706), .ZN(n1712) );
  IND4D1BWP12T U2597 ( .A1(n1720), .B1(n1718), .B2(n1749), .B3(n1740), .ZN(
        n1711) );
  OA21D1BWP12T U2598 ( .A1(n1709), .A2(n1749), .B(n1708), .Z(n1710) );
  ND3D1BWP12T U2599 ( .A1(n1712), .A2(n1711), .A3(n1710), .ZN(n2195) );
  AN2XD2BWP12T U2600 ( .A1(n1749), .A2(n1740), .Z(n1726) );
  INVD1BWP12T U2601 ( .I(n1726), .ZN(n1714) );
  TPAOI21D2BWP12T U2602 ( .A1(write1_in[27]), .A2(n2920), .B(n1713), .ZN(n1723) );
  TPNR2D1BWP12T U2603 ( .A1(n1723), .A2(n2919), .ZN(n1719) );
  CKND2D1BWP12T U2604 ( .A1(n1714), .A2(n1719), .ZN(n1730) );
  INVD1BWP12T U2605 ( .I(n1723), .ZN(n1738) );
  CKND0BWP12T U2606 ( .I(pc_out[27]), .ZN(n1716) );
  ND2XD0BWP12T U2607 ( .A1(next_pc_in[27]), .A2(n1488), .ZN(n1715) );
  OAI21D0BWP12T U2608 ( .A1(n2924), .A2(n1716), .B(n1715), .ZN(n1717) );
  AO21D1BWP12T U2609 ( .A1(n1718), .A2(n1738), .B(n1717), .Z(n1722) );
  ND3D1BWP12T U2610 ( .A1(n1739), .A2(n1723), .A3(n2914), .ZN(n1724) );
  INR2D1BWP12T U2611 ( .A1(n1725), .B1(n1724), .ZN(n1727) );
  ND2D1BWP12T U2612 ( .A1(n1727), .A2(n1726), .ZN(n1728) );
  ND3D1BWP12T U2613 ( .A1(n1730), .A2(n1729), .A3(n1728), .ZN(n2196) );
  NR2D1BWP12T U2614 ( .A1(write1_in[27]), .A2(n2916), .ZN(n1734) );
  AOI21D0BWP12T U2615 ( .A1(n2916), .A2(n1731), .B(n2919), .ZN(n1732) );
  CKND2D2BWP12T U2616 ( .A1(n1739), .A2(n1732), .ZN(n1733) );
  TPNR3D2BWP12T U2617 ( .A1(n1735), .A2(n1734), .A3(n1733), .ZN(n1736) );
  ND3D1BWP12T U2618 ( .A1(n1736), .A2(n1741), .A3(n2912), .ZN(n1747) );
  TPAOI21D0BWP12T U2619 ( .A1(next_pc_in[28]), .A2(n1488), .B(n1737), .ZN(
        n1746) );
  CKND2D1BWP12T U2620 ( .A1(n1738), .A2(n2912), .ZN(n1744) );
  CKND2D1BWP12T U2621 ( .A1(n1740), .A2(n1739), .ZN(n1743) );
  NR2D1BWP12T U2622 ( .A1(n1741), .A2(n2919), .ZN(n1742) );
  OAI21D1BWP12T U2623 ( .A1(n1744), .A2(n1743), .B(n1742), .ZN(n1745) );
  ND3D1BWP12T U2624 ( .A1(n1747), .A2(n1746), .A3(n1745), .ZN(n2197) );
  XNR2XD1BWP12T U2625 ( .A1(n1749), .A2(n1748), .ZN(n1753) );
  TPNR2D0BWP12T U2626 ( .A1(n2924), .A2(n1750), .ZN(n1751) );
  AOI21D1BWP12T U2627 ( .A1(next_pc_in[22]), .A2(n1488), .B(n1751), .ZN(n1752)
         );
  OAI21D1BWP12T U2628 ( .A1(n1753), .A2(n2919), .B(n1752), .ZN(n2191) );
  AOI22D1BWP12T U2629 ( .A1(n2795), .A2(r0[31]), .B1(n2791), .B2(r4[31]), .ZN(
        n1755) );
  AOI22D1BWP12T U2630 ( .A1(tmp1[31]), .A2(n2820), .B1(n2819), .B2(r9[31]), 
        .ZN(n1754) );
  OA211D1BWP12T U2631 ( .A1(n1756), .A2(n2789), .B(n1755), .C(n1754), .Z(n1764) );
  AOI22D1BWP12T U2632 ( .A1(n2808), .A2(r11[31]), .B1(n2807), .B2(n[2937]), 
        .ZN(n1760) );
  AOI22D1BWP12T U2633 ( .A1(r3[31]), .A2(n2810), .B1(n2809), .B2(r5[31]), .ZN(
        n1759) );
  AOI22D1BWP12T U2634 ( .A1(n2812), .A2(r7[31]), .B1(n2811), .B2(pc_out[31]), 
        .ZN(n1758) );
  AOI22D1BWP12T U2635 ( .A1(n2814), .A2(r1[31]), .B1(n2813), .B2(r12[31]), 
        .ZN(n1757) );
  AN4XD1BWP12T U2636 ( .A1(n1760), .A2(n1759), .A3(n1758), .A4(n1757), .Z(
        n1763) );
  AOI22D1BWP12T U2637 ( .A1(n2892), .A2(r8[31]), .B1(n2891), .B2(lr[31]), .ZN(
        n1762) );
  AOI22D1BWP12T U2638 ( .A1(r6[31]), .A2(n2894), .B1(n2893), .B2(r10[31]), 
        .ZN(n1761) );
  ND4D1BWP12T U2639 ( .A1(n1764), .A2(n1763), .A3(n1762), .A4(n1761), .ZN(
        regA_out[31]) );
  AOI22D1BWP12T U2640 ( .A1(r1[30]), .A2(n118), .B1(n2761), .B2(r12[30]), .ZN(
        n1768) );
  AOI22D1BWP12T U2641 ( .A1(r3[30]), .A2(n2763), .B1(n2762), .B2(lr[30]), .ZN(
        n1767) );
  AOI22D1BWP12T U2642 ( .A1(r8[30]), .A2(n2765), .B1(n2764), .B2(n[2938]), 
        .ZN(n1766) );
  AOI22D1BWP12T U2643 ( .A1(pc_out[30]), .A2(n2767), .B1(n2766), .B2(r6[30]), 
        .ZN(n1765) );
  AN4XD1BWP12T U2644 ( .A1(n1768), .A2(n1767), .A3(n1766), .A4(n1765), .Z(
        n1775) );
  AOI22D1BWP12T U2645 ( .A1(tmp1[30]), .A2(n2746), .B1(n2135), .B2(
        immediate2_in[30]), .ZN(n1771) );
  AOI22D1BWP12T U2646 ( .A1(r9[30]), .A2(n105), .B1(n2753), .B2(r4[30]), .ZN(
        n1770) );
  AOI22D1BWP12T U2647 ( .A1(r11[30]), .A2(n2755), .B1(n2650), .B2(r0[30]), 
        .ZN(n1769) );
  AN3XD1BWP12T U2648 ( .A1(n1771), .A2(n1770), .A3(n1769), .Z(n1774) );
  AOI22D1BWP12T U2649 ( .A1(r5[30]), .A2(n2748), .B1(n2747), .B2(r10[30]), 
        .ZN(n1773) );
  AOI22D1BWP12T U2650 ( .A1(r7[30]), .A2(n2750), .B1(n2749), .B2(r2[30]), .ZN(
        n1772) );
  ND4D1BWP12T U2651 ( .A1(n1775), .A2(n1774), .A3(n1773), .A4(n1772), .ZN(
        regB_out[30]) );
  INVD1BWP12T U2652 ( .I(r2[29]), .ZN(n1778) );
  AOI22D1BWP12T U2653 ( .A1(r4[29]), .A2(n2791), .B1(n2795), .B2(r0[29]), .ZN(
        n1777) );
  AOI22D1BWP12T U2654 ( .A1(tmp1[29]), .A2(n2820), .B1(n2819), .B2(r9[29]), 
        .ZN(n1776) );
  OA211D1BWP12T U2655 ( .A1(n1778), .A2(n2789), .B(n1777), .C(n1776), .Z(n1787) );
  AOI22D1BWP12T U2656 ( .A1(n2808), .A2(r11[29]), .B1(n2807), .B2(n[2939]), 
        .ZN(n1782) );
  AOI22D1BWP12T U2657 ( .A1(r3[29]), .A2(n2810), .B1(n2809), .B2(r5[29]), .ZN(
        n1781) );
  AOI22D1BWP12T U2658 ( .A1(n2812), .A2(r7[29]), .B1(n2776), .B2(pc_out[29]), 
        .ZN(n1780) );
  AOI22D1BWP12T U2659 ( .A1(n2814), .A2(r1[29]), .B1(n2708), .B2(r12[29]), 
        .ZN(n1779) );
  AN4XD1BWP12T U2660 ( .A1(n1782), .A2(n1781), .A3(n1780), .A4(n1779), .Z(
        n1786) );
  AOI22D1BWP12T U2661 ( .A1(n2892), .A2(r8[29]), .B1(n2891), .B2(lr[29]), .ZN(
        n1784) );
  AOI22D1BWP12T U2662 ( .A1(r6[29]), .A2(n2894), .B1(n2893), .B2(r10[29]), 
        .ZN(n1783) );
  AN2XD1BWP12T U2663 ( .A1(n1784), .A2(n1783), .Z(n1785) );
  ND3D1BWP12T U2664 ( .A1(n1787), .A2(n1786), .A3(n1785), .ZN(regA_out[29]) );
  INVD1BWP12T U2665 ( .I(r2[28]), .ZN(n1790) );
  AOI22D1BWP12T U2666 ( .A1(n2791), .A2(r4[28]), .B1(n2795), .B2(r0[28]), .ZN(
        n1789) );
  AOI22D1BWP12T U2667 ( .A1(tmp1[28]), .A2(n2820), .B1(n2819), .B2(r9[28]), 
        .ZN(n1788) );
  OA211D1BWP12T U2668 ( .A1(n1790), .A2(n2789), .B(n1789), .C(n1788), .Z(n1799) );
  AOI22D1BWP12T U2669 ( .A1(n2808), .A2(r11[28]), .B1(n2807), .B2(n[2940]), 
        .ZN(n1795) );
  AOI22D1BWP12T U2670 ( .A1(r7[28]), .A2(n2812), .B1(n2811), .B2(pc_out[28]), 
        .ZN(n1794) );
  AOI22D1BWP12T U2671 ( .A1(r3[28]), .A2(n2810), .B1(n2809), .B2(r5[28]), .ZN(
        n1793) );
  INVD1BWP12T U2672 ( .I(r12[28]), .ZN(n1791) );
  AN4XD1BWP12T U2673 ( .A1(n1795), .A2(n1794), .A3(n1793), .A4(n1792), .Z(
        n1798) );
  AOI22D1BWP12T U2674 ( .A1(n2892), .A2(r8[28]), .B1(n2891), .B2(lr[28]), .ZN(
        n1797) );
  AOI22D1BWP12T U2675 ( .A1(n2894), .A2(r6[28]), .B1(n2893), .B2(r10[28]), 
        .ZN(n1796) );
  ND4D1BWP12T U2676 ( .A1(n1799), .A2(n1798), .A3(n1797), .A4(n1796), .ZN(
        regA_out[28]) );
  AOI22D1BWP12T U2677 ( .A1(r1[27]), .A2(n118), .B1(n2761), .B2(r12[27]), .ZN(
        n1803) );
  AOI22D1BWP12T U2678 ( .A1(r3[27]), .A2(n2763), .B1(n2762), .B2(lr[27]), .ZN(
        n1802) );
  AOI22D1BWP12T U2679 ( .A1(r8[27]), .A2(n2765), .B1(n2764), .B2(n[2941]), 
        .ZN(n1801) );
  AOI22D1BWP12T U2680 ( .A1(pc_out[27]), .A2(n2767), .B1(n2766), .B2(r6[27]), 
        .ZN(n1800) );
  AN4XD1BWP12T U2681 ( .A1(n1803), .A2(n1802), .A3(n1801), .A4(n1800), .Z(
        n1810) );
  AOI22D1BWP12T U2682 ( .A1(tmp1[27]), .A2(n2746), .B1(n2745), .B2(
        immediate2_in[27]), .ZN(n1806) );
  AOI22D1BWP12T U2683 ( .A1(r9[27]), .A2(n105), .B1(n2753), .B2(r4[27]), .ZN(
        n1805) );
  AOI22D1BWP12T U2684 ( .A1(r11[27]), .A2(n2755), .B1(n2650), .B2(r0[27]), 
        .ZN(n1804) );
  AN3XD1BWP12T U2685 ( .A1(n1806), .A2(n1805), .A3(n1804), .Z(n1809) );
  AOI22D1BWP12T U2686 ( .A1(r5[27]), .A2(n2748), .B1(n2747), .B2(r10[27]), 
        .ZN(n1808) );
  AOI22D1BWP12T U2687 ( .A1(r7[27]), .A2(n2750), .B1(n2749), .B2(r2[27]), .ZN(
        n1807) );
  ND4D1BWP12T U2688 ( .A1(n1810), .A2(n1809), .A3(n1808), .A4(n1807), .ZN(
        regB_out[27]) );
  AOI22D1BWP12T U2689 ( .A1(r1[26]), .A2(n118), .B1(n2761), .B2(r12[26]), .ZN(
        n1814) );
  AOI22D1BWP12T U2690 ( .A1(r3[26]), .A2(n2763), .B1(n2762), .B2(lr[26]), .ZN(
        n1813) );
  AOI22D1BWP12T U2691 ( .A1(r8[26]), .A2(n2765), .B1(n2764), .B2(n[2942]), 
        .ZN(n1812) );
  AOI22D1BWP12T U2692 ( .A1(pc_out[26]), .A2(n2767), .B1(n2766), .B2(r6[26]), 
        .ZN(n1811) );
  AN4XD1BWP12T U2693 ( .A1(n1814), .A2(n1813), .A3(n1812), .A4(n1811), .Z(
        n1821) );
  AOI22D1BWP12T U2694 ( .A1(tmp1[26]), .A2(n2746), .B1(n2730), .B2(
        immediate2_in[26]), .ZN(n1817) );
  AOI22D1BWP12T U2695 ( .A1(r9[26]), .A2(n105), .B1(n2753), .B2(r4[26]), .ZN(
        n1816) );
  AOI22D1BWP12T U2696 ( .A1(r11[26]), .A2(n2755), .B1(n2754), .B2(r0[26]), 
        .ZN(n1815) );
  AN3XD1BWP12T U2697 ( .A1(n1817), .A2(n1816), .A3(n1815), .Z(n1820) );
  AOI22D1BWP12T U2698 ( .A1(r5[26]), .A2(n2748), .B1(n2747), .B2(r10[26]), 
        .ZN(n1819) );
  AOI22D1BWP12T U2699 ( .A1(r7[26]), .A2(n2750), .B1(n2749), .B2(r2[26]), .ZN(
        n1818) );
  ND4D1BWP12T U2700 ( .A1(n1821), .A2(n1820), .A3(n1819), .A4(n1818), .ZN(
        regB_out[26]) );
  AOI22D1BWP12T U2701 ( .A1(n2808), .A2(r11[0]), .B1(n2807), .B2(n[2968]), 
        .ZN(n1825) );
  AOI22D1BWP12T U2702 ( .A1(r3[0]), .A2(n2810), .B1(n2809), .B2(r5[0]), .ZN(
        n1824) );
  AOI22D1BWP12T U2703 ( .A1(n2812), .A2(r7[0]), .B1(n2776), .B2(pc_out[0]), 
        .ZN(n1823) );
  AOI22D1BWP12T U2704 ( .A1(n2814), .A2(r1[0]), .B1(n2708), .B2(r12[0]), .ZN(
        n1822) );
  AN4XD1BWP12T U2705 ( .A1(n1825), .A2(n1824), .A3(n1823), .A4(n1822), .Z(
        n1838) );
  AOI22D1BWP12T U2706 ( .A1(tmp1[0]), .A2(n2820), .B1(n2819), .B2(r9[0]), .ZN(
        n1826) );
  IOA21D1BWP12T U2707 ( .A1(r2[0]), .A2(n2890), .B(n1826), .ZN(n1836) );
  INVD1BWP12T U2708 ( .I(r8[0]), .ZN(n1827) );
  OAI22D1BWP12T U2709 ( .A1(n2825), .A2(n1828), .B1(n1827), .B2(n2822), .ZN(
        n1835) );
  INVD1BWP12T U2710 ( .I(r6[0]), .ZN(n1829) );
  OAI22D1BWP12T U2711 ( .A1(n2829), .A2(n1830), .B1(n1829), .B2(n2826), .ZN(
        n1834) );
  INVD1BWP12T U2712 ( .I(r4[0]), .ZN(n1832) );
  INVD1BWP12T U2713 ( .I(r0[0]), .ZN(n1831) );
  OAI22D1BWP12T U2714 ( .A1(n2887), .A2(n1832), .B1(n1831), .B2(n2884), .ZN(
        n1833) );
  NR4D0BWP12T U2715 ( .A1(n1836), .A2(n1835), .A3(n1834), .A4(n1833), .ZN(
        n1837) );
  ND2D1BWP12T U2716 ( .A1(n1838), .A2(n1837), .ZN(regA_out[0]) );
  OAI22D1BWP12T U2717 ( .A1(n2030), .A2(n2664), .B1(n2663), .B2(n2048), .ZN(
        n1845) );
  INVD1BWP12T U2718 ( .I(tmp1[21]), .ZN(n2041) );
  MOAI22D0BWP12T U2719 ( .A1(n2041), .A2(n2666), .B1(n2135), .B2(
        immediate2_in[21]), .ZN(n1844) );
  AOI22D1BWP12T U2720 ( .A1(r9[21]), .A2(n105), .B1(n2753), .B2(r4[21]), .ZN(
        n1840) );
  AOI22D1BWP12T U2721 ( .A1(r11[21]), .A2(n2755), .B1(n2733), .B2(r0[21]), 
        .ZN(n1839) );
  ND2D1BWP12T U2722 ( .A1(n1840), .A2(n1839), .ZN(n1843) );
  OAI22D1BWP12T U2723 ( .A1(n2673), .A2(n2033), .B1(n2671), .B2(n1841), .ZN(
        n1842) );
  NR4D0BWP12T U2724 ( .A1(n1845), .A2(n1844), .A3(n1843), .A4(n1842), .ZN(
        n1851) );
  OAI22D1BWP12T U2725 ( .A1(n2035), .A2(n2680), .B1(n2679), .B2(n2036), .ZN(
        n1849) );
  OAI22D1BWP12T U2726 ( .A1(n2029), .A2(n2684), .B1(n2683), .B2(n2050), .ZN(
        n1848) );
  OAI22D1BWP12T U2727 ( .A1(n2689), .A2(n2049), .B1(n2687), .B2(n2032), .ZN(
        n1847) );
  INVD1BWP12T U2728 ( .I(pc_out[21]), .ZN(n2034) );
  OAI22D1BWP12T U2729 ( .A1(n2693), .A2(n2034), .B1(n2691), .B2(n2047), .ZN(
        n1846) );
  NR4D0BWP12T U2730 ( .A1(n1849), .A2(n1848), .A3(n1847), .A4(n1846), .ZN(
        n1850) );
  ND2D1BWP12T U2731 ( .A1(n1851), .A2(n1850), .ZN(regB_out[21]) );
  INVD1BWP12T U2732 ( .I(n[2964]), .ZN(n2019) );
  NR2XD0BWP12T U2733 ( .A1(n1854), .A2(readA_sel[1]), .ZN(n1857) );
  INVD1BWP12T U2734 ( .I(tmp1[4]), .ZN(n2006) );
  NR2D1BWP12T U2735 ( .A1(n2880), .A2(n2006), .ZN(n1858) );
  INR3D0BWP12T U2736 ( .A1(n1861), .B1(n1860), .B2(n1859), .ZN(n1872) );
  NR2D1BWP12T U2737 ( .A1(n2860), .A2(n2018), .ZN(n1862) );
  RCIAO21D0BWP12T U2738 ( .A1(n2863), .A2(n2005), .B(n1862), .ZN(n1870) );
  ND2D1BWP12T U2739 ( .A1(n2813), .A2(r12[4]), .ZN(n1863) );
  IOA21D1BWP12T U2740 ( .A1(n2814), .A2(r1[4]), .B(n1863), .ZN(n1869) );
  NR2D1BWP12T U2741 ( .A1(n2822), .A2(n2020), .ZN(n1864) );
  AOI21D0BWP12T U2742 ( .A1(n2891), .A2(lr[4]), .B(n1864), .ZN(n1867) );
  NR2D1BWP12T U2743 ( .A1(n2826), .A2(n2021), .ZN(n1865) );
  TPAOI21D0BWP12T U2744 ( .A1(n2893), .A2(r10[4]), .B(n1865), .ZN(n1866) );
  CKND2D1BWP12T U2745 ( .A1(n1867), .A2(n1866), .ZN(n1868) );
  INR3XD0BWP12T U2746 ( .A1(n1870), .B1(n1869), .B2(n1868), .ZN(n1871) );
  ND2D1BWP12T U2747 ( .A1(n1872), .A2(n1871), .ZN(regA_out[4]) );
  NR2D1BWP12T U2748 ( .A1(n2880), .A2(n1875), .ZN(n1876) );
  INR3D0BWP12T U2749 ( .A1(n1880), .B1(n1879), .B2(n1878), .ZN(n1892) );
  CKND2D1BWP12T U2750 ( .A1(n2807), .A2(n[2966]), .ZN(n1882) );
  OAI21D1BWP12T U2751 ( .A1(n2864), .A2(n1883), .B(n1882), .ZN(n1889) );
  ND2D1BWP12T U2752 ( .A1(n1887), .A2(n1886), .ZN(n1888) );
  INR3D0BWP12T U2753 ( .A1(n1890), .B1(n1889), .B2(n1888), .ZN(n1891) );
  ND2D1BWP12T U2754 ( .A1(n1892), .A2(n1891), .ZN(regA_out[2]) );
  INVD1BWP12T U2755 ( .I(r2[26]), .ZN(n1895) );
  AOI22D1BWP12T U2756 ( .A1(r0[26]), .A2(n2795), .B1(n2791), .B2(r4[26]), .ZN(
        n1894) );
  AOI22D1BWP12T U2757 ( .A1(tmp1[26]), .A2(n2820), .B1(n2819), .B2(r9[26]), 
        .ZN(n1893) );
  OA211D1BWP12T U2758 ( .A1(n1895), .A2(n2789), .B(n1894), .C(n1893), .Z(n1903) );
  AOI22D1BWP12T U2759 ( .A1(n2808), .A2(r11[26]), .B1(n2807), .B2(n[2942]), 
        .ZN(n1899) );
  AOI22D1BWP12T U2760 ( .A1(r3[26]), .A2(n2810), .B1(n2809), .B2(r5[26]), .ZN(
        n1898) );
  AOI22D1BWP12T U2761 ( .A1(n2812), .A2(r7[26]), .B1(n2811), .B2(pc_out[26]), 
        .ZN(n1897) );
  AOI22D1BWP12T U2762 ( .A1(n2814), .A2(r1[26]), .B1(n2813), .B2(r12[26]), 
        .ZN(n1896) );
  AN4XD1BWP12T U2763 ( .A1(n1899), .A2(n1898), .A3(n1897), .A4(n1896), .Z(
        n1902) );
  AOI22D1BWP12T U2764 ( .A1(n2892), .A2(r8[26]), .B1(n2891), .B2(lr[26]), .ZN(
        n1901) );
  AOI22D1BWP12T U2765 ( .A1(r6[26]), .A2(n2894), .B1(n2893), .B2(r10[26]), 
        .ZN(n1900) );
  ND4D1BWP12T U2766 ( .A1(n1903), .A2(n1902), .A3(n1901), .A4(n1900), .ZN(
        regA_out[26]) );
  AOI22D1BWP12T U2767 ( .A1(tmp1[13]), .A2(n2746), .B1(n2730), .B2(
        immediate2_in[13]), .ZN(n1910) );
  AOI22D1BWP12T U2768 ( .A1(r5[13]), .A2(n2748), .B1(n2747), .B2(r10[13]), 
        .ZN(n1905) );
  AOI22D1BWP12T U2769 ( .A1(r7[13]), .A2(n2750), .B1(n2749), .B2(r2[13]), .ZN(
        n1904) );
  ND2D1BWP12T U2770 ( .A1(n1905), .A2(n1904), .ZN(n1909) );
  AOI22D1BWP12T U2771 ( .A1(r9[13]), .A2(n105), .B1(n2753), .B2(r4[13]), .ZN(
        n1907) );
  AOI22D1BWP12T U2772 ( .A1(r11[13]), .A2(n2755), .B1(n2733), .B2(r0[13]), 
        .ZN(n1906) );
  ND2D1BWP12T U2773 ( .A1(n1907), .A2(n1906), .ZN(n1908) );
  INR3XD0BWP12T U2774 ( .A1(n1910), .B1(n1909), .B2(n1908), .ZN(n1916) );
  AOI22D1BWP12T U2775 ( .A1(r1[13]), .A2(n118), .B1(n2761), .B2(r12[13]), .ZN(
        n1914) );
  AOI22D1BWP12T U2776 ( .A1(r3[13]), .A2(n2763), .B1(n2762), .B2(lr[13]), .ZN(
        n1913) );
  AOI22D1BWP12T U2777 ( .A1(r8[13]), .A2(n2765), .B1(n2764), .B2(n[2955]), 
        .ZN(n1912) );
  AOI22D1BWP12T U2778 ( .A1(pc_out[13]), .A2(n2767), .B1(n2766), .B2(r6[13]), 
        .ZN(n1911) );
  AN4XD1BWP12T U2779 ( .A1(n1914), .A2(n1913), .A3(n1912), .A4(n1911), .Z(
        n1915) );
  ND2D1BWP12T U2780 ( .A1(n1916), .A2(n1915), .ZN(regB_out[13]) );
  OAI22D1BWP12T U2781 ( .A1(n1918), .A2(n2664), .B1(n2663), .B2(n1917), .ZN(
        n1927) );
  MOAI22D0BWP12T U2782 ( .A1(n1919), .A2(n2666), .B1(n2135), .B2(
        immediate2_in[11]), .ZN(n1926) );
  AOI22D1BWP12T U2783 ( .A1(r9[11]), .A2(n105), .B1(n2753), .B2(r4[11]), .ZN(
        n1921) );
  AOI22D1BWP12T U2784 ( .A1(r11[11]), .A2(n2755), .B1(n2733), .B2(r0[11]), 
        .ZN(n1920) );
  ND2D1BWP12T U2785 ( .A1(n1921), .A2(n1920), .ZN(n1925) );
  OAI22D1BWP12T U2786 ( .A1(n2673), .A2(n1923), .B1(n2671), .B2(n1922), .ZN(
        n1924) );
  NR4D0BWP12T U2787 ( .A1(n1927), .A2(n1926), .A3(n1925), .A4(n1924), .ZN(
        n1941) );
  OAI22D1BWP12T U2788 ( .A1(n1931), .A2(n2684), .B1(n2683), .B2(n1930), .ZN(
        n1938) );
  OAI22D1BWP12T U2789 ( .A1(n2689), .A2(n1933), .B1(n2687), .B2(n1932), .ZN(
        n1937) );
  INVD1BWP12T U2790 ( .I(pc_out[11]), .ZN(n1935) );
  OAI22D1BWP12T U2791 ( .A1(n2693), .A2(n1935), .B1(n2691), .B2(n1934), .ZN(
        n1936) );
  NR4D0BWP12T U2792 ( .A1(n1939), .A2(n1938), .A3(n1937), .A4(n1936), .ZN(
        n1940) );
  ND2D1BWP12T U2793 ( .A1(n1941), .A2(n1940), .ZN(regB_out[11]) );
  NR2D1BWP12T U2794 ( .A1(n1943), .A2(n1942), .ZN(n1944) );
  RCAOI21D0BWP12T U2795 ( .A1(n2891), .A2(lr[12]), .B(n1944), .ZN(n1956) );
  CKND2D1BWP12T U2796 ( .A1(n2893), .A2(r10[12]), .ZN(n1945) );
  TPOAI21D0BWP12T U2797 ( .A1(n2826), .A2(n1946), .B(n1945), .ZN(n1955) );
  NR2D1BWP12T U2798 ( .A1(n2880), .A2(n1947), .ZN(n1948) );
  AOI21D1BWP12T U2799 ( .A1(n2819), .A2(r9[12]), .B(n1948), .ZN(n1953) );
  TPND2D0BWP12T U2800 ( .A1(n2890), .A2(r2[12]), .ZN(n1952) );
  NR2D1BWP12T U2801 ( .A1(n2884), .A2(n1949), .ZN(n1950) );
  TPAOI21D0BWP12T U2802 ( .A1(n2791), .A2(r4[12]), .B(n1950), .ZN(n1951) );
  ND3D1BWP12T U2803 ( .A1(n1953), .A2(n1952), .A3(n1951), .ZN(n1954) );
  INR3D0BWP12T U2804 ( .A1(n1956), .B1(n1955), .B2(n1954), .ZN(n1971) );
  NR2D1BWP12T U2805 ( .A1(n2868), .A2(n1957), .ZN(n1958) );
  AOI21D1BWP12T U2806 ( .A1(n2776), .A2(pc_out[12]), .B(n1958), .ZN(n1969) );
  CKND2D1BWP12T U2807 ( .A1(n2807), .A2(n[2956]), .ZN(n1959) );
  OAI21D1BWP12T U2808 ( .A1(n2864), .A2(n1960), .B(n1959), .ZN(n1968) );
  NR2D1BWP12T U2809 ( .A1(n2860), .A2(n1961), .ZN(n1962) );
  AOI21D1BWP12T U2810 ( .A1(n2809), .A2(r5[12]), .B(n1962), .ZN(n1966) );
  NR2D1BWP12T U2811 ( .A1(n2872), .A2(n1963), .ZN(n1964) );
  AOI21D1BWP12T U2812 ( .A1(n2813), .A2(r12[12]), .B(n1964), .ZN(n1965) );
  ND2D1BWP12T U2813 ( .A1(n1966), .A2(n1965), .ZN(n1967) );
  INR3D0BWP12T U2814 ( .A1(n1969), .B1(n1968), .B2(n1967), .ZN(n1970) );
  ND2D1BWP12T U2815 ( .A1(n1971), .A2(n1970), .ZN(regA_out[12]) );
  OAI22D1BWP12T U2816 ( .A1(n2863), .A2(n2057), .B1(n2070), .B2(n2860), .ZN(
        n1976) );
  OAI22D0BWP12T U2817 ( .A1(n2867), .A2(n2071), .B1(n1972), .B2(n2864), .ZN(
        n1975) );
  INVD1BWP12T U2818 ( .I(pc_out[20]), .ZN(n2074) );
  OAI22D1BWP12T U2819 ( .A1(n2871), .A2(n2074), .B1(n2062), .B2(n2868), .ZN(
        n1974) );
  OAI22D1BWP12T U2820 ( .A1(n2851), .A2(n2067), .B1(n2068), .B2(n2872), .ZN(
        n1973) );
  NR4D0BWP12T U2821 ( .A1(n1976), .A2(n1975), .A3(n1974), .A4(n1973), .ZN(
        n1986) );
  INVD1BWP12T U2822 ( .I(tmp1[20]), .ZN(n2058) );
  OAI22D1BWP12T U2823 ( .A1(n2883), .A2(n1977), .B1(n2058), .B2(n2880), .ZN(
        n1981) );
  OAI22D1BWP12T U2824 ( .A1(n2887), .A2(n1979), .B1(n1978), .B2(n2884), .ZN(
        n1980) );
  AOI211D1BWP12T U2825 ( .A1(r2[20]), .A2(n2890), .B(n1981), .C(n1980), .ZN(
        n1985) );
  OAI22D1BWP12T U2826 ( .A1(n2829), .A2(n2056), .B1(n2073), .B2(n2826), .ZN(
        n1983) );
  OAI22D1BWP12T U2827 ( .A1(n2825), .A2(n2069), .B1(n2072), .B2(n2822), .ZN(
        n1982) );
  NR2D1BWP12T U2828 ( .A1(n1983), .A2(n1982), .ZN(n1984) );
  ND3D1BWP12T U2829 ( .A1(n1986), .A2(n1985), .A3(n1984), .ZN(regA_out[20]) );
  AOI22D1BWP12T U2830 ( .A1(n2808), .A2(r11[18]), .B1(n2807), .B2(n[2950]), 
        .ZN(n1990) );
  AOI22D1BWP12T U2831 ( .A1(r3[18]), .A2(n2810), .B1(n2809), .B2(r5[18]), .ZN(
        n1989) );
  AOI22D1BWP12T U2832 ( .A1(n2812), .A2(r7[18]), .B1(n2811), .B2(pc_out[18]), 
        .ZN(n1988) );
  AOI22D1BWP12T U2833 ( .A1(n2814), .A2(r1[18]), .B1(n2708), .B2(r12[18]), 
        .ZN(n1987) );
  AN4XD1BWP12T U2834 ( .A1(n1990), .A2(n1989), .A3(n1988), .A4(n1987), .Z(
        n2003) );
  AOI22D1BWP12T U2835 ( .A1(tmp1[18]), .A2(n2820), .B1(n2819), .B2(r9[18]), 
        .ZN(n1991) );
  IOA21D1BWP12T U2836 ( .A1(r2[18]), .A2(n2890), .B(n1991), .ZN(n2001) );
  INVD1BWP12T U2837 ( .I(lr[18]), .ZN(n1993) );
  OAI22D1BWP12T U2838 ( .A1(n2825), .A2(n1993), .B1(n1992), .B2(n2822), .ZN(
        n2000) );
  INVD1BWP12T U2839 ( .I(r10[18]), .ZN(n1995) );
  INVD1BWP12T U2840 ( .I(r6[18]), .ZN(n1994) );
  OAI22D1BWP12T U2841 ( .A1(n2829), .A2(n1995), .B1(n1994), .B2(n2826), .ZN(
        n1999) );
  INVD1BWP12T U2842 ( .I(r4[18]), .ZN(n1997) );
  INVD1BWP12T U2843 ( .I(r0[18]), .ZN(n1996) );
  OAI22D1BWP12T U2844 ( .A1(n2887), .A2(n1997), .B1(n1996), .B2(n2884), .ZN(
        n1998) );
  NR4D0BWP12T U2845 ( .A1(n2001), .A2(n2000), .A3(n1999), .A4(n1998), .ZN(
        n2002) );
  OAI22D1BWP12T U2846 ( .A1(n2005), .A2(n2664), .B1(n2663), .B2(n2004), .ZN(
        n2014) );
  MOAI22D0BWP12T U2847 ( .A1(n2006), .A2(n2666), .B1(n2135), .B2(
        immediate2_in[4]), .ZN(n2013) );
  AOI22D1BWP12T U2848 ( .A1(r9[4]), .A2(n105), .B1(n2753), .B2(r4[4]), .ZN(
        n2008) );
  AOI22D1BWP12T U2849 ( .A1(r11[4]), .A2(n2755), .B1(n2733), .B2(r0[4]), .ZN(
        n2007) );
  ND2D1BWP12T U2850 ( .A1(n2008), .A2(n2007), .ZN(n2012) );
  OAI22D1BWP12T U2851 ( .A1(n2673), .A2(n2010), .B1(n2671), .B2(n2009), .ZN(
        n2011) );
  NR4D0BWP12T U2852 ( .A1(n2014), .A2(n2013), .A3(n2012), .A4(n2011), .ZN(
        n2028) );
  OAI22D1BWP12T U2853 ( .A1(n2016), .A2(n2680), .B1(n2679), .B2(n2015), .ZN(
        n2026) );
  OAI22D1BWP12T U2854 ( .A1(n2018), .A2(n2684), .B1(n2683), .B2(n2017), .ZN(
        n2025) );
  OAI22D1BWP12T U2855 ( .A1(n2689), .A2(n2020), .B1(n2687), .B2(n2019), .ZN(
        n2024) );
  OAI22D1BWP12T U2856 ( .A1(n2693), .A2(n2022), .B1(n2691), .B2(n2021), .ZN(
        n2023) );
  NR4D0BWP12T U2857 ( .A1(n2026), .A2(n2025), .A3(n2024), .A4(n2023), .ZN(
        n2027) );
  ND2D1BWP12T U2858 ( .A1(n2028), .A2(n2027), .ZN(regB_out[4]) );
  OAI22D1BWP12T U2859 ( .A1(n2863), .A2(n2030), .B1(n2029), .B2(n2860), .ZN(
        n2040) );
  OAI22D0BWP12T U2860 ( .A1(n2867), .A2(n2032), .B1(n2031), .B2(n2864), .ZN(
        n2039) );
  OAI22D1BWP12T U2861 ( .A1(n2871), .A2(n2034), .B1(n2033), .B2(n2868), .ZN(
        n2038) );
  OAI22D1BWP12T U2862 ( .A1(n2851), .A2(n2036), .B1(n2035), .B2(n2872), .ZN(
        n2037) );
  NR4D0BWP12T U2863 ( .A1(n2040), .A2(n2039), .A3(n2038), .A4(n2037), .ZN(
        n2055) );
  OAI22D1BWP12T U2864 ( .A1(n2883), .A2(n2042), .B1(n2041), .B2(n2880), .ZN(
        n2046) );
  OAI22D1BWP12T U2865 ( .A1(n2887), .A2(n2044), .B1(n2043), .B2(n2884), .ZN(
        n2045) );
  AOI211D1BWP12T U2866 ( .A1(r2[21]), .A2(n2890), .B(n2046), .C(n2045), .ZN(
        n2054) );
  OAI22D1BWP12T U2867 ( .A1(n2829), .A2(n2048), .B1(n2047), .B2(n2826), .ZN(
        n2052) );
  OAI22D1BWP12T U2868 ( .A1(n2825), .A2(n2050), .B1(n2049), .B2(n2822), .ZN(
        n2051) );
  NR2D1BWP12T U2869 ( .A1(n2052), .A2(n2051), .ZN(n2053) );
  ND3D1BWP12T U2870 ( .A1(n2055), .A2(n2054), .A3(n2053), .ZN(regA_out[21]) );
  OAI22D1BWP12T U2871 ( .A1(n2057), .A2(n2664), .B1(n2663), .B2(n2056), .ZN(
        n2066) );
  MOAI22D0BWP12T U2872 ( .A1(n2058), .A2(n2666), .B1(n2745), .B2(
        immediate2_in[20]), .ZN(n2065) );
  AOI22D1BWP12T U2873 ( .A1(r9[20]), .A2(n105), .B1(n2753), .B2(r4[20]), .ZN(
        n2060) );
  AOI22D1BWP12T U2874 ( .A1(r11[20]), .A2(n2755), .B1(n2650), .B2(r0[20]), 
        .ZN(n2059) );
  ND2D1BWP12T U2875 ( .A1(n2060), .A2(n2059), .ZN(n2064) );
  OAI22D1BWP12T U2876 ( .A1(n2673), .A2(n2062), .B1(n2671), .B2(n2061), .ZN(
        n2063) );
  NR4D0BWP12T U2877 ( .A1(n2066), .A2(n2065), .A3(n2064), .A4(n2063), .ZN(
        n2080) );
  OAI22D1BWP12T U2878 ( .A1(n2068), .A2(n2680), .B1(n2679), .B2(n2067), .ZN(
        n2078) );
  OAI22D1BWP12T U2879 ( .A1(n2070), .A2(n2684), .B1(n2683), .B2(n2069), .ZN(
        n2077) );
  OAI22D1BWP12T U2880 ( .A1(n2689), .A2(n2072), .B1(n2687), .B2(n2071), .ZN(
        n2076) );
  OAI22D1BWP12T U2881 ( .A1(n2693), .A2(n2074), .B1(n2691), .B2(n2073), .ZN(
        n2075) );
  NR4D0BWP12T U2882 ( .A1(n2078), .A2(n2077), .A3(n2076), .A4(n2075), .ZN(
        n2079) );
  ND2D1BWP12T U2883 ( .A1(n2080), .A2(n2079), .ZN(regB_out[20]) );
  OAI22D1BWP12T U2884 ( .A1(n2863), .A2(n2082), .B1(n2081), .B2(n2860), .ZN(
        n2092) );
  OAI22D0BWP12T U2885 ( .A1(n2867), .A2(n2084), .B1(n2083), .B2(n2864), .ZN(
        n2091) );
  OAI22D1BWP12T U2886 ( .A1(n2871), .A2(n2086), .B1(n2085), .B2(n2868), .ZN(
        n2090) );
  OAI22D1BWP12T U2887 ( .A1(n2875), .A2(n2088), .B1(n2087), .B2(n2872), .ZN(
        n2089) );
  NR4D0BWP12T U2888 ( .A1(n2092), .A2(n2091), .A3(n2090), .A4(n2089), .ZN(
        n2107) );
  OAI22D1BWP12T U2889 ( .A1(n2883), .A2(n2094), .B1(n2093), .B2(n2880), .ZN(
        n2098) );
  OAI22D1BWP12T U2890 ( .A1(n2887), .A2(n2096), .B1(n2095), .B2(n2884), .ZN(
        n2097) );
  AOI211D1BWP12T U2891 ( .A1(r2[6]), .A2(n2890), .B(n2098), .C(n2097), .ZN(
        n2106) );
  OAI22D1BWP12T U2892 ( .A1(n2829), .A2(n2100), .B1(n2099), .B2(n2826), .ZN(
        n2104) );
  OAI22D1BWP12T U2893 ( .A1(n2825), .A2(n2102), .B1(n2101), .B2(n2822), .ZN(
        n2103) );
  NR2D1BWP12T U2894 ( .A1(n2104), .A2(n2103), .ZN(n2105) );
  ND3D1BWP12T U2895 ( .A1(n2107), .A2(n2106), .A3(n2105), .ZN(regA_out[6]) );
  OAI22D1BWP12T U2896 ( .A1(n2863), .A2(n2109), .B1(n2108), .B2(n2860), .ZN(
        n2119) );
  OAI22D1BWP12T U2897 ( .A1(n2867), .A2(n2111), .B1(n2110), .B2(n2864), .ZN(
        n2118) );
  OAI22D1BWP12T U2898 ( .A1(n2871), .A2(n2113), .B1(n2112), .B2(n2868), .ZN(
        n2117) );
  OAI22D1BWP12T U2899 ( .A1(n2851), .A2(n2115), .B1(n2114), .B2(n2872), .ZN(
        n2116) );
  NR4D0BWP12T U2900 ( .A1(n2119), .A2(n2118), .A3(n2117), .A4(n2116), .ZN(
        n2134) );
  OAI22D1BWP12T U2901 ( .A1(n2883), .A2(n2121), .B1(n2120), .B2(n2880), .ZN(
        n2125) );
  OAI22D1BWP12T U2902 ( .A1(n2887), .A2(n2123), .B1(n2122), .B2(n2884), .ZN(
        n2124) );
  RCAOI211D0BWP12T U2903 ( .A1(r2[5]), .A2(n2890), .B(n2125), .C(n2124), .ZN(
        n2133) );
  OAI22D1BWP12T U2904 ( .A1(n2829), .A2(n2127), .B1(n2126), .B2(n2826), .ZN(
        n2131) );
  OAI22D1BWP12T U2905 ( .A1(n2825), .A2(n2129), .B1(n2128), .B2(n2822), .ZN(
        n2130) );
  NR2D1BWP12T U2906 ( .A1(n2131), .A2(n2130), .ZN(n2132) );
  ND3D1BWP12T U2907 ( .A1(n2134), .A2(n2133), .A3(n2132), .ZN(regA_out[5]) );
  AOI22D1BWP12T U2908 ( .A1(tmp1[18]), .A2(n2746), .B1(n2135), .B2(
        immediate2_in[18]), .ZN(n2655) );
  AOI22D1BWP12T U2909 ( .A1(r5[18]), .A2(n2748), .B1(n2747), .B2(r10[18]), 
        .ZN(n2649) );
  AOI22D1BWP12T U2910 ( .A1(r7[18]), .A2(n2750), .B1(n2749), .B2(r2[18]), .ZN(
        n2137) );
  ND2D1BWP12T U2911 ( .A1(n2649), .A2(n2137), .ZN(n2654) );
  AOI22D1BWP12T U2912 ( .A1(r9[18]), .A2(n105), .B1(n2753), .B2(r4[18]), .ZN(
        n2652) );
  AOI22D1BWP12T U2913 ( .A1(r11[18]), .A2(n2755), .B1(n2650), .B2(r0[18]), 
        .ZN(n2651) );
  ND2D1BWP12T U2914 ( .A1(n2652), .A2(n2651), .ZN(n2653) );
  INR3XD0BWP12T U2915 ( .A1(n2655), .B1(n2654), .B2(n2653), .ZN(n2661) );
  AOI22D1BWP12T U2916 ( .A1(r1[18]), .A2(n118), .B1(n2761), .B2(r12[18]), .ZN(
        n2659) );
  AOI22D1BWP12T U2917 ( .A1(r3[18]), .A2(n2763), .B1(n2762), .B2(lr[18]), .ZN(
        n2658) );
  AOI22D1BWP12T U2918 ( .A1(r8[18]), .A2(n2765), .B1(n2764), .B2(n[2950]), 
        .ZN(n2657) );
  AOI22D1BWP12T U2919 ( .A1(pc_out[18]), .A2(n2767), .B1(n2766), .B2(r6[18]), 
        .ZN(n2656) );
  AN4XD1BWP12T U2920 ( .A1(n2659), .A2(n2658), .A3(n2657), .A4(n2656), .Z(
        n2660) );
  ND2D1BWP12T U2921 ( .A1(n2661), .A2(n2660), .ZN(regB_out[18]) );
  OAI22D1BWP12T U2922 ( .A1(n2665), .A2(n2664), .B1(n2663), .B2(n2662), .ZN(
        n2677) );
  MOAI22D0BWP12T U2923 ( .A1(n2667), .A2(n2666), .B1(n2730), .B2(
        immediate2_in[17]), .ZN(n2676) );
  AOI22D1BWP12T U2924 ( .A1(r9[17]), .A2(n105), .B1(n2753), .B2(r4[17]), .ZN(
        n2669) );
  AOI22D1BWP12T U2925 ( .A1(r11[17]), .A2(n2755), .B1(n2754), .B2(r0[17]), 
        .ZN(n2668) );
  ND2D1BWP12T U2926 ( .A1(n2669), .A2(n2668), .ZN(n2675) );
  OAI22D1BWP12T U2927 ( .A1(n2673), .A2(n2672), .B1(n2671), .B2(n2670), .ZN(
        n2674) );
  OAI22D1BWP12T U2928 ( .A1(n2681), .A2(n2680), .B1(n2679), .B2(n2678), .ZN(
        n2697) );
  OAI22D1BWP12T U2929 ( .A1(n2685), .A2(n2684), .B1(n2683), .B2(n2682), .ZN(
        n2696) );
  OAI22D1BWP12T U2930 ( .A1(n2689), .A2(n2688), .B1(n2687), .B2(n2686), .ZN(
        n2695) );
  INVD0BWP12T U2931 ( .I(pc_out[17]), .ZN(n2692) );
  OAI22D1BWP12T U2932 ( .A1(n2693), .A2(n2692), .B1(n2691), .B2(n2690), .ZN(
        n2694) );
  NR4D0BWP12T U2933 ( .A1(n2697), .A2(n2696), .A3(n2695), .A4(n2694), .ZN(
        n2698) );
  ND2D1BWP12T U2934 ( .A1(n2699), .A2(n2698), .ZN(regB_out[17]) );
  NR2D1BWP12T U2935 ( .A1(n2868), .A2(n2700), .ZN(n2701) );
  AOI21D1BWP12T U2936 ( .A1(n2776), .A2(pc_out[8]), .B(n2701), .ZN(n2713) );
  ND2D1BWP12T U2937 ( .A1(n2807), .A2(n[2960]), .ZN(n2702) );
  OAI21D1BWP12T U2938 ( .A1(n2864), .A2(n2703), .B(n2702), .ZN(n2712) );
  NR2D1BWP12T U2939 ( .A1(n2860), .A2(n2704), .ZN(n2705) );
  AOI21D1BWP12T U2940 ( .A1(n2809), .A2(r5[8]), .B(n2705), .ZN(n2710) );
  NR2D1BWP12T U2941 ( .A1(n2872), .A2(n2706), .ZN(n2707) );
  AOI21D1BWP12T U2942 ( .A1(n2708), .A2(r12[8]), .B(n2707), .ZN(n2709) );
  ND2D1BWP12T U2943 ( .A1(n2710), .A2(n2709), .ZN(n2711) );
  INR3D0BWP12T U2944 ( .A1(n2713), .B1(n2712), .B2(n2711), .ZN(n2729) );
  NR2D1BWP12T U2945 ( .A1(n2884), .A2(n2714), .ZN(n2715) );
  AOI21D1BWP12T U2946 ( .A1(n2791), .A2(r4[8]), .B(n2715), .ZN(n2727) );
  NR2D1BWP12T U2947 ( .A1(n2880), .A2(n2716), .ZN(n2717) );
  AOI21D1BWP12T U2948 ( .A1(n2819), .A2(r9[8]), .B(n2717), .ZN(n2718) );
  IOA21D1BWP12T U2949 ( .A1(n2890), .A2(r2[8]), .B(n2718), .ZN(n2726) );
  NR2D1BWP12T U2950 ( .A1(n2822), .A2(n2719), .ZN(n2720) );
  AOI21D0BWP12T U2951 ( .A1(n2891), .A2(lr[8]), .B(n2720), .ZN(n2724) );
  NR2D1BWP12T U2952 ( .A1(n2826), .A2(n2721), .ZN(n2722) );
  TPAOI21D0BWP12T U2953 ( .A1(n2893), .A2(r10[8]), .B(n2722), .ZN(n2723) );
  CKND2D1BWP12T U2954 ( .A1(n2724), .A2(n2723), .ZN(n2725) );
  INR3D0BWP12T U2955 ( .A1(n2727), .B1(n2726), .B2(n2725), .ZN(n2728) );
  ND2D1BWP12T U2956 ( .A1(n2729), .A2(n2728), .ZN(regA_out[8]) );
  AOI22D1BWP12T U2957 ( .A1(tmp1[16]), .A2(n2746), .B1(n2730), .B2(
        immediate2_in[16]), .ZN(n2738) );
  AOI22D1BWP12T U2958 ( .A1(r5[16]), .A2(n2748), .B1(n2747), .B2(r10[16]), 
        .ZN(n2732) );
  AOI22D1BWP12T U2959 ( .A1(r7[16]), .A2(n2750), .B1(n2749), .B2(r2[16]), .ZN(
        n2731) );
  ND2D1BWP12T U2960 ( .A1(n2732), .A2(n2731), .ZN(n2737) );
  AOI22D1BWP12T U2961 ( .A1(r9[16]), .A2(n105), .B1(n2753), .B2(r4[16]), .ZN(
        n2735) );
  AOI22D1BWP12T U2962 ( .A1(r11[16]), .A2(n2755), .B1(n2733), .B2(r0[16]), 
        .ZN(n2734) );
  ND2D1BWP12T U2963 ( .A1(n2735), .A2(n2734), .ZN(n2736) );
  INR3XD0BWP12T U2964 ( .A1(n2738), .B1(n2737), .B2(n2736), .ZN(n2744) );
  AOI22D1BWP12T U2965 ( .A1(r1[16]), .A2(n118), .B1(n2761), .B2(r12[16]), .ZN(
        n2742) );
  AOI22D1BWP12T U2966 ( .A1(r3[16]), .A2(n2763), .B1(n2762), .B2(lr[16]), .ZN(
        n2741) );
  AOI22D1BWP12T U2967 ( .A1(r8[16]), .A2(n2765), .B1(n2764), .B2(n[2952]), 
        .ZN(n2740) );
  AOI22D1BWP12T U2968 ( .A1(pc_out[16]), .A2(n2767), .B1(n2766), .B2(r6[16]), 
        .ZN(n2739) );
  AN4XD1BWP12T U2969 ( .A1(n2742), .A2(n2741), .A3(n2740), .A4(n2739), .Z(
        n2743) );
  ND2D1BWP12T U2970 ( .A1(n2744), .A2(n2743), .ZN(regB_out[16]) );
  AOI22D1BWP12T U2971 ( .A1(tmp1[15]), .A2(n2746), .B1(n2745), .B2(
        immediate2_in[15]), .ZN(n2760) );
  AOI22D1BWP12T U2972 ( .A1(r5[15]), .A2(n2748), .B1(n2747), .B2(r10[15]), 
        .ZN(n2752) );
  AOI22D1BWP12T U2973 ( .A1(r7[15]), .A2(n2750), .B1(n2749), .B2(r2[15]), .ZN(
        n2751) );
  ND2D1BWP12T U2974 ( .A1(n2752), .A2(n2751), .ZN(n2759) );
  AOI22D1BWP12T U2975 ( .A1(r9[15]), .A2(n105), .B1(n2753), .B2(r4[15]), .ZN(
        n2757) );
  AOI22D1BWP12T U2976 ( .A1(r11[15]), .A2(n2755), .B1(n2754), .B2(r0[15]), 
        .ZN(n2756) );
  ND2D1BWP12T U2977 ( .A1(n2757), .A2(n2756), .ZN(n2758) );
  INR3XD0BWP12T U2978 ( .A1(n2760), .B1(n2759), .B2(n2758), .ZN(n2773) );
  AOI22D1BWP12T U2979 ( .A1(r1[15]), .A2(n118), .B1(n2761), .B2(r12[15]), .ZN(
        n2771) );
  AOI22D1BWP12T U2980 ( .A1(r3[15]), .A2(n2763), .B1(n2762), .B2(lr[15]), .ZN(
        n2770) );
  AOI22D1BWP12T U2981 ( .A1(r8[15]), .A2(n2765), .B1(n2764), .B2(n[2953]), 
        .ZN(n2769) );
  AOI22D1BWP12T U2982 ( .A1(pc_out[15]), .A2(n2767), .B1(n2766), .B2(r6[15]), 
        .ZN(n2768) );
  AN4XD1BWP12T U2983 ( .A1(n2771), .A2(n2770), .A3(n2769), .A4(n2768), .Z(
        n2772) );
  ND2D1BWP12T U2984 ( .A1(n2773), .A2(n2772), .ZN(regB_out[15]) );
  NR2D1BWP12T U2985 ( .A1(n2868), .A2(n2774), .ZN(n2775) );
  AOI21D1BWP12T U2986 ( .A1(n2776), .A2(pc_out[10]), .B(n2775), .ZN(n2787) );
  ND2D1BWP12T U2987 ( .A1(n2807), .A2(n[2958]), .ZN(n2777) );
  OAI21D1BWP12T U2988 ( .A1(n2864), .A2(n2778), .B(n2777), .ZN(n2786) );
  NR2D1BWP12T U2989 ( .A1(n2860), .A2(n2779), .ZN(n2780) );
  AOI21D1BWP12T U2990 ( .A1(n2809), .A2(r5[10]), .B(n2780), .ZN(n2784) );
  NR2D1BWP12T U2991 ( .A1(n2872), .A2(n2781), .ZN(n2782) );
  AOI21D1BWP12T U2992 ( .A1(n2813), .A2(r12[10]), .B(n2782), .ZN(n2783) );
  ND2D1BWP12T U2993 ( .A1(n2784), .A2(n2783), .ZN(n2785) );
  INR3D0BWP12T U2994 ( .A1(n2787), .B1(n2786), .B2(n2785), .ZN(n2806) );
  NR2D1BWP12T U2995 ( .A1(n2789), .A2(n2788), .ZN(n2790) );
  AOI21D1BWP12T U2996 ( .A1(n2791), .A2(r4[10]), .B(n2790), .ZN(n2804) );
  NR2D1BWP12T U2997 ( .A1(n2880), .A2(n2792), .ZN(n2793) );
  AOI21D1BWP12T U2998 ( .A1(n2819), .A2(r9[10]), .B(n2793), .ZN(n2794) );
  IOA21D1BWP12T U2999 ( .A1(r0[10]), .A2(n2795), .B(n2794), .ZN(n2803) );
  NR2D1BWP12T U3000 ( .A1(n2822), .A2(n2796), .ZN(n2797) );
  AOI21D0BWP12T U3001 ( .A1(n2891), .A2(lr[10]), .B(n2797), .ZN(n2801) );
  NR2D1BWP12T U3002 ( .A1(n2826), .A2(n2798), .ZN(n2799) );
  TPAOI21D0BWP12T U3003 ( .A1(n2893), .A2(r10[10]), .B(n2799), .ZN(n2800) );
  CKND2D1BWP12T U3004 ( .A1(n2801), .A2(n2800), .ZN(n2802) );
  INR3D0BWP12T U3005 ( .A1(n2804), .B1(n2803), .B2(n2802), .ZN(n2805) );
  ND2D1BWP12T U3006 ( .A1(n2806), .A2(n2805), .ZN(regA_out[10]) );
  AOI22D1BWP12T U3007 ( .A1(n2808), .A2(r11[25]), .B1(n2807), .B2(n[2943]), 
        .ZN(n2818) );
  AOI22D1BWP12T U3008 ( .A1(r3[25]), .A2(n2810), .B1(n2809), .B2(r5[25]), .ZN(
        n2817) );
  AOI22D1BWP12T U3009 ( .A1(n2812), .A2(r7[25]), .B1(n2811), .B2(pc_out[25]), 
        .ZN(n2816) );
  AOI22D1BWP12T U3010 ( .A1(n2814), .A2(r1[25]), .B1(n2813), .B2(r12[25]), 
        .ZN(n2815) );
  AN4XD1BWP12T U3011 ( .A1(n2818), .A2(n2817), .A3(n2816), .A4(n2815), .Z(
        n2837) );
  AOI22D1BWP12T U3012 ( .A1(tmp1[25]), .A2(n2820), .B1(n2819), .B2(r9[25]), 
        .ZN(n2821) );
  IOA21D1BWP12T U3013 ( .A1(r2[25]), .A2(n2890), .B(n2821), .ZN(n2835) );
  INVD1BWP12T U3014 ( .I(lr[25]), .ZN(n2824) );
  OAI22D1BWP12T U3015 ( .A1(n2825), .A2(n2824), .B1(n2823), .B2(n2822), .ZN(
        n2834) );
  INVD1BWP12T U3016 ( .I(r10[25]), .ZN(n2828) );
  INVD1BWP12T U3017 ( .I(r6[25]), .ZN(n2827) );
  OAI22D1BWP12T U3018 ( .A1(n2829), .A2(n2828), .B1(n2827), .B2(n2826), .ZN(
        n2833) );
  INVD1BWP12T U3019 ( .I(r4[25]), .ZN(n2831) );
  INVD1BWP12T U3020 ( .I(r0[25]), .ZN(n2830) );
  OAI22D1BWP12T U3021 ( .A1(n2887), .A2(n2831), .B1(n2830), .B2(n2884), .ZN(
        n2832) );
  NR4D0BWP12T U3022 ( .A1(n2835), .A2(n2834), .A3(n2833), .A4(n2832), .ZN(
        n2836) );
  ND2D1BWP12T U3023 ( .A1(n2837), .A2(n2836), .ZN(regA_out[25]) );
  INVD1BWP12T U3024 ( .I(r9[24]), .ZN(n2839) );
  OAI22D1BWP12T U3025 ( .A1(n2883), .A2(n2839), .B1(n2838), .B2(n2880), .ZN(
        n2843) );
  INVD1BWP12T U3026 ( .I(r4[24]), .ZN(n2841) );
  INVD1BWP12T U3027 ( .I(r0[24]), .ZN(n2840) );
  OAI22D1BWP12T U3028 ( .A1(n2887), .A2(n2841), .B1(n2840), .B2(n2884), .ZN(
        n2842) );
  AOI211D1BWP12T U3029 ( .A1(r2[24]), .A2(n2890), .B(n2843), .C(n2842), .ZN(
        n2859) );
  INVD1BWP12T U3030 ( .I(r3[24]), .ZN(n2844) );
  OAI22D1BWP12T U3031 ( .A1(n2863), .A2(n2845), .B1(n2844), .B2(n2860), .ZN(
        n2855) );
  INVD1BWP12T U3032 ( .I(r11[24]), .ZN(n2846) );
  OAI22D0BWP12T U3033 ( .A1(n2867), .A2(n2847), .B1(n2846), .B2(n2864), .ZN(
        n2854) );
  INVD1BWP12T U3034 ( .I(pc_out[24]), .ZN(n2901) );
  OAI22D1BWP12T U3035 ( .A1(n2871), .A2(n2901), .B1(n2848), .B2(n2868), .ZN(
        n2853) );
  INVD1BWP12T U3036 ( .I(r1[24]), .ZN(n2849) );
  OAI22D1BWP12T U3037 ( .A1(n2851), .A2(n2850), .B1(n2849), .B2(n2872), .ZN(
        n2852) );
  NR4D0BWP12T U3038 ( .A1(n2855), .A2(n2854), .A3(n2853), .A4(n2852), .ZN(
        n2858) );
  AOI22D1BWP12T U3039 ( .A1(n2892), .A2(r8[24]), .B1(n2891), .B2(lr[24]), .ZN(
        n2857) );
  AOI22D1BWP12T U3040 ( .A1(r6[24]), .A2(n2894), .B1(n2893), .B2(r10[24]), 
        .ZN(n2856) );
  ND4D1BWP12T U3041 ( .A1(n2859), .A2(n2858), .A3(n2857), .A4(n2856), .ZN(
        regA_out[24]) );
  INVD1BWP12T U3042 ( .I(r3[23]), .ZN(n2861) );
  OAI22D1BWP12T U3043 ( .A1(n2863), .A2(n2862), .B1(n2861), .B2(n2860), .ZN(
        n2879) );
  INVD1BWP12T U3044 ( .I(n[2945]), .ZN(n2866) );
  OAI22D0BWP12T U3045 ( .A1(n2867), .A2(n2866), .B1(n2865), .B2(n2864), .ZN(
        n2878) );
  INVD1BWP12T U3046 ( .I(pc_out[23]), .ZN(n2870) );
  OAI22D1BWP12T U3047 ( .A1(n2871), .A2(n2870), .B1(n2869), .B2(n2868), .ZN(
        n2877) );
  INVD1BWP12T U3048 ( .I(r12[23]), .ZN(n2874) );
  INVD1BWP12T U3049 ( .I(r1[23]), .ZN(n2873) );
  OAI22D1BWP12T U3050 ( .A1(n2875), .A2(n2874), .B1(n2873), .B2(n2872), .ZN(
        n2876) );
  NR4D0BWP12T U3051 ( .A1(n2879), .A2(n2878), .A3(n2877), .A4(n2876), .ZN(
        n2898) );
  INVD1BWP12T U3052 ( .I(r9[23]), .ZN(n2882) );
  OAI22D1BWP12T U3053 ( .A1(n2883), .A2(n2882), .B1(n2881), .B2(n2880), .ZN(
        n2889) );
  INVD1BWP12T U3054 ( .I(r4[23]), .ZN(n2886) );
  INVD1BWP12T U3055 ( .I(r0[23]), .ZN(n2885) );
  OAI22D1BWP12T U3056 ( .A1(n2887), .A2(n2886), .B1(n2885), .B2(n2884), .ZN(
        n2888) );
  AOI211D1BWP12T U3057 ( .A1(r2[23]), .A2(n2890), .B(n2889), .C(n2888), .ZN(
        n2897) );
  AOI22D1BWP12T U3058 ( .A1(n2892), .A2(r8[23]), .B1(n2891), .B2(lr[23]), .ZN(
        n2896) );
  AOI22D1BWP12T U3059 ( .A1(r6[23]), .A2(n2894), .B1(n2893), .B2(r10[23]), 
        .ZN(n2895) );
  ND4D1BWP12T U3060 ( .A1(n2898), .A2(n2897), .A3(n2896), .A4(n2895), .ZN(
        regA_out[23]) );
  TPND3D0BWP12T U3061 ( .A1(n2900), .A2(n2906), .A3(n2914), .ZN(n2899) );
  NR2XD0BWP12T U3062 ( .A1(n2905), .A2(n2899), .ZN(n2909) );
  TPNR2D0BWP12T U3063 ( .A1(n2900), .A2(n2919), .ZN(n2904) );
  CKND1BWP12T U3064 ( .I(n2906), .ZN(n2903) );
  AOI21D1BWP12T U3065 ( .A1(n2904), .A2(n2903), .B(n2902), .ZN(n2908) );
  IND3D1BWP12T U3066 ( .A1(n2906), .B1(n2914), .B2(n2905), .ZN(n2907) );
  IND3D1BWP12T U3067 ( .A1(n2909), .B1(n2908), .B2(n2907), .ZN(n2193) );
  AO21D0BWP12T U3068 ( .A1(write1_in[28]), .A2(n2920), .B(n2910), .Z(n2913) );
  ND3D2BWP12T U3069 ( .A1(n2913), .A2(n2912), .A3(n2911), .ZN(n2935) );
  INR2D1BWP12T U3070 ( .A1(n2914), .B1(n2931), .ZN(n2934) );
  INVD2BWP12T U3071 ( .I(n2935), .ZN(n2932) );
  AOI21D0BWP12T U3072 ( .A1(n2916), .A2(n2915), .B(n2919), .ZN(n2917) );
  OA21XD0BWP12T U3073 ( .A1(write1_in[29]), .A2(n2918), .B(n2917), .Z(n2930)
         );
  IAO21D0BWP12T U3074 ( .A1(n2922), .A2(n2920), .B(n2919), .ZN(n2921) );
  OAI21D1BWP12T U3075 ( .A1(write1_in[30]), .A2(n2922), .B(n2921), .ZN(n2928)
         );
  TPNR2D0BWP12T U3076 ( .A1(n2924), .A2(n2923), .ZN(n2925) );
  AOI21D1BWP12T U3077 ( .A1(next_pc_in[30]), .A2(n1488), .B(n2925), .ZN(n2926)
         );
  OAI21D1BWP12T U3078 ( .A1(n2928), .A2(n2927), .B(n2926), .ZN(n2929) );
  TPAOI31D1BWP12T U3079 ( .A1(n2932), .A2(n2931), .A3(n2930), .B(n2929), .ZN(
        n2933) );
  IOA21D1BWP12T U3080 ( .A1(n2935), .A2(n2934), .B(n2933), .ZN(n2199) );
endmodule


module ALU_VARIABLE ( a, b, op, c_in, result, c_out, z, n, v );
  input [31:0] a;
  input [31:0] b;
  input [3:0] op;
  output [31:0] result;
  input c_in;
  output c_out, z, n, v;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218;

  OAI22D1BWP12T U3 ( .A1(n2130), .A2(n817), .B1(n754), .B2(n829), .ZN(n824) );
  TPND2D1BWP12T U4 ( .A1(n2003), .A2(n1516), .ZN(n2005) );
  XNR2D1BWP12T U5 ( .A1(n1977), .A2(n3938), .ZN(n1252) );
  INVD1BWP12T U6 ( .I(n1421), .ZN(n3135) );
  AOI21D1BWP12T U7 ( .A1(n2227), .A2(n2225), .B(n1726), .ZN(n3508) );
  CKBD1BWP12T U8 ( .I(b[27]), .Z(n3942) );
  IND2D1BWP12T U9 ( .A1(n1469), .B1(n1242), .ZN(n1254) );
  FA1D0BWP12T U10 ( .A(n768), .B(n767), .CI(n766), .CO(n792), .S(n770) );
  OAI22D1BWP12T U11 ( .A1(n2088), .A2(n816), .B1(n2086), .B2(n815), .ZN(n825)
         );
  INVD2BWP12T U12 ( .I(n3911), .ZN(n4089) );
  XNR2D1BWP12T U13 ( .A1(n1977), .A2(n3942), .ZN(n1592) );
  HA1D0BWP12T U14 ( .A(n1887), .B(n1886), .CO(n1993), .S(n1914) );
  OAI22D1BWP12T U15 ( .A1(n2023), .A2(n1343), .B1(n2021), .B2(n1525), .ZN(
        n1529) );
  FA1D0BWP12T U16 ( .A(n1638), .B(n1637), .CI(n1636), .CO(n1885), .S(n1634) );
  CKBD1BWP12T U17 ( .I(n1911), .Z(n2100) );
  FA1D0BWP12T U18 ( .A(n1899), .B(n1898), .CI(n1897), .CO(n1972), .S(n1904) );
  OAI22D1BWP12T U19 ( .A1(n2130), .A2(n829), .B1(n754), .B2(n867), .ZN(n881)
         );
  OAI22D1BWP12T U20 ( .A1(n2019), .A2(n888), .B1(n1282), .B2(n2018), .ZN(n1384) );
  OAI22D1BWP12T U21 ( .A1(n2079), .A2(n1184), .B1(n2077), .B2(n1371), .ZN(
        n1369) );
  FA1D0BWP12T U22 ( .A(n1366), .B(n1365), .CI(n1364), .CO(n1556), .S(n1352) );
  FA1D0BWP12T U23 ( .A(n1667), .B(n1666), .CI(n1665), .CO(n1922), .S(n1658) );
  FA1D0BWP12T U24 ( .A(n1559), .B(n1558), .CI(n1557), .CO(n1601), .S(n1615) );
  OAI22D1BWP12T U25 ( .A1(n2083), .A2(n1294), .B1(n2080), .B2(n1293), .ZN(
        n1404) );
  OAI22D1BWP12T U26 ( .A1(n2072), .A2(n1296), .B1(n2070), .B2(n1295), .ZN(
        n1403) );
  OAI22D1BWP12T U27 ( .A1(n2127), .A2(n1166), .B1(n2125), .B2(n1173), .ZN(
        n1220) );
  CKBD1BWP12T U28 ( .I(n3916), .Z(n1962) );
  FA1D0BWP12T U29 ( .A(n1922), .B(n1921), .CI(n1920), .CO(n1935), .S(n1862) );
  FA1D0BWP12T U30 ( .A(n2054), .B(n2053), .CI(n2052), .CO(n2096), .S(n2040) );
  FA1D0BWP12T U31 ( .A(n2048), .B(n2047), .CI(n2046), .CO(n2149), .S(n2151) );
  ND2D1BWP12T U32 ( .A1(n1394), .A2(n1393), .ZN(n1446) );
  MUX2D1BWP12T U33 ( .I0(n4075), .I1(n4081), .S(b[0]), .Z(n2823) );
  INVD1BWP12T U34 ( .I(n338), .ZN(n718) );
  OAI22D1BWP12T U35 ( .A1(n2127), .A2(n1156), .B1(n2125), .B2(n1166), .ZN(
        n1177) );
  INR2D1BWP12T U36 ( .A1(n1979), .B1(n2077), .ZN(n1300) );
  OAI22D1BWP12T U37 ( .A1(n2019), .A2(n1281), .B1(n1252), .B2(n2018), .ZN(
        n1301) );
  FA1D0BWP12T U38 ( .A(n1206), .B(n1205), .CI(n1204), .CO(n1333), .S(n1228) );
  OAI21D1BWP12T U39 ( .A1(n1688), .A2(n1687), .B(n1686), .ZN(n1690) );
  XOR3D1BWP12T U40 ( .A1(n1484), .A2(n1483), .A3(n1482), .Z(n1485) );
  INVD1BWP12T U41 ( .I(n3942), .ZN(n3851) );
  CKBD1BWP12T U42 ( .I(b[28]), .Z(n3944) );
  INVD1BWP12T U43 ( .I(n2641), .ZN(n2949) );
  XNR2D1BWP12T U44 ( .A1(n1517), .A2(n4082), .ZN(n817) );
  OAI22D1BWP12T U45 ( .A1(n1110), .A2(n787), .B1(n789), .B2(n2018), .ZN(n797)
         );
  OAI22D1BWP12T U46 ( .A1(n2072), .A2(n788), .B1(n2070), .B2(n828), .ZN(n795)
         );
  FA1D0BWP12T U47 ( .A(n1245), .B(n1244), .CI(n1243), .CO(n1225), .S(n1260) );
  OAI22D1BWP12T U48 ( .A1(n2079), .A2(n1155), .B1(n2077), .B2(n1154), .ZN(
        n1244) );
  NR2D1BWP12T U49 ( .A1(n1498), .A2(n1497), .ZN(n3089) );
  HA1D0BWP12T U50 ( .A(n725), .B(n724), .CO(n749), .S(n734) );
  OAI22D1BWP12T U51 ( .A1(n2009), .A2(n719), .B1(n764), .B2(n2006), .ZN(n758)
         );
  ND2D1BWP12T U52 ( .A1(n1927), .A2(n1926), .ZN(n2746) );
  OAI21D1BWP12T U53 ( .A1(n2694), .A2(n2844), .B(n2695), .ZN(n2742) );
  ND2D1BWP12T U54 ( .A1(n1692), .A2(n1691), .ZN(n2739) );
  INVD1BWP12T U55 ( .I(n4089), .ZN(n3395) );
  INR2D1BWP12T U56 ( .A1(b[0]), .B1(n3780), .ZN(n2632) );
  ND2D1BWP12T U57 ( .A1(n1502), .A2(n1501), .ZN(n3046) );
  OAI21D1BWP12T U58 ( .A1(n3508), .A2(n3506), .B(n3507), .ZN(n3001) );
  INVD1BWP12T U59 ( .I(n4076), .ZN(n3896) );
  BUFFD2BWP12T U60 ( .I(a[26]), .Z(n4076) );
  ND2D1BWP12T U61 ( .A1(n3505), .A2(n4173), .ZN(n2218) );
  INVD1BWP12T U62 ( .I(n2470), .ZN(n2463) );
  OAI21D1BWP12T U63 ( .A1(n3120), .A2(n3118), .B(n3123), .ZN(n3057) );
  NR3D1BWP12T U64 ( .A1(n539), .A2(n538), .A3(n537), .ZN(n550) );
  AOI21D1BWP12T U65 ( .A1(n2847), .A2(n2845), .B(n2693), .ZN(n2698) );
  FA1D0BWP12T U66 ( .A(n3395), .B(n2207), .CI(n3394), .CO(n3396), .S(n3609) );
  XOR2D1BWP12T U67 ( .A1(n3134), .A2(n896), .Z(n3435) );
  AOI21D1BWP12T U68 ( .A1(n3134), .A2(n317), .B(n3133), .ZN(n3139) );
  AO21D1BWP12T U69 ( .A1(n3450), .A2(n140), .B(n1782), .Z(result[29]) );
  INVD1BWP12T U70 ( .I(b[5]), .ZN(n3842) );
  DEL025D1BWP12T U71 ( .I(b[18]), .Z(n3951) );
  DEL025D1BWP12T U72 ( .I(b[21]), .Z(n3939) );
  OAI21D1BWP12T U73 ( .A1(n1323), .A2(n1262), .B(n1261), .ZN(n1271) );
  AOI21D1BWP12T U74 ( .A1(n3057), .A2(n3056), .B(n2238), .ZN(n2233) );
  INVD1BWP12T U75 ( .I(a[31]), .ZN(n3911) );
  INVD1BWP12T U76 ( .I(n4078), .ZN(n3876) );
  XNR2D1BWP12T U77 ( .A1(n4044), .A2(n2629), .ZN(n3300) );
  IOA21D1BWP12T U78 ( .A1(n3444), .A2(n4171), .B(n3329), .ZN(result[21]) );
  RCOAI21D1BWP12T U79 ( .A1(n2178), .A2(n3407), .B(n2177), .ZN(v) );
  CKBD1BWP12T U80 ( .I(result[31]), .Z(n) );
  AO21D1BWP12T U81 ( .A1(n3420), .A2(n4171), .B(n2843), .Z(result[9]) );
  CKBD1BWP12T U82 ( .I(n340), .Z(n1110) );
  ND2D1BWP12T U83 ( .A1(n468), .A2(n467), .ZN(n2795) );
  INVD2BWP12T U84 ( .I(n3840), .ZN(n3929) );
  INVD1BWP12T U85 ( .I(n3916), .ZN(n582) );
  INVD3BWP12T U86 ( .I(n2668), .ZN(n4067) );
  BUFFD2BWP12T U87 ( .I(a[6]), .Z(n4083) );
  INVD1BWP12T U88 ( .I(n3928), .ZN(n1909) );
  BUFFD2BWP12T U89 ( .I(a[8]), .Z(n4062) );
  INVD1BWP12T U90 ( .I(n3957), .ZN(n1959) );
  INVD1BWP12T U91 ( .I(n3933), .ZN(n3833) );
  INVD2BWP12T U92 ( .I(n3832), .ZN(n3928) );
  ND2D1BWP12T U93 ( .A1(n372), .A2(n371), .ZN(n2363) );
  TPNR2D1BWP12T U94 ( .A1(n691), .A2(n690), .ZN(n2367) );
  CKND2D2BWP12T U95 ( .A1(n348), .A2(n347), .ZN(n1986) );
  INVD1BWP12T U96 ( .I(n2281), .ZN(n777) );
  XOR3D1BWP12T U97 ( .A1(n841), .A2(n840), .A3(n839), .Z(n846) );
  INVD1BWP12T U98 ( .I(n3950), .ZN(n3829) );
  INVD1BWP12T U99 ( .I(n3931), .ZN(n3830) );
  INVD1BWP12T U100 ( .I(n3930), .ZN(n3827) );
  INVD1BWP12T U101 ( .I(n3949), .ZN(n3828) );
  INVD1BWP12T U102 ( .I(n4191), .ZN(n3821) );
  INVD1BWP12T U103 ( .I(n3952), .ZN(n3826) );
  INVD1BWP12T U104 ( .I(n3951), .ZN(n3819) );
  BUFFD2BWP12T U105 ( .I(b[12]), .Z(n3950) );
  BUFFD2BWP12T U106 ( .I(a[12]), .Z(n4078) );
  INVD1BWP12T U107 ( .I(n4061), .ZN(n3877) );
  INVD1BWP12T U108 ( .I(n3487), .ZN(n3276) );
  INVD1BWP12T U109 ( .I(n3938), .ZN(n3817) );
  INR2D1BWP12T U110 ( .A1(n1741), .B1(n3579), .ZN(n2236) );
  BUFFD2BWP12T U111 ( .I(b[24]), .Z(n3918) );
  OR2XD1BWP12T U112 ( .A1(n3921), .A2(n3922), .Z(n2955) );
  NR2D1BWP12T U113 ( .A1(n3886), .A2(n3916), .ZN(n3242) );
  INVD1BWP12T U114 ( .I(n1724), .ZN(n3519) );
  INVD3BWP12T U115 ( .I(n3922), .ZN(n4044) );
  TPNR2D1BWP12T U116 ( .A1(n3170), .A2(n3300), .ZN(n4179) );
  INVD1BWP12T U117 ( .I(n2667), .ZN(n4182) );
  INR2D1BWP12T U118 ( .A1(n4182), .B1(n3910), .ZN(n4184) );
  INVD1BWP12T U119 ( .I(n4181), .ZN(n4185) );
  INVD1BWP12T U120 ( .I(n4183), .ZN(n4187) );
  INVD1BWP12T U121 ( .I(n4163), .ZN(n4201) );
  OAI22D1BWP12T U122 ( .A1(n2019), .A2(n404), .B1(n412), .B2(n2018), .ZN(n416)
         );
  RCOAI21D1BWP12T U123 ( .A1(n2279), .A2(n3407), .B(n2278), .ZN(result[24]) );
  XNR2D1BWP12T U124 ( .A1(n1977), .A2(n1189), .ZN(n385) );
  OAI22D1BWP12T U125 ( .A1(n2072), .A2(n351), .B1(n2070), .B2(n362), .ZN(n367)
         );
  INR2D1BWP12T U126 ( .A1(n370), .B1(n372), .ZN(n689) );
  INVD1BWP12T U127 ( .I(n3921), .ZN(n583) );
  INVD1BWP12T U128 ( .I(n3920), .ZN(n588) );
  INVD1BWP12T U129 ( .I(n3929), .ZN(n594) );
  INVD1BWP12T U130 ( .I(n3927), .ZN(n589) );
  OAI22D1BWP12T U131 ( .A1(n2072), .A2(n673), .B1(n2070), .B2(n701), .ZN(n721)
         );
  OAI22D1BWP12T U132 ( .A1(n2009), .A2(n678), .B1(n713), .B2(n2006), .ZN(n727)
         );
  OAI22D1BWP12T U133 ( .A1(n2088), .A2(n697), .B1(n2086), .B2(n710), .ZN(n715)
         );
  OAI22D1BWP12T U134 ( .A1(n2083), .A2(n700), .B1(n717), .B2(n2080), .ZN(n706)
         );
  NR2D1BWP12T U135 ( .A1(n3930), .A2(a[14]), .ZN(n2910) );
  AOI21D1BWP12T U136 ( .A1(n3098), .A2(n3097), .B(n1725), .ZN(n3052) );
  AN2D1BWP12T U137 ( .A1(n319), .A2(n3452), .Z(n2223) );
  FA1D0BWP12T U138 ( .A(n425), .B(n424), .CI(n423), .CO(n428), .S(n410) );
  HA1D0BWP12T U139 ( .A(n388), .B(n387), .CO(n389), .S(n383) );
  INVD2BWP12T U140 ( .I(n3443), .ZN(n2279) );
  CKND0BWP12T U141 ( .I(n4044), .ZN(n1) );
  MAOI22D0BWP12T U142 ( .A1(n2388), .A2(n1), .B1(n3356), .B2(n2420), .ZN(n2)
         );
  OAI211D0BWP12T U143 ( .A1(n2955), .A2(n2414), .B(n3841), .C(n2), .ZN(n2404)
         );
  CKND2D0BWP12T U144 ( .A1(n2912), .A2(n2905), .ZN(n3) );
  CKND0BWP12T U145 ( .I(n2910), .ZN(n4) );
  AOI32D0BWP12T U146 ( .A1(n2907), .A2(n4), .A3(n2962), .B1(n2908), .B2(n4), 
        .ZN(n5) );
  IND4D0BWP12T U147 ( .A1(n3388), .B1(n2907), .B2(n2958), .B3(n4), .ZN(n6) );
  ND3D0BWP12T U148 ( .A1(n2909), .A2(n5), .A3(n6), .ZN(n7) );
  MOAI22D0BWP12T U149 ( .A1(n3), .A2(n7), .B1(n3), .B2(n7), .ZN(n3566) );
  CKND2D0BWP12T U150 ( .A1(n3249), .A2(n3013), .ZN(n8) );
  MOAI22D0BWP12T U151 ( .A1(n3012), .A2(n8), .B1(n3919), .B2(n3371), .ZN(n9)
         );
  OAI22D0BWP12T U152 ( .A1(n3786), .A2(n3015), .B1(n3784), .B2(n3014), .ZN(n10) );
  OAI22D0BWP12T U153 ( .A1(n3782), .A2(n3017), .B1(n3780), .B2(n3016), .ZN(n11) );
  OAI32D0BWP12T U154 ( .A1(n9), .A2(n10), .A3(n11), .B1(n3788), .B2(n9), .ZN(
        n12) );
  CKND2D0BWP12T U155 ( .A1(n3986), .A2(n12), .ZN(n3812) );
  OAI21D0BWP12T U156 ( .A1(n2318), .A2(n3379), .B(n2319), .ZN(n13) );
  CKND2D0BWP12T U157 ( .A1(n2380), .A2(n2382), .ZN(n14) );
  MOAI22D0BWP12T U158 ( .A1(n13), .A2(n14), .B1(n13), .B2(n14), .ZN(n4098) );
  OAI21D0BWP12T U159 ( .A1(n2656), .A2(n2657), .B(n2655), .ZN(n15) );
  CKND2D0BWP12T U160 ( .A1(n2659), .A2(n2679), .ZN(n16) );
  MOAI22D0BWP12T U161 ( .A1(n15), .A2(n16), .B1(n15), .B2(n16), .ZN(n3482) );
  CKND0BWP12T U162 ( .I(n3939), .ZN(n17) );
  OAI32D0BWP12T U163 ( .A1(n17), .A2(n4182), .A3(a[21]), .B1(n4181), .B2(n17), 
        .ZN(n18) );
  AOI22D0BWP12T U164 ( .A1(n3939), .A2(n2664), .B1(n4184), .B2(n17), .ZN(n19)
         );
  CKND0BWP12T U165 ( .I(n3864), .ZN(n20) );
  CKND0BWP12T U166 ( .I(n2205), .ZN(n21) );
  OAI32D0BWP12T U167 ( .A1(n3864), .A2(n4185), .A3(n19), .B1(n20), .B2(n21), 
        .ZN(n22) );
  MAOI22D0BWP12T U168 ( .A1(n3723), .A2(n3289), .B1(n3290), .B2(n4034), .ZN(
        n23) );
  AOI22D0BWP12T U169 ( .A1(n3617), .A2(n4203), .B1(n4163), .B2(n3671), .ZN(n24) );
  OA211D0BWP12T U170 ( .A1(n3796), .A2(n3773), .B(n23), .C(n24), .Z(n25) );
  IND4D0BWP12T U171 ( .A1(n18), .B1(n4193), .B2(n22), .B3(n25), .ZN(n3327) );
  CKND2D0BWP12T U172 ( .A1(n1712), .A2(n1709), .ZN(n26) );
  NR2D0BWP12T U173 ( .A1(n1708), .A2(n3140), .ZN(n27) );
  CKND0BWP12T U174 ( .I(n3519), .ZN(n28) );
  AOI32D0BWP12T U175 ( .A1(n3510), .A2(n27), .A3(n28), .B1(n3516), .B2(n27), 
        .ZN(n29) );
  OAI211D0BWP12T U176 ( .A1(n1708), .A2(n3143), .B(n3189), .C(n29), .ZN(n30)
         );
  MOAI22D0BWP12T U177 ( .A1(n26), .A2(n30), .B1(n26), .B2(n30), .ZN(n3526) );
  OAI22D0BWP12T U178 ( .A1(n2520), .A2(n2949), .B1(n2519), .B2(n2948), .ZN(n31) );
  IAO21D0BWP12T U179 ( .A1(n2525), .A2(n2955), .B(n31), .ZN(n32) );
  OA211D0BWP12T U180 ( .A1(n2524), .A2(n3356), .B(n3841), .C(n32), .Z(n561) );
  MAOI22D0BWP12T U181 ( .A1(n3921), .A2(n3713), .B1(n3921), .B2(n3712), .ZN(
        n33) );
  NR2D0BWP12T U182 ( .A1(n3702), .A2(n3701), .ZN(n34) );
  NR2D0BWP12T U183 ( .A1(n3704), .A2(n3783), .ZN(n35) );
  OAI22D0BWP12T U184 ( .A1(n3703), .A2(n3785), .B1(n3705), .B2(n3787), .ZN(n36) );
  AOI211D0BWP12T U185 ( .A1(n3707), .A2(n3706), .B(n35), .C(n36), .ZN(n37) );
  ND3D0BWP12T U186 ( .A1(n4175), .A2(n3709), .A3(n3708), .ZN(n38) );
  OAI211D0BWP12T U187 ( .A1(n3711), .A2(n37), .B(n3710), .C(n38), .ZN(n39) );
  OAI22D0BWP12T U188 ( .A1(n3767), .A2(n33), .B1(n34), .B2(n39), .ZN(n4162) );
  CKND2D0BWP12T U189 ( .A1(n3375), .A2(n3377), .ZN(n40) );
  CKND2D0BWP12T U190 ( .A1(n3378), .A2(n3377), .ZN(n41) );
  OAI211D0BWP12T U191 ( .A1(n3379), .A2(n40), .B(n3376), .C(n41), .ZN(n42) );
  CKND2D0BWP12T U192 ( .A1(n3389), .A2(n3390), .ZN(n43) );
  MOAI22D0BWP12T U193 ( .A1(n42), .A2(n43), .B1(n42), .B2(n43), .ZN(n4124) );
  NR4D0BWP12T U194 ( .A1(n3481), .A2(n3482), .A3(n3480), .A4(n3479), .ZN(n44)
         );
  NR4D0BWP12T U195 ( .A1(n3477), .A2(n3483), .A3(n3478), .A4(n3476), .ZN(n45)
         );
  IND3D0BWP12T U196 ( .A1(n3484), .B1(n44), .B2(n45), .ZN(n46) );
  NR4D0BWP12T U197 ( .A1(n3492), .A2(n3493), .A3(n4174), .A4(n46), .ZN(n47) );
  NR4D0BWP12T U198 ( .A1(n3475), .A2(n3474), .A3(n3473), .A4(n3472), .ZN(n48)
         );
  NR4D0BWP12T U199 ( .A1(n3471), .A2(n3470), .A3(n3469), .A4(n3468), .ZN(n49)
         );
  NR4D0BWP12T U200 ( .A1(n3467), .A2(n3466), .A3(n3465), .A4(n3464), .ZN(n50)
         );
  ND4D0BWP12T U201 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(n51) );
  OR4D0BWP12T U202 ( .A1(n3498), .A2(n4168), .A3(n3497), .A4(n51), .Z(n52) );
  OR4D0BWP12T U203 ( .A1(n3499), .A2(n3501), .A3(n3500), .A4(n52), .Z(n3502)
         );
  CKND2D0BWP12T U204 ( .A1(n3145), .A2(n3144), .ZN(n53) );
  NR2D0BWP12T U205 ( .A1(n3142), .A2(n3140), .ZN(n54) );
  CKND0BWP12T U206 ( .I(n3519), .ZN(n55) );
  AOI32D0BWP12T U207 ( .A1(n3510), .A2(n54), .A3(n55), .B1(n3516), .B2(n54), 
        .ZN(n56) );
  OAI211D0BWP12T U208 ( .A1(n3142), .A2(n3143), .B(n3141), .C(n56), .ZN(n57)
         );
  MOAI22D0BWP12T U209 ( .A1(n53), .A2(n57), .B1(n53), .B2(n57), .ZN(n3525) );
  INR3D0BWP12T U210 ( .A1(n3351), .B1(n4078), .B2(n2977), .ZN(n58) );
  MOAI22D0BWP12T U211 ( .A1(a[13]), .A2(n58), .B1(a[13]), .B2(n58), .ZN(n3633)
         );
  OAI21D0BWP12T U212 ( .A1(n3157), .A2(n3579), .B(n3158), .ZN(n59) );
  CKND2D0BWP12T U213 ( .A1(n3159), .A2(n3160), .ZN(n60) );
  MOAI22D0BWP12T U214 ( .A1(n59), .A2(n60), .B1(n59), .B2(n60), .ZN(n3568) );
  CKND0BWP12T U215 ( .I(n3694), .ZN(n61) );
  OAI222D0BWP12T U216 ( .A1(n3704), .A2(n3017), .B1(n3005), .B2(n3016), .C1(
        n3705), .C2(n3015), .ZN(n62) );
  NR2D0BWP12T U217 ( .A1(n3703), .A2(n3014), .ZN(n63) );
  OAI21D0BWP12T U218 ( .A1(n63), .A2(n62), .B(n4179), .ZN(n64) );
  OAI211D0BWP12T U219 ( .A1(n3007), .A2(n3006), .B(n3710), .C(n64), .ZN(n65)
         );
  AOI21D0BWP12T U220 ( .A1(n3170), .A2(n61), .B(n65), .ZN(n3715) );
  CKND0BWP12T U221 ( .I(n3379), .ZN(n66) );
  AOI21D0BWP12T U222 ( .A1(n3375), .A2(n66), .B(n3378), .ZN(n67) );
  CKND2D0BWP12T U223 ( .A1(n3376), .A2(n3377), .ZN(n68) );
  MAOI22D0BWP12T U224 ( .A1(n67), .A2(n68), .B1(n67), .B2(n68), .ZN(n4125) );
  INR2D0BWP12T U225 ( .A1(n2935), .B1(n3345), .ZN(n69) );
  OAI32D0BWP12T U226 ( .A1(n2936), .A2(n69), .A3(n2938), .B1(n2937), .B2(n2936), .ZN(n70) );
  CKND2D0BWP12T U227 ( .A1(n2940), .A2(n2932), .ZN(n71) );
  MAOI22D0BWP12T U228 ( .A1(n70), .A2(n71), .B1(n70), .B2(n71), .ZN(n3464) );
  CKND0BWP12T U229 ( .I(n4152), .ZN(n72) );
  CKND0BWP12T U230 ( .I(n4159), .ZN(n73) );
  CKND0BWP12T U231 ( .I(b[25]), .ZN(n74) );
  OAI32D0BWP12T U232 ( .A1(n74), .A2(n4182), .A3(n4157), .B1(n4181), .B2(n74), 
        .ZN(n75) );
  CKND0BWP12T U233 ( .I(n4154), .ZN(n76) );
  AOI22D0BWP12T U234 ( .A1(n4155), .A2(n4195), .B1(n4203), .B2(n4156), .ZN(n77) );
  AOI22D0BWP12T U235 ( .A1(b[25]), .A2(n2664), .B1(n4184), .B2(n74), .ZN(n78)
         );
  CKND0BWP12T U236 ( .I(n4160), .ZN(n79) );
  CKND0BWP12T U237 ( .I(n2205), .ZN(n80) );
  OAI32D0BWP12T U238 ( .A1(n4160), .A2(n4185), .A3(n78), .B1(n79), .B2(n80), 
        .ZN(n81) );
  OAI211D0BWP12T U239 ( .A1(n4161), .A2(n76), .B(n77), .C(n81), .ZN(n82) );
  AOI211D0BWP12T U240 ( .A1(n4158), .A2(n73), .B(n75), .C(n82), .ZN(n83) );
  AOI22D0BWP12T U241 ( .A1(n4162), .A2(n4163), .B1(n4206), .B2(n4153), .ZN(n84) );
  OAI211D0BWP12T U242 ( .A1(n4164), .A2(n72), .B(n83), .C(n84), .ZN(n4165) );
  AN4D0BWP12T U243 ( .A1(n3681), .A2(n3679), .A3(n3682), .A4(n3680), .Z(n85)
         );
  IND4D0BWP12T U244 ( .A1(n3683), .B1(n3684), .B2(n4014), .B3(n85), .ZN(n3999)
         );
  OA22D0BWP12T U245 ( .A1(n2955), .A2(n2950), .B1(n3356), .B2(n3712), .Z(n2495) );
  IIND4D0BWP12T U246 ( .A1(n2977), .A2(n2917), .B1(n3873), .B2(n3351), .ZN(n86) );
  MAOI22D0BWP12T U247 ( .A1(n4082), .A2(n86), .B1(n4082), .B2(n86), .ZN(n3631)
         );
  CKND0BWP12T U248 ( .I(n3579), .ZN(n87) );
  AN3D0BWP12T U249 ( .A1(n87), .A2(n3302), .A3(n3122), .Z(n88) );
  AOI211D0BWP12T U250 ( .A1(n3122), .A2(n3306), .B(n3121), .C(n88), .ZN(n89)
         );
  CKND2D0BWP12T U251 ( .A1(n3123), .A2(n3124), .ZN(n90) );
  MAOI22D0BWP12T U252 ( .A1(n89), .A2(n90), .B1(n89), .B2(n90), .ZN(n3570) );
  CKND2D0BWP12T U253 ( .A1(n622), .A2(n624), .ZN(n91) );
  AOI21D0BWP12T U254 ( .A1(n2535), .A2(n2498), .B(n2497), .ZN(n92) );
  OAI21D0BWP12T U255 ( .A1(n2499), .A2(n92), .B(n2500), .ZN(n93) );
  MOAI22D0BWP12T U256 ( .A1(n91), .A2(n93), .B1(n91), .B2(n93), .ZN(n4106) );
  CKND0BWP12T U257 ( .I(n3582), .ZN(n94) );
  AOI22D0BWP12T U258 ( .A1(n4210), .A2(n4100), .B1(n3567), .B2(n94), .ZN(n95)
         );
  MOAI22D0BWP12T U259 ( .A1(n3290), .A2(n4033), .B1(n3629), .B2(n4203), .ZN(
        n96) );
  OAI21D0BWP12T U260 ( .A1(a[19]), .A2(n4182), .B(n4181), .ZN(n97) );
  NR2D0BWP12T U261 ( .A1(n3166), .A2(n4185), .ZN(n98) );
  MUX2ND0BWP12T U262 ( .I0(n98), .I1(n2205), .S(n3866), .ZN(n99) );
  AOI211D0BWP12T U263 ( .A1(b[19]), .A2(n97), .B(n3216), .C(n99), .ZN(n100) );
  CKND2D0BWP12T U264 ( .A1(n3725), .A2(n3289), .ZN(n101) );
  OAI211D0BWP12T U265 ( .A1(n3798), .A2(n3773), .B(n100), .C(n101), .ZN(n102)
         );
  AOI211D0BWP12T U266 ( .A1(n3696), .A2(n4163), .B(n96), .C(n102), .ZN(n103)
         );
  CKND2D0BWP12T U267 ( .A1(n95), .A2(n103), .ZN(n3174) );
  CKND2D0BWP12T U268 ( .A1(n4067), .A2(n2632), .ZN(n104) );
  AOI31D0BWP12T U269 ( .A1(n2584), .A2(n2583), .A3(n104), .B(n3922), .ZN(n105)
         );
  OAI222D0BWP12T U270 ( .A1(n3356), .A2(n2585), .B1(n2812), .B2(n2949), .C1(
        n2951), .C2(n2948), .ZN(n106) );
  NR2D0BWP12T U271 ( .A1(n105), .A2(n106), .ZN(n3719) );
  IND2D0BWP12T U272 ( .A1(n3172), .B1(n3293), .ZN(n107) );
  MAOI22D0BWP12T U273 ( .A1(a[18]), .A2(n107), .B1(a[18]), .B2(n107), .ZN(
        n3610) );
  CKND0BWP12T U274 ( .I(n3160), .ZN(n108) );
  OA21D0BWP12T U275 ( .A1(n3158), .A2(n108), .B(n3159), .Z(n109) );
  OAI31D0BWP12T U276 ( .A1(n3579), .A2(n3157), .A3(n108), .B(n109), .ZN(n110)
         );
  CKND2D0BWP12T U277 ( .A1(n3162), .A2(n3154), .ZN(n111) );
  MOAI22D0BWP12T U278 ( .A1(n110), .A2(n111), .B1(n110), .B2(n111), .ZN(n3567)
         );
  MAOI22D0BWP12T U279 ( .A1(n4210), .A2(n4099), .B1(n4052), .B2(n3029), .ZN(
        n112) );
  OAI21D0BWP12T U280 ( .A1(n4069), .A2(n4182), .B(n4181), .ZN(n113) );
  MAOI22D0BWP12T U281 ( .A1(n3938), .A2(n113), .B1(n3799), .B2(n3773), .ZN(
        n114) );
  CKND0BWP12T U282 ( .I(n2205), .ZN(n115) );
  CKND0BWP12T U283 ( .I(n3865), .ZN(n116) );
  OAI32D0BWP12T U284 ( .A1(n3865), .A2(n4185), .A3(n1841), .B1(n115), .B2(n116), .ZN(n117) );
  OA211D0BWP12T U285 ( .A1(n3669), .A2(n4201), .B(n114), .C(n117), .Z(n118) );
  AOI22D0BWP12T U286 ( .A1(n3724), .A2(n3289), .B1(n3628), .B2(n4203), .ZN(
        n119) );
  AOI22D0BWP12T U287 ( .A1(n3475), .A2(n4173), .B1(n4206), .B2(n3572), .ZN(
        n120) );
  ND4D0BWP12T U288 ( .A1(n112), .A2(n118), .A3(n119), .A4(n120), .ZN(n1842) );
  CKND2D0BWP12T U289 ( .A1(n1856), .A2(n1857), .ZN(n121) );
  MAOI22D0BWP12T U290 ( .A1(b[0]), .A2(n121), .B1(b[0]), .B2(n121), .ZN(n3480)
         );
  CKND2D0BWP12T U291 ( .A1(n3096), .A2(n3097), .ZN(n122) );
  MOAI22D0BWP12T U292 ( .A1(n3098), .A2(n122), .B1(n3098), .B2(n122), .ZN(
        n3548) );
  CKND0BWP12T U293 ( .I(n3478), .ZN(n123) );
  OAI22D0BWP12T U294 ( .A1(n3479), .A2(n123), .B1(n2675), .B2(n3076), .ZN(n124) );
  AOI22D0BWP12T U295 ( .A1(n3929), .A2(n1027), .B1(n3587), .B2(n4206), .ZN(
        n125) );
  MUX2ND0BWP12T U296 ( .I0(n1029), .I1(n3366), .S(n3891), .ZN(n126) );
  OAI211D0BWP12T U297 ( .A1(n2480), .A2(n3064), .B(n125), .C(n126), .ZN(n127)
         );
  AO211D0BWP12T U298 ( .A1(n3540), .A2(n4215), .B(n124), .C(n127), .Z(n1053)
         );
  AOI22D0BWP12T U299 ( .A1(n3245), .A2(n2768), .B1(n3242), .B2(n2767), .ZN(
        n128) );
  IND2D0BWP12T U300 ( .A1(n2769), .B1(n3238), .ZN(n129) );
  OAI211D0BWP12T U301 ( .A1(a[29]), .A2(n2770), .B(n128), .C(n129), .ZN(n130)
         );
  CKND0BWP12T U302 ( .I(n3658), .ZN(n131) );
  AOI211D0BWP12T U303 ( .A1(n3788), .A2(n130), .B(n3655), .C(n131), .ZN(n132)
         );
  AOI22D0BWP12T U304 ( .A1(n2779), .A2(n2778), .B1(n3249), .B2(n3102), .ZN(
        n133) );
  OAI211D0BWP12T U305 ( .A1(n2780), .A2(n3754), .B(n132), .C(n133), .ZN(n3775)
         );
  CKND2D0BWP12T U306 ( .A1(n4187), .A2(n3293), .ZN(n134) );
  MAOI22D0BWP12T U307 ( .A1(a[17]), .A2(n134), .B1(a[17]), .B2(n134), .ZN(
        n3611) );
  OAI21D0BWP12T U308 ( .A1(n2401), .A2(n3388), .B(n2400), .ZN(n135) );
  CKND2D0BWP12T U309 ( .A1(n2959), .A2(n2961), .ZN(n136) );
  MOAI22D0BWP12T U310 ( .A1(n135), .A2(n136), .B1(n135), .B2(n136), .ZN(n3576)
         );
  OA222D0BWP12T U311 ( .A1(n2955), .A2(n633), .B1(n3356), .B2(n636), .C1(n3357), .C2(n2949), .Z(n137) );
  OA211D0BWP12T U312 ( .A1(n2301), .A2(n2948), .B(n3841), .C(n137), .Z(n3718)
         );
  CKND2D0BWP12T U313 ( .A1(n3485), .A2(n2902), .ZN(n138) );
  MOAI22D0BWP12T U314 ( .A1(n3276), .A2(n138), .B1(n3276), .B2(n138), .ZN(
        n3474) );
  CKND2D0BWP12T U315 ( .A1(n3507), .A2(n3495), .ZN(n139) );
  MAOI22D0BWP12T U316 ( .A1(n3508), .A2(n139), .B1(n3508), .B2(n139), .ZN(
        n4166) );
  CKND0BWP12T U317 ( .I(n3407), .ZN(n140) );
  AN3D0BWP12T U318 ( .A1(n141), .A2(n568), .A3(op[0]), .Z(n2667) );
  CKND0BWP12T U319 ( .I(op[3]), .ZN(n141) );
  NR4D0BWP12T U320 ( .A1(n3615), .A2(n3614), .A3(n3616), .A4(n3613), .ZN(n142)
         );
  NR4D0BWP12T U321 ( .A1(n3610), .A2(n3617), .A3(n3612), .A4(n3611), .ZN(n143)
         );
  ND3D0BWP12T U322 ( .A1(n320), .A2(n142), .A3(n143), .ZN(n3640) );
  NR2D0BWP12T U323 ( .A1(n3058), .A2(n3059), .ZN(n144) );
  CKND2D0BWP12T U324 ( .A1(n3060), .A2(n3056), .ZN(n145) );
  MAOI22D0BWP12T U325 ( .A1(n144), .A2(n145), .B1(n144), .B2(n145), .ZN(n3571)
         );
  INR3D0BWP12T U326 ( .A1(n3351), .B1(n4061), .B2(n3350), .ZN(n146) );
  MOAI22D0BWP12T U327 ( .A1(n4060), .A2(n146), .B1(n4060), .B2(n146), .ZN(
        n3627) );
  NR2D0BWP12T U328 ( .A1(n3841), .A2(n4158), .ZN(n147) );
  MAOI22D0BWP12T U329 ( .A1(n3702), .A2(n3701), .B1(n2837), .B2(n147), .ZN(
        n3743) );
  OAI21D0BWP12T U330 ( .A1(n1083), .A2(n3379), .B(n1082), .ZN(n148) );
  CKND2D0BWP12T U331 ( .A1(n1085), .A2(n1086), .ZN(n149) );
  MOAI22D0BWP12T U332 ( .A1(n148), .A2(n149), .B1(n148), .B2(n149), .ZN(n4126)
         );
  CKND0BWP12T U333 ( .I(n3566), .ZN(n150) );
  MUX2ND0BWP12T U334 ( .I0(n2915), .I1(n2205), .S(n3874), .ZN(n151) );
  AOI21D0BWP12T U335 ( .A1(n4195), .A2(n3760), .B(n151), .ZN(n152) );
  OAI21D0BWP12T U336 ( .A1(n4185), .A2(n2916), .B(n3949), .ZN(n153) );
  OAI211D0BWP12T U337 ( .A1(n3582), .A2(n150), .B(n152), .C(n153), .ZN(n154)
         );
  AOI22D0BWP12T U338 ( .A1(n4011), .A2(n4024), .B1(n4116), .B2(n4210), .ZN(
        n155) );
  CKND0BWP12T U339 ( .I(n3735), .ZN(n156) );
  OAI21D0BWP12T U340 ( .A1(n3988), .A2(n156), .B(n2921), .ZN(n157) );
  OAI211D0BWP12T U341 ( .A1(n4201), .A2(n3728), .B(n155), .C(n157), .ZN(n158)
         );
  AOI211D0BWP12T U342 ( .A1(n4203), .A2(n3631), .B(n154), .C(n158), .ZN(n2923)
         );
  CKND2D0BWP12T U343 ( .A1(n2999), .A2(n3000), .ZN(n159) );
  MOAI22D0BWP12T U344 ( .A1(n3001), .A2(n159), .B1(n3001), .B2(n159), .ZN(
        n3555) );
  CKND0BWP12T U345 ( .I(n3563), .ZN(n160) );
  CKND2D0BWP12T U346 ( .A1(n4173), .A2(n3504), .ZN(n161) );
  OAI211D0BWP12T U347 ( .A1(n3532), .A2(n160), .B(n2790), .C(n161), .ZN(n162)
         );
  AO21D1BWP12T U348 ( .A1(n3403), .A2(n4171), .B(n162), .Z(result[30]) );
  INR2D0BWP12T U349 ( .A1(n2935), .B1(n3345), .ZN(n163) );
  OAI32D0BWP12T U350 ( .A1(n2373), .A2(n163), .A3(n2938), .B1(n316), .B2(n2373), .ZN(n164) );
  CKND2D0BWP12T U351 ( .A1(n2379), .A2(n2376), .ZN(n165) );
  MAOI22D0BWP12T U352 ( .A1(n164), .A2(n165), .B1(n164), .B2(n165), .ZN(n3465)
         );
  AOI22D0BWP12T U353 ( .A1(n4206), .A2(n3580), .B1(n4106), .B2(n4210), .ZN(
        n166) );
  CKND0BWP12T U354 ( .I(n3479), .ZN(n167) );
  AOI22D0BWP12T U355 ( .A1(n4203), .A2(n3620), .B1(n3476), .B2(n167), .ZN(n168) );
  OAI211D0BWP12T U356 ( .A1(n3972), .A2(n2834), .B(n166), .C(n168), .ZN(n657)
         );
  OA222D0BWP12T U357 ( .A1(n3782), .A2(n1832), .B1(n1831), .B2(n3886), .C1(
        n1833), .C2(n3780), .Z(n3752) );
  IND2D0BWP12T U358 ( .A1(n3655), .B1(n3774), .ZN(n169) );
  NR2D0BWP12T U359 ( .A1(n3767), .A2(n3012), .ZN(n170) );
  AO222D0BWP12T U360 ( .A1(n169), .A2(n3765), .B1(n3013), .B2(n170), .C1(n3011), .C2(n3249), .Z(n3803) );
  INR3D0BWP12T U361 ( .A1(n3293), .B1(a[18]), .B2(n3172), .ZN(n171) );
  MOAI22D0BWP12T U362 ( .A1(n3173), .A2(n171), .B1(n3173), .B2(n171), .ZN(
        n3629) );
  CKND2D0BWP12T U363 ( .A1(n3386), .A2(n3390), .ZN(n172) );
  CKND2D0BWP12T U364 ( .A1(n3387), .A2(n3390), .ZN(n173) );
  OAI211D0BWP12T U365 ( .A1(n3388), .A2(n172), .B(n3389), .C(n173), .ZN(n174)
         );
  CKND2D0BWP12T U366 ( .A1(n929), .A2(n2382), .ZN(n175) );
  MOAI22D0BWP12T U367 ( .A1(n174), .A2(n175), .B1(n174), .B2(n175), .ZN(n3577)
         );
  AOI21D0BWP12T U368 ( .A1(n2535), .A2(n2498), .B(n2497), .ZN(n176) );
  CKND2D0BWP12T U369 ( .A1(n2500), .A2(n2493), .ZN(n177) );
  MAOI22D0BWP12T U370 ( .A1(n176), .A2(n177), .B1(n176), .B2(n177), .ZN(n4107)
         );
  AOI21D0BWP12T U371 ( .A1(n3276), .A2(n3147), .B(n3146), .ZN(n178) );
  CKND2D0BWP12T U372 ( .A1(n3149), .A2(n3145), .ZN(n179) );
  MAOI22D0BWP12T U373 ( .A1(n178), .A2(n179), .B1(n178), .B2(n179), .ZN(n3468)
         );
  INR2D0BWP12T U374 ( .A1(n2372), .B1(n3519), .ZN(n180) );
  OAI32D0BWP12T U375 ( .A1(n2373), .A2(n180), .A3(n2374), .B1(n316), .B2(n2373), .ZN(n181) );
  CKND2D0BWP12T U376 ( .A1(n2375), .A2(n2376), .ZN(n182) );
  MAOI22D0BWP12T U377 ( .A1(n181), .A2(n182), .B1(n181), .B2(n182), .ZN(n3527)
         );
  AN2D0BWP12T U378 ( .A1(n601), .A2(n570), .Z(n3910) );
  AO222D0BWP12T U379 ( .A1(n2586), .A2(n3242), .B1(n3238), .B2(n2824), .C1(
        n3241), .C2(n2823), .Z(n2478) );
  CKND2D0BWP12T U380 ( .A1(n3880), .A2(n3351), .ZN(n183) );
  MAOI22D0BWP12T U381 ( .A1(n4063), .A2(n183), .B1(n4063), .B2(n183), .ZN(
        n3624) );
  IOA21D0BWP12T U382 ( .A1(n3713), .A2(n2641), .B(n2495), .ZN(n3723) );
  OA21D0BWP12T U383 ( .A1(b[0]), .A2(n4066), .B(n2605), .Z(n3583) );
  CKND2D0BWP12T U384 ( .A1(n2926), .A2(n2927), .ZN(n184) );
  MAOI22D1BWP12T U385 ( .A1(n2928), .A2(n184), .B1(n2928), .B2(n184), .ZN(
        n3426) );
  AOI22D0BWP12T U386 ( .A1(n4206), .A2(n3568), .B1(n4210), .B2(n4101), .ZN(
        n185) );
  CKND0BWP12T U387 ( .I(n3951), .ZN(n186) );
  OAI32D0BWP12T U388 ( .A1(n186), .A2(a[18]), .A3(n4182), .B1(n4181), .B2(n186), .ZN(n187) );
  AOI211D0BWP12T U389 ( .A1(n3610), .A2(n4203), .B(n187), .C(n997), .ZN(n188)
         );
  OAI21D0BWP12T U390 ( .A1(n3803), .A2(n3773), .B(n188), .ZN(n189) );
  OAI22D0BWP12T U391 ( .A1(n3744), .A2(n4201), .B1(n4041), .B2(n3029), .ZN(
        n190) );
  AOI211D0BWP12T U392 ( .A1(n3992), .A2(n3019), .B(n189), .C(n190), .ZN(n191)
         );
  CKND2D0BWP12T U393 ( .A1(n4173), .A2(n3469), .ZN(n192) );
  ND3D0BWP12T U394 ( .A1(n185), .A2(n191), .A3(n192), .ZN(n998) );
  CKND2D0BWP12T U395 ( .A1(n3126), .A2(n3097), .ZN(n193) );
  MAOI22D0BWP12T U396 ( .A1(n3127), .A2(n193), .B1(n3127), .B2(n193), .ZN(
        n3473) );
  CKND0BWP12T U397 ( .I(n3519), .ZN(n194) );
  AOI21D0BWP12T U398 ( .A1(n2372), .A2(n194), .B(n2374), .ZN(n195) );
  CKND2D0BWP12T U399 ( .A1(n898), .A2(n316), .ZN(n196) );
  MAOI22D0BWP12T U400 ( .A1(n195), .A2(n196), .B1(n195), .B2(n196), .ZN(n3528)
         );
  IND3D0BWP12T U401 ( .A1(op[1]), .B1(op[0]), .B2(n197), .ZN(n4164) );
  CKND0BWP12T U402 ( .I(n563), .ZN(n197) );
  IAO21D0BWP12T U403 ( .A1(n2462), .A2(n3911), .B(n2304), .ZN(n961) );
  MOAI22D0BWP12T U404 ( .A1(n3922), .A2(n3165), .B1(n3922), .B2(n3756), .ZN(
        n3751) );
  IND2D0BWP12T U405 ( .A1(n3350), .B1(n3351), .ZN(n198) );
  MAOI22D0BWP12T U406 ( .A1(n4061), .A2(n198), .B1(n4061), .B2(n198), .ZN(
        n3622) );
  CKND2D0BWP12T U407 ( .A1(n1082), .A2(n1045), .ZN(n199) );
  MAOI22D0BWP12T U408 ( .A1(n3379), .A2(n199), .B1(n3379), .B2(n199), .ZN(
        n4112) );
  CKND2D0BWP12T U409 ( .A1(n2492), .A2(n2493), .ZN(n200) );
  IOA21D0BWP12T U410 ( .A1(n2490), .A2(n2439), .B(n2489), .ZN(n201) );
  MOAI22D0BWP12T U411 ( .A1(n200), .A2(n201), .B1(n200), .B2(n201), .ZN(n3581)
         );
  OAI21D0BWP12T U412 ( .A1(n2800), .A2(n3519), .B(n2799), .ZN(n202) );
  CKND2D0BWP12T U413 ( .A1(n2802), .A2(n3341), .ZN(n203) );
  MOAI22D0BWP12T U414 ( .A1(n202), .A2(n203), .B1(n202), .B2(n203), .ZN(n3530)
         );
  CKND2D0BWP12T U415 ( .A1(n1056), .A2(n2793), .ZN(n204) );
  MAOI22D0BWP12T U416 ( .A1(n2791), .A2(n204), .B1(n2791), .B2(n204), .ZN(
        n3418) );
  CKND0BWP12T U417 ( .I(n3407), .ZN(n205) );
  AOI22D0BWP12T U418 ( .A1(n3408), .A2(n205), .B1(n4206), .B2(n3583), .ZN(n206) );
  AOI22D0BWP12T U419 ( .A1(b[0]), .A2(n4185), .B1(n2018), .B2(n3366), .ZN(n207) );
  CKND0BWP12T U420 ( .I(b[0]), .ZN(n208) );
  AOI22D0BWP12T U421 ( .A1(b[0]), .A2(n2664), .B1(n4184), .B2(n208), .ZN(n209)
         );
  OAI31D0BWP12T U422 ( .A1(n4185), .A2(n4203), .A3(n209), .B(n4066), .ZN(n210)
         );
  OAI211D0BWP12T U423 ( .A1(n3674), .A2(n2592), .B(n207), .C(n210), .ZN(n211)
         );
  AOI222D0BWP12T U424 ( .A1(n3748), .A2(n1860), .B1(n4103), .B2(n4210), .C1(
        n3480), .C2(n4173), .ZN(n212) );
  OAI21D0BWP12T U425 ( .A1(n4018), .A2(n2423), .B(n4011), .ZN(n213) );
  OAI211D0BWP12T U426 ( .A1(n3974), .A2(n2834), .B(n212), .C(n213), .ZN(n214)
         );
  AOI211D0BWP12T U427 ( .A1(n4215), .A2(n3533), .B(n211), .C(n214), .ZN(n215)
         );
  OAI211D0BWP12T U428 ( .A1(n4182), .A2(n3887), .B(n206), .C(n215), .ZN(n216)
         );
  AO21D0BWP12T U429 ( .A1(n4163), .A2(n3677), .B(n216), .Z(result[0]) );
  NR3D0BWP12T U430 ( .A1(n4070), .A2(n3107), .A3(n3067), .ZN(n217) );
  MOAI22D0BWP12T U431 ( .A1(a[23]), .A2(n217), .B1(a[23]), .B2(n217), .ZN(
        n3623) );
  MOAI22D0BWP12T U432 ( .A1(n2547), .A2(n3687), .B1(n2547), .B2(n3167), .ZN(
        n3693) );
  AOI21D0BWP12T U433 ( .A1(n2490), .A2(n1010), .B(n1012), .ZN(n218) );
  CKND2D0BWP12T U434 ( .A1(n1013), .A2(n624), .ZN(n219) );
  MAOI22D0BWP12T U435 ( .A1(n218), .A2(n219), .B1(n218), .B2(n219), .ZN(n3580)
         );
  CKND2D0BWP12T U436 ( .A1(n2438), .A2(n2439), .ZN(n220) );
  IOA21D0BWP12T U437 ( .A1(n2535), .A2(n2534), .B(n2533), .ZN(n221) );
  MOAI22D0BWP12T U438 ( .A1(n220), .A2(n221), .B1(n220), .B2(n221), .ZN(n4109)
         );
  OAI21D0BWP12T U439 ( .A1(n3334), .A2(n3519), .B(n3333), .ZN(n222) );
  CKND2D0BWP12T U440 ( .A1(n3336), .A2(n3337), .ZN(n223) );
  MOAI22D0BWP12T U441 ( .A1(n222), .A2(n223), .B1(n222), .B2(n223), .ZN(n3529)
         );
  OAI21D0BWP12T U442 ( .A1(n1058), .A2(n3345), .B(n1057), .ZN(n224) );
  CKND2D0BWP12T U443 ( .A1(n1060), .A2(n1061), .ZN(n225) );
  MOAI22D0BWP12T U444 ( .A1(n224), .A2(n225), .B1(n224), .B2(n225), .ZN(n3493)
         );
  MOAI22D0BWP12T U445 ( .A1(a[19]), .A2(n3930), .B1(a[19]), .B2(n3930), .ZN(
        n226) );
  OAI22D0BWP12T U446 ( .A1(n2127), .A2(n2126), .B1(n2125), .B2(n226), .ZN(
        n2135) );
  OAI22D0BWP12T U447 ( .A1(n2470), .A2(n3898), .B1(n2471), .B2(n4160), .ZN(
        n227) );
  OAI22D0BWP12T U448 ( .A1(n2469), .A2(n3863), .B1(n2468), .B2(n3896), .ZN(
        n228) );
  NR2D0BWP12T U449 ( .A1(n227), .A2(n228), .ZN(n2519) );
  CKND0BWP12T U450 ( .I(n3886), .ZN(n229) );
  CKND0BWP12T U451 ( .I(n641), .ZN(n230) );
  AOI221D0BWP12T U452 ( .A1(n1005), .A2(n3886), .B1(n3911), .B2(n229), .C(n230), .ZN(n2523) );
  INR3D0BWP12T U453 ( .A1(n3293), .B1(n3107), .B2(n3291), .ZN(n231) );
  MOAI22D0BWP12T U454 ( .A1(n4070), .A2(n231), .B1(n4070), .B2(n231), .ZN(
        n3612) );
  INR3D0BWP12T U455 ( .A1(n3890), .B1(n1046), .B2(n2479), .ZN(n232) );
  MOAI22D0BWP12T U456 ( .A1(n4084), .A2(n232), .B1(n4084), .B2(n232), .ZN(
        n3630) );
  CKND2D0BWP12T U457 ( .A1(n2489), .A2(n2439), .ZN(n233) );
  MOAI22D0BWP12T U458 ( .A1(n2490), .A2(n233), .B1(n2490), .B2(n233), .ZN(
        n3588) );
  CKND2D0BWP12T U459 ( .A1(n2533), .A2(n2534), .ZN(n234) );
  MOAI22D0BWP12T U460 ( .A1(n2535), .A2(n234), .B1(n2535), .B2(n234), .ZN(
        n4108) );
  AOI222D0BWP12T U461 ( .A1(n4067), .A2(n2630), .B1(n3885), .B2(n2633), .C1(
        n581), .C2(n2632), .ZN(n235) );
  MAOI22D0BWP12T U462 ( .A1(n2579), .A2(n2418), .B1(n2414), .B2(n2948), .ZN(
        n236) );
  OAI21D0BWP12T U463 ( .A1(b[3]), .A2(n235), .B(n236), .ZN(n237) );
  AOI211D0BWP12T U464 ( .A1(n2641), .A2(n2413), .B(n3748), .C(n237), .ZN(n3674) );
  CKND2D0BWP12T U465 ( .A1(n2363), .A2(n2365), .ZN(n238) );
  MOAI22D0BWP12T U466 ( .A1(n2366), .A2(n238), .B1(n2366), .B2(n238), .ZN(
        n3425) );
  CKND2D0BWP12T U467 ( .A1(n2799), .A2(n1061), .ZN(n239) );
  MAOI22D0BWP12T U468 ( .A1(n3519), .A2(n239), .B1(n3519), .B2(n239), .ZN(
        n3541) );
  AOI21D0BWP12T U469 ( .A1(n2539), .A2(n2508), .B(n2507), .ZN(n240) );
  CKND2D0BWP12T U470 ( .A1(n2510), .A2(n2511), .ZN(n241) );
  MAOI22D0BWP12T U471 ( .A1(n240), .A2(n241), .B1(n240), .B2(n241), .ZN(n3477)
         );
  OAI211D0BWP12T U472 ( .A1(n3479), .A2(n3382), .B(n3381), .C(n3380), .ZN(n242) );
  AOI22D0BWP12T U473 ( .A1(n3973), .A2(n3982), .B1(n4206), .B2(n3591), .ZN(
        n243) );
  AOI22D0BWP12T U474 ( .A1(n4058), .A2(n4011), .B1(n3529), .B2(n4215), .ZN(
        n244) );
  CKND2D0BWP12T U475 ( .A1(n243), .A2(n244), .ZN(n245) );
  AO211D1BWP12T U476 ( .A1(n4171), .A2(n3423), .B(n242), .C(n245), .Z(
        result[10]) );
  MAOI22D0BWP12T U477 ( .A1(n1189), .A2(n3897), .B1(n1189), .B2(n3897), .ZN(
        n1906) );
  MAOI22D0BWP12T U478 ( .A1(n3820), .A2(n2463), .B1(n2468), .B2(n3865), .ZN(
        n246) );
  CKND2D0BWP12T U479 ( .A1(n2462), .A2(a[17]), .ZN(n247) );
  OAI211D0BWP12T U480 ( .A1(n2471), .A2(n3866), .B(n246), .C(n247), .ZN(n2577)
         );
  AN2D0BWP12T U481 ( .A1(n2634), .A2(n2633), .Z(n2635) );
  MAOI222D0BWP12T U482 ( .A(n1448), .B(n248), .C(n249), .ZN(n1452) );
  CKND0BWP12T U483 ( .I(n1446), .ZN(n248) );
  CKND0BWP12T U484 ( .I(n1447), .ZN(n249) );
  IOA21D0BWP12T U485 ( .A1(n965), .A2(n2641), .B(n978), .ZN(n979) );
  CKND0BWP12T U486 ( .I(n3065), .ZN(n250) );
  OAI21D0BWP12T U487 ( .A1(n3921), .A2(n3030), .B(n250), .ZN(n251) );
  AO21D0BWP12T U488 ( .A1(n2427), .A2(n251), .B(n4046), .Z(n4052) );
  NR2D0BWP12T U489 ( .A1(n4064), .A2(n2245), .ZN(n252) );
  CKND2D0BWP12T U490 ( .A1(n3293), .A2(n252), .ZN(n253) );
  CKND0BWP12T U491 ( .I(n3618), .ZN(n254) );
  NR2D0BWP12T U492 ( .A1(n253), .A2(n254), .ZN(n3009) );
  MAOI22D0BWP12T U493 ( .A1(n253), .A2(n254), .B1(n253), .B2(n254), .ZN(n4156)
         );
  CKND0BWP12T U494 ( .I(n3353), .ZN(n255) );
  CKND0BWP12T U495 ( .I(n2525), .ZN(n256) );
  AOI21D0BWP12T U496 ( .A1(n2579), .A2(n256), .B(n3919), .ZN(n257) );
  OAI21D0BWP12T U497 ( .A1(n2526), .A2(n255), .B(n257), .ZN(n258) );
  AOI21D0BWP12T U498 ( .A1(b[3]), .A2(n2919), .B(n258), .ZN(n3726) );
  OAI21D0BWP12T U499 ( .A1(n2660), .A2(n2663), .B(n2661), .ZN(n259) );
  CKND2D0BWP12T U500 ( .A1(n2532), .A2(n2534), .ZN(n260) );
  MAOI22D0BWP12T U501 ( .A1(n259), .A2(n260), .B1(n259), .B2(n260), .ZN(n322)
         );
  OR4XD1BWP12T U502 ( .A1(n3938), .A2(b[19]), .A3(n3939), .A4(n3951), .Z(n542)
         );
  CKND2D0BWP12T U503 ( .A1(n1859), .A2(n1857), .ZN(n261) );
  MOAI22D0BWP12T U504 ( .A1(b[0]), .A2(n261), .B1(b[0]), .B2(n261), .ZN(n4103)
         );
  CKND2D0BWP12T U505 ( .A1(n3330), .A2(n3331), .ZN(n262) );
  MOAI22D0BWP12T U506 ( .A1(n3332), .A2(n262), .B1(n3332), .B2(n262), .ZN(
        n3423) );
  CKND0BWP12T U507 ( .I(n3345), .ZN(n263) );
  AOI21D0BWP12T U508 ( .A1(n3338), .A2(n263), .B(n3342), .ZN(n264) );
  CKND2D0BWP12T U509 ( .A1(n3339), .A2(n3341), .ZN(n265) );
  MAOI22D0BWP12T U510 ( .A1(n264), .A2(n265), .B1(n264), .B2(n265), .ZN(n3492)
         );
  IOA21D0BWP12T U511 ( .A1(n4210), .A2(n4126), .B(n1087), .ZN(n266) );
  AO21D0BWP12T U512 ( .A1(n4203), .A2(n3634), .B(n266), .Z(n1106) );
  AOI21D0BWP12T U513 ( .A1(n2504), .A2(n1030), .B(n1032), .ZN(n267) );
  CKND2D0BWP12T U514 ( .A1(n1033), .A2(n610), .ZN(n268) );
  MAOI22D0BWP12T U515 ( .A1(n267), .A2(n268), .B1(n267), .B2(n268), .ZN(n3536)
         );
  CKND0BWP12T U516 ( .I(n3528), .ZN(n269) );
  OAI211D0BWP12T U517 ( .A1(n3532), .A2(n269), .B(n603), .C(n602), .ZN(n270)
         );
  AO21D1BWP12T U518 ( .A1(n4171), .A2(n3425), .B(n270), .Z(result[11]) );
  AOI22D0BWP12T U519 ( .A1(n4173), .A2(n3477), .B1(n3537), .B2(n4215), .ZN(
        n271) );
  ND4D1BWP12T U520 ( .A1(n2512), .A2(n2513), .A3(n271), .A4(n2514), .ZN(n272)
         );
  AO21D1BWP12T U521 ( .A1(n3412), .A2(n4171), .B(n272), .Z(result[5]) );
  OA21D0BWP12T U522 ( .A1(n2471), .A2(n3911), .B(n2621), .Z(n3682) );
  AOI22D0BWP12T U523 ( .A1(n4081), .A2(n2632), .B1(n3885), .B2(n2582), .ZN(
        n273) );
  AOI21D0BWP12T U524 ( .A1(n2527), .A2(n273), .B(b[3]), .ZN(n274) );
  OAI22D0BWP12T U525 ( .A1(n2524), .A2(n2948), .B1(n2525), .B2(n2949), .ZN(
        n275) );
  OAI21D0BWP12T U526 ( .A1(n3356), .A2(n2526), .B(n3841), .ZN(n276) );
  NR3D0BWP12T U527 ( .A1(n274), .A2(n275), .A3(n276), .ZN(n2573) );
  OAI21D0BWP12T U528 ( .A1(n2683), .A2(n2684), .B(n2682), .ZN(n277) );
  CKND2D0BWP12T U529 ( .A1(n2686), .A2(n2662), .ZN(n278) );
  MOAI22D0BWP12T U530 ( .A1(n277), .A2(n278), .B1(n277), .B2(n278), .ZN(n4105)
         );
  OR4XD1BWP12T U531 ( .A1(n4191), .A2(n3949), .A3(n3952), .A4(n3930), .Z(n547)
         );
  CKND2D0BWP12T U532 ( .A1(n3261), .A2(n3262), .ZN(n279) );
  MOAI22D0BWP12T U533 ( .A1(n3263), .A2(n279), .B1(n3263), .B2(n279), .ZN(
        n3444) );
  NR2D0BWP12T U534 ( .A1(n3399), .A2(n3660), .ZN(n280) );
  AOI211D0BWP12T U535 ( .A1(n3399), .A2(n3660), .B(n3613), .C(n280), .ZN(n2176) );
  CKND2D0BWP12T U536 ( .A1(n3053), .A2(n3054), .ZN(n281) );
  MOAI22D0BWP12T U537 ( .A1(n3055), .A2(n281), .B1(n3055), .B2(n281), .ZN(
        n3498) );
  CKND2D0BWP12T U538 ( .A1(n2391), .A2(n3351), .ZN(n282) );
  MAOI22D0BWP12T U539 ( .A1(n4078), .A2(n282), .B1(n4078), .B2(n282), .ZN(
        n3626) );
  OAI21D0BWP12T U540 ( .A1(n2817), .A2(n3388), .B(n2816), .ZN(n283) );
  CKND2D0BWP12T U541 ( .A1(n2819), .A2(n3377), .ZN(n284) );
  MOAI22D0BWP12T U542 ( .A1(n283), .A2(n284), .B1(n283), .B2(n284), .ZN(n3592)
         );
  CKND2D0BWP12T U543 ( .A1(n2506), .A2(n2511), .ZN(n285) );
  IOA21D0BWP12T U544 ( .A1(n2504), .A2(n2503), .B(n2502), .ZN(n286) );
  MOAI22D0BWP12T U545 ( .A1(n285), .A2(n286), .B1(n285), .B2(n286), .ZN(n3537)
         );
  IND2D0BWP12T U546 ( .A1(n2410), .B1(n2411), .ZN(n287) );
  MAOI22D0BWP12T U547 ( .A1(n2412), .A2(n287), .B1(n2412), .B2(n287), .ZN(
        n3414) );
  CKND0BWP12T U548 ( .I(n3853), .ZN(n288) );
  OAI222D1BWP12T U549 ( .A1(n288), .A2(n1065), .B1(n2468), .B2(a[29]), .C1(
        n4065), .C2(n2471), .ZN(n965) );
  MOAI22D0BWP12T U550 ( .A1(n4089), .A2(n3921), .B1(n4089), .B2(n3921), .ZN(
        n289) );
  OAI22D0BWP12T U551 ( .A1(n2103), .A2(n2104), .B1(n2102), .B2(n289), .ZN(
        n2105) );
  OAI21D0BWP12T U552 ( .A1(n1328), .A2(n1329), .B(n1326), .ZN(n1327) );
  CKND0BWP12T U553 ( .I(n4068), .ZN(n290) );
  MAOI22D0BWP12T U554 ( .A1(n2632), .A2(n290), .B1(n4081), .B2(n2631), .ZN(
        n2637) );
  MOAI22D0BWP12T U555 ( .A1(a[21]), .A2(n1979), .B1(a[21]), .B2(n1979), .ZN(
        n291) );
  OAI22D1BWP12T U556 ( .A1(n2079), .A2(n291), .B1(n2077), .B2(n1155), .ZN(
        n1286) );
  AN2XD2BWP12T U557 ( .A1(n1450), .A2(n1451), .Z(n3136) );
  INR2D0BWP12T U558 ( .A1(n2241), .B1(n2238), .ZN(n1742) );
  IOA21D0BWP12T U559 ( .A1(n2461), .A2(n3922), .B(n2495), .ZN(n3288) );
  OA21D0BWP12T U560 ( .A1(n2598), .A2(n2597), .B(n2599), .Z(n3406) );
  IOA21D0BWP12T U561 ( .A1(a[23]), .A2(n3943), .B(n3056), .ZN(n292) );
  MOAI22D0BWP12T U562 ( .A1(n3057), .A2(n292), .B1(n3057), .B2(n292), .ZN(
        n4134) );
  MOAI22D0BWP12T U563 ( .A1(n2547), .A2(n3004), .B1(n2547), .B2(n3003), .ZN(
        n3694) );
  NR2D0BWP12T U564 ( .A1(n1046), .A2(n2479), .ZN(n293) );
  MOAI22D0BWP12T U565 ( .A1(n4083), .A2(n293), .B1(n4083), .B2(n293), .ZN(
        n3620) );
  CKND2D0BWP12T U566 ( .A1(n2661), .A2(n2662), .ZN(n294) );
  MAOI22D0BWP12T U567 ( .A1(n2663), .A2(n294), .B1(n2663), .B2(n294), .ZN(
        n3585) );
  IAO21D0BWP12T U568 ( .A1(n3919), .A2(n512), .B(n2491), .ZN(n1010) );
  AO22D0BWP12T U569 ( .A1(n4113), .A2(n4210), .B1(n4206), .B2(n3573), .Z(n3326) );
  INR2D0BWP12T U570 ( .A1(n2941), .B1(n3379), .ZN(n295) );
  OAI32D0BWP12T U571 ( .A1(n2942), .A2(n295), .A3(n2944), .B1(n2943), .B2(
        n2942), .ZN(n296) );
  CKND2D0BWP12T U572 ( .A1(n2946), .A2(n2967), .ZN(n297) );
  MAOI22D0BWP12T U573 ( .A1(n296), .A2(n297), .B1(n296), .B2(n297), .ZN(n4096)
         );
  CKND2D0BWP12T U574 ( .A1(n2446), .A2(n2503), .ZN(n298) );
  IOA21D0BWP12T U575 ( .A1(n2539), .A2(n2537), .B(n2536), .ZN(n299) );
  MOAI22D0BWP12T U576 ( .A1(n298), .A2(n299), .B1(n298), .B2(n299), .ZN(n3483)
         );
  IND2D1BWP12T U577 ( .A1(n4084), .B1(n3880), .ZN(n347) );
  IND2XD2BWP12T U578 ( .A1(b[0]), .B1(n3916), .ZN(n2471) );
  NR2D0BWP12T U579 ( .A1(n2245), .A2(n3619), .ZN(n300) );
  MOAI22D0BWP12T U580 ( .A1(n4064), .A2(n300), .B1(n4064), .B2(n300), .ZN(
        n3641) );
  OAI21D0BWP12T U581 ( .A1(n1532), .A2(n1531), .B(n1530), .ZN(n1534) );
  MOAI22D0BWP12T U582 ( .A1(a[29]), .A2(n2098), .B1(a[29]), .B2(n2098), .ZN(
        n301) );
  OAI22D0BWP12T U583 ( .A1(n2100), .A2(n2101), .B1(n2099), .B2(n301), .ZN(
        n2106) );
  OAI21D0BWP12T U584 ( .A1(n1478), .A2(n1479), .B(n1477), .ZN(n1481) );
  OAI21D0BWP12T U585 ( .A1(n1211), .A2(n1212), .B(n1210), .ZN(n1214) );
  IOA21D0BWP12T U586 ( .A1(n3323), .A2(n3315), .B(n3322), .ZN(n1731) );
  OA21D0BWP12T U587 ( .A1(b[0]), .A2(n581), .B(n3887), .Z(n2586) );
  AOI222D0BWP12T U588 ( .A1(n3229), .A2(n3230), .B1(n3228), .B2(n3227), .C1(
        n3231), .C2(n2821), .ZN(n302) );
  IOA21D0BWP12T U589 ( .A1(n3707), .A2(n3226), .B(n302), .ZN(n3062) );
  CKND2D0BWP12T U590 ( .A1(n2542), .A2(n2672), .ZN(n303) );
  MAOI22D0BWP12T U591 ( .A1(n4068), .A2(n303), .B1(n4068), .B2(n303), .ZN(
        n3615) );
  OAI21D0BWP12T U592 ( .A1(n1241), .A2(n1240), .B(n1239), .ZN(n1135) );
  IND2D0BWP12T U593 ( .A1(n1783), .B1(n3134), .ZN(n1785) );
  OA32D0BWP12T U594 ( .A1(n2973), .A2(n2955), .A3(n3682), .B1(n3919), .B2(
        n2973), .Z(n3966) );
  IND2D0BWP12T U595 ( .A1(n2889), .B1(n2890), .ZN(n2892) );
  IND2D0BWP12T U596 ( .A1(n651), .B1(n3986), .ZN(n3372) );
  IOA21D0BWP12T U597 ( .A1(n2582), .A2(n3027), .B(n3066), .ZN(n1047) );
  NR2D0BWP12T U598 ( .A1(n4081), .A2(n2479), .ZN(n304) );
  MOAI22D0BWP12T U599 ( .A1(n4075), .A2(n304), .B1(n4075), .B2(n304), .ZN(
        n3621) );
  CKND2D0BWP12T U600 ( .A1(n2646), .A2(n2647), .ZN(n305) );
  MOAI22D0BWP12T U601 ( .A1(n2648), .A2(n305), .B1(n2648), .B2(n305), .ZN(
        n3411) );
  IND2D0BWP12T U602 ( .A1(n4081), .B1(n2634), .ZN(n1046) );
  CKND2D0BWP12T U603 ( .A1(n3494), .A2(n3495), .ZN(n306) );
  MOAI22D0BWP12T U604 ( .A1(n3496), .A2(n306), .B1(n3496), .B2(n306), .ZN(
        n4168) );
  CKND0BWP12T U605 ( .I(n3388), .ZN(n307) );
  AOI21D0BWP12T U606 ( .A1(n3386), .A2(n307), .B(n3387), .ZN(n308) );
  CKND2D0BWP12T U607 ( .A1(n3389), .A2(n3390), .ZN(n309) );
  MAOI22D0BWP12T U608 ( .A1(n308), .A2(n309), .B1(n308), .B2(n309), .ZN(n3591)
         );
  CKND2D0BWP12T U609 ( .A1(n2502), .A2(n2503), .ZN(n310) );
  MOAI22D0BWP12T U610 ( .A1(n2504), .A2(n310), .B1(n2504), .B2(n310), .ZN(
        n3542) );
  MAOI222D0BWP12T U611 ( .A(n446), .B(n447), .C(n445), .ZN(n311) );
  CKND0BWP12T U612 ( .I(n311), .ZN(n465) );
  IND4D0BWP12T U613 ( .A1(n3107), .B1(n3863), .B2(n3862), .B3(n3106), .ZN(
        n2245) );
  CKND0BWP12T U614 ( .I(n3396), .ZN(n312) );
  AOI222D0BWP12T U615 ( .A1(n312), .A2(n4206), .B1(n4210), .B2(n3398), .C1(
        n3399), .C2(n4203), .ZN(n3400) );
  IND2D0BWP12T U616 ( .A1(n4063), .B1(n3880), .ZN(n3350) );
  NR2D0BWP12T U617 ( .A1(n1740), .A2(n1817), .ZN(n3058) );
  IAO21D0BWP12T U618 ( .A1(n3841), .A2(n4089), .B(n3655), .ZN(n4036) );
  CKND2D0BWP12T U619 ( .A1(n2241), .A2(n2242), .ZN(n313) );
  MAOI22D0BWP12T U620 ( .A1(n2233), .A2(n313), .B1(n2233), .B2(n313), .ZN(
        n4133) );
  OAI22D0BWP12T U621 ( .A1(n3886), .A2(n983), .B1(n3782), .B2(n1833), .ZN(n314) );
  OAI22D0BWP12T U622 ( .A1(n3780), .A2(n1838), .B1(n3786), .B2(n966), .ZN(n315) );
  NR2D0BWP12T U623 ( .A1(n314), .A2(n315), .ZN(n3754) );
  FA1D2BWP12T U624 ( .A(a[29]), .B(n2169), .CI(n2166), .CO(n2789), .S(n3503)
         );
  FA1D2BWP12T U625 ( .A(n3395), .B(b[31]), .CI(n2179), .CO(n2170), .S(n3562)
         );
  RCAOI21D1BWP12T U626 ( .A1(n1724), .A2(n1723), .B(n1722), .ZN(n3267) );
  TPND2D3BWP12T U627 ( .A1(n2021), .A2(n1185), .ZN(n2023) );
  TPAOI21D2BWP12T U628 ( .A1(n1455), .A2(n3134), .B(n1454), .ZN(n3043) );
  CKND2D2BWP12T U629 ( .A1(n1498), .A2(n1497), .ZN(n3261) );
  TPND2D2BWP12T U630 ( .A1(n1500), .A2(n1499), .ZN(n3092) );
  BUFFD2BWP12T U631 ( .I(b[3]), .Z(n1189) );
  TPND2D3BWP12T U632 ( .A1(n3451), .A2(n4171), .ZN(n2222) );
  HA1D0BWP12T U633 ( .A(n3899), .B(n2752), .CO(n2165), .S(n3662) );
  FA1D2BWP12T U634 ( .A(n3848), .B(a[30]), .CI(n2789), .CO(n2217), .S(n3504)
         );
  OAI22D1BWP12T U635 ( .A1(n2469), .A2(n3899), .B1(n2470), .B2(n3911), .ZN(
        n2304) );
  INVD3BWP12T U636 ( .I(a[9]), .ZN(n3879) );
  TPAOI21D2BWP12T U637 ( .A1(n2792), .A2(n2796), .B(n469), .ZN(n470) );
  INVD9BWP12T U638 ( .I(n3891), .ZN(n4084) );
  FA1D2BWP12T U639 ( .A(n1319), .B(n1318), .CI(n1317), .CO(n1461), .S(n1440)
         );
  OAI22D1BWP12T U640 ( .A1(n2127), .A2(n1313), .B1(n2125), .B2(n1236), .ZN(
        n1319) );
  INR2D2BWP12T U641 ( .A1(n2469), .B1(n2454), .ZN(n527) );
  TPOAI21D1BWP12T U642 ( .A1(n3267), .A2(n3264), .B(n3265), .ZN(n3098) );
  ND2D4BWP12T U643 ( .A1(n2222), .A2(n2221), .ZN(result[31]) );
  XNR2D1BWP12T U644 ( .A1(n2064), .A2(n1190), .ZN(n1341) );
  ND2XD8BWP12T U645 ( .A1(n754), .A2(n753), .ZN(n2130) );
  TPAOI21D2BWP12T U646 ( .A1(n3044), .A2(n321), .B(n1503), .ZN(n1504) );
  TPND2D2BWP12T U647 ( .A1(n2362), .A2(n2361), .ZN(result[14]) );
  CKND0BWP12T U648 ( .I(n2791), .ZN(n2794) );
  TPOAI21D1BWP12T U649 ( .A1(n2791), .A2(n471), .B(n470), .ZN(n3332) );
  XNR2XD2BWP12T U650 ( .A1(n1004), .A2(n1003), .ZN(n3415) );
  TPAOI21D2BWP12T U651 ( .A1(n1004), .A2(n1002), .B(n430), .ZN(n2791) );
  FA1D2BWP12T U652 ( .A(n397), .B(n396), .CI(n395), .CO(n398), .S(n390) );
  INVD3BWP12T U653 ( .I(n3897), .ZN(n4077) );
  INVD3BWP12T U654 ( .I(a[14]), .ZN(n3873) );
  TPND2D2BWP12T U655 ( .A1(n1931), .A2(n1930), .ZN(n2163) );
  TPOAI22D2BWP12T U656 ( .A1(n2068), .A2(n1191), .B1(n1341), .B2(n2065), .ZN(
        n1356) );
  INVD3BWP12T U657 ( .I(n3300), .ZN(n2547) );
  INVD1BWP12T U658 ( .I(a[21]), .ZN(n3864) );
  NR2D0BWP12T U659 ( .A1(n3833), .A2(n4060), .ZN(n912) );
  BUFFD2BWP12T U660 ( .I(a[0]), .Z(n4066) );
  INVD3BWP12T U661 ( .I(n4066), .ZN(n2018) );
  INVD4BWP12T U662 ( .I(n4160), .ZN(n4157) );
  CKBD1BWP12T U663 ( .I(n500), .Z(n499) );
  AO21D2BWP12T U664 ( .A1(n4170), .A2(n4171), .B(n4169), .Z(result[25]) );
  INVD1BWP12T U665 ( .I(n3407), .ZN(n4171) );
  ND2D1BWP12T U666 ( .A1(n523), .A2(n483), .ZN(n3407) );
  INVD1BWP12T U667 ( .I(a[30]), .ZN(n3899) );
  OR2XD1BWP12T U668 ( .A1(n3833), .A2(n4060), .Z(n316) );
  OR2XD1BWP12T U669 ( .A1(n895), .A2(n894), .Z(n317) );
  INVD1BWP12T U670 ( .I(n3454), .ZN(n2993) );
  INVD1BWP12T U671 ( .I(a[17]), .ZN(n3868) );
  OR2XD1BWP12T U672 ( .A1(n3817), .A2(n4069), .Z(n1801) );
  OR2XD1BWP12T U673 ( .A1(n3827), .A2(a[14]), .Z(n2291) );
  OR2XD1BWP12T U674 ( .A1(n3829), .A2(n4078), .Z(n2376) );
  OR2XD1BWP12T U675 ( .A1(n399), .A2(n398), .Z(n318) );
  INVD2BWP12T U676 ( .I(a[27]), .ZN(n3897) );
  OR2XD1BWP12T U677 ( .A1(n1714), .A2(n1713), .Z(n3145) );
  OR2XD1BWP12T U678 ( .A1(n3830), .A2(n905), .Z(n2932) );
  OR2XD1BWP12T U679 ( .A1(n1508), .A2(n1507), .Z(n319) );
  XNR2D1BWP12T U680 ( .A1(n2479), .A2(n4081), .ZN(n320) );
  INVD4BWP12T U681 ( .I(a[13]), .ZN(n989) );
  OR2XD1BWP12T U682 ( .A1(n3819), .A2(n3820), .Z(n1712) );
  OR2D2BWP12T U683 ( .A1(n1502), .A2(n1501), .Z(n321) );
  NR2D1BWP12T U684 ( .A1(n4075), .A2(n3920), .ZN(n2499) );
  INVD1BWP12T U685 ( .I(a[19]), .ZN(n1312) );
  INVD8BWP12T U686 ( .I(n3892), .ZN(n4075) );
  CKBD1BWP12T U687 ( .I(a[19]), .Z(n3173) );
  INVD1BWP12T U688 ( .I(n4066), .ZN(n324) );
  INVD3BWP12T U689 ( .I(a[1]), .ZN(n323) );
  INVD9BWP12T U690 ( .I(n323), .ZN(n1977) );
  TPND2D2BWP12T U691 ( .A1(n324), .A2(n1977), .ZN(n340) );
  BUFFD8BWP12T U692 ( .I(n340), .Z(n2019) );
  INVD1BWP12T U693 ( .I(b[8]), .ZN(n3832) );
  XNR2D1BWP12T U694 ( .A1(n1977), .A2(n3928), .ZN(n330) );
  INVD1BWP12T U695 ( .I(b[9]), .ZN(n3838) );
  INVD4BWP12T U696 ( .I(n3838), .ZN(n3957) );
  XNR2XD2BWP12T U697 ( .A1(n1977), .A2(n3957), .ZN(n341) );
  OAI22D1BWP12T U698 ( .A1(n2019), .A2(n330), .B1(n341), .B2(n2018), .ZN(n344)
         );
  INVD3BWP12T U699 ( .I(a[5]), .ZN(n3892) );
  INVD2BWP12T U700 ( .I(a[4]), .ZN(n3893) );
  CKND8BWP12T U701 ( .I(n3893), .ZN(n4081) );
  INVD3BWP12T U702 ( .I(n4081), .ZN(n325) );
  XNR2XD4BWP12T U703 ( .A1(n4075), .A2(n325), .ZN(n327) );
  BUFFXD8BWP12T U704 ( .I(a[3]), .Z(n4068) );
  BUFFXD6BWP12T U705 ( .I(a[3]), .Z(n331) );
  ND2D8BWP12T U706 ( .A1(n4081), .A2(n331), .ZN(n326) );
  TPOAI21D8BWP12T U707 ( .A1(n4068), .A2(n4081), .B(n326), .ZN(n2080) );
  ND2XD8BWP12T U708 ( .A1(n327), .A2(n2080), .ZN(n2083) );
  BUFFD2BWP12T U709 ( .I(b[4]), .Z(n328) );
  INVD6BWP12T U710 ( .I(n328), .ZN(n338) );
  XNR2D1BWP12T U711 ( .A1(n4075), .A2(n718), .ZN(n441) );
  INVD3BWP12T U712 ( .I(n3842), .ZN(n3920) );
  XNR2D1BWP12T U713 ( .A1(n4075), .A2(n3920), .ZN(n337) );
  TPOAI22D1BWP12T U714 ( .A1(n2083), .A2(n441), .B1(n337), .B2(n2080), .ZN(
        n343) );
  XNR2XD8BWP12T U715 ( .A1(n4075), .A2(n4083), .ZN(n2011) );
  INVD4BWP12T U716 ( .I(a[7]), .ZN(n3891) );
  XOR2D2BWP12T U717 ( .A1(n4084), .A2(n4083), .Z(n329) );
  ND2XD8BWP12T U718 ( .A1(n2011), .A2(n329), .ZN(n2013) );
  INVD4BWP12T U719 ( .I(b[2]), .ZN(n3886) );
  INVD15BWP12T U720 ( .I(n3886), .ZN(n3921) );
  XNR2XD1BWP12T U721 ( .A1(n3921), .A2(n4084), .ZN(n439) );
  XNR2D1BWP12T U722 ( .A1(b[3]), .A2(n4084), .ZN(n339) );
  OAI22D1BWP12T U723 ( .A1(n2013), .A2(n439), .B1(n2011), .B2(n339), .ZN(n459)
         );
  INVD1BWP12T U724 ( .I(b[7]), .ZN(n3840) );
  XNR2D1BWP12T U725 ( .A1(n3929), .A2(n1977), .ZN(n411) );
  OAI22D1BWP12T U726 ( .A1(n2019), .A2(n411), .B1(n330), .B2(n2018), .ZN(n438)
         );
  BUFFXD8BWP12T U727 ( .I(b[0]), .Z(n1979) );
  ND2D1BWP12T U728 ( .A1(n4062), .A2(n4084), .ZN(n348) );
  INVD3BWP12T U729 ( .I(n4062), .ZN(n3880) );
  INR2D1BWP12T U730 ( .A1(n1979), .B1(n1986), .ZN(n437) );
  INVD1BWP12T U731 ( .I(a[2]), .ZN(n2668) );
  XNR2XD8BWP12T U732 ( .A1(n4067), .A2(n1977), .ZN(n334) );
  BUFFXD6BWP12T U733 ( .I(n334), .Z(n333) );
  XOR2XD2BWP12T U734 ( .A1(n4067), .A2(n331), .Z(n332) );
  ND2XD8BWP12T U735 ( .A1(n333), .A2(n332), .ZN(n2072) );
  XNR2D1BWP12T U736 ( .A1(n4068), .A2(n3920), .ZN(n417) );
  BUFFXD8BWP12T U737 ( .I(n334), .Z(n2070) );
  INVD1BWP12T U738 ( .I(b[6]), .ZN(n3839) );
  INVD3BWP12T U739 ( .I(n3839), .ZN(n3927) );
  XNR2D1BWP12T U740 ( .A1(n4068), .A2(n3927), .ZN(n352) );
  OAI22D1BWP12T U741 ( .A1(n2072), .A2(n417), .B1(n2070), .B2(n352), .ZN(n436)
         );
  ND2D3BWP12T U742 ( .A1(n348), .A2(n347), .ZN(n336) );
  INVD12BWP12T U743 ( .I(n3879), .ZN(n4063) );
  XOR2D2BWP12T U744 ( .A1(n4062), .A2(n4063), .Z(n335) );
  CKND2D8BWP12T U745 ( .A1(n336), .A2(n335), .ZN(n2027) );
  INVD2BWP12T U746 ( .I(b[1]), .ZN(n3853) );
  INVD8BWP12T U747 ( .I(n3853), .ZN(n3916) );
  BUFFXD8BWP12T U748 ( .I(n3916), .Z(n1517) );
  XNR2D1BWP12T U749 ( .A1(n1517), .A2(n4063), .ZN(n349) );
  XNR2XD1BWP12T U750 ( .A1(n3921), .A2(n4063), .ZN(n364) );
  OAI22D1BWP12T U751 ( .A1(n2027), .A2(n349), .B1(n1986), .B2(n364), .ZN(n358)
         );
  XNR2D1BWP12T U752 ( .A1(n4075), .A2(n3927), .ZN(n359) );
  OAI22D1BWP12T U753 ( .A1(n2083), .A2(n337), .B1(n359), .B2(n2080), .ZN(n357)
         );
  INVD8BWP12T U754 ( .I(n338), .ZN(n2098) );
  XNR2XD1BWP12T U755 ( .A1(n2098), .A2(n4084), .ZN(n363) );
  OAI22D1BWP12T U756 ( .A1(n2013), .A2(n339), .B1(n2011), .B2(n363), .ZN(n356)
         );
  INVD1BWP12T U757 ( .I(b[10]), .ZN(n3831) );
  INVD3BWP12T U758 ( .I(n3831), .ZN(n3932) );
  XNR2D1BWP12T U759 ( .A1(n1977), .A2(n3932), .ZN(n365) );
  TPOAI22D1BWP12T U760 ( .A1(n1110), .A2(n341), .B1(n365), .B2(n2018), .ZN(
        n369) );
  BUFFD3BWP12T U761 ( .I(a[10]), .Z(n4061) );
  XNR2XD8BWP12T U762 ( .A1(n4063), .A2(n4061), .ZN(n342) );
  BUFFXD12BWP12T U763 ( .I(n342), .Z(n2006) );
  INR2D2BWP12T U764 ( .A1(n1979), .B1(n2006), .ZN(n368) );
  XNR2D1BWP12T U765 ( .A1(n4068), .A2(n3929), .ZN(n351) );
  XNR2D1BWP12T U766 ( .A1(n4068), .A2(n3928), .ZN(n362) );
  HA1D1BWP12T U767 ( .A(n344), .B(n343), .CO(n354), .S(n460) );
  INVD1BWP12T U768 ( .I(n4063), .ZN(n346) );
  IND2D1BWP12T U769 ( .A1(b[0]), .B1(n595), .ZN(n345) );
  TPOAI22D1BWP12T U770 ( .A1(n2027), .A2(n346), .B1(n1986), .B2(n345), .ZN(
        n450) );
  XNR2D1BWP12T U771 ( .A1(n1979), .A2(n4063), .ZN(n350) );
  CKND2D2BWP12T U772 ( .A1(n348), .A2(n347), .ZN(n2025) );
  TPOAI22D1BWP12T U773 ( .A1(n2027), .A2(n350), .B1(n2025), .B2(n349), .ZN(
        n449) );
  OAI22D1BWP12T U774 ( .A1(n2072), .A2(n352), .B1(n2070), .B2(n351), .ZN(n448)
         );
  INVD1BWP12T U775 ( .I(n371), .ZN(n370) );
  FA1D1BWP12T U776 ( .A(n355), .B(n354), .CI(n353), .CO(n688), .S(n472) );
  FA1D0BWP12T U777 ( .A(n358), .B(n357), .CI(n356), .CO(n687), .S(n473) );
  XNR2D1BWP12T U778 ( .A1(n4075), .A2(n3929), .ZN(n677) );
  OAI22D1BWP12T U779 ( .A1(n2083), .A2(n359), .B1(n677), .B2(n2080), .ZN(n676)
         );
  DCCKND4BWP12T U780 ( .I(a[11]), .ZN(n3878) );
  INVD9BWP12T U781 ( .I(n3878), .ZN(n4060) );
  XOR2D2BWP12T U782 ( .A1(n4060), .A2(n4061), .Z(n360) );
  ND2XD16BWP12T U783 ( .A1(n360), .A2(n2006), .ZN(n2009) );
  XNR2XD1BWP12T U784 ( .A1(n4060), .A2(n1979), .ZN(n361) );
  XNR2D1BWP12T U785 ( .A1(n4060), .A2(n1517), .ZN(n678) );
  TPOAI22D1BWP12T U786 ( .A1(n2009), .A2(n361), .B1(n678), .B2(n2006), .ZN(
        n675) );
  BUFFD6BWP12T U787 ( .I(a[3]), .Z(n3885) );
  XNR2D1BWP12T U788 ( .A1(n3885), .A2(n3957), .ZN(n673) );
  OAI22D1BWP12T U789 ( .A1(n2072), .A2(n362), .B1(n2070), .B2(n673), .ZN(n674)
         );
  XNR2D1BWP12T U790 ( .A1(n4084), .A2(n3920), .ZN(n679) );
  OAI22D1BWP12T U791 ( .A1(n2013), .A2(n363), .B1(n2011), .B2(n679), .ZN(n681)
         );
  BUFFXD8BWP12T U792 ( .I(b[3]), .Z(n3922) );
  XNR2XD1BWP12T U793 ( .A1(n3922), .A2(n4063), .ZN(n671) );
  TPOAI22D1BWP12T U794 ( .A1(n2027), .A2(n364), .B1(n2025), .B2(n671), .ZN(
        n682) );
  BUFFD2BWP12T U795 ( .I(b[11]), .Z(n3933) );
  XNR2D1BWP12T U796 ( .A1(n1977), .A2(n3933), .ZN(n672) );
  OAI22D1BWP12T U797 ( .A1(n2019), .A2(n365), .B1(n672), .B2(n2018), .ZN(n670)
         );
  INVD1BWP12T U798 ( .I(n4060), .ZN(n987) );
  IND2D0BWP12T U799 ( .A1(b[0]), .B1(n4060), .ZN(n366) );
  TPOAI22D1BWP12T U800 ( .A1(n2009), .A2(n987), .B1(n2006), .B2(n366), .ZN(
        n669) );
  XOR3D2BWP12T U801 ( .A1(n681), .A2(n682), .A3(n680), .Z(n665) );
  FA1D2BWP12T U802 ( .A(n369), .B(n368), .CI(n367), .CO(n664), .S(n355) );
  XOR3D2BWP12T U803 ( .A1(n663), .A2(n665), .A3(n664), .Z(n686) );
  INVD1BWP12T U804 ( .I(n689), .ZN(n2365) );
  XNR2D1BWP12T U805 ( .A1(n3921), .A2(n1977), .ZN(n376) );
  OAI22D1BWP12T U806 ( .A1(n2019), .A2(n376), .B1(n385), .B2(n2018), .ZN(n388)
         );
  XNR2XD1BWP12T U807 ( .A1(n1979), .A2(n4068), .ZN(n373) );
  XNR2D1BWP12T U808 ( .A1(n1517), .A2(n3885), .ZN(n386) );
  OAI22D1BWP12T U809 ( .A1(n2072), .A2(n373), .B1(n2070), .B2(n386), .ZN(n387)
         );
  INVD0BWP12T U810 ( .I(n4068), .ZN(n375) );
  IND2D0BWP12T U811 ( .A1(b[0]), .B1(n3885), .ZN(n374) );
  OAI22D1BWP12T U812 ( .A1(n2072), .A2(n375), .B1(n2070), .B2(n374), .ZN(n382)
         );
  OR2D2BWP12T U813 ( .A1(n383), .A2(n382), .Z(n2516) );
  XNR2D1BWP12T U814 ( .A1(n1517), .A2(n1977), .ZN(n377) );
  OAI22D1BWP12T U815 ( .A1(n2019), .A2(n377), .B1(n376), .B2(n2018), .ZN(n380)
         );
  INR2D1BWP12T U816 ( .A1(n1979), .B1(n2070), .ZN(n379) );
  OR2XD1BWP12T U817 ( .A1(n380), .A2(n379), .Z(n2647) );
  OAI22D1BWP12T U818 ( .A1(n2019), .A2(n1979), .B1(n377), .B2(n2018), .ZN(
        n2598) );
  IND2D1BWP12T U819 ( .A1(b[0]), .B1(n1977), .ZN(n378) );
  ND2D1BWP12T U820 ( .A1(n2019), .A2(n378), .ZN(n2597) );
  ND2D1BWP12T U821 ( .A1(n2598), .A2(n2597), .ZN(n2599) );
  INVD1BWP12T U822 ( .I(n2599), .ZN(n2648) );
  ND2D1BWP12T U823 ( .A1(n380), .A2(n379), .ZN(n2646) );
  INVD1BWP12T U824 ( .I(n2646), .ZN(n381) );
  AO21D1BWP12T U825 ( .A1(n2647), .A2(n2648), .B(n381), .Z(n2517) );
  ND2D1BWP12T U826 ( .A1(n383), .A2(n382), .ZN(n2515) );
  INVD1BWP12T U827 ( .I(n2515), .ZN(n384) );
  AOI21D1BWP12T U828 ( .A1(n2516), .A2(n2517), .B(n384), .ZN(n2412) );
  XNR2D1BWP12T U829 ( .A1(n2098), .A2(n1977), .ZN(n393) );
  OAI22D1BWP12T U830 ( .A1(n393), .A2(n2018), .B1(n2019), .B2(n385), .ZN(n397)
         );
  INR2D1BWP12T U831 ( .A1(n1979), .B1(n2080), .ZN(n396) );
  XNR2XD1BWP12T U832 ( .A1(n3921), .A2(n3885), .ZN(n391) );
  OAI22D1BWP12T U833 ( .A1(n2072), .A2(n386), .B1(n2070), .B2(n391), .ZN(n395)
         );
  NR2D1BWP12T U834 ( .A1(n390), .A2(n389), .ZN(n2410) );
  ND2D1BWP12T U835 ( .A1(n390), .A2(n389), .ZN(n2411) );
  OAI21D1BWP12T U836 ( .A1(n2412), .A2(n2410), .B(n2411), .ZN(n2452) );
  XNR2XD1BWP12T U837 ( .A1(n3922), .A2(n3885), .ZN(n405) );
  OAI22D1BWP12T U838 ( .A1(n2072), .A2(n391), .B1(n2070), .B2(n405), .ZN(n408)
         );
  XNR2D1BWP12T U839 ( .A1(n4075), .A2(n1979), .ZN(n392) );
  XNR2D1BWP12T U840 ( .A1(n4075), .A2(n1517), .ZN(n403) );
  OAI22D1BWP12T U841 ( .A1(n2083), .A2(n392), .B1(n403), .B2(n2080), .ZN(n407)
         );
  XNR2D1BWP12T U842 ( .A1(n3920), .A2(n1977), .ZN(n404) );
  OAI22D1BWP12T U843 ( .A1(n2019), .A2(n393), .B1(n404), .B2(n2018), .ZN(n402)
         );
  IND2XD1BWP12T U844 ( .A1(b[0]), .B1(n4075), .ZN(n394) );
  OAI22D1BWP12T U845 ( .A1(n2083), .A2(n2634), .B1(n2080), .B2(n394), .ZN(n401) );
  ND2D1BWP12T U846 ( .A1(n399), .A2(n398), .ZN(n2451) );
  INVD1BWP12T U847 ( .I(n2451), .ZN(n400) );
  AOI21D1BWP12T U848 ( .A1(n2452), .A2(n318), .B(n400), .ZN(n607) );
  HA1D1BWP12T U849 ( .A(n402), .B(n401), .CO(n425), .S(n406) );
  XNR2D1BWP12T U850 ( .A1(n4075), .A2(n3921), .ZN(n413) );
  OAI22D1BWP12T U851 ( .A1(n2083), .A2(n403), .B1(n413), .B2(n2080), .ZN(n424)
         );
  XNR2D1BWP12T U852 ( .A1(n3927), .A2(n1977), .ZN(n412) );
  INR2D1BWP12T U853 ( .A1(n1979), .B1(n2011), .ZN(n415) );
  XNR2XD1BWP12T U854 ( .A1(n2098), .A2(n4068), .ZN(n418) );
  OAI22D1BWP12T U855 ( .A1(n2072), .A2(n405), .B1(n2070), .B2(n418), .ZN(n414)
         );
  FA1D0BWP12T U856 ( .A(n408), .B(n407), .CI(n406), .CO(n409), .S(n399) );
  NR2D1BWP12T U857 ( .A1(n410), .A2(n409), .ZN(n604) );
  ND2D1BWP12T U858 ( .A1(n410), .A2(n409), .ZN(n605) );
  OAI21D1BWP12T U859 ( .A1(n607), .A2(n604), .B(n605), .ZN(n1004) );
  OAI22D1BWP12T U860 ( .A1(n2019), .A2(n412), .B1(n411), .B2(n2018), .ZN(n444)
         );
  XNR2D1BWP12T U861 ( .A1(n4075), .A2(n3922), .ZN(n442) );
  OAI22D1BWP12T U862 ( .A1(n2083), .A2(n413), .B1(n442), .B2(n2080), .ZN(n443)
         );
  INVD1BWP12T U863 ( .I(n446), .ZN(n422) );
  FA1D1BWP12T U864 ( .A(n416), .B(n415), .CI(n414), .CO(n447), .S(n423) );
  OAI22D1BWP12T U865 ( .A1(n2072), .A2(n418), .B1(n2070), .B2(n417), .ZN(n431)
         );
  XNR2D1BWP12T U866 ( .A1(n1979), .A2(n4084), .ZN(n419) );
  XNR2D1BWP12T U867 ( .A1(n1517), .A2(n4084), .ZN(n440) );
  OAI22D1BWP12T U868 ( .A1(n2013), .A2(n419), .B1(n2011), .B2(n440), .ZN(n433)
         );
  INVD0BWP12T U869 ( .I(n4084), .ZN(n421) );
  IND2D0BWP12T U870 ( .A1(b[0]), .B1(n4084), .ZN(n420) );
  OAI22D1BWP12T U871 ( .A1(n2013), .A2(n421), .B1(n2011), .B2(n420), .ZN(n432)
         );
  XOR3D1BWP12T U872 ( .A1(n431), .A2(n433), .A3(n432), .Z(n445) );
  XNR3D1BWP12T U873 ( .A1(n422), .A2(n447), .A3(n445), .ZN(n429) );
  INVD1BWP12T U874 ( .I(n429), .ZN(n427) );
  INVD1BWP12T U875 ( .I(n428), .ZN(n426) );
  ND2D1BWP12T U876 ( .A1(n427), .A2(n426), .ZN(n1002) );
  ND2D1BWP12T U877 ( .A1(n429), .A2(n428), .ZN(n1001) );
  INVD1BWP12T U878 ( .I(n1001), .ZN(n430) );
  OAI21D1BWP12T U879 ( .A1(n433), .A2(n432), .B(n431), .ZN(n435) );
  CKND2D1BWP12T U880 ( .A1(n433), .A2(n432), .ZN(n434) );
  ND2D1BWP12T U881 ( .A1(n435), .A2(n434), .ZN(n463) );
  FA1D1BWP12T U882 ( .A(n438), .B(n437), .CI(n436), .CO(n458), .S(n462) );
  OAI22D1BWP12T U883 ( .A1(n2013), .A2(n440), .B1(n2011), .B2(n439), .ZN(n454)
         );
  OAI22D1BWP12T U884 ( .A1(n2083), .A2(n442), .B1(n441), .B2(n2080), .ZN(n455)
         );
  HA1D1BWP12T U885 ( .A(n444), .B(n443), .CO(n453), .S(n446) );
  XOR3D1BWP12T U886 ( .A1(n454), .A2(n455), .A3(n453), .Z(n461) );
  OR2D2BWP12T U887 ( .A1(n466), .A2(n465), .Z(n2793) );
  FA1D1BWP12T U888 ( .A(n450), .B(n449), .CI(n448), .CO(n353), .S(n477) );
  INVD1BWP12T U889 ( .I(n454), .ZN(n451) );
  IND2XD1BWP12T U890 ( .A1(n455), .B1(n451), .ZN(n452) );
  ND2D1BWP12T U891 ( .A1(n453), .A2(n452), .ZN(n457) );
  CKND2D1BWP12T U892 ( .A1(n455), .A2(n454), .ZN(n456) );
  ND2D1BWP12T U893 ( .A1(n457), .A2(n456), .ZN(n476) );
  FA1D1BWP12T U894 ( .A(n460), .B(n459), .CI(n458), .CO(n474), .S(n475) );
  FA1D1BWP12T U895 ( .A(n463), .B(n462), .CI(n461), .CO(n467), .S(n466) );
  TPNR2D1BWP12T U896 ( .A1(n468), .A2(n467), .ZN(n464) );
  INVD1P75BWP12T U897 ( .I(n464), .ZN(n2796) );
  CKND2D1BWP12T U898 ( .A1(n2793), .A2(n2796), .ZN(n471) );
  ND2D1BWP12T U899 ( .A1(n466), .A2(n465), .ZN(n1056) );
  INVD1BWP12T U900 ( .I(n1056), .ZN(n2792) );
  INVD1BWP12T U901 ( .I(n2795), .ZN(n469) );
  FA1D1BWP12T U902 ( .A(n474), .B(n473), .CI(n472), .CO(n371), .S(n481) );
  INVD1BWP12T U903 ( .I(n481), .ZN(n479) );
  FA1D1BWP12T U904 ( .A(n477), .B(n476), .CI(n475), .CO(n480), .S(n468) );
  INVD1BWP12T U905 ( .I(n480), .ZN(n478) );
  ND2D1BWP12T U906 ( .A1(n479), .A2(n478), .ZN(n3331) );
  ND2D1BWP12T U907 ( .A1(n481), .A2(n480), .ZN(n3330) );
  INVD1BWP12T U908 ( .I(n3330), .ZN(n482) );
  TPAOI21D1BWP12T U909 ( .A1(n3332), .A2(n3331), .B(n482), .ZN(n694) );
  INVD1BWP12T U910 ( .I(n694), .ZN(n2366) );
  ND2D1BWP12T U911 ( .A1(op[3]), .A2(op[0]), .ZN(n573) );
  INVD1BWP12T U912 ( .I(n573), .ZN(n523) );
  INR2D1BWP12T U913 ( .A1(op[2]), .B1(op[1]), .ZN(n483) );
  INVD1BWP12T U914 ( .I(b[0]), .ZN(n1854) );
  NR2XD0BWP12T U915 ( .A1(n1854), .A2(n4066), .ZN(n2590) );
  CKND0BWP12T U916 ( .I(a[1]), .ZN(n484) );
  INVD1BWP12T U917 ( .I(n484), .ZN(n581) );
  NR2D1BWP12T U918 ( .A1(n582), .A2(n496), .ZN(n2587) );
  ND2D1BWP12T U919 ( .A1(n582), .A2(n581), .ZN(n2588) );
  OAI21D1BWP12T U920 ( .A1(n2590), .A2(n2587), .B(n2588), .ZN(n2559) );
  INVD1BWP12T U921 ( .I(n3885), .ZN(n485) );
  INVD1BWP12T U922 ( .I(b[3]), .ZN(n486) );
  INR2D1BWP12T U923 ( .A1(n485), .B1(n486), .ZN(n2560) );
  NR2D1BWP12T U924 ( .A1(n583), .A2(n4067), .ZN(n2677) );
  NR2D1BWP12T U925 ( .A1(n2560), .A2(n2677), .ZN(n488) );
  CKND2D1BWP12T U926 ( .A1(n583), .A2(n4067), .ZN(n2678) );
  ND2D1BWP12T U927 ( .A1(n486), .A2(n4068), .ZN(n2561) );
  OAI21D1BWP12T U928 ( .A1(n2560), .A2(n2678), .B(n2561), .ZN(n487) );
  AOI21D1BWP12T U929 ( .A1(n2559), .A2(n488), .B(n487), .ZN(n609) );
  BUFFD2BWP12T U930 ( .I(b[4]), .Z(n500) );
  NR2D1BWP12T U931 ( .A1(n3841), .A2(n4081), .ZN(n2447) );
  NR2D1BWP12T U932 ( .A1(n588), .A2(n4075), .ZN(n2505) );
  NR2D1BWP12T U933 ( .A1(n2447), .A2(n2505), .ZN(n1030) );
  NR2D1BWP12T U934 ( .A1(n594), .A2(n4084), .ZN(n1038) );
  NR2D1BWP12T U935 ( .A1(n589), .A2(n4083), .ZN(n1034) );
  NR2D1BWP12T U936 ( .A1(n1038), .A2(n1034), .ZN(n490) );
  CKND2D1BWP12T U937 ( .A1(n1030), .A2(n490), .ZN(n492) );
  ND2D1BWP12T U938 ( .A1(n3841), .A2(n4081), .ZN(n2502) );
  CKND2D1BWP12T U939 ( .A1(n588), .A2(n4075), .ZN(n2506) );
  OAI21D1BWP12T U940 ( .A1(n2502), .A2(n2505), .B(n2506), .ZN(n1032) );
  CKND2D1BWP12T U941 ( .A1(n589), .A2(n4083), .ZN(n1033) );
  ND2D1BWP12T U942 ( .A1(n594), .A2(n4084), .ZN(n1039) );
  OAI21D1BWP12T U943 ( .A1(n1038), .A2(n1033), .B(n1039), .ZN(n489) );
  AOI21D1BWP12T U944 ( .A1(n1032), .A2(n490), .B(n489), .ZN(n491) );
  OAI21D1BWP12T U945 ( .A1(n609), .A2(n492), .B(n491), .ZN(n1724) );
  INVD1BWP12T U946 ( .I(n3957), .ZN(n493) );
  NR2D1BWP12T U947 ( .A1(n493), .A2(n4063), .ZN(n2801) );
  NR2D1BWP12T U948 ( .A1(n1909), .A2(n4062), .ZN(n2800) );
  NR2D1BWP12T U949 ( .A1(n2801), .A2(n2800), .ZN(n897) );
  INVD0BWP12T U950 ( .I(n897), .ZN(n3334) );
  INVD2P3BWP12T U951 ( .I(n3932), .ZN(n2063) );
  NR2D1BWP12T U952 ( .A1(n2063), .A2(n4061), .ZN(n3335) );
  NR2XD0BWP12T U953 ( .A1(n3334), .A2(n3335), .ZN(n2372) );
  CKND2D1BWP12T U954 ( .A1(n1909), .A2(n4062), .ZN(n2799) );
  ND2D1BWP12T U955 ( .A1(n493), .A2(n4063), .ZN(n2802) );
  OAI21D1BWP12T U956 ( .A1(n2801), .A2(n2799), .B(n2802), .ZN(n903) );
  INVD1BWP12T U957 ( .I(n903), .ZN(n3333) );
  ND2D1BWP12T U958 ( .A1(n2063), .A2(n4061), .ZN(n3336) );
  OAI21D1BWP12T U959 ( .A1(n3333), .A2(n3335), .B(n3336), .ZN(n2374) );
  CKND2D1BWP12T U960 ( .A1(n3833), .A2(n4060), .ZN(n898) );
  INVD0BWP12T U961 ( .I(op[0]), .ZN(n494) );
  IND2XD1BWP12T U962 ( .A1(op[2]), .B1(op[1]), .ZN(n518) );
  INR2D1BWP12T U963 ( .A1(n494), .B1(n518), .ZN(n566) );
  ND2D1BWP12T U964 ( .A1(n566), .A2(op[3]), .ZN(n3532) );
  INR2D1BWP12T U965 ( .A1(op[2]), .B1(op[3]), .ZN(n600) );
  INVD1BWP12T U966 ( .I(n600), .ZN(n563) );
  INVD2BWP12T U967 ( .I(n4164), .ZN(n4210) );
  NR2D1BWP12T U968 ( .A1(n3921), .A2(n4067), .ZN(n2685) );
  BUFFXD0BWP12T U969 ( .I(a[1]), .Z(n496) );
  NR2D1BWP12T U970 ( .A1(n3916), .A2(n496), .ZN(n2683) );
  TPNR2D0BWP12T U971 ( .A1(n2685), .A2(n2683), .ZN(n498) );
  CKND1BWP12T U972 ( .I(b[0]), .ZN(n495) );
  NR2D1BWP12T U973 ( .A1(n4066), .A2(c_in), .ZN(n1858) );
  CKND2D1BWP12T U974 ( .A1(n4066), .A2(c_in), .ZN(n1859) );
  OAI21D1BWP12T U975 ( .A1(n495), .A2(n1858), .B(n1859), .ZN(n2600) );
  CKND2D1BWP12T U976 ( .A1(n3916), .A2(n496), .ZN(n2682) );
  ND2D1BWP12T U977 ( .A1(n3921), .A2(n4067), .ZN(n2686) );
  OAI21D1BWP12T U978 ( .A1(n2685), .A2(n2682), .B(n2686), .ZN(n497) );
  AOI21D1BWP12T U979 ( .A1(n498), .A2(n2600), .B(n497), .ZN(n620) );
  NR2D1BWP12T U980 ( .A1(b[3]), .A2(n4068), .ZN(n2436) );
  CKBD1BWP12T U981 ( .I(n4081), .Z(n501) );
  NR2D1BWP12T U982 ( .A1(n499), .A2(n501), .ZN(n2437) );
  NR2D1BWP12T U983 ( .A1(n2436), .A2(n2437), .ZN(n2498) );
  NR2D1BWP12T U984 ( .A1(n3927), .A2(n4083), .ZN(n621) );
  NR2D1BWP12T U985 ( .A1(n2499), .A2(n621), .ZN(n503) );
  CKND2D1BWP12T U986 ( .A1(n2498), .A2(n503), .ZN(n505) );
  CKND2D1BWP12T U987 ( .A1(b[3]), .A2(n4068), .ZN(n2533) );
  BUFFXD4BWP12T U988 ( .I(n500), .Z(n3919) );
  CKND2D1BWP12T U989 ( .A1(n3919), .A2(n501), .ZN(n2438) );
  OAI21D1BWP12T U990 ( .A1(n2437), .A2(n2533), .B(n2438), .ZN(n2497) );
  CKND2D1BWP12T U991 ( .A1(n4075), .A2(n3920), .ZN(n2500) );
  CKND2D1BWP12T U992 ( .A1(n3927), .A2(n4083), .ZN(n622) );
  OAI21D1BWP12T U993 ( .A1(n621), .A2(n2500), .B(n622), .ZN(n502) );
  AOI21D1BWP12T U994 ( .A1(n2497), .A2(n503), .B(n502), .ZN(n504) );
  OAI21D1BWP12T U995 ( .A1(n620), .A2(n505), .B(n504), .ZN(n952) );
  INVD1BWP12T U996 ( .I(n952), .ZN(n3379) );
  NR2D1BWP12T U997 ( .A1(n4084), .A2(n3929), .ZN(n1083) );
  NR2D1BWP12T U998 ( .A1(n3928), .A2(n4062), .ZN(n1084) );
  NR2D1BWP12T U999 ( .A1(n1083), .A2(n1084), .ZN(n3375) );
  CKBD1BWP12T U1000 ( .I(n4063), .Z(n506) );
  NR2D1BWP12T U1001 ( .A1(n506), .A2(n3957), .ZN(n2804) );
  NR2D1BWP12T U1002 ( .A1(n3932), .A2(n4061), .ZN(n928) );
  NR2D1BWP12T U1003 ( .A1(n2804), .A2(n928), .ZN(n508) );
  ND2D1BWP12T U1004 ( .A1(n3375), .A2(n508), .ZN(n2318) );
  ND2D1BWP12T U1005 ( .A1(n4084), .A2(n3929), .ZN(n1082) );
  CKND2D1BWP12T U1006 ( .A1(n3928), .A2(n4062), .ZN(n1085) );
  OAI21D1BWP12T U1007 ( .A1(n1084), .A2(n1082), .B(n1085), .ZN(n3378) );
  ND2D1BWP12T U1008 ( .A1(n506), .A2(n3957), .ZN(n3376) );
  ND2D1BWP12T U1009 ( .A1(n3932), .A2(n4061), .ZN(n3389) );
  OAI21D1BWP12T U1010 ( .A1(n928), .A2(n3376), .B(n3389), .ZN(n507) );
  AOI21D1BWP12T U1011 ( .A1(n508), .A2(n3378), .B(n507), .ZN(n2319) );
  NR2D1BWP12T U1012 ( .A1(n4060), .A2(n3933), .ZN(n944) );
  INVD1BWP12T U1013 ( .I(n944), .ZN(n2382) );
  CKND2D1BWP12T U1014 ( .A1(n4060), .A2(n3933), .ZN(n2380) );
  CKND2D1BWP12T U1015 ( .A1(b[0]), .A2(n4066), .ZN(n2605) );
  NR2D1BWP12T U1016 ( .A1(n1962), .A2(n496), .ZN(n2602) );
  CKND2D1BWP12T U1017 ( .A1(n1962), .A2(n496), .ZN(n2603) );
  OAI21D1BWP12T U1018 ( .A1(n2605), .A2(n2602), .B(n2603), .ZN(n2530) );
  NR2D1BWP12T U1019 ( .A1(b[3]), .A2(n4068), .ZN(n2531) );
  CKBD1BWP12T U1020 ( .I(n4067), .Z(n509) );
  NR2D1BWP12T U1021 ( .A1(n3921), .A2(n509), .ZN(n2660) );
  NR2D1BWP12T U1022 ( .A1(n2531), .A2(n2660), .ZN(n511) );
  CKND2D1BWP12T U1023 ( .A1(n3921), .A2(n509), .ZN(n2661) );
  CKND2D1BWP12T U1024 ( .A1(n3922), .A2(n3885), .ZN(n2532) );
  OAI21D1BWP12T U1025 ( .A1(n2531), .A2(n2661), .B(n2532), .ZN(n510) );
  AOI21D1BWP12T U1026 ( .A1(n2530), .A2(n511), .B(n510), .ZN(n623) );
  CKBD1BWP12T U1027 ( .I(n4081), .Z(n512) );
  NR2D1BWP12T U1028 ( .A1(n4075), .A2(n3920), .ZN(n2491) );
  NR2D1BWP12T U1029 ( .A1(n4084), .A2(n3929), .ZN(n1018) );
  NR2D1BWP12T U1030 ( .A1(n3927), .A2(n4083), .ZN(n1014) );
  NR2D1BWP12T U1031 ( .A1(n1018), .A2(n1014), .ZN(n514) );
  ND2D1BWP12T U1032 ( .A1(n1010), .A2(n514), .ZN(n516) );
  CKND2D1BWP12T U1033 ( .A1(n3919), .A2(n512), .ZN(n2489) );
  CKND2D1BWP12T U1034 ( .A1(n4075), .A2(n3920), .ZN(n2492) );
  OAI21D1BWP12T U1035 ( .A1(n2491), .A2(n2489), .B(n2492), .ZN(n1012) );
  CKND2D1BWP12T U1036 ( .A1(n3927), .A2(n4083), .ZN(n1013) );
  CKND2D1BWP12T U1037 ( .A1(n4084), .A2(n3929), .ZN(n1019) );
  OAI21D1BWP12T U1038 ( .A1(n1018), .A2(n1013), .B(n1019), .ZN(n513) );
  AOI21D1BWP12T U1039 ( .A1(n1012), .A2(n514), .B(n513), .ZN(n515) );
  TPOAI21D1BWP12T U1040 ( .A1(n623), .A2(n516), .B(n515), .ZN(n941) );
  INVD1BWP12T U1041 ( .I(n941), .ZN(n3388) );
  CKBD1BWP12T U1042 ( .I(n4063), .Z(n517) );
  NR2D1BWP12T U1043 ( .A1(n517), .A2(n3957), .ZN(n2818) );
  NR2D1BWP12T U1044 ( .A1(n3928), .A2(n4062), .ZN(n2817) );
  NR2D1BWP12T U1045 ( .A1(n2818), .A2(n2817), .ZN(n3386) );
  INVD1BWP12T U1046 ( .I(n928), .ZN(n3390) );
  CKND2D1BWP12T U1047 ( .A1(n3928), .A2(n4062), .ZN(n2816) );
  CKND2D1BWP12T U1048 ( .A1(n517), .A2(n3957), .ZN(n2819) );
  OAI21D1BWP12T U1049 ( .A1(n2818), .A2(n2816), .B(n2819), .ZN(n3387) );
  NR2D1BWP12T U1050 ( .A1(n4060), .A2(n3933), .ZN(n930) );
  CKND2D1BWP12T U1051 ( .A1(n4060), .A2(n3933), .ZN(n929) );
  NR2D2BWP12T U1052 ( .A1(n518), .A2(n573), .ZN(n4206) );
  INVD1BWP12T U1053 ( .I(n4083), .ZN(n3890) );
  ND2D1BWP12T U1054 ( .A1(n421), .A2(n3890), .ZN(n519) );
  NR2D1BWP12T U1055 ( .A1(n1046), .A2(n519), .ZN(n522) );
  INVD1BWP12T U1056 ( .I(n4068), .ZN(n520) );
  INVD1BWP12T U1057 ( .I(n4067), .ZN(n2542) );
  ND2D1BWP12T U1058 ( .A1(n520), .A2(n2542), .ZN(n521) );
  ND2D1BWP12T U1059 ( .A1(n484), .A2(n2018), .ZN(n2541) );
  NR2D1BWP12T U1060 ( .A1(n521), .A2(n2541), .ZN(n625) );
  ND2D1BWP12T U1061 ( .A1(n522), .A2(n625), .ZN(n993) );
  INVD1BWP12T U1062 ( .I(n993), .ZN(n3351) );
  TPNR2D0BWP12T U1063 ( .A1(op[2]), .A2(op[1]), .ZN(n568) );
  ND2D1BWP12T U1064 ( .A1(n523), .A2(n568), .ZN(n3613) );
  INVD2BWP12T U1065 ( .I(n3613), .ZN(n4203) );
  INVD1BWP12T U1066 ( .I(n3886), .ZN(n524) );
  NR2D1BWP12T U1067 ( .A1(n524), .A2(b[0]), .ZN(n525) );
  ND2D2BWP12T U1068 ( .A1(n582), .A2(n525), .ZN(n2629) );
  ND2D1BWP12T U1069 ( .A1(b[3]), .A2(n3919), .ZN(n2780) );
  INVD1BWP12T U1070 ( .I(n2780), .ZN(n526) );
  AOI21D2BWP12T U1071 ( .A1(n2629), .A2(n3919), .B(n526), .ZN(n3170) );
  CKND2D1BWP12T U1072 ( .A1(op[0]), .A2(op[1]), .ZN(n551) );
  INR2D2BWP12T U1073 ( .A1(n600), .B1(n551), .ZN(n4163) );
  NR2D1BWP12T U1074 ( .A1(n3170), .A2(n4201), .ZN(n3361) );
  TPNR2D3BWP12T U1075 ( .A1(n3916), .A2(b[0]), .ZN(n2462) );
  INVD3BWP12T U1076 ( .I(n2462), .ZN(n2469) );
  ND2XD3BWP12T U1077 ( .A1(n2469), .A2(n3921), .ZN(n641) );
  CKND2D2BWP12T U1078 ( .A1(n641), .A2(n2629), .ZN(n967) );
  ND2D3BWP12T U1079 ( .A1(n3916), .A2(b[0]), .ZN(n2468) );
  INVD1P75BWP12T U1080 ( .I(n2468), .ZN(n2454) );
  INVD1P75BWP12T U1081 ( .I(n527), .ZN(n640) );
  INVD2BWP12T U1082 ( .I(n640), .ZN(n1088) );
  ND2D1BWP12T U1083 ( .A1(n967), .A2(n1088), .ZN(n970) );
  INVD1BWP12T U1084 ( .I(n970), .ZN(n2806) );
  CKND2D1BWP12T U1085 ( .A1(b[0]), .A2(n2018), .ZN(n3887) );
  INVD2BWP12T U1086 ( .I(n967), .ZN(n1089) );
  NR2XD3BWP12T U1087 ( .A1(n1089), .A2(n1088), .ZN(n3707) );
  MUX2D1BWP12T U1088 ( .I0(n4068), .I1(n4067), .S(b[0]), .Z(n2824) );
  AOI22D1BWP12T U1089 ( .A1(n2806), .A2(n2586), .B1(n3707), .B2(n2824), .ZN(
        n3687) );
  MUX2XD0BWP12T U1090 ( .I0(n3879), .I1(n3880), .S(b[0]), .Z(n2807) );
  INVD1BWP12T U1091 ( .I(n2807), .ZN(n2821) );
  INR2D2BWP12T U1092 ( .A1(n640), .B1(n967), .ZN(n3229) );
  INVD2BWP12T U1093 ( .I(n3229), .ZN(n3703) );
  MUX2D1BWP12T U1094 ( .I0(n4084), .I1(n4083), .S(b[0]), .Z(n2822) );
  OAI22D1BWP12T U1095 ( .A1(n970), .A2(n2821), .B1(n3703), .B2(n2822), .ZN(
        n530) );
  INVD2BWP12T U1096 ( .I(n3707), .ZN(n3005) );
  MUX2XD0BWP12T U1097 ( .I0(n3878), .I1(n3877), .S(b[0]), .Z(n3244) );
  INVD1BWP12T U1098 ( .I(n3244), .ZN(n3230) );
  INVD1BWP12T U1099 ( .I(n641), .ZN(n528) );
  NR2D2BWP12T U1100 ( .A1(n640), .A2(n528), .ZN(n3231) );
  INVD1BWP12T U1101 ( .I(n3231), .ZN(n3705) );
  OAI22D1BWP12T U1102 ( .A1(n3005), .A2(n3230), .B1(n2823), .B2(n3705), .ZN(
        n529) );
  NR2D1BWP12T U1103 ( .A1(n530), .A2(n529), .ZN(n3167) );
  AOI22D1BWP12T U1104 ( .A1(n3627), .A2(n4203), .B1(n3361), .B2(n3693), .ZN(
        n531) );
  IOA21D1BWP12T U1105 ( .A1(n3577), .A2(n4206), .B(n531), .ZN(n580) );
  NR2D1BWP12T U1106 ( .A1(n3957), .A2(n3928), .ZN(n533) );
  NR2D1BWP12T U1107 ( .A1(n3929), .A2(n3927), .ZN(n532) );
  ND2D1BWP12T U1108 ( .A1(n533), .A2(n532), .ZN(n539) );
  NR2XD0BWP12T U1109 ( .A1(b[29]), .A2(b[28]), .ZN(n535) );
  BUFFD2BWP12T U1110 ( .I(b[26]), .Z(n3917) );
  NR2XD0BWP12T U1111 ( .A1(n3942), .A2(n3917), .ZN(n534) );
  ND2D1BWP12T U1112 ( .A1(n535), .A2(n534), .ZN(n538) );
  BUFFD2BWP12T U1113 ( .I(b[30]), .Z(n3940) );
  NR2XD0BWP12T U1114 ( .A1(b[31]), .A2(n3940), .ZN(n536) );
  CKND2D1BWP12T U1115 ( .A1(n536), .A2(n3842), .ZN(n537) );
  NR2XD0BWP12T U1116 ( .A1(b[25]), .A2(n3918), .ZN(n541) );
  BUFFD2BWP12T U1117 ( .I(b[23]), .Z(n3943) );
  BUFFD2BWP12T U1118 ( .I(b[22]), .Z(n3941) );
  NR2D1BWP12T U1119 ( .A1(n3943), .A2(n3941), .ZN(n540) );
  CKND2D1BWP12T U1120 ( .A1(n541), .A2(n540), .ZN(n543) );
  BUFFD2BWP12T U1121 ( .I(b[20]), .Z(n3938) );
  NR2XD0BWP12T U1122 ( .A1(n543), .A2(n542), .ZN(n549) );
  BUFFD2BWP12T U1123 ( .I(b[17]), .Z(n3952) );
  BUFFD2BWP12T U1124 ( .I(b[16]), .Z(n4191) );
  BUFFD2BWP12T U1125 ( .I(b[15]), .Z(n3949) );
  BUFFD2BWP12T U1126 ( .I(b[14]), .Z(n3930) );
  BUFFD2BWP12T U1127 ( .I(b[13]), .Z(n3931) );
  NR2D1BWP12T U1128 ( .A1(n3931), .A2(n3950), .ZN(n545) );
  NR2D1BWP12T U1129 ( .A1(n3933), .A2(n3932), .ZN(n544) );
  ND2D1BWP12T U1130 ( .A1(n545), .A2(n544), .ZN(n546) );
  NR2XD0BWP12T U1131 ( .A1(n547), .A2(n546), .ZN(n548) );
  ND3D2BWP12T U1132 ( .A1(n550), .A2(n549), .A3(n548), .ZN(n3655) );
  INVD2BWP12T U1133 ( .I(n3655), .ZN(n650) );
  NR3D1BWP12T U1134 ( .A1(n551), .A2(op[3]), .A3(op[2]), .ZN(n3973) );
  ND2D1BWP12T U1135 ( .A1(n650), .A2(n3973), .ZN(n2978) );
  CKND2D1BWP12T U1136 ( .A1(n2978), .A2(n4201), .ZN(n2921) );
  INVD1BWP12T U1137 ( .I(n2921), .ZN(n2529) );
  INVD1P75BWP12T U1138 ( .I(n2471), .ZN(n1845) );
  IND2D4BWP12T U1139 ( .A1(n3916), .B1(b[0]), .ZN(n2470) );
  BUFFD6BWP12T U1140 ( .I(a[28]), .Z(n4065) );
  AOI22D1BWP12T U1141 ( .A1(n1845), .A2(a[29]), .B1(n2463), .B2(n4065), .ZN(
        n553) );
  AOI22D1BWP12T U1142 ( .A1(n2454), .A2(a[30]), .B1(n2462), .B2(n4077), .ZN(
        n552) );
  ND2D1BWP12T U1143 ( .A1(n553), .A2(n552), .ZN(n2570) );
  INVD1BWP12T U1144 ( .I(n2570), .ZN(n1005) );
  CKND2D1BWP12T U1145 ( .A1(n2523), .A2(n4044), .ZN(n3994) );
  INVD1BWP12T U1146 ( .I(a[23]), .ZN(n3863) );
  CKND3BWP12T U1147 ( .I(a[25]), .ZN(n4160) );
  BUFFD6BWP12T U1148 ( .I(a[24]), .Z(n4064) );
  INVD2BWP12T U1149 ( .I(n4064), .ZN(n3898) );
  ND2D1BWP12T U1150 ( .A1(b[3]), .A2(n3921), .ZN(n2948) );
  INVD1BWP12T U1151 ( .I(a[19]), .ZN(n3866) );
  BUFFD2BWP12T U1152 ( .I(a[22]), .Z(n4070) );
  INVD1BWP12T U1153 ( .I(n4070), .ZN(n3862) );
  OAI22D0BWP12T U1154 ( .A1(n2469), .A2(n3866), .B1(n2468), .B2(n3862), .ZN(
        n555) );
  BUFFD2BWP12T U1155 ( .I(a[20]), .Z(n4069) );
  INVD1BWP12T U1156 ( .I(n4069), .ZN(n3865) );
  OAI22D1BWP12T U1157 ( .A1(n3864), .A2(n2471), .B1(n2470), .B2(n3865), .ZN(
        n554) );
  NR2D1BWP12T U1158 ( .A1(n555), .A2(n554), .ZN(n2520) );
  TPNR2D3BWP12T U1159 ( .A1(n4044), .A2(n3921), .ZN(n2641) );
  OAI22D0BWP12T U1160 ( .A1(n2469), .A2(n3878), .B1(n2468), .B2(n3873), .ZN(
        n557) );
  CKND0BWP12T U1161 ( .I(a[13]), .ZN(n3875) );
  OAI22D1BWP12T U1162 ( .A1(n2471), .A2(n3875), .B1(n2470), .B2(n3876), .ZN(
        n556) );
  NR2D1BWP12T U1163 ( .A1(n557), .A2(n556), .ZN(n2525) );
  INVD2BWP12T U1164 ( .I(b[4]), .ZN(n3841) );
  INVD4BWP12T U1165 ( .I(a[15]), .ZN(n3874) );
  BUFFD2BWP12T U1166 ( .I(a[18]), .Z(n3820) );
  INVD1BWP12T U1167 ( .I(n3820), .ZN(n3867) );
  OAI22D1BWP12T U1168 ( .A1(n2469), .A2(n3874), .B1(n2468), .B2(n3867), .ZN(
        n559) );
  BUFFD6BWP12T U1169 ( .I(a[16]), .Z(n4183) );
  OAI22D1BWP12T U1170 ( .A1(n2471), .A2(n3868), .B1(n2470), .B2(n4187), .ZN(
        n558) );
  NR2D1BWP12T U1171 ( .A1(n559), .A2(n558), .ZN(n2524) );
  IND2D1BWP12T U1172 ( .A1(n1189), .B1(n3921), .ZN(n3356) );
  AO21D0BWP12T U1173 ( .A1(n3994), .A2(n3919), .B(n561), .Z(n3734) );
  INVD1BWP12T U1174 ( .I(n2955), .ZN(n3353) );
  CKND2D0BWP12T U1175 ( .A1(n2570), .A2(n3353), .ZN(n560) );
  ND2D1BWP12T U1176 ( .A1(n3922), .A2(n4089), .ZN(n2970) );
  OAI211D0BWP12T U1177 ( .A1(n3356), .A2(n3911), .B(n560), .C(n2970), .ZN(
        n2869) );
  BUFFD6BWP12T U1178 ( .I(n650), .Z(n3986) );
  ND2D4BWP12T U1179 ( .A1(n650), .A2(n3841), .ZN(n3765) );
  CKND4BWP12T U1180 ( .I(n3765), .ZN(n3997) );
  AOI21D0BWP12T U1181 ( .A1(n2869), .A2(n3986), .B(n3997), .ZN(n562) );
  ND2D2BWP12T U1182 ( .A1(n3655), .A2(n4089), .ZN(n3384) );
  OAI21D0BWP12T U1183 ( .A1(n562), .A2(n561), .B(n3384), .ZN(n4016) );
  NR2D1BWP12T U1184 ( .A1(op[0]), .A2(op[1]), .ZN(n2202) );
  INR2D2BWP12T U1185 ( .A1(n2202), .B1(n563), .ZN(n4011) );
  CKND2D0BWP12T U1186 ( .A1(n4016), .A2(n4011), .ZN(n578) );
  ND2D1BWP12T U1187 ( .A1(n3916), .A2(n3921), .ZN(n3786) );
  OR2D2BWP12T U1188 ( .A1(n3921), .A2(n3916), .Z(n3780) );
  INVD1BWP12T U1189 ( .I(n3780), .ZN(n3241) );
  IND2XD2BWP12T U1190 ( .A1(n3921), .B1(n3916), .ZN(n3782) );
  INVD1BWP12T U1191 ( .I(n3782), .ZN(n3238) );
  AOI22D0BWP12T U1192 ( .A1(n3241), .A2(n3244), .B1(n2807), .B2(n3238), .ZN(
        n565) );
  INVD1BWP12T U1193 ( .I(n2822), .ZN(n2805) );
  TPND2D0BWP12T U1194 ( .A1(n2805), .A2(n3242), .ZN(n564) );
  OAI211D1BWP12T U1195 ( .A1(n2823), .A2(n3786), .B(n565), .C(n564), .ZN(n3165) );
  INVD1BWP12T U1196 ( .I(n2824), .ZN(n2808) );
  INVD1BWP12T U1197 ( .I(n2586), .ZN(n2595) );
  OAI22D1BWP12T U1198 ( .A1(n2808), .A2(n3780), .B1(n2595), .B2(n3782), .ZN(
        n3756) );
  INVD0BWP12T U1199 ( .I(op[3]), .ZN(n567) );
  ND2D1BWP12T U1200 ( .A1(n566), .A2(n567), .ZN(n3773) );
  INVD1BWP12T U1201 ( .I(n3773), .ZN(n4195) );
  CKND2D1BWP12T U1202 ( .A1(n3841), .A2(n4195), .ZN(n651) );
  INVD1BWP12T U1203 ( .I(n3372), .ZN(n1860) );
  INR2D1BWP12T U1204 ( .A1(op[2]), .B1(n567), .ZN(n570) );
  ND2D1BWP12T U1205 ( .A1(n570), .A2(n2202), .ZN(n4181) );
  NR2D0BWP12T U1206 ( .A1(n4060), .A2(n4182), .ZN(n569) );
  OA21XD0BWP12T U1207 ( .A1(n4185), .A2(n569), .B(n3933), .Z(n576) );
  INR2D1BWP12T U1208 ( .A1(op[1]), .B1(op[0]), .ZN(n601) );
  CKND0BWP12T U1209 ( .I(op[2]), .ZN(n2201) );
  TPND2D0BWP12T U1210 ( .A1(n2202), .A2(n2201), .ZN(n2664) );
  INVD1BWP12T U1211 ( .I(n2664), .ZN(n3363) );
  MUX2ND0BWP12T U1212 ( .I0(n4184), .I1(n2664), .S(n3933), .ZN(n571) );
  NR2D0BWP12T U1213 ( .A1(n571), .A2(n4185), .ZN(n574) );
  CKND2D0BWP12T U1214 ( .A1(op[2]), .A2(op[1]), .ZN(n572) );
  NR2D1BWP12T U1215 ( .A1(n573), .A2(n572), .ZN(n3366) );
  INVD1BWP12T U1216 ( .I(n3366), .ZN(n2205) );
  MUX2ND0BWP12T U1217 ( .I0(n574), .I1(n2205), .S(n3878), .ZN(n575) );
  AOI211D1BWP12T U1218 ( .A1(n3751), .A2(n1860), .B(n576), .C(n575), .ZN(n577)
         );
  OAI211D1BWP12T U1219 ( .A1(n2529), .A2(n3734), .B(n578), .C(n577), .ZN(n579)
         );
  RCAOI211D0BWP12T U1220 ( .A1(n4210), .A2(n4098), .B(n580), .C(n579), .ZN(
        n603) );
  NR2D1BWP12T U1221 ( .A1(n583), .A2(n4067), .ZN(n2658) );
  NR2D1BWP12T U1222 ( .A1(n582), .A2(n581), .ZN(n2656) );
  NR2D1BWP12T U1223 ( .A1(n2658), .A2(n2656), .ZN(n585) );
  NR2D1BWP12T U1224 ( .A1(n4066), .A2(c_in), .ZN(n1855) );
  CKND2D1BWP12T U1225 ( .A1(n4066), .A2(c_in), .ZN(n1856) );
  OAI21D1BWP12T U1226 ( .A1(b[0]), .A2(n1855), .B(n1856), .ZN(n2593) );
  CKND2D1BWP12T U1227 ( .A1(n582), .A2(n581), .ZN(n2655) );
  CKND2D1BWP12T U1228 ( .A1(n583), .A2(n4067), .ZN(n2659) );
  OAI21D1BWP12T U1229 ( .A1(n2658), .A2(n2655), .B(n2659), .ZN(n584) );
  AOI21D1BWP12T U1230 ( .A1(n585), .A2(n2593), .B(n584), .ZN(n611) );
  INVD1BWP12T U1231 ( .I(n3922), .ZN(n586) );
  NR2D1BWP12T U1232 ( .A1(n586), .A2(n3885), .ZN(n2444) );
  CKBD1BWP12T U1233 ( .I(n4081), .Z(n587) );
  NR2D1BWP12T U1234 ( .A1(n3841), .A2(n587), .ZN(n2445) );
  NR2D1BWP12T U1235 ( .A1(n2444), .A2(n2445), .ZN(n2508) );
  NR2D1BWP12T U1236 ( .A1(n588), .A2(n4075), .ZN(n2509) );
  NR2D1BWP12T U1237 ( .A1(n589), .A2(n4083), .ZN(n616) );
  NR2D1BWP12T U1238 ( .A1(n2509), .A2(n616), .ZN(n591) );
  CKND2D1BWP12T U1239 ( .A1(n2508), .A2(n591), .ZN(n593) );
  ND2D1BWP12T U1240 ( .A1(n586), .A2(n4068), .ZN(n2536) );
  ND2D1BWP12T U1241 ( .A1(n3841), .A2(n587), .ZN(n2446) );
  OAI21D1BWP12T U1242 ( .A1(n2445), .A2(n2536), .B(n2446), .ZN(n2507) );
  CKND2D1BWP12T U1243 ( .A1(n588), .A2(n4075), .ZN(n2510) );
  CKND2D1BWP12T U1244 ( .A1(n589), .A2(n4083), .ZN(n617) );
  OAI21D1BWP12T U1245 ( .A1(n616), .A2(n2510), .B(n617), .ZN(n590) );
  AOI21D1BWP12T U1246 ( .A1(n2507), .A2(n591), .B(n590), .ZN(n592) );
  OAI21D1BWP12T U1247 ( .A1(n611), .A2(n593), .B(n592), .ZN(n920) );
  INVD1BWP12T U1248 ( .I(n920), .ZN(n3345) );
  NR2D1BWP12T U1249 ( .A1(n594), .A2(n4084), .ZN(n1058) );
  NR2D1BWP12T U1250 ( .A1(n1909), .A2(n4062), .ZN(n1059) );
  NR2D1BWP12T U1251 ( .A1(n1058), .A2(n1059), .ZN(n3338) );
  CKBD1BWP12T U1252 ( .I(n4063), .Z(n595) );
  NR2D1BWP12T U1253 ( .A1(n1959), .A2(n595), .ZN(n2803) );
  NR2D1BWP12T U1254 ( .A1(n2063), .A2(n4061), .ZN(n3346) );
  NR2D1BWP12T U1255 ( .A1(n2803), .A2(n3346), .ZN(n597) );
  ND2D1BWP12T U1256 ( .A1(n3338), .A2(n597), .ZN(n2346) );
  ND2D1BWP12T U1257 ( .A1(n594), .A2(n4084), .ZN(n1057) );
  CKND2D1BWP12T U1258 ( .A1(n1909), .A2(n4062), .ZN(n1060) );
  OAI21D1BWP12T U1259 ( .A1(n1059), .A2(n1057), .B(n1060), .ZN(n3342) );
  ND2D1BWP12T U1260 ( .A1(n1959), .A2(n595), .ZN(n3339) );
  CKND2D1BWP12T U1261 ( .A1(n2063), .A2(n4061), .ZN(n3347) );
  OAI21D1BWP12T U1262 ( .A1(n3346), .A2(n3339), .B(n3347), .ZN(n596) );
  RCAOI21D1BWP12T U1263 ( .A1(n597), .A2(n3342), .B(n596), .ZN(n2347) );
  OAI21D1BWP12T U1264 ( .A1(n3345), .A2(n2346), .B(n2347), .ZN(n599) );
  ND2D1BWP12T U1265 ( .A1(n3833), .A2(n4060), .ZN(n2377) );
  ND2D1BWP12T U1266 ( .A1(n316), .A2(n2377), .ZN(n598) );
  XNR2XD1BWP12T U1267 ( .A1(n599), .A2(n598), .ZN(n3466) );
  ND2D1BWP12T U1268 ( .A1(n601), .A2(n600), .ZN(n3479) );
  INVD2BWP12T U1269 ( .I(n3479), .ZN(n4173) );
  CKND2D1BWP12T U1270 ( .A1(n3466), .A2(n4173), .ZN(n602) );
  INVD0BWP12T U1271 ( .I(n604), .ZN(n606) );
  CKND2D1BWP12T U1272 ( .A1(n606), .A2(n605), .ZN(n608) );
  XOR2XD1BWP12T U1273 ( .A1(n608), .A2(n607), .Z(n3417) );
  INVD1BWP12T U1274 ( .I(n3417), .ZN(n662) );
  INVD2BWP12T U1275 ( .I(n3532), .ZN(n4215) );
  INVD1BWP12T U1276 ( .I(n609), .ZN(n2504) );
  CKND0BWP12T U1277 ( .I(n1034), .ZN(n610) );
  INVD1BWP12T U1278 ( .I(n611), .ZN(n2539) );
  CKND0BWP12T U1279 ( .I(n2508), .ZN(n612) );
  NR2D0BWP12T U1280 ( .A1(n612), .A2(n2509), .ZN(n615) );
  CKND0BWP12T U1281 ( .I(n2507), .ZN(n613) );
  OAI21D0BWP12T U1282 ( .A1(n613), .A2(n2509), .B(n2510), .ZN(n614) );
  AOI21D1BWP12T U1283 ( .A1(n2539), .A2(n615), .B(n614), .ZN(n619) );
  CKND2D0BWP12T U1284 ( .A1(n610), .A2(n617), .ZN(n618) );
  XOR2XD1BWP12T U1285 ( .A1(n619), .A2(n618), .Z(n3476) );
  INVD1BWP12T U1286 ( .I(n620), .ZN(n2535) );
  INVD1BWP12T U1287 ( .I(n623), .ZN(n2490) );
  INVD0BWP12T U1288 ( .I(n1014), .ZN(n624) );
  INVD1BWP12T U1289 ( .I(n625), .ZN(n2479) );
  OAI22D1BWP12T U1290 ( .A1(n2469), .A2(n3862), .B1(n2468), .B2(n4160), .ZN(
        n627) );
  OAI22D1BWP12T U1291 ( .A1(n2471), .A2(n3898), .B1(n2470), .B2(n3863), .ZN(
        n626) );
  NR2D1BWP12T U1292 ( .A1(n627), .A2(n626), .ZN(n962) );
  INVD1BWP12T U1293 ( .I(n962), .ZN(n2299) );
  MUX2D1BWP12T U1294 ( .I0(n4076), .I1(n4077), .S(b[0]), .Z(n1065) );
  INVD1BWP12T U1295 ( .I(n965), .ZN(n3026) );
  INVD1BWP12T U1296 ( .I(n3356), .ZN(n2579) );
  AOI22D1BWP12T U1297 ( .A1(n2299), .A2(n3353), .B1(n3026), .B2(n2579), .ZN(
        n658) );
  TPND2D0BWP12T U1298 ( .A1(n2304), .A2(n2641), .ZN(n628) );
  ND2D1BWP12T U1299 ( .A1(n658), .A2(n628), .ZN(n3683) );
  OAI22D1BWP12T U1300 ( .A1(n2469), .A2(n3873), .B1(n2468), .B2(n3868), .ZN(
        n630) );
  OAI22D1BWP12T U1301 ( .A1(n2471), .A2(n4187), .B1(n2470), .B2(n3874), .ZN(
        n629) );
  NR2D1BWP12T U1302 ( .A1(n630), .A2(n629), .ZN(n3357) );
  AOI22D1BWP12T U1303 ( .A1(n1845), .A2(n4062), .B1(n2463), .B2(n4084), .ZN(
        n632) );
  AOI22D1BWP12T U1304 ( .A1(n2454), .A2(n4063), .B1(n2462), .B2(n4083), .ZN(
        n631) );
  ND2D1BWP12T U1305 ( .A1(n632), .A2(n631), .ZN(n2628) );
  CKND1BWP12T U1306 ( .I(n2628), .ZN(n633) );
  OAI22D0BWP12T U1307 ( .A1(n2469), .A2(n4061), .B1(a[13]), .B2(n2468), .ZN(
        n635) );
  OAI22D1BWP12T U1308 ( .A1(n4078), .A2(n2471), .B1(n2470), .B2(n4060), .ZN(
        n634) );
  NR2D1BWP12T U1309 ( .A1(n635), .A2(n634), .ZN(n3354) );
  CKND0BWP12T U1310 ( .I(n3354), .ZN(n636) );
  OAI22D1BWP12T U1311 ( .A1(n2469), .A2(n3867), .B1(n2468), .B2(n3864), .ZN(
        n638) );
  OAI22D1BWP12T U1312 ( .A1(n2471), .A2(n3865), .B1(n2470), .B2(n3866), .ZN(
        n637) );
  NR2D1BWP12T U1313 ( .A1(n638), .A2(n637), .ZN(n2301) );
  INVD0BWP12T U1314 ( .I(n3718), .ZN(n639) );
  OAI211D1BWP12T U1315 ( .A1(n3841), .A2(n3683), .B(n639), .C(n3986), .ZN(
        n3972) );
  INVD1BWP12T U1316 ( .I(n3973), .ZN(n2834) );
  NR2D1BWP12T U1317 ( .A1(n3919), .A2(n4201), .ZN(n3360) );
  AOI21D0BWP12T U1318 ( .A1(n4163), .A2(n3683), .B(n3360), .ZN(n655) );
  OAI21D0BWP12T U1319 ( .A1(n4083), .A2(n4182), .B(n4181), .ZN(n649) );
  MUX2D1BWP12T U1320 ( .I0(n4067), .I1(n581), .S(b[0]), .Z(n1832) );
  INVD1BWP12T U1321 ( .I(n1832), .ZN(n652) );
  MUX2D1BWP12T U1322 ( .I0(n4083), .I1(n4075), .S(b[0]), .Z(n1838) );
  CKND2D1BWP12T U1323 ( .A1(n3707), .A2(n1838), .ZN(n643) );
  CKND2D1BWP12T U1324 ( .A1(n1845), .A2(n4066), .ZN(n981) );
  INVD1BWP12T U1325 ( .I(n981), .ZN(n966) );
  TPNR2D2BWP12T U1326 ( .A1(n641), .A2(n640), .ZN(n3227) );
  CKMUX2D1BWP12T U1327 ( .I0(n4081), .I1(n3885), .S(b[0]), .Z(n1833) );
  AOI22D1BWP12T U1328 ( .A1(n1089), .A2(n966), .B1(n3227), .B2(n1833), .ZN(
        n642) );
  OAI211D1BWP12T U1329 ( .A1(n3703), .A2(n652), .B(n643), .C(n642), .ZN(n3100)
         );
  INVD1BWP12T U1330 ( .I(n3100), .ZN(n3688) );
  NR2D0BWP12T U1331 ( .A1(n3170), .A2(n4201), .ZN(n644) );
  ND2D1BWP12T U1332 ( .A1(n2547), .A2(n644), .ZN(n2480) );
  NR2D1BWP12T U1333 ( .A1(n3688), .A2(n2480), .ZN(n648) );
  MUX2ND0BWP12T U1334 ( .I0(n4184), .I1(n2664), .S(n3927), .ZN(n645) );
  NR2XD0BWP12T U1335 ( .A1(n645), .A2(n4185), .ZN(n646) );
  MUX2NXD0BWP12T U1336 ( .I0(n646), .I1(n2205), .S(n3890), .ZN(n647) );
  AOI211D1BWP12T U1337 ( .A1(n3927), .A2(n649), .B(n648), .C(n647), .ZN(n654)
         );
  IND3D4BWP12T U1338 ( .A1(n651), .B1(n4044), .B2(n650), .ZN(n2675) );
  INVD1BWP12T U1339 ( .I(n2675), .ZN(n2596) );
  ND2D1BWP12T U1340 ( .A1(n981), .A2(n652), .ZN(n983) );
  ND2D1BWP12T U1341 ( .A1(n2596), .A2(n3754), .ZN(n653) );
  OAI211D1BWP12T U1342 ( .A1(n3718), .A2(n655), .B(n654), .C(n653), .ZN(n656)
         );
  AOI211D1BWP12T U1343 ( .A1(n4215), .A2(n3536), .B(n657), .C(n656), .ZN(n661)
         );
  INVD1BWP12T U1344 ( .I(n961), .ZN(n3025) );
  MUX2NXD0BWP12T U1345 ( .I0(n3025), .I1(n4089), .S(n3921), .ZN(n2314) );
  OAI21D1BWP12T U1346 ( .A1(n2314), .A2(n4044), .B(n658), .ZN(n4038) );
  AOI21D1BWP12T U1347 ( .A1(n4038), .A2(n3986), .B(n3997), .ZN(n659) );
  OAI21D1BWP12T U1348 ( .A1(n659), .A2(n3718), .B(n3384), .ZN(n4031) );
  ND2D1BWP12T U1349 ( .A1(n4031), .A2(n4011), .ZN(n660) );
  OAI211D1BWP12T U1350 ( .A1(n3407), .A2(n662), .B(n661), .C(n660), .ZN(
        result[6]) );
  ND2D1BWP12T U1351 ( .A1(n663), .A2(n665), .ZN(n668) );
  CKND2D1BWP12T U1352 ( .A1(n663), .A2(n664), .ZN(n667) );
  CKND2D1BWP12T U1353 ( .A1(n665), .A2(n664), .ZN(n666) );
  ND3D1BWP12T U1354 ( .A1(n668), .A2(n667), .A3(n666), .ZN(n745) );
  HA1D0BWP12T U1355 ( .A(n670), .B(n669), .CO(n704), .S(n680) );
  XNR2XD1BWP12T U1356 ( .A1(n2098), .A2(n4063), .ZN(n695) );
  OAI22D1BWP12T U1357 ( .A1(n2027), .A2(n671), .B1(n2025), .B2(n695), .ZN(n703) );
  XNR2D1BWP12T U1358 ( .A1(n1977), .A2(n3950), .ZN(n712) );
  OAI22D1BWP12T U1359 ( .A1(n2019), .A2(n672), .B1(n712), .B2(n2018), .ZN(n723) );
  XNR2XD8BWP12T U1360 ( .A1(n4060), .A2(n4078), .ZN(n2086) );
  INR2D1BWP12T U1361 ( .A1(n1979), .B1(n2086), .ZN(n722) );
  XNR2D1BWP12T U1362 ( .A1(n4068), .A2(n3932), .ZN(n701) );
  FA1D1BWP12T U1363 ( .A(n676), .B(n675), .CI(n674), .CO(n731), .S(n663) );
  XNR2D1BWP12T U1364 ( .A1(n4075), .A2(n3928), .ZN(n700) );
  OAI22D1BWP12T U1365 ( .A1(n2083), .A2(n677), .B1(n700), .B2(n2080), .ZN(n728) );
  XNR2D1BWP12T U1366 ( .A1(n4060), .A2(n3921), .ZN(n713) );
  XNR2D1BWP12T U1367 ( .A1(n4084), .A2(n3927), .ZN(n698) );
  OAI22D1BWP12T U1368 ( .A1(n2013), .A2(n679), .B1(n2011), .B2(n698), .ZN(n726) );
  OAI21D0BWP12T U1369 ( .A1(n682), .A2(n681), .B(n680), .ZN(n684) );
  CKND2D1BWP12T U1370 ( .A1(n682), .A2(n681), .ZN(n683) );
  ND2D1BWP12T U1371 ( .A1(n684), .A2(n683), .ZN(n729) );
  INVD1BWP12T U1372 ( .I(n729), .ZN(n685) );
  XNR3XD4BWP12T U1373 ( .A1(n731), .A2(n732), .A3(n685), .ZN(n743) );
  FA1D2BWP12T U1374 ( .A(n688), .B(n687), .CI(n686), .CO(n690), .S(n372) );
  OR2D2BWP12T U1375 ( .A1(n2367), .A2(n689), .Z(n693) );
  ND2D1BWP12T U1376 ( .A1(n691), .A2(n690), .ZN(n2368) );
  OA21D1BWP12T U1377 ( .A1(n2367), .A2(n2363), .B(n2368), .Z(n692) );
  TPOAI21D1BWP12T U1378 ( .A1(n694), .A2(n693), .B(n692), .ZN(n2890) );
  XNR2D1BWP12T U1379 ( .A1(n4063), .A2(n3920), .ZN(n709) );
  TPOAI22D1BWP12T U1380 ( .A1(n2027), .A2(n695), .B1(n1986), .B2(n709), .ZN(
        n716) );
  INVD15BWP12T U1381 ( .I(n989), .ZN(n2084) );
  XOR2D2BWP12T U1382 ( .A1(n2084), .A2(n4078), .Z(n696) );
  ND2D4BWP12T U1383 ( .A1(n2086), .A2(n696), .ZN(n2088) );
  XNR2D1BWP12T U1384 ( .A1(n1979), .A2(n2084), .ZN(n697) );
  XNR2D1BWP12T U1385 ( .A1(n1517), .A2(n2084), .ZN(n710) );
  XNR2D1BWP12T U1386 ( .A1(n4084), .A2(n3929), .ZN(n720) );
  OAI22D1BWP12T U1387 ( .A1(n2013), .A2(n698), .B1(n2011), .B2(n720), .ZN(n714) );
  IND2XD1BWP12T U1388 ( .A1(b[0]), .B1(n2084), .ZN(n699) );
  OAI22D1BWP12T U1389 ( .A1(n2088), .A2(n3875), .B1(n2086), .B2(n699), .ZN(
        n707) );
  XNR2D1BWP12T U1390 ( .A1(n4075), .A2(n3957), .ZN(n717) );
  XNR2D1BWP12T U1391 ( .A1(n3885), .A2(n3933), .ZN(n708) );
  OAI22D1BWP12T U1392 ( .A1(n2072), .A2(n701), .B1(n2070), .B2(n708), .ZN(n705) );
  FA1D1BWP12T U1393 ( .A(n704), .B(n703), .CI(n702), .CO(n736), .S(n744) );
  FA1D2BWP12T U1394 ( .A(n707), .B(n706), .CI(n705), .CO(n771), .S(n737) );
  XNR2D1BWP12T U1395 ( .A1(n1977), .A2(n3931), .ZN(n711) );
  XNR2D1BWP12T U1396 ( .A1(n1977), .A2(n3930), .ZN(n763) );
  OAI22D1BWP12T U1397 ( .A1(n2019), .A2(n711), .B1(n763), .B2(n2018), .ZN(n768) );
  XNR2XD8BWP12T U1398 ( .A1(a[14]), .A2(n2084), .ZN(n754) );
  INR2D1BWP12T U1399 ( .A1(n1979), .B1(n754), .ZN(n767) );
  XNR2D1BWP12T U1400 ( .A1(n4068), .A2(n3950), .ZN(n762) );
  OAI22D1BWP12T U1401 ( .A1(n2072), .A2(n708), .B1(n2070), .B2(n762), .ZN(n766) );
  XNR2D1BWP12T U1402 ( .A1(n4063), .A2(n3927), .ZN(n765) );
  TPOAI22D1BWP12T U1403 ( .A1(n2027), .A2(n709), .B1(n1986), .B2(n765), .ZN(
        n751) );
  XNR2XD1BWP12T U1404 ( .A1(n3921), .A2(n2084), .ZN(n752) );
  TPOAI22D1BWP12T U1405 ( .A1(n2088), .A2(n710), .B1(n2086), .B2(n752), .ZN(
        n750) );
  OAI22D1BWP12T U1406 ( .A1(n2019), .A2(n712), .B1(n711), .B2(n2018), .ZN(n725) );
  XNR2D1BWP12T U1407 ( .A1(n4060), .A2(n3922), .ZN(n719) );
  OAI22D1BWP12T U1408 ( .A1(n2009), .A2(n713), .B1(n719), .B2(n2006), .ZN(n724) );
  FA1D1BWP12T U1409 ( .A(n716), .B(n715), .CI(n714), .CO(n748), .S(n738) );
  XNR2D1BWP12T U1410 ( .A1(n4075), .A2(n3932), .ZN(n761) );
  OAI22D1BWP12T U1411 ( .A1(n2083), .A2(n717), .B1(n761), .B2(n2080), .ZN(n759) );
  XNR2D1BWP12T U1412 ( .A1(n4060), .A2(n718), .ZN(n764) );
  XNR2D1BWP12T U1413 ( .A1(n4084), .A2(n3928), .ZN(n756) );
  OAI22D1BWP12T U1414 ( .A1(n2013), .A2(n720), .B1(n2011), .B2(n756), .ZN(n757) );
  FA1D1BWP12T U1415 ( .A(n723), .B(n722), .CI(n721), .CO(n735), .S(n702) );
  FA1D2BWP12T U1416 ( .A(n728), .B(n727), .CI(n726), .CO(n733), .S(n732) );
  INVD1BWP12T U1417 ( .I(n2282), .ZN(n739) );
  OAI21D1BWP12T U1418 ( .A1(n731), .A2(n732), .B(n729), .ZN(n730) );
  IOA21D1BWP12T U1419 ( .A1(n732), .A2(n731), .B(n730), .ZN(n742) );
  FA1D1BWP12T U1420 ( .A(n735), .B(n734), .CI(n733), .CO(n746), .S(n741) );
  FA1D1BWP12T U1421 ( .A(n738), .B(n737), .CI(n736), .CO(n774), .S(n740) );
  TPND2D2BWP12T U1422 ( .A1(n739), .A2(n777), .ZN(n2284) );
  FA1D1BWP12T U1423 ( .A(n742), .B(n741), .CI(n740), .CO(n2281), .S(n776) );
  FA1D1BWP12T U1424 ( .A(n745), .B(n744), .CI(n743), .CO(n775), .S(n691) );
  NR2D1BWP12T U1425 ( .A1(n776), .A2(n775), .ZN(n2280) );
  INVD1BWP12T U1426 ( .I(n2280), .ZN(n2927) );
  CKND2D2BWP12T U1427 ( .A1(n2284), .A2(n2927), .ZN(n2889) );
  FA1D2BWP12T U1428 ( .A(n748), .B(n747), .CI(n746), .CO(n850), .S(n772) );
  FA1D1BWP12T U1429 ( .A(n751), .B(n750), .CI(n749), .CO(n805), .S(n769) );
  XNR2D1BWP12T U1430 ( .A1(n3922), .A2(n2084), .ZN(n816) );
  OAI22D1BWP12T U1431 ( .A1(n2088), .A2(n752), .B1(n2086), .B2(n816), .ZN(n811) );
  INVD12BWP12T U1432 ( .I(n3874), .ZN(n4082) );
  XNR2D1BWP12T U1433 ( .A1(n3873), .A2(n4082), .ZN(n753) );
  INVD8BWP12T U1434 ( .I(n4082), .ZN(n990) );
  IND2XD1BWP12T U1435 ( .A1(b[0]), .B1(n4082), .ZN(n755) );
  TPOAI22D1BWP12T U1436 ( .A1(n2130), .A2(n990), .B1(n754), .B2(n755), .ZN(
        n810) );
  XNR2D1BWP12T U1437 ( .A1(n4084), .A2(n3957), .ZN(n786) );
  OAI22D1BWP12T U1438 ( .A1(n2013), .A2(n756), .B1(n2011), .B2(n786), .ZN(n809) );
  FA1D0BWP12T U1439 ( .A(n759), .B(n758), .CI(n757), .CO(n803), .S(n747) );
  XNR2D1BWP12T U1440 ( .A1(n1979), .A2(n4082), .ZN(n760) );
  OAI22D1BWP12T U1441 ( .A1(n2130), .A2(n760), .B1(n754), .B2(n817), .ZN(n802)
         );
  XNR2D1BWP12T U1442 ( .A1(n4075), .A2(n3933), .ZN(n784) );
  OAI22D1BWP12T U1443 ( .A1(n2083), .A2(n761), .B1(n784), .B2(n2080), .ZN(n801) );
  XNR2D1BWP12T U1444 ( .A1(n4068), .A2(n3931), .ZN(n788) );
  OAI22D1BWP12T U1445 ( .A1(n2072), .A2(n762), .B1(n2070), .B2(n788), .ZN(n800) );
  XNR2D1BWP12T U1446 ( .A1(n1977), .A2(n3949), .ZN(n787) );
  OAI22D1BWP12T U1447 ( .A1(n2019), .A2(n763), .B1(n787), .B2(n2018), .ZN(n799) );
  XNR2D1BWP12T U1448 ( .A1(n4060), .A2(n3920), .ZN(n785) );
  OAI22D1BWP12T U1449 ( .A1(n2009), .A2(n764), .B1(n785), .B2(n2006), .ZN(n798) );
  XNR2D1BWP12T U1450 ( .A1(n4063), .A2(n3929), .ZN(n819) );
  OAI22D1BWP12T U1451 ( .A1(n2027), .A2(n765), .B1(n2025), .B2(n819), .ZN(n793) );
  FA1D2BWP12T U1452 ( .A(n771), .B(n770), .CI(n769), .CO(n833), .S(n773) );
  XOR3D2BWP12T U1453 ( .A1(n837), .A2(n838), .A3(n833), .Z(n848) );
  FA1D2BWP12T U1454 ( .A(n774), .B(n773), .CI(n772), .CO(n780), .S(n2282) );
  TPNR2D2BWP12T U1455 ( .A1(n781), .A2(n780), .ZN(n2893) );
  TPNR2D1BWP12T U1456 ( .A1(n2889), .A2(n2893), .ZN(n783) );
  CKND2D2BWP12T U1457 ( .A1(n776), .A2(n775), .ZN(n2926) );
  NR2D1BWP12T U1458 ( .A1(n2926), .A2(n777), .ZN(n779) );
  ND2D1BWP12T U1459 ( .A1(n2926), .A2(n777), .ZN(n778) );
  OAI21D1BWP12T U1460 ( .A1(n779), .A2(n2282), .B(n778), .ZN(n2891) );
  ND2D1BWP12T U1461 ( .A1(n781), .A2(n780), .ZN(n2894) );
  TPOAI21D1BWP12T U1462 ( .A1(n2891), .A2(n2893), .B(n2894), .ZN(n782) );
  TPAOI21D2BWP12T U1463 ( .A1(n2890), .A2(n783), .B(n782), .ZN(n3430) );
  XNR2D1BWP12T U1464 ( .A1(n4075), .A2(n3950), .ZN(n830) );
  OAI22D1BWP12T U1465 ( .A1(n2083), .A2(n784), .B1(n830), .B2(n2080), .ZN(n814) );
  XNR2D1BWP12T U1466 ( .A1(n4060), .A2(n3927), .ZN(n826) );
  OAI22D1BWP12T U1467 ( .A1(n2009), .A2(n785), .B1(n826), .B2(n2006), .ZN(n813) );
  XNR2D1BWP12T U1468 ( .A1(n4084), .A2(n3932), .ZN(n831) );
  OAI22D1BWP12T U1469 ( .A1(n2013), .A2(n786), .B1(n2011), .B2(n831), .ZN(n812) );
  XNR2D1BWP12T U1470 ( .A1(n1977), .A2(n4191), .ZN(n789) );
  XOR2XD8BWP12T U1471 ( .A1(n990), .A2(n4183), .Z(n2059) );
  INVD1BWP12T U1472 ( .I(n1979), .ZN(n1593) );
  NR2D1BWP12T U1473 ( .A1(n2059), .A2(n1593), .ZN(n796) );
  XNR2D1BWP12T U1474 ( .A1(n4068), .A2(n3930), .ZN(n828) );
  XNR2D1BWP12T U1475 ( .A1(n4063), .A2(n3928), .ZN(n818) );
  XNR2D1BWP12T U1476 ( .A1(n4063), .A2(n3957), .ZN(n869) );
  TPOAI22D1BWP12T U1477 ( .A1(n2027), .A2(n818), .B1(n2025), .B2(n869), .ZN(
        n884) );
  XNR2XD1BWP12T U1478 ( .A1(n2098), .A2(n2084), .ZN(n815) );
  XNR2D1BWP12T U1479 ( .A1(n2084), .A2(n3920), .ZN(n887) );
  OAI22D1BWP12T U1480 ( .A1(n2088), .A2(n815), .B1(n2086), .B2(n887), .ZN(n883) );
  XNR2D1BWP12T U1481 ( .A1(n1977), .A2(n3952), .ZN(n888) );
  OAI22D1BWP12T U1482 ( .A1(n2019), .A2(n789), .B1(n888), .B2(n2018), .ZN(n886) );
  INVD8BWP12T U1483 ( .I(a[17]), .ZN(n1339) );
  XNR2XD2BWP12T U1484 ( .A1(n1339), .A2(n4183), .ZN(n790) );
  TPND2D3BWP12T U1485 ( .A1(n2059), .A2(n790), .ZN(n2062) );
  BUFFXD12BWP12T U1486 ( .I(n2059), .Z(n1648) );
  INVD8BWP12T U1487 ( .I(n1339), .ZN(n2058) );
  IND2XD1BWP12T U1488 ( .A1(b[0]), .B1(n2058), .ZN(n791) );
  TPOAI22D1BWP12T U1489 ( .A1(n2062), .A2(n1339), .B1(n1648), .B2(n791), .ZN(
        n885) );
  INVD1BWP12T U1490 ( .I(n892), .ZN(n832) );
  FA1D2BWP12T U1491 ( .A(n794), .B(n793), .CI(n792), .CO(n844), .S(n838) );
  FA1D2BWP12T U1492 ( .A(n797), .B(n796), .CI(n795), .CO(n877), .S(n808) );
  HA1D1BWP12T U1493 ( .A(n799), .B(n798), .CO(n807), .S(n794) );
  FA1D2BWP12T U1494 ( .A(n802), .B(n801), .CI(n800), .CO(n806), .S(n837) );
  FA1D1BWP12T U1495 ( .A(n805), .B(n804), .CI(n803), .CO(n842), .S(n849) );
  FA1D1BWP12T U1496 ( .A(n808), .B(n807), .CI(n806), .CO(n857), .S(n843) );
  FA1D1BWP12T U1497 ( .A(n811), .B(n810), .CI(n809), .CO(n840), .S(n804) );
  FA1D1BWP12T U1498 ( .A(n814), .B(n813), .CI(n812), .CO(n878), .S(n841) );
  NR2D1BWP12T U1499 ( .A1(n840), .A2(n841), .ZN(n822) );
  XNR2XD1BWP12T U1500 ( .A1(n3921), .A2(n4082), .ZN(n829) );
  OAI22D1BWP12T U1501 ( .A1(n2027), .A2(n819), .B1(n2025), .B2(n818), .ZN(n823) );
  INVD1BWP12T U1502 ( .I(n839), .ZN(n821) );
  CKND2D1BWP12T U1503 ( .A1(n840), .A2(n841), .ZN(n820) );
  OAI21D1BWP12T U1504 ( .A1(n822), .A2(n821), .B(n820), .ZN(n858) );
  FA1D2BWP12T U1505 ( .A(n825), .B(n824), .CI(n823), .CO(n870), .S(n839) );
  XNR2D1BWP12T U1506 ( .A1(n4060), .A2(n3929), .ZN(n861) );
  OAI22D1BWP12T U1507 ( .A1(n2009), .A2(n826), .B1(n861), .B2(n2006), .ZN(n866) );
  BUFFXD4BWP12T U1508 ( .I(n2062), .Z(n1650) );
  XNR2D1BWP12T U1509 ( .A1(n2058), .A2(n1979), .ZN(n827) );
  XNR2D1BWP12T U1510 ( .A1(n2058), .A2(n1517), .ZN(n862) );
  TPOAI22D1BWP12T U1511 ( .A1(n1650), .A2(n827), .B1(n862), .B2(n1648), .ZN(
        n865) );
  XNR2D0BWP12T U1512 ( .A1(n4068), .A2(n3949), .ZN(n889) );
  OAI22D1BWP12T U1513 ( .A1(n2072), .A2(n828), .B1(n2070), .B2(n889), .ZN(n864) );
  XNR2D1BWP12T U1514 ( .A1(n1189), .A2(n4082), .ZN(n867) );
  XNR2XD1BWP12T U1515 ( .A1(n4075), .A2(n3931), .ZN(n868) );
  OAI22D1BWP12T U1516 ( .A1(n2083), .A2(n830), .B1(n868), .B2(n2080), .ZN(n880) );
  XNR2D1BWP12T U1517 ( .A1(n4084), .A2(n3933), .ZN(n863) );
  OAI22D1BWP12T U1518 ( .A1(n2013), .A2(n831), .B1(n2011), .B2(n863), .ZN(n879) );
  XOR3D2BWP12T U1519 ( .A1(n870), .A2(n872), .A3(n871), .Z(n856) );
  XOR3D2BWP12T U1520 ( .A1(n857), .A2(n858), .A3(n856), .Z(n890) );
  XNR3XD4BWP12T U1521 ( .A1(n832), .A2(n893), .A3(n890), .ZN(n3180) );
  INVD1BWP12T U1522 ( .I(n838), .ZN(n835) );
  INVD1BWP12T U1523 ( .I(n837), .ZN(n834) );
  IOA21D1BWP12T U1524 ( .A1(n835), .A2(n834), .B(n833), .ZN(n836) );
  IOA21D1BWP12T U1525 ( .A1(n838), .A2(n837), .B(n836), .ZN(n847) );
  FA1D1BWP12T U1526 ( .A(n844), .B(n843), .CI(n842), .CO(n893), .S(n845) );
  OR2XD4BWP12T U1527 ( .A1(n3180), .A2(n3179), .Z(n3182) );
  FA1D1BWP12T U1528 ( .A(n847), .B(n846), .CI(n845), .CO(n3179), .S(n852) );
  FA1D1BWP12T U1529 ( .A(n850), .B(n849), .CI(n848), .CO(n851), .S(n781) );
  OR2D2BWP12T U1530 ( .A1(n852), .A2(n851), .Z(n3428) );
  ND2D1BWP12T U1531 ( .A1(n3182), .A2(n3428), .ZN(n855) );
  ND2D1BWP12T U1532 ( .A1(n852), .A2(n851), .ZN(n3427) );
  INVD1BWP12T U1533 ( .I(n3427), .ZN(n3177) );
  AN2XD2BWP12T U1534 ( .A1(n3180), .A2(n3179), .Z(n853) );
  TPAOI21D2BWP12T U1535 ( .A1(n3182), .A2(n3177), .B(n853), .ZN(n854) );
  TPOAI21D2BWP12T U1536 ( .A1(n3430), .A2(n855), .B(n854), .ZN(n3134) );
  OAI21D1BWP12T U1537 ( .A1(n857), .A2(n858), .B(n856), .ZN(n860) );
  CKND2D1BWP12T U1538 ( .A1(n858), .A2(n857), .ZN(n859) );
  ND2D1BWP12T U1539 ( .A1(n860), .A2(n859), .ZN(n1420) );
  XNR2D1BWP12T U1540 ( .A1(n4060), .A2(n3928), .ZN(n1292) );
  OAI22D1BWP12T U1541 ( .A1(n2009), .A2(n861), .B1(n1292), .B2(n2006), .ZN(
        n1389) );
  XNR2D1BWP12T U1542 ( .A1(n2058), .A2(n3921), .ZN(n1284) );
  TPOAI22D1BWP12T U1543 ( .A1(n1650), .A2(n862), .B1(n1284), .B2(n1648), .ZN(
        n1388) );
  XNR2D1BWP12T U1544 ( .A1(n4084), .A2(n3950), .ZN(n1316) );
  OAI22D1BWP12T U1545 ( .A1(n2013), .A2(n863), .B1(n2011), .B2(n1316), .ZN(
        n1387) );
  FA1D2BWP12T U1546 ( .A(n866), .B(n865), .CI(n864), .CO(n1415), .S(n872) );
  XNR2XD1BWP12T U1547 ( .A1(n2098), .A2(n4082), .ZN(n1411) );
  OAI22D1BWP12T U1548 ( .A1(n2130), .A2(n867), .B1(n754), .B2(n1411), .ZN(
        n1407) );
  XNR2D1BWP12T U1549 ( .A1(n4075), .A2(n3930), .ZN(n1294) );
  OAI22D1BWP12T U1550 ( .A1(n2083), .A2(n868), .B1(n1294), .B2(n2080), .ZN(
        n1406) );
  XNR2XD1BWP12T U1551 ( .A1(n506), .A2(n3932), .ZN(n1413) );
  OAI22D1BWP12T U1552 ( .A1(n2027), .A2(n869), .B1(n1986), .B2(n1413), .ZN(
        n1405) );
  ND2D1BWP12T U1553 ( .A1(n870), .A2(n872), .ZN(n875) );
  ND2D1BWP12T U1554 ( .A1(n870), .A2(n871), .ZN(n874) );
  ND2D1BWP12T U1555 ( .A1(n872), .A2(n871), .ZN(n873) );
  ND3D1BWP12T U1556 ( .A1(n875), .A2(n874), .A3(n873), .ZN(n1392) );
  FA1D2BWP12T U1557 ( .A(n878), .B(n877), .CI(n876), .CO(n1391), .S(n892) );
  FA1D1BWP12T U1558 ( .A(n881), .B(n880), .CI(n879), .CO(n1399), .S(n871) );
  FA1D1BWP12T U1559 ( .A(n884), .B(n883), .CI(n882), .CO(n1400), .S(n876) );
  HA1D1BWP12T U1560 ( .A(n886), .B(n885), .CO(n1378), .S(n882) );
  XNR2D1BWP12T U1561 ( .A1(n2084), .A2(n3927), .ZN(n1409) );
  OAI22D1BWP12T U1562 ( .A1(n2088), .A2(n887), .B1(n2086), .B2(n1409), .ZN(
        n1377) );
  XNR2D1BWP12T U1563 ( .A1(n1977), .A2(n3951), .ZN(n1282) );
  XNR2XD8BWP12T U1564 ( .A1(n2058), .A2(n3820), .ZN(n2125) );
  INR2D1BWP12T U1565 ( .A1(n1979), .B1(n2125), .ZN(n1383) );
  XNR2D1BWP12T U1566 ( .A1(n3885), .A2(n4191), .ZN(n1296) );
  OAI22D1BWP12T U1567 ( .A1(n2072), .A2(n889), .B1(n2070), .B2(n1296), .ZN(
        n1382) );
  XOR3D1BWP12T U1568 ( .A1(n1399), .A2(n1400), .A3(n1395), .Z(n1390) );
  XOR3D2BWP12T U1569 ( .A1(n1392), .A2(n1391), .A3(n1390), .Z(n1418) );
  OAI21D1BWP12T U1570 ( .A1(n892), .A2(n893), .B(n890), .ZN(n891) );
  IOA21D1BWP12T U1571 ( .A1(n893), .A2(n892), .B(n891), .ZN(n894) );
  CKND2D2BWP12T U1572 ( .A1(n895), .A2(n894), .ZN(n1449) );
  AN2XD1BWP12T U1573 ( .A1(n317), .A2(n1449), .Z(n896) );
  INVD1BWP12T U1574 ( .I(n3435), .ZN(n1000) );
  BUFFXD0BWP12T U1575 ( .I(a[13]), .Z(n905) );
  ND2D1BWP12T U1576 ( .A1(n2932), .A2(n2291), .ZN(n3509) );
  CKBD1BWP12T U1577 ( .I(n4082), .Z(n907) );
  NR2D1BWP12T U1578 ( .A1(n3828), .A2(n907), .ZN(n3512) );
  INVD1BWP12T U1579 ( .I(n3512), .ZN(n2902) );
  OR2XD1BWP12T U1580 ( .A1(n3821), .A2(n4183), .Z(n3521) );
  ND2D1BWP12T U1581 ( .A1(n2902), .A2(n3521), .ZN(n910) );
  NR2D1BWP12T U1582 ( .A1(n3509), .A2(n910), .ZN(n3186) );
  INVD1BWP12T U1583 ( .I(n3186), .ZN(n3140) );
  CKBD1BWP12T U1584 ( .I(a[17]), .Z(n911) );
  NR2D1BWP12T U1585 ( .A1(n3826), .A2(n911), .ZN(n1708) );
  ND2D1BWP12T U1586 ( .A1(n316), .A2(n2376), .ZN(n901) );
  NR2D1BWP12T U1587 ( .A1(n901), .A2(n3335), .ZN(n904) );
  ND2D1BWP12T U1588 ( .A1(n904), .A2(n897), .ZN(n2930) );
  INVD1BWP12T U1589 ( .I(n2930), .ZN(n3510) );
  INVD1BWP12T U1590 ( .I(n898), .ZN(n2373) );
  CKND2D1BWP12T U1591 ( .A1(n3829), .A2(n4078), .ZN(n2375) );
  INVD1BWP12T U1592 ( .I(n2375), .ZN(n899) );
  AOI21D1BWP12T U1593 ( .A1(n2376), .A2(n2373), .B(n899), .ZN(n900) );
  OAI21D1BWP12T U1594 ( .A1(n901), .A2(n3336), .B(n900), .ZN(n902) );
  AOI21D1BWP12T U1595 ( .A1(n904), .A2(n903), .B(n902), .ZN(n2929) );
  INVD1BWP12T U1596 ( .I(n2929), .ZN(n3516) );
  ND2D1BWP12T U1597 ( .A1(n3830), .A2(n905), .ZN(n2931) );
  INVD1BWP12T U1598 ( .I(n2931), .ZN(n2287) );
  CKND2D1BWP12T U1599 ( .A1(n3827), .A2(a[14]), .ZN(n2290) );
  INVD1BWP12T U1600 ( .I(n2290), .ZN(n906) );
  AOI21D1BWP12T U1601 ( .A1(n2291), .A2(n2287), .B(n906), .ZN(n3513) );
  ND2D1BWP12T U1602 ( .A1(n3828), .A2(n907), .ZN(n3511) );
  ND2D1BWP12T U1603 ( .A1(n3821), .A2(n4183), .ZN(n3520) );
  INVD1BWP12T U1604 ( .I(n3520), .ZN(n908) );
  AOI21D1BWP12T U1605 ( .A1(n3521), .A2(n922), .B(n908), .ZN(n909) );
  OAI21D1BWP12T U1606 ( .A1(n3513), .A2(n910), .B(n909), .ZN(n3185) );
  INVD1BWP12T U1607 ( .I(n3185), .ZN(n3143) );
  ND2D1BWP12T U1608 ( .A1(n3826), .A2(n911), .ZN(n3189) );
  CKND2D1BWP12T U1609 ( .A1(n3819), .A2(n3820), .ZN(n1709) );
  NR2D1BWP12T U1610 ( .A1(n3829), .A2(n4078), .ZN(n2378) );
  NR2D1BWP12T U1611 ( .A1(n912), .A2(n2378), .ZN(n2937) );
  CKBD1BWP12T U1612 ( .I(a[13]), .Z(n913) );
  NR2D1BWP12T U1613 ( .A1(n3830), .A2(n913), .ZN(n2939) );
  NR2D1BWP12T U1614 ( .A1(n3827), .A2(a[14]), .ZN(n2353) );
  NR2D1BWP12T U1615 ( .A1(n2939), .A2(n2353), .ZN(n915) );
  ND2D1BWP12T U1616 ( .A1(n2937), .A2(n915), .ZN(n917) );
  NR2D1BWP12T U1617 ( .A1(n2346), .A2(n917), .ZN(n919) );
  CKND2D1BWP12T U1618 ( .A1(n3829), .A2(n4078), .ZN(n2379) );
  OAI21D1BWP12T U1619 ( .A1(n2378), .A2(n2377), .B(n2379), .ZN(n2936) );
  ND2D1BWP12T U1620 ( .A1(n3830), .A2(n913), .ZN(n2940) );
  CKND2D1BWP12T U1621 ( .A1(n3827), .A2(a[14]), .ZN(n2354) );
  OAI21D1BWP12T U1622 ( .A1(n2353), .A2(n2940), .B(n2354), .ZN(n914) );
  AOI21D1BWP12T U1623 ( .A1(n915), .A2(n2936), .B(n914), .ZN(n916) );
  OAI21D1BWP12T U1624 ( .A1(n2347), .A2(n917), .B(n916), .ZN(n918) );
  AOI21D1BWP12T U1625 ( .A1(n920), .A2(n919), .B(n918), .ZN(n3487) );
  CKBD1BWP12T U1626 ( .I(n4082), .Z(n921) );
  NR2D1BWP12T U1627 ( .A1(n3828), .A2(n921), .ZN(n3486) );
  OR2XD1BWP12T U1628 ( .A1(n3821), .A2(n4183), .Z(n3489) );
  ND2D1BWP12T U1629 ( .A1(n2902), .A2(n3489), .ZN(n3193) );
  CKBD1BWP12T U1630 ( .I(a[17]), .Z(n923) );
  NR2D1BWP12T U1631 ( .A1(n3826), .A2(n923), .ZN(n3197) );
  NR2D0BWP12T U1632 ( .A1(n3193), .A2(n3197), .ZN(n925) );
  ND2D1BWP12T U1633 ( .A1(n3828), .A2(n921), .ZN(n3485) );
  INVD0BWP12T U1634 ( .I(n3485), .ZN(n922) );
  ND2D1BWP12T U1635 ( .A1(n3821), .A2(n4183), .ZN(n3488) );
  AOI21D1BWP12T U1636 ( .A1(n3489), .A2(n922), .B(n908), .ZN(n3194) );
  ND2D1BWP12T U1637 ( .A1(n3826), .A2(n923), .ZN(n3198) );
  TPOAI21D0BWP12T U1638 ( .A1(n3194), .A2(n3197), .B(n3198), .ZN(n924) );
  AOI21D1BWP12T U1639 ( .A1(n3276), .A2(n925), .B(n924), .ZN(n927) );
  NR2D1BWP12T U1640 ( .A1(n3819), .A2(a[18]), .ZN(n1696) );
  ND2D1BWP12T U1641 ( .A1(n3819), .A2(a[18]), .ZN(n1695) );
  ND2D1BWP12T U1642 ( .A1(n1712), .A2(n1695), .ZN(n926) );
  XOR2XD1BWP12T U1643 ( .A1(n927), .A2(n926), .Z(n3469) );
  NR2D1BWP12T U1644 ( .A1(n930), .A2(n928), .ZN(n932) );
  ND2D1BWP12T U1645 ( .A1(n3386), .A2(n932), .ZN(n2401) );
  CKBD1BWP12T U1646 ( .I(a[13]), .Z(n933) );
  NR2D1BWP12T U1647 ( .A1(n933), .A2(n3931), .ZN(n2965) );
  NR2D1BWP12T U1648 ( .A1(n3950), .A2(n4078), .ZN(n2385) );
  NR2D1BWP12T U1649 ( .A1(n2965), .A2(n2385), .ZN(n2907) );
  CKBD1BWP12T U1650 ( .I(n4082), .Z(n934) );
  NR2D1BWP12T U1651 ( .A1(n934), .A2(n3949), .ZN(n2911) );
  NR2D1BWP12T U1652 ( .A1(n2911), .A2(n2910), .ZN(n936) );
  ND2D1BWP12T U1653 ( .A1(n2907), .A2(n936), .ZN(n938) );
  NR2D1BWP12T U1654 ( .A1(n2401), .A2(n938), .ZN(n940) );
  OAI21D1BWP12T U1655 ( .A1(n930), .A2(n3389), .B(n929), .ZN(n931) );
  AOI21D1BWP12T U1656 ( .A1(n932), .A2(n3387), .B(n931), .ZN(n2400) );
  ND2D1BWP12T U1657 ( .A1(n3950), .A2(n4078), .ZN(n2959) );
  CKND2D1BWP12T U1658 ( .A1(n933), .A2(n3931), .ZN(n2966) );
  OAI21D1BWP12T U1659 ( .A1(n2965), .A2(n2959), .B(n2966), .ZN(n2908) );
  ND2D1BWP12T U1660 ( .A1(n3930), .A2(a[14]), .ZN(n2909) );
  CKND2D1BWP12T U1661 ( .A1(n934), .A2(n3949), .ZN(n2912) );
  TPOAI21D0BWP12T U1662 ( .A1(n2911), .A2(n2909), .B(n2912), .ZN(n935) );
  TPAOI21D0BWP12T U1663 ( .A1(n936), .A2(n2908), .B(n935), .ZN(n937) );
  OAI21D1BWP12T U1664 ( .A1(n2400), .A2(n938), .B(n937), .ZN(n939) );
  TPAOI21D2BWP12T U1665 ( .A1(n941), .A2(n940), .B(n939), .ZN(n3579) );
  BUFFD1BWP12T U1666 ( .I(a[17]), .Z(n942) );
  OR2XD1BWP12T U1667 ( .A1(n942), .A2(n3952), .Z(n3203) );
  NR2D1BWP12T U1668 ( .A1(n4191), .A2(n4183), .ZN(n3201) );
  ND2D1BWP12T U1669 ( .A1(n3203), .A2(n4121), .ZN(n3157) );
  ND2D1BWP12T U1670 ( .A1(n4191), .A2(n4183), .ZN(n4120) );
  INVD1BWP12T U1671 ( .I(n4120), .ZN(n954) );
  CKND2D1BWP12T U1672 ( .A1(n942), .A2(n3952), .ZN(n3202) );
  INVD1BWP12T U1673 ( .I(n3202), .ZN(n943) );
  AOI21D1BWP12T U1674 ( .A1(n3203), .A2(n954), .B(n943), .ZN(n3158) );
  NR2D1BWP12T U1675 ( .A1(n3951), .A2(n3820), .ZN(n1737) );
  INVD1BWP12T U1676 ( .I(n1737), .ZN(n3160) );
  ND2D1BWP12T U1677 ( .A1(n3951), .A2(n3820), .ZN(n3159) );
  NR2D1BWP12T U1678 ( .A1(n944), .A2(n2385), .ZN(n2943) );
  CKBD1BWP12T U1679 ( .I(a[13]), .Z(n945) );
  NR2D1BWP12T U1680 ( .A1(n945), .A2(n3931), .ZN(n2945) );
  NR2D1BWP12T U1681 ( .A1(n2945), .A2(n2910), .ZN(n947) );
  ND2D1BWP12T U1682 ( .A1(n2943), .A2(n947), .ZN(n949) );
  NR2D1BWP12T U1683 ( .A1(n2318), .A2(n949), .ZN(n951) );
  OAI21D1BWP12T U1684 ( .A1(n2385), .A2(n2380), .B(n2959), .ZN(n2942) );
  CKND2D1BWP12T U1685 ( .A1(n945), .A2(n3931), .ZN(n2946) );
  OAI21D1BWP12T U1686 ( .A1(n2910), .A2(n2946), .B(n2909), .ZN(n946) );
  TPAOI21D0BWP12T U1687 ( .A1(n947), .A2(n2942), .B(n946), .ZN(n948) );
  OAI21D1BWP12T U1688 ( .A1(n2319), .A2(n949), .B(n948), .ZN(n950) );
  AOI21D1BWP12T U1689 ( .A1(n952), .A2(n951), .B(n950), .ZN(n4119) );
  INVD1P75BWP12T U1690 ( .I(n4119), .ZN(n3321) );
  CKBD1BWP12T U1691 ( .I(n4082), .Z(n953) );
  NR2D1BWP12T U1692 ( .A1(n953), .A2(n3949), .ZN(n4118) );
  INVD1BWP12T U1693 ( .I(n4118), .ZN(n2905) );
  OR2XD1BWP12T U1694 ( .A1(n4191), .A2(n4183), .Z(n4121) );
  ND2D1BWP12T U1695 ( .A1(n2905), .A2(n4121), .ZN(n3206) );
  CKBD1BWP12T U1696 ( .I(a[17]), .Z(n956) );
  NR2D1BWP12T U1697 ( .A1(n956), .A2(n3952), .ZN(n3210) );
  NR2D0BWP12T U1698 ( .A1(n3206), .A2(n3210), .ZN(n958) );
  CKND2D1BWP12T U1699 ( .A1(n953), .A2(n3949), .ZN(n4117) );
  INVD1BWP12T U1700 ( .I(n4117), .ZN(n955) );
  AOI21D1BWP12T U1701 ( .A1(n4121), .A2(n955), .B(n954), .ZN(n3207) );
  ND2D1BWP12T U1702 ( .A1(n956), .A2(n3952), .ZN(n3211) );
  TPOAI21D0BWP12T U1703 ( .A1(n3207), .A2(n3210), .B(n3211), .ZN(n957) );
  AOI21D1BWP12T U1704 ( .A1(n3321), .A2(n958), .B(n957), .ZN(n960) );
  CKND2D1BWP12T U1705 ( .A1(n3160), .A2(n3159), .ZN(n959) );
  XOR2XD1BWP12T U1706 ( .A1(n960), .A2(n959), .Z(n4101) );
  INVD1BWP12T U1707 ( .I(n2948), .ZN(n1072) );
  CKND2D1BWP12T U1708 ( .A1(n961), .A2(n1072), .ZN(n963) );
  MUX2D1BWP12T U1709 ( .I0(n2301), .I1(n962), .S(n3921), .Z(n3352) );
  CKND2D1BWP12T U1710 ( .A1(n3352), .A2(n4044), .ZN(n978) );
  INR2D1BWP12T U1711 ( .A1(n963), .B1(n979), .ZN(n2649) );
  INVD1BWP12T U1712 ( .I(n2649), .ZN(n964) );
  INVD0BWP12T U1713 ( .I(n4036), .ZN(n4013) );
  ND2D1BWP12T U1714 ( .A1(n3765), .A2(n4089), .ZN(n2920) );
  OA21D1BWP12T U1715 ( .A1(n964), .A2(n4013), .B(n2920), .Z(n4041) );
  INVD1BWP12T U1716 ( .I(n4011), .ZN(n3029) );
  INVD1BWP12T U1717 ( .I(n2304), .ZN(n3679) );
  MUX2D1BWP12T U1718 ( .I0(n3679), .I1(n965), .S(n3886), .Z(n3018) );
  OR2XD1BWP12T U1719 ( .A1(b[3]), .A2(n3919), .Z(n3767) );
  OAI21D0BWP12T U1720 ( .A1(n3018), .A2(n3919), .B(n3767), .ZN(n977) );
  CKND2D0BWP12T U1721 ( .A1(n967), .A2(n966), .ZN(n969) );
  INVD1BWP12T U1722 ( .I(n983), .ZN(n968) );
  AOI21D1BWP12T U1723 ( .A1(n3005), .A2(n969), .B(n968), .ZN(n2654) );
  INVD1BWP12T U1724 ( .I(n2654), .ZN(n3004) );
  MUX2XD0BWP12T U1725 ( .I0(n3880), .I1(n3891), .S(b[0]), .Z(n2333) );
  INVD1BWP12T U1726 ( .I(n2333), .ZN(n2294) );
  MUX2XD0BWP12T U1727 ( .I0(n3877), .I1(n3879), .S(b[0]), .Z(n2330) );
  INVD1BWP12T U1728 ( .I(n2330), .ZN(n2255) );
  OAI22D1BWP12T U1729 ( .A1(n2294), .A2(n970), .B1(n3005), .B2(n2255), .ZN(
        n972) );
  OAI22D1BWP12T U1730 ( .A1(n3703), .A2(n1838), .B1(n1833), .B2(n3705), .ZN(
        n971) );
  NR2D1BWP12T U1731 ( .A1(n972), .A2(n971), .ZN(n3003) );
  MUX2XD0BWP12T U1732 ( .I0(n3820), .I1(a[17]), .S(b[0]), .Z(n2258) );
  INVD1BWP12T U1733 ( .I(n2258), .ZN(n2772) );
  MUX2XD0BWP12T U1734 ( .I0(a[14]), .I1(a[13]), .S(b[0]), .Z(n2296) );
  TPNR2D0BWP12T U1735 ( .A1(n3703), .A2(n2296), .ZN(n974) );
  MUX2XD0BWP12T U1736 ( .I0(n3876), .I1(n3878), .S(b[0]), .Z(n2332) );
  INVD1BWP12T U1737 ( .I(n2332), .ZN(n2295) );
  INVD1P75BWP12T U1738 ( .I(n3227), .ZN(n3704) );
  MUX2XD0BWP12T U1739 ( .I0(n4187), .I1(n3874), .S(b[0]), .Z(n2775) );
  INVD1BWP12T U1740 ( .I(n2775), .ZN(n2756) );
  TPOAI22D0BWP12T U1741 ( .A1(n3705), .A2(n2295), .B1(n3704), .B2(n2756), .ZN(
        n973) );
  AOI211D1BWP12T U1742 ( .A1(n3707), .A2(n2772), .B(n974), .C(n973), .ZN(n3007) );
  INVD2BWP12T U1743 ( .I(n4179), .ZN(n3711) );
  OAI22D0BWP12T U1744 ( .A1(n3003), .A2(n2547), .B1(n3007), .B2(n3711), .ZN(
        n975) );
  ND2D1BWP12T U1745 ( .A1(n3300), .A2(n3170), .ZN(n2760) );
  NR2D1BWP12T U1746 ( .A1(n2629), .A2(n3767), .ZN(n2771) );
  INVD1BWP12T U1747 ( .I(n2771), .ZN(n3710) );
  ND2D1BWP12T U1748 ( .A1(n2760), .A2(n3710), .ZN(n3298) );
  AOI211D0BWP12T U1749 ( .A1(n3170), .A2(n3004), .B(n975), .C(n3298), .ZN(n976) );
  AOI21D1BWP12T U1750 ( .A1(n978), .A2(n977), .B(n976), .ZN(n3744) );
  TPND2D0BWP12T U1751 ( .A1(n3679), .A2(n1072), .ZN(n980) );
  INR2D1BWP12T U1752 ( .A1(n980), .B1(n979), .ZN(n3992) );
  NR2D1BWP12T U1753 ( .A1(n3765), .A2(n2834), .ZN(n3019) );
  OAI21D0BWP12T U1754 ( .A1(n981), .A2(n3921), .B(n3780), .ZN(n982) );
  ND2D1BWP12T U1755 ( .A1(n983), .A2(n982), .ZN(n3010) );
  NR2D0BWP12T U1756 ( .A1(n3010), .A2(b[3]), .ZN(n3774) );
  INVD1BWP12T U1757 ( .I(n3786), .ZN(n3245) );
  INVD1BWP12T U1758 ( .I(n1833), .ZN(n1827) );
  CKND0BWP12T U1759 ( .I(n1838), .ZN(n984) );
  AOI22D1BWP12T U1760 ( .A1(n3245), .A2(n1827), .B1(n984), .B2(n3242), .ZN(
        n986) );
  AOI22D0BWP12T U1761 ( .A1(n3241), .A2(n2330), .B1(n2333), .B2(n3238), .ZN(
        n985) );
  ND2D1BWP12T U1762 ( .A1(n986), .A2(n985), .ZN(n3011) );
  NR2D1BWP12T U1763 ( .A1(n4044), .A2(n3919), .ZN(n3249) );
  INVD1BWP12T U1764 ( .I(n2296), .ZN(n2331) );
  INVD1BWP12T U1765 ( .I(n3242), .ZN(n3784) );
  OAI22D0BWP12T U1766 ( .A1(n3786), .A2(n2332), .B1(n2331), .B2(n3784), .ZN(
        n3012) );
  AOI22D0BWP12T U1767 ( .A1(n3241), .A2(n2258), .B1(n2756), .B2(n3238), .ZN(
        n3013) );
  ND2D1BWP12T U1768 ( .A1(n987), .A2(n3877), .ZN(n988) );
  NR2D1BWP12T U1769 ( .A1(n3350), .A2(n988), .ZN(n2391) );
  ND2D1BWP12T U1770 ( .A1(n989), .A2(n3876), .ZN(n2917) );
  ND2D1BWP12T U1771 ( .A1(n990), .A2(n3873), .ZN(n991) );
  NR2D1BWP12T U1772 ( .A1(n2917), .A2(n991), .ZN(n992) );
  ND2D1BWP12T U1773 ( .A1(n2391), .A2(n992), .ZN(n994) );
  NR2D1BWP12T U1774 ( .A1(n994), .A2(n993), .ZN(n3293) );
  ND2D1BWP12T U1775 ( .A1(n1339), .A2(n4187), .ZN(n3172) );
  MUX2ND0BWP12T U1776 ( .I0(n4184), .I1(n2664), .S(n3951), .ZN(n995) );
  NR2XD0BWP12T U1777 ( .A1(n995), .A2(n4185), .ZN(n996) );
  MUX2ND0BWP12T U1778 ( .I0(n996), .I1(n2205), .S(n3867), .ZN(n997) );
  AOI21D1BWP12T U1779 ( .A1(n3526), .A2(n4215), .B(n998), .ZN(n999) );
  OAI21D4BWP12T U1780 ( .A1(n1000), .A2(n3407), .B(n999), .ZN(result[18]) );
  CKND2D1BWP12T U1781 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  CKND2D1BWP12T U1782 ( .A1(n3415), .A2(n4171), .ZN(n1055) );
  MUX2NXD0BWP12T U1783 ( .I0(n2519), .I1(n1005), .S(n3921), .ZN(n2918) );
  CKND2D1BWP12T U1784 ( .A1(n2918), .A2(n4044), .ZN(n3066) );
  CKND1BWP12T U1785 ( .I(n2629), .ZN(n2582) );
  INVD1BWP12T U1786 ( .I(n2970), .ZN(n3027) );
  CKND2D0BWP12T U1787 ( .A1(n1047), .A2(n3986), .ZN(n1008) );
  MUX2NXD0BWP12T U1788 ( .I0(n2524), .I1(n2520), .S(n3921), .ZN(n2919) );
  OAI22D1BWP12T U1789 ( .A1(n2469), .A2(n3891), .B1(n2468), .B2(n3877), .ZN(
        n1007) );
  OAI22D1BWP12T U1790 ( .A1(n2471), .A2(n3879), .B1(n2470), .B2(n3880), .ZN(
        n1006) );
  NR2D1BWP12T U1791 ( .A1(n1007), .A2(n1006), .ZN(n2526) );
  AOI21D0BWP12T U1792 ( .A1(n1008), .A2(n3765), .B(n3726), .ZN(n3985) );
  CKND2D0BWP12T U1793 ( .A1(n1040), .A2(n1057), .ZN(n1009) );
  XOR2XD1BWP12T U1794 ( .A1(n3345), .A2(n1009), .Z(n3478) );
  CKND0BWP12T U1795 ( .I(n1010), .ZN(n1011) );
  NR2D0BWP12T U1796 ( .A1(n1011), .A2(n1014), .ZN(n1017) );
  CKND0BWP12T U1797 ( .I(n1012), .ZN(n1015) );
  OAI21D0BWP12T U1798 ( .A1(n1015), .A2(n1014), .B(n1013), .ZN(n1016) );
  AOI21D1BWP12T U1799 ( .A1(n2490), .A2(n1017), .B(n1016), .ZN(n1021) );
  CKND2D0BWP12T U1800 ( .A1(n1045), .A2(n1019), .ZN(n1020) );
  XOR2XD1BWP12T U1801 ( .A1(n1021), .A2(n1020), .Z(n3587) );
  TPOAI22D0BWP12T U1802 ( .A1(n2586), .A2(n3786), .B1(n2823), .B2(n3782), .ZN(
        n1023) );
  OAI22D1BWP12T U1803 ( .A1(n2824), .A2(n3784), .B1(n2822), .B2(n3780), .ZN(
        n1022) );
  NR2D1BWP12T U1804 ( .A1(n1023), .A2(n1022), .ZN(n3753) );
  INVD1BWP12T U1805 ( .I(n3753), .ZN(n3076) );
  TPND2D0BWP12T U1806 ( .A1(n3229), .A2(n2824), .ZN(n1026) );
  AOI22D1BWP12T U1807 ( .A1(n2823), .A2(n3227), .B1(n3231), .B2(n2586), .ZN(
        n1025) );
  CKND2D1BWP12T U1808 ( .A1(n3707), .A2(n2822), .ZN(n1024) );
  ND3D1BWP12T U1809 ( .A1(n1026), .A2(n1025), .A3(n1024), .ZN(n3686) );
  INVD1BWP12T U1810 ( .I(n3686), .ZN(n3064) );
  OAI21D0BWP12T U1811 ( .A1(n4084), .A2(n4182), .B(n4181), .ZN(n1027) );
  INVD1BWP12T U1812 ( .I(n4184), .ZN(n3364) );
  MUX2ND0BWP12T U1813 ( .I0(n3364), .I1(n3363), .S(n3929), .ZN(n1028) );
  CKND2D0BWP12T U1814 ( .A1(n1028), .A2(n4181), .ZN(n1029) );
  CKND0BWP12T U1815 ( .I(n1030), .ZN(n1031) );
  NR2D0BWP12T U1816 ( .A1(n1031), .A2(n1034), .ZN(n1037) );
  CKND0BWP12T U1817 ( .I(n1032), .ZN(n1035) );
  TPOAI21D0BWP12T U1818 ( .A1(n1035), .A2(n1034), .B(n1033), .ZN(n1036) );
  AOI21D1BWP12T U1819 ( .A1(n2504), .A2(n1037), .B(n1036), .ZN(n1042) );
  CKND0BWP12T U1820 ( .I(n1038), .ZN(n1040) );
  TPND2D0BWP12T U1821 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XOR2XD1BWP12T U1822 ( .A1(n1042), .A2(n1041), .Z(n3540) );
  OAI21D0BWP12T U1823 ( .A1(n2918), .A2(n3841), .B(n2780), .ZN(n1043) );
  AOI211D0BWP12T U1824 ( .A1(n2970), .A2(n1043), .B(n3726), .C(n3655), .ZN(
        n1044) );
  INVD1BWP12T U1825 ( .I(n3384), .ZN(n2423) );
  NR2D0BWP12T U1826 ( .A1(n1044), .A2(n2423), .ZN(n4026) );
  CKND0BWP12T U1827 ( .I(n1083), .ZN(n1045) );
  RCAOI22D0BWP12T U1828 ( .A1(n4210), .A2(n4112), .B1(n3630), .B2(n4203), .ZN(
        n1051) );
  INVD1BWP12T U1829 ( .I(n1047), .ZN(n3684) );
  TPNR2D0BWP12T U1830 ( .A1(n3684), .A2(n4201), .ZN(n1049) );
  INVD1BWP12T U1831 ( .I(n3726), .ZN(n1048) );
  TPOAI21D0BWP12T U1832 ( .A1(n1049), .A2(n3360), .B(n1048), .ZN(n1050) );
  OAI211D1BWP12T U1833 ( .A1(n4026), .A2(n3029), .B(n1051), .C(n1050), .ZN(
        n1052) );
  AOI211D1BWP12T U1834 ( .A1(n3985), .A2(n3973), .B(n1053), .C(n1052), .ZN(
        n1054) );
  ND2D1BWP12T U1835 ( .A1(n1055), .A2(n1054), .ZN(result[7]) );
  INVD0BWP12T U1836 ( .I(n2800), .ZN(n1061) );
  XNR2XD1BWP12T U1837 ( .A1(n3351), .A2(n4062), .ZN(n3634) );
  CKND2D1BWP12T U1838 ( .A1(n1086), .A2(n2816), .ZN(n1062) );
  XOR2XD1BWP12T U1839 ( .A1(n3388), .A2(n1062), .Z(n3589) );
  INVD8BWP12T U1840 ( .I(n4065), .ZN(n3895) );
  OAI22D1BWP12T U1841 ( .A1(n2469), .A2(n3895), .B1(n3911), .B2(n2468), .ZN(
        n1064) );
  CKND1BWP12T U1842 ( .I(a[29]), .ZN(n3894) );
  OAI22D1BWP12T U1843 ( .A1(n2471), .A2(n3899), .B1(n2470), .B2(n3894), .ZN(
        n1063) );
  NR2D1BWP12T U1844 ( .A1(n1064), .A2(n1063), .ZN(n3681) );
  INVD1BWP12T U1845 ( .I(n3681), .ZN(n2402) );
  ND2D0BWP12T U1846 ( .A1(n1065), .A2(n3916), .ZN(n1067) );
  AOI22D1BWP12T U1847 ( .A1(n2463), .A2(n4157), .B1(n2462), .B2(n4064), .ZN(
        n1066) );
  ND2D1BWP12T U1848 ( .A1(n1067), .A2(n1066), .ZN(n1852) );
  AOI22D1BWP12T U1849 ( .A1(n2579), .A2(n2402), .B1(n1852), .B2(n3353), .ZN(
        n4014) );
  OAI21D0BWP12T U1850 ( .A1(n4014), .A2(n3655), .B(n3765), .ZN(n1081) );
  OAI22D1BWP12T U1851 ( .A1(n2469), .A2(n3865), .B1(n2471), .B2(n3862), .ZN(
        n1069) );
  OAI22D1BWP12T U1852 ( .A1(n2470), .A2(n3864), .B1(n2468), .B2(n3863), .ZN(
        n1068) );
  NR2D1BWP12T U1853 ( .A1(n1069), .A2(n1068), .ZN(n1849) );
  INVD1BWP12T U1854 ( .I(n1849), .ZN(n1815) );
  OAI22D1BWP12T U1855 ( .A1(n2469), .A2(n4062), .B1(n4060), .B2(n2468), .ZN(
        n1071) );
  OAI22D1BWP12T U1856 ( .A1(n4061), .A2(n2471), .B1(n2470), .B2(n4063), .ZN(
        n1070) );
  NR2D1BWP12T U1857 ( .A1(n1071), .A2(n1070), .ZN(n2413) );
  AOI22D1BWP12T U1858 ( .A1(n1072), .A2(n1815), .B1(n2413), .B2(n3353), .ZN(
        n1080) );
  OAI22D1BWP12T U1859 ( .A1(n2469), .A2(n3876), .B1(n2468), .B2(n3874), .ZN(
        n1074) );
  OAI22D1BWP12T U1860 ( .A1(n2471), .A2(n3873), .B1(n2470), .B2(n3875), .ZN(
        n1073) );
  NR2D1BWP12T U1861 ( .A1(n1074), .A2(n1073), .ZN(n2414) );
  OAI21D0BWP12T U1862 ( .A1(n2414), .A2(n3356), .B(n3841), .ZN(n1078) );
  OAI22D1BWP12T U1863 ( .A1(n2469), .A2(n4187), .B1(n2470), .B2(n3868), .ZN(
        n1076) );
  OAI22D1BWP12T U1864 ( .A1(n2471), .A2(n3867), .B1(n2468), .B2(n3866), .ZN(
        n1075) );
  NR2D1BWP12T U1865 ( .A1(n1076), .A2(n1075), .ZN(n2420) );
  TPNR2D0BWP12T U1866 ( .A1(n2420), .A2(n2949), .ZN(n1077) );
  NR2XD0BWP12T U1867 ( .A1(n1078), .A2(n1077), .ZN(n1079) );
  ND2D1BWP12T U1868 ( .A1(n1080), .A2(n1079), .ZN(n1101) );
  ND2D1BWP12T U1869 ( .A1(n1081), .A2(n1101), .ZN(n3978) );
  MAOI22D0BWP12T U1870 ( .A1(n3589), .A2(n4206), .B1(n3978), .B2(n2834), .ZN(
        n1087) );
  INVD0BWP12T U1871 ( .I(n1084), .ZN(n1086) );
  CKND2D0BWP12T U1872 ( .A1(n4014), .A2(n3919), .ZN(n1092) );
  NR2D1BWP12T U1873 ( .A1(n2547), .A2(n3170), .ZN(n4175) );
  CKND2D1BWP12T U1874 ( .A1(n2462), .A2(n4066), .ZN(n1848) );
  INVD1BWP12T U1875 ( .I(n1848), .ZN(n1831) );
  CKND2D1BWP12T U1876 ( .A1(n1831), .A2(n3886), .ZN(n3772) );
  INVD1BWP12T U1877 ( .I(n3772), .ZN(n4178) );
  AOI22D1BWP12T U1878 ( .A1(n3229), .A2(n1833), .B1(n2806), .B2(n1838), .ZN(
        n1091) );
  ND3D0BWP12T U1879 ( .A1(n1089), .A2(n1088), .A3(n1832), .ZN(n1090) );
  OAI211D1BWP12T U1880 ( .A1(n2333), .A2(n3005), .B(n1091), .C(n1090), .ZN(
        n4176) );
  AOI222D1BWP12T U1881 ( .A1(n1092), .A2(n1101), .B1(n4175), .B2(n4178), .C1(
        n4176), .C2(n4179), .ZN(n3665) );
  OAI21D0BWP12T U1882 ( .A1(n4062), .A2(n4182), .B(n4181), .ZN(n1100) );
  OAI22D1BWP12T U1883 ( .A1(n1838), .A2(n3782), .B1(n2294), .B2(n3780), .ZN(
        n1094) );
  TPNR2D0BWP12T U1884 ( .A1(n1832), .A2(n3786), .ZN(n1093) );
  AOI211D1BWP12T U1885 ( .A1(n3242), .A2(n1827), .B(n1094), .C(n1093), .ZN(
        n3769) );
  INVD1BWP12T U1886 ( .I(n3769), .ZN(n2264) );
  MUX2ND0BWP12T U1887 ( .I0(n2264), .I1(n3772), .S(n3922), .ZN(n1095) );
  ND2D1BWP12T U1888 ( .A1(n1095), .A2(n3997), .ZN(n3806) );
  NR2D1BWP12T U1889 ( .A1(n3806), .A2(n3773), .ZN(n1099) );
  MUX2ND0BWP12T U1890 ( .I0(n4184), .I1(n2664), .S(n3928), .ZN(n1096) );
  NR2XD0BWP12T U1891 ( .A1(n1096), .A2(n4185), .ZN(n1097) );
  MUX2NXD0BWP12T U1892 ( .I0(n1097), .I1(n2205), .S(n3880), .ZN(n1098) );
  AOI211D1BWP12T U1893 ( .A1(n3928), .A2(n1100), .B(n1099), .C(n1098), .ZN(
        n1104) );
  CKND0BWP12T U1894 ( .I(n1101), .ZN(n1102) );
  OAI211D1BWP12T U1895 ( .A1(n1102), .A2(n2970), .B(n3978), .C(n3384), .ZN(
        n4022) );
  CKND2D1BWP12T U1896 ( .A1(n4022), .A2(n4011), .ZN(n1103) );
  OAI211D1BWP12T U1897 ( .A1(n3665), .A2(n4201), .B(n1104), .C(n1103), .ZN(
        n1105) );
  AOI211D1BWP12T U1898 ( .A1(n4215), .A2(n3541), .B(n1106), .C(n1105), .ZN(
        n1107) );
  IOA21D1BWP12T U1899 ( .A1(n4173), .A2(n3493), .B(n1107), .ZN(n1108) );
  AO21D1BWP12T U1900 ( .A1(n3418), .A2(n4171), .B(n1108), .Z(result[8]) );
  XNR2D1BWP12T U1901 ( .A1(n1977), .A2(n3941), .ZN(n1115) );
  XNR2D1BWP12T U1902 ( .A1(n1977), .A2(n3943), .ZN(n1109) );
  OAI22D1BWP12T U1903 ( .A1(n2019), .A2(n1115), .B1(n1109), .B2(n2018), .ZN(
        n1113) );
  XNR2D1BWP12T U1904 ( .A1(n2058), .A2(n3927), .ZN(n1114) );
  XNR2D1BWP12T U1905 ( .A1(n2058), .A2(n3929), .ZN(n1179) );
  TPOAI22D1BWP12T U1906 ( .A1(n1650), .A2(n1114), .B1(n1179), .B2(n1648), .ZN(
        n1112) );
  XNR2D1BWP12T U1907 ( .A1(n4082), .A2(n3957), .ZN(n1111) );
  XNR2D1BWP12T U1908 ( .A1(n4082), .A2(n3932), .ZN(n1172) );
  OAI22D1BWP12T U1909 ( .A1(n2130), .A2(n1111), .B1(n754), .B2(n1172), .ZN(
        n1208) );
  XNR2D1BWP12T U1910 ( .A1(n1977), .A2(n3918), .ZN(n1202) );
  OAI22D1BWP12T U1911 ( .A1(n1110), .A2(n1109), .B1(n1202), .B2(n2018), .ZN(
        n1201) );
  INVD4BWP12T U1912 ( .I(a[23]), .ZN(n2064) );
  XNR2XD4BWP12T U1913 ( .A1(n2064), .A2(n3898), .ZN(n2021) );
  INR2D2BWP12T U1914 ( .A1(n1979), .B1(n2021), .ZN(n1200) );
  XNR2D1BWP12T U1915 ( .A1(n3885), .A2(n3939), .ZN(n1151) );
  XNR2D1BWP12T U1916 ( .A1(n3885), .A2(n3941), .ZN(n1192) );
  OAI22D1BWP12T U1917 ( .A1(n2072), .A2(n1151), .B1(n2070), .B2(n1192), .ZN(
        n1199) );
  XNR2D1BWP12T U1918 ( .A1(n2084), .A2(n3932), .ZN(n1125) );
  XNR2D1BWP12T U1919 ( .A1(n2084), .A2(n3933), .ZN(n1168) );
  OAI22D1BWP12T U1920 ( .A1(n2088), .A2(n1125), .B1(n2086), .B2(n1168), .ZN(
        n1118) );
  XNR2D1BWP12T U1921 ( .A1(n4082), .A2(n3928), .ZN(n1123) );
  OAI22D1BWP12T U1922 ( .A1(n2130), .A2(n1123), .B1(n754), .B2(n1111), .ZN(
        n1117) );
  HA1D1BWP12T U1923 ( .A(n1113), .B(n1112), .CO(n1209), .S(n1116) );
  XNR2D1BWP12T U1924 ( .A1(n4060), .A2(n3933), .ZN(n1127) );
  XNR2D1BWP12T U1925 ( .A1(n4060), .A2(n3950), .ZN(n1121) );
  OAI22D1BWP12T U1926 ( .A1(n2009), .A2(n1127), .B1(n1121), .B2(n2006), .ZN(
        n1141) );
  XNR2D1BWP12T U1927 ( .A1(n2058), .A2(n3920), .ZN(n1133) );
  TPOAI22D1BWP12T U1928 ( .A1(n1650), .A2(n1133), .B1(n1114), .B2(n1648), .ZN(
        n1140) );
  XNR2D1BWP12T U1929 ( .A1(n4084), .A2(n3949), .ZN(n1142) );
  XNR2D1BWP12T U1930 ( .A1(n4084), .A2(n4191), .ZN(n1122) );
  OAI22D1BWP12T U1931 ( .A1(n2013), .A2(n1142), .B1(n2011), .B2(n1122), .ZN(
        n1139) );
  XNR2D1BWP12T U1932 ( .A1(n1977), .A2(n3939), .ZN(n1132) );
  OAI22D1BWP12T U1933 ( .A1(n2019), .A2(n1132), .B1(n1115), .B2(n2018), .ZN(
        n1131) );
  XNR2XD8BWP12T U1934 ( .A1(n4070), .A2(a[21]), .ZN(n2065) );
  INR2D1BWP12T U1935 ( .A1(n1979), .B1(n2065), .ZN(n1130) );
  XNR2D0BWP12T U1936 ( .A1(n3885), .A2(b[19]), .ZN(n1128) );
  XNR2D1BWP12T U1937 ( .A1(n4068), .A2(n3938), .ZN(n1152) );
  OAI22D1BWP12T U1938 ( .A1(n2072), .A2(n1128), .B1(n2070), .B2(n1152), .ZN(
        n1129) );
  FA1D0BWP12T U1939 ( .A(n1118), .B(n1117), .CI(n1116), .CO(n1197), .S(n1136)
         );
  OAI21D1BWP12T U1940 ( .A1(n1138), .A2(n1137), .B(n1136), .ZN(n1119) );
  IOA21D1BWP12T U1941 ( .A1(n1137), .A2(n1138), .B(n1119), .ZN(n1196) );
  XNR2XD8BWP12T U1942 ( .A1(n4069), .A2(a[19]), .ZN(n2077) );
  XOR2XD2BWP12T U1943 ( .A1(n4069), .A2(a[21]), .Z(n1120) );
  ND2XD16BWP12T U1944 ( .A1(n2077), .A2(n1120), .ZN(n2079) );
  XNR2D1BWP12T U1945 ( .A1(n3921), .A2(a[21]), .ZN(n1154) );
  XNR2D1BWP12T U1946 ( .A1(n3922), .A2(a[21]), .ZN(n1169) );
  OAI22D1BWP12T U1947 ( .A1(n2079), .A2(n1154), .B1(n2077), .B2(n1169), .ZN(
        n1211) );
  XNR2XD1BWP12T U1948 ( .A1(n4060), .A2(n3931), .ZN(n1170) );
  OAI22D1BWP12T U1949 ( .A1(n2009), .A2(n1121), .B1(n1170), .B2(n2006), .ZN(
        n1212) );
  XNR2D1BWP12T U1950 ( .A1(n4084), .A2(n3952), .ZN(n1180) );
  OAI22D1BWP12T U1951 ( .A1(n2013), .A2(n1122), .B1(n2011), .B2(n1180), .ZN(
        n1210) );
  XOR3D2BWP12T U1952 ( .A1(n1211), .A2(n1212), .A3(n1210), .Z(n1257) );
  XNR2D1BWP12T U1953 ( .A1(n4082), .A2(n3929), .ZN(n1234) );
  TPOAI22D1BWP12T U1954 ( .A1(n2130), .A2(n1234), .B1(n754), .B2(n1123), .ZN(
        n1145) );
  XOR2XD8BWP12T U1955 ( .A1(n3820), .A2(a[19]), .Z(n1124) );
  ND2XD8BWP12T U1956 ( .A1(n2125), .A2(n1124), .ZN(n2127) );
  XNR2D1BWP12T U1957 ( .A1(n3922), .A2(a[19]), .ZN(n1235) );
  XNR2D1BWP12T U1958 ( .A1(n2098), .A2(a[19]), .ZN(n1156) );
  TPOAI22D2BWP12T U1959 ( .A1(n2127), .A2(n1235), .B1(n2125), .B2(n1156), .ZN(
        n1144) );
  XNR2D1BWP12T U1960 ( .A1(n2084), .A2(n3957), .ZN(n1251) );
  OAI22D1BWP12T U1961 ( .A1(n2088), .A2(n1251), .B1(n2086), .B2(n1125), .ZN(
        n1143) );
  IND2XD1BWP12T U1962 ( .A1(b[0]), .B1(a[21]), .ZN(n1126) );
  TPOAI22D2BWP12T U1963 ( .A1(n2079), .A2(n1746), .B1(n2077), .B2(n1126), .ZN(
        n1278) );
  XNR2D1BWP12T U1964 ( .A1(n4060), .A2(n3932), .ZN(n1231) );
  OAI22D1BWP12T U1965 ( .A1(n2009), .A2(n1231), .B1(n1127), .B2(n2006), .ZN(
        n1277) );
  XNR2D1BWP12T U1966 ( .A1(n3885), .A2(n3951), .ZN(n1253) );
  OAI22D1BWP12T U1967 ( .A1(n2072), .A2(n1253), .B1(n2070), .B2(n1128), .ZN(
        n1276) );
  FA1D2BWP12T U1968 ( .A(n1131), .B(n1130), .CI(n1129), .CO(n1138), .S(n1240)
         );
  OAI22D1BWP12T U1969 ( .A1(n2019), .A2(n1252), .B1(n1132), .B2(n2018), .ZN(
        n1250) );
  XNR2D1BWP12T U1970 ( .A1(n2058), .A2(n2098), .ZN(n1232) );
  OAI22D2BWP12T U1971 ( .A1(n1650), .A2(n1232), .B1(n1133), .B2(n1648), .ZN(
        n1249) );
  ND2D1BWP12T U1972 ( .A1(n1240), .A2(n1241), .ZN(n1134) );
  TPND2D1BWP12T U1973 ( .A1(n1135), .A2(n1134), .ZN(n1255) );
  INVD1BWP12T U1974 ( .I(n1267), .ZN(n1164) );
  INVD1BWP12T U1975 ( .I(n1268), .ZN(n1163) );
  XOR3D1BWP12T U1976 ( .A1(n1138), .A2(n1137), .A3(n1136), .Z(n1322) );
  CKND1BWP12T U1977 ( .I(n1322), .ZN(n1160) );
  FA1D2BWP12T U1978 ( .A(n1141), .B(n1140), .CI(n1139), .CO(n1137), .S(n1272)
         );
  XNR2XD1BWP12T U1979 ( .A1(n4075), .A2(n4191), .ZN(n1230) );
  XNR2D1BWP12T U1980 ( .A1(n4075), .A2(n3952), .ZN(n1153) );
  OAI22D1BWP12T U1981 ( .A1(n2083), .A2(n1230), .B1(n1153), .B2(n2080), .ZN(
        n1287) );
  XNR2D1BWP12T U1982 ( .A1(n1517), .A2(a[21]), .ZN(n1155) );
  XNR2D1BWP12T U1983 ( .A1(n4084), .A2(n3930), .ZN(n1233) );
  OAI22D1BWP12T U1984 ( .A1(n2013), .A2(n1233), .B1(n2011), .B2(n1142), .ZN(
        n1285) );
  ND2D1BWP12T U1985 ( .A1(n1272), .A2(n1275), .ZN(n1147) );
  FA1D1BWP12T U1986 ( .A(n1145), .B(n1144), .CI(n1143), .CO(n1256), .S(n1274)
         );
  OAI21D1BWP12T U1987 ( .A1(n1272), .A2(n1275), .B(n1274), .ZN(n1146) );
  ND2D1BWP12T U1988 ( .A1(n1147), .A2(n1146), .ZN(n1321) );
  CKND1BWP12T U1989 ( .I(n1321), .ZN(n1159) );
  XNR2D1BWP12T U1990 ( .A1(n2064), .A2(n4070), .ZN(n1148) );
  ND2D4BWP12T U1991 ( .A1(n2065), .A2(n1148), .ZN(n2068) );
  XNR2D0BWP12T U1992 ( .A1(n1979), .A2(a[23]), .ZN(n1149) );
  XNR2D1BWP12T U1993 ( .A1(n1517), .A2(a[23]), .ZN(n1178) );
  OAI22D1BWP12T U1994 ( .A1(n2068), .A2(n1149), .B1(n1178), .B2(n2065), .ZN(
        n1217) );
  OR2XD1BWP12T U1995 ( .A1(b[0]), .A2(n2064), .Z(n1150) );
  OAI22D1BWP12T U1996 ( .A1(n2068), .A2(n2064), .B1(n2065), .B2(n1150), .ZN(
        n1216) );
  OAI22D1BWP12T U1997 ( .A1(n2072), .A2(n1152), .B1(n2070), .B2(n1151), .ZN(
        n1215) );
  XNR2XD1BWP12T U1998 ( .A1(n4075), .A2(n3951), .ZN(n1157) );
  OAI22D1BWP12T U1999 ( .A1(n2083), .A2(n1153), .B1(n1157), .B2(n2080), .ZN(
        n1245) );
  XNR2XD1BWP12T U2000 ( .A1(n595), .A2(n3931), .ZN(n1237) );
  XNR2D1BWP12T U2001 ( .A1(n4063), .A2(n3930), .ZN(n1158) );
  OAI22D1BWP12T U2002 ( .A1(n2027), .A2(n1237), .B1(n1986), .B2(n1158), .ZN(
        n1243) );
  XNR2D1BWP12T U2003 ( .A1(a[19]), .A2(n3920), .ZN(n1166) );
  XNR2XD1BWP12T U2004 ( .A1(n4075), .A2(b[19]), .ZN(n1167) );
  OAI22D1BWP12T U2005 ( .A1(n2083), .A2(n1157), .B1(n1167), .B2(n2080), .ZN(
        n1176) );
  XNR2XD1BWP12T U2006 ( .A1(n4063), .A2(n3949), .ZN(n1171) );
  OAI22D1BWP12T U2007 ( .A1(n2027), .A2(n1158), .B1(n1986), .B2(n1171), .ZN(
        n1175) );
  IOA21D1BWP12T U2008 ( .A1(n1160), .A2(n1159), .B(n1320), .ZN(n1162) );
  CKND2D1BWP12T U2009 ( .A1(n1321), .A2(n1322), .ZN(n1161) );
  ND2D1BWP12T U2010 ( .A1(n1162), .A2(n1161), .ZN(n1266) );
  IOA21D1BWP12T U2011 ( .A1(n1164), .A2(n1163), .B(n1266), .ZN(n1165) );
  IOA21D1BWP12T U2012 ( .A1(n1268), .A2(n1267), .B(n1165), .ZN(n1375) );
  XNR2D1BWP12T U2013 ( .A1(n1699), .A2(n3927), .ZN(n1173) );
  XNR2XD1BWP12T U2014 ( .A1(n4075), .A2(n3938), .ZN(n1193) );
  OAI22D1BWP12T U2015 ( .A1(n2083), .A2(n1167), .B1(n1193), .B2(n2080), .ZN(
        n1219) );
  XNR2D1BWP12T U2016 ( .A1(n2084), .A2(n3950), .ZN(n1174) );
  OAI22D1BWP12T U2017 ( .A1(n2088), .A2(n1168), .B1(n2086), .B2(n1174), .ZN(
        n1218) );
  XNR2XD1BWP12T U2018 ( .A1(n2098), .A2(a[21]), .ZN(n1184) );
  OAI22D1BWP12T U2019 ( .A1(n2079), .A2(n1169), .B1(n2077), .B2(n1184), .ZN(
        n1183) );
  XNR2D1BWP12T U2020 ( .A1(n4060), .A2(n3930), .ZN(n1188) );
  OAI22D1BWP12T U2021 ( .A1(n2009), .A2(n1170), .B1(n1188), .B2(n2006), .ZN(
        n1182) );
  XNR2XD1BWP12T U2022 ( .A1(n4063), .A2(n4191), .ZN(n1187) );
  OAI22D1BWP12T U2023 ( .A1(n2027), .A2(n1171), .B1(n1986), .B2(n1187), .ZN(
        n1181) );
  XNR2D1BWP12T U2024 ( .A1(n4082), .A2(n3933), .ZN(n1360) );
  TPOAI22D1BWP12T U2025 ( .A1(n2130), .A2(n1172), .B1(n754), .B2(n1360), .ZN(
        n1338) );
  XNR2D1BWP12T U2026 ( .A1(n1699), .A2(n3929), .ZN(n1361) );
  OAI22D1BWP12T U2027 ( .A1(n2127), .A2(n1173), .B1(n2125), .B2(n1361), .ZN(
        n1337) );
  XNR2D0BWP12T U2028 ( .A1(n2084), .A2(n3931), .ZN(n1372) );
  OAI22D1BWP12T U2029 ( .A1(n2088), .A2(n1174), .B1(n2086), .B2(n1372), .ZN(
        n1336) );
  FA1D0BWP12T U2030 ( .A(n1177), .B(n1176), .CI(n1175), .CO(n1229), .S(n1224)
         );
  XOR2XD1BWP12T U2031 ( .A1(n3921), .A2(n2064), .Z(n1191) );
  OAI22D1BWP12T U2032 ( .A1(n2068), .A2(n1178), .B1(n1191), .B2(n2065), .ZN(
        n1206) );
  XNR2D1BWP12T U2033 ( .A1(n2058), .A2(n3928), .ZN(n1203) );
  OAI22D1BWP12T U2034 ( .A1(n2062), .A2(n1179), .B1(n1203), .B2(n1648), .ZN(
        n1205) );
  XNR2XD1BWP12T U2035 ( .A1(n4084), .A2(n3951), .ZN(n1195) );
  OAI22D1BWP12T U2036 ( .A1(n2013), .A2(n1180), .B1(n2011), .B2(n1195), .ZN(
        n1204) );
  FA1D2BWP12T U2037 ( .A(n1183), .B(n1182), .CI(n1181), .CO(n1331), .S(n1227)
         );
  XNR2D1BWP12T U2038 ( .A1(a[21]), .A2(n3920), .ZN(n1371) );
  CKXOR2D1BWP12T U2039 ( .A1(n4157), .A2(n4064), .Z(n1185) );
  IND2D0BWP12T U2040 ( .A1(b[0]), .B1(n4157), .ZN(n1186) );
  OAI22D1BWP12T U2041 ( .A1(n2023), .A2(n3618), .B1(n2021), .B2(n1186), .ZN(
        n1368) );
  XNR2D1BWP12T U2042 ( .A1(n4063), .A2(n3952), .ZN(n1345) );
  OAI22D1BWP12T U2043 ( .A1(n2027), .A2(n1187), .B1(n1986), .B2(n1345), .ZN(
        n1367) );
  XNR2D1BWP12T U2044 ( .A1(n4060), .A2(n3949), .ZN(n1344) );
  OAI22D1BWP12T U2045 ( .A1(n2009), .A2(n1188), .B1(n1344), .B2(n2006), .ZN(
        n1357) );
  CKND1BWP12T U2046 ( .I(n1189), .ZN(n1190) );
  XNR2D1BWP12T U2047 ( .A1(n3885), .A2(n3943), .ZN(n1359) );
  OAI22D1BWP12T U2048 ( .A1(n2072), .A2(n1192), .B1(n2070), .B2(n1359), .ZN(
        n1355) );
  XNR2XD1BWP12T U2049 ( .A1(n4075), .A2(n3939), .ZN(n1370) );
  OAI22D1BWP12T U2050 ( .A1(n2083), .A2(n1193), .B1(n1370), .B2(n2080), .ZN(
        n1366) );
  XNR2XD1BWP12T U2051 ( .A1(n1979), .A2(n4157), .ZN(n1194) );
  XNR2D1BWP12T U2052 ( .A1(n1517), .A2(n4157), .ZN(n1343) );
  OAI22D1BWP12T U2053 ( .A1(n2023), .A2(n1194), .B1(n2021), .B2(n1343), .ZN(
        n1365) );
  XNR2XD1BWP12T U2054 ( .A1(n4084), .A2(b[19]), .ZN(n1342) );
  OAI22D1BWP12T U2055 ( .A1(n2013), .A2(n1195), .B1(n2011), .B2(n1342), .ZN(
        n1364) );
  FA1D2BWP12T U2056 ( .A(n1198), .B(n1197), .CI(n1196), .CO(n1328), .S(n1268)
         );
  FA1D0BWP12T U2057 ( .A(n1201), .B(n1200), .CI(n1199), .CO(n1335), .S(n1207)
         );
  XNR2D1BWP12T U2058 ( .A1(n1977), .A2(b[25]), .ZN(n1358) );
  OAI22D1BWP12T U2059 ( .A1(n2019), .A2(n1202), .B1(n1358), .B2(n2018), .ZN(
        n1363) );
  XNR2D1BWP12T U2060 ( .A1(n1339), .A2(n1959), .ZN(n1340) );
  OAI22D1BWP12T U2061 ( .A1(n1650), .A2(n1203), .B1(n1340), .B2(n1648), .ZN(
        n1362) );
  FA1D1BWP12T U2062 ( .A(n1209), .B(n1208), .CI(n1207), .CO(n1347), .S(n1198)
         );
  ND2D1BWP12T U2063 ( .A1(n1212), .A2(n1211), .ZN(n1213) );
  ND2D1BWP12T U2064 ( .A1(n1214), .A2(n1213), .ZN(n1223) );
  FA1D1BWP12T U2065 ( .A(n1217), .B(n1216), .CI(n1215), .CO(n1222), .S(n1226)
         );
  FA1D1BWP12T U2066 ( .A(n1220), .B(n1219), .CI(n1218), .CO(n1332), .S(n1221)
         );
  FA1D1BWP12T U2067 ( .A(n1223), .B(n1222), .CI(n1221), .CO(n1346), .S(n1265)
         );
  FA1D1BWP12T U2068 ( .A(n1226), .B(n1225), .CI(n1224), .CO(n1264), .S(n1320)
         );
  FA1D1BWP12T U2069 ( .A(n1229), .B(n1228), .CI(n1227), .CO(n1350), .S(n1263)
         );
  XOR3D2BWP12T U2070 ( .A1(n1328), .A2(n1329), .A3(n1326), .Z(n1373) );
  XNR2D1BWP12T U2071 ( .A1(n1517), .A2(a[19]), .ZN(n1313) );
  XNR2D1BWP12T U2072 ( .A1(n3921), .A2(a[19]), .ZN(n1236) );
  XNR2XD1BWP12T U2073 ( .A1(n4075), .A2(n3949), .ZN(n1293) );
  OAI22D1BWP12T U2074 ( .A1(n2083), .A2(n1293), .B1(n1230), .B2(n2080), .ZN(
        n1318) );
  XNR2D1BWP12T U2075 ( .A1(n4063), .A2(n3933), .ZN(n1412) );
  XNR2D1BWP12T U2076 ( .A1(n4063), .A2(n3950), .ZN(n1238) );
  OAI22D1BWP12T U2077 ( .A1(n2027), .A2(n1412), .B1(n2025), .B2(n1238), .ZN(
        n1317) );
  XNR2D1BWP12T U2078 ( .A1(n4060), .A2(n3957), .ZN(n1291) );
  OAI22D1BWP12T U2079 ( .A1(n2009), .A2(n1291), .B1(n1231), .B2(n2006), .ZN(
        n1310) );
  XNR2D1BWP12T U2080 ( .A1(n2058), .A2(n3922), .ZN(n1283) );
  TPOAI22D1BWP12T U2081 ( .A1(n1650), .A2(n1283), .B1(n1232), .B2(n1648), .ZN(
        n1309) );
  XNR2D1BWP12T U2082 ( .A1(n4084), .A2(n3931), .ZN(n1315) );
  OAI22D1BWP12T U2083 ( .A1(n2013), .A2(n1315), .B1(n2011), .B2(n1233), .ZN(
        n1308) );
  XNR2D1BWP12T U2084 ( .A1(n4082), .A2(n3927), .ZN(n1280) );
  OAI22D1BWP12T U2085 ( .A1(n2130), .A2(n1280), .B1(n754), .B2(n1234), .ZN(
        n1248) );
  OAI22D1BWP12T U2086 ( .A1(n2127), .A2(n1236), .B1(n2125), .B2(n1235), .ZN(
        n1247) );
  OAI22D1BWP12T U2087 ( .A1(n2027), .A2(n1238), .B1(n2025), .B2(n1237), .ZN(
        n1246) );
  XOR3D1BWP12T U2088 ( .A1(n1241), .A2(n1240), .A3(n1239), .Z(n1470) );
  CKND1BWP12T U2089 ( .I(n1470), .ZN(n1242) );
  FA1D0BWP12T U2090 ( .A(n1248), .B(n1247), .CI(n1246), .CO(n1259), .S(n1459)
         );
  HA1D1BWP12T U2091 ( .A(n1250), .B(n1249), .CO(n1241), .S(n1307) );
  XNR2D1BWP12T U2092 ( .A1(n2084), .A2(n3928), .ZN(n1279) );
  OAI22D1BWP12T U2093 ( .A1(n2088), .A2(n1279), .B1(n2086), .B2(n1251), .ZN(
        n1306) );
  XNR2D1BWP12T U2094 ( .A1(n1977), .A2(b[19]), .ZN(n1281) );
  XNR2D1BWP12T U2095 ( .A1(n3885), .A2(n3952), .ZN(n1295) );
  OAI22D1BWP12T U2096 ( .A1(n2072), .A2(n1295), .B1(n2070), .B2(n1253), .ZN(
        n1299) );
  AOI22D1BWP12T U2097 ( .A1(n1254), .A2(n1468), .B1(n1470), .B2(n1469), .ZN(
        n1323) );
  FA1D2BWP12T U2098 ( .A(n1257), .B(n1256), .CI(n1255), .CO(n1267), .S(n1324)
         );
  FA1D1BWP12T U2099 ( .A(n1260), .B(n1259), .CI(n1258), .CO(n1325), .S(n1468)
         );
  NR2D1BWP12T U2100 ( .A1(n1324), .A2(n1325), .ZN(n1262) );
  ND2D1BWP12T U2101 ( .A1(n1324), .A2(n1325), .ZN(n1261) );
  FA1D1BWP12T U2102 ( .A(n1265), .B(n1264), .CI(n1263), .CO(n1326), .S(n1270)
         );
  XOR3D2BWP12T U2103 ( .A1(n1268), .A2(n1267), .A3(n1266), .Z(n1269) );
  TPNR2D1BWP12T U2104 ( .A1(n1510), .A2(n1509), .ZN(n1511) );
  INVD1BWP12T U2105 ( .I(n1511), .ZN(n3456) );
  FA1D1BWP12T U2106 ( .A(n1271), .B(n1270), .CI(n1269), .CO(n1509), .S(n1508)
         );
  INVD1BWP12T U2107 ( .I(n1272), .ZN(n1273) );
  XNR3XD4BWP12T U2108 ( .A1(n1275), .A2(n1274), .A3(n1273), .ZN(n1473) );
  FA1D2BWP12T U2109 ( .A(n1278), .B(n1277), .CI(n1276), .CO(n1239), .S(n1458)
         );
  XNR2D1BWP12T U2110 ( .A1(n2084), .A2(n3929), .ZN(n1408) );
  OAI22D1BWP12T U2111 ( .A1(n2088), .A2(n1408), .B1(n2086), .B2(n1279), .ZN(
        n1290) );
  XNR2D1BWP12T U2112 ( .A1(n4082), .A2(n3920), .ZN(n1410) );
  OAI22D1BWP12T U2113 ( .A1(n2130), .A2(n1410), .B1(n754), .B2(n1280), .ZN(
        n1289) );
  OAI22D1BWP12T U2114 ( .A1(n2019), .A2(n1282), .B1(n1281), .B2(n2018), .ZN(
        n1386) );
  OAI22D1BWP12T U2115 ( .A1(n1650), .A2(n1284), .B1(n1283), .B2(n1648), .ZN(
        n1385) );
  FA1D2BWP12T U2116 ( .A(n1287), .B(n1286), .CI(n1285), .CO(n1275), .S(n1456)
         );
  FA1D2BWP12T U2117 ( .A(n1290), .B(n1289), .CI(n1288), .CO(n1457), .S(n1437)
         );
  INVD1BWP12T U2118 ( .I(n1437), .ZN(n1304) );
  OAI22D1BWP12T U2119 ( .A1(n2009), .A2(n1292), .B1(n1291), .B2(n2006), .ZN(
        n1401) );
  OAI21D1BWP12T U2120 ( .A1(n1401), .A2(n1404), .B(n1403), .ZN(n1298) );
  CKND2D1BWP12T U2121 ( .A1(n1401), .A2(n1404), .ZN(n1297) );
  ND2D1BWP12T U2122 ( .A1(n1298), .A2(n1297), .ZN(n1438) );
  FA1D0BWP12T U2123 ( .A(n1301), .B(n1300), .CI(n1299), .CO(n1305), .S(n1439)
         );
  NR2D1BWP12T U2124 ( .A1(n1438), .A2(n1439), .ZN(n1303) );
  ND2D1BWP12T U2125 ( .A1(n1438), .A2(n1439), .ZN(n1302) );
  OAI21D1BWP12T U2126 ( .A1(n1304), .A2(n1303), .B(n1302), .ZN(n1476) );
  FA1D1BWP12T U2127 ( .A(n1307), .B(n1306), .CI(n1305), .CO(n1258), .S(n1475)
         );
  FA1D1BWP12T U2128 ( .A(n1310), .B(n1309), .CI(n1308), .CO(n1460), .S(n1442)
         );
  IND2XD1BWP12T U2129 ( .A1(b[0]), .B1(n3173), .ZN(n1311) );
  TPOAI22D1BWP12T U2130 ( .A1(n2127), .A2(n1312), .B1(n2125), .B2(n1311), .ZN(
        n1381) );
  XNR2D1BWP12T U2131 ( .A1(n1979), .A2(n1730), .ZN(n1314) );
  OAI22D1BWP12T U2132 ( .A1(n2127), .A2(n1314), .B1(n2125), .B2(n1313), .ZN(
        n1380) );
  OAI22D1BWP12T U2133 ( .A1(n2013), .A2(n1316), .B1(n2011), .B2(n1315), .ZN(
        n1379) );
  XOR3D2BWP12T U2134 ( .A1(n1322), .A2(n1321), .A3(n1320), .Z(n1492) );
  XNR3D1BWP12T U2135 ( .A1(n1325), .A2(n1324), .A3(n1323), .ZN(n1491) );
  TPND2D1BWP12T U2136 ( .A1(n3456), .A2(n319), .ZN(n2992) );
  IOA21D1BWP12T U2137 ( .A1(n1329), .A2(n1328), .B(n1327), .ZN(n1625) );
  FA1D1BWP12T U2138 ( .A(n1332), .B(n1331), .CI(n1330), .CO(n1605), .S(n1351)
         );
  FA1D1BWP12T U2139 ( .A(n1335), .B(n1334), .CI(n1333), .CO(n1604), .S(n1348)
         );
  FA1D1BWP12T U2140 ( .A(n1338), .B(n1337), .CI(n1336), .CO(n1550), .S(n1330)
         );
  XNR2D1BWP12T U2141 ( .A1(n1339), .A2(n2063), .ZN(n1569) );
  OAI22D1BWP12T U2142 ( .A1(n2062), .A2(n1340), .B1(n1569), .B2(n2059), .ZN(
        n1531) );
  XOR2XD1BWP12T U2143 ( .A1(n2098), .A2(n2064), .Z(n1519) );
  TPOAI22D1BWP12T U2144 ( .A1(n1341), .A2(n2068), .B1(n1519), .B2(n2065), .ZN(
        n1532) );
  XNR2D1BWP12T U2145 ( .A1(n4084), .A2(n3938), .ZN(n1566) );
  OAI22D1BWP12T U2146 ( .A1(n2013), .A2(n1342), .B1(n2011), .B2(n1566), .ZN(
        n1530) );
  XOR3D1BWP12T U2147 ( .A1(n1531), .A2(n1532), .A3(n1530), .Z(n1549) );
  XNR2XD1BWP12T U2148 ( .A1(n3921), .A2(n4157), .ZN(n1525) );
  XNR2XD1BWP12T U2149 ( .A1(n4060), .A2(n4191), .ZN(n1563) );
  OAI22D1BWP12T U2150 ( .A1(n2009), .A2(n1344), .B1(n1563), .B2(n2006), .ZN(
        n1528) );
  XNR2D0BWP12T U2151 ( .A1(n4063), .A2(n3951), .ZN(n1526) );
  OAI22D1BWP12T U2152 ( .A1(n2027), .A2(n1345), .B1(n1986), .B2(n1526), .ZN(
        n1527) );
  FA1D2BWP12T U2153 ( .A(n1348), .B(n1347), .CI(n1346), .CO(n1612), .S(n1329)
         );
  FA1D2BWP12T U2154 ( .A(n1351), .B(n1350), .CI(n1349), .CO(n1613), .S(n1374)
         );
  FA1D0BWP12T U2155 ( .A(n1354), .B(n1353), .CI(n1352), .CO(n1616), .S(n1349)
         );
  FA1D1BWP12T U2156 ( .A(n1357), .B(n1356), .CI(n1355), .CO(n1559), .S(n1353)
         );
  XNR2D1BWP12T U2157 ( .A1(n1977), .A2(n3917), .ZN(n1567) );
  OAI22D1BWP12T U2158 ( .A1(n2019), .A2(n1358), .B1(n1567), .B2(n2018), .ZN(
        n1573) );
  XNR2XD4BWP12T U2159 ( .A1(n4076), .A2(n4157), .ZN(n2003) );
  INR2D1BWP12T U2160 ( .A1(n1979), .B1(n2003), .ZN(n1572) );
  XNR2D0BWP12T U2161 ( .A1(n3885), .A2(n3918), .ZN(n1520) );
  OAI22D1BWP12T U2162 ( .A1(n2072), .A2(n1359), .B1(n2070), .B2(n1520), .ZN(
        n1571) );
  XNR2D1BWP12T U2163 ( .A1(n4082), .A2(n3950), .ZN(n1570) );
  OAI22D1BWP12T U2164 ( .A1(n2130), .A2(n1360), .B1(n754), .B2(n1570), .ZN(
        n1562) );
  XNR2D1BWP12T U2165 ( .A1(n1730), .A2(n3928), .ZN(n1535) );
  OAI22D1BWP12T U2166 ( .A1(n2127), .A2(n1361), .B1(n2125), .B2(n1535), .ZN(
        n1561) );
  HA1D1BWP12T U2167 ( .A(n1363), .B(n1362), .CO(n1560), .S(n1334) );
  FA1D0BWP12T U2168 ( .A(n1369), .B(n1368), .CI(n1367), .CO(n1555), .S(n1354)
         );
  XNR2XD1BWP12T U2169 ( .A1(n4075), .A2(n3941), .ZN(n1524) );
  OAI22D1BWP12T U2170 ( .A1(n2083), .A2(n1370), .B1(n1524), .B2(n2080), .ZN(
        n1523) );
  XNR2D1BWP12T U2171 ( .A1(n1735), .A2(n3927), .ZN(n1536) );
  OAI22D1BWP12T U2172 ( .A1(n2079), .A2(n1371), .B1(n2077), .B2(n1536), .ZN(
        n1522) );
  XNR2XD1BWP12T U2173 ( .A1(n2084), .A2(n3930), .ZN(n1537) );
  OAI22D1BWP12T U2174 ( .A1(n2088), .A2(n1372), .B1(n2086), .B2(n1537), .ZN(
        n1521) );
  XOR3D2BWP12T U2175 ( .A1(n1612), .A2(n1613), .A3(n1610), .Z(n1623) );
  FA1D1BWP12T U2176 ( .A(n1375), .B(n1374), .CI(n1373), .CO(n1512), .S(n1510)
         );
  TPNR2D2BWP12T U2177 ( .A1(n1513), .A2(n1512), .ZN(n2994) );
  TPNR2D1BWP12T U2178 ( .A1(n2992), .A2(n2994), .ZN(n1506) );
  FA1D1BWP12T U2179 ( .A(n1378), .B(n1377), .CI(n1376), .CO(n1445), .S(n1395)
         );
  FA1D1BWP12T U2180 ( .A(n1381), .B(n1380), .CI(n1379), .CO(n1441), .S(n1444)
         );
  FA1D2BWP12T U2181 ( .A(n1384), .B(n1383), .CI(n1382), .CO(n1430), .S(n1376)
         );
  HA1D1BWP12T U2182 ( .A(n1386), .B(n1385), .CO(n1288), .S(n1429) );
  FA1D1BWP12T U2183 ( .A(n1389), .B(n1388), .CI(n1387), .CO(n1428), .S(n1416)
         );
  OAI21D1BWP12T U2184 ( .A1(n1392), .A2(n1391), .B(n1390), .ZN(n1394) );
  ND2D1BWP12T U2185 ( .A1(n1392), .A2(n1391), .ZN(n1393) );
  CKND1BWP12T U2186 ( .I(n1399), .ZN(n1397) );
  CKND1BWP12T U2187 ( .I(n1400), .ZN(n1396) );
  IOA21D1BWP12T U2188 ( .A1(n1397), .A2(n1396), .B(n1395), .ZN(n1398) );
  IOA21D1BWP12T U2189 ( .A1(n1400), .A2(n1399), .B(n1398), .ZN(n1423) );
  INVD1BWP12T U2190 ( .I(n1401), .ZN(n1402) );
  XNR3XD4BWP12T U2191 ( .A1(n1404), .A2(n1403), .A3(n1402), .ZN(n1436) );
  FA1D1BWP12T U2192 ( .A(n1407), .B(n1406), .CI(n1405), .CO(n1435), .S(n1414)
         );
  OAI22D1BWP12T U2193 ( .A1(n2088), .A2(n1409), .B1(n2086), .B2(n1408), .ZN(
        n1433) );
  OAI22D1BWP12T U2194 ( .A1(n2130), .A2(n1411), .B1(n754), .B2(n1410), .ZN(
        n1432) );
  OAI22D1BWP12T U2195 ( .A1(n2027), .A2(n1413), .B1(n2025), .B2(n1412), .ZN(
        n1431) );
  FA1D1BWP12T U2196 ( .A(n1416), .B(n1415), .CI(n1414), .CO(n1424), .S(n1419)
         );
  INVD1BWP12T U2197 ( .I(n1424), .ZN(n1417) );
  XOR3XD4BWP12T U2198 ( .A1(n1423), .A2(n1422), .A3(n1417), .Z(n1448) );
  XNR3XD4BWP12T U2199 ( .A1(n1447), .A2(n1446), .A3(n1448), .ZN(n1450) );
  FA1D1BWP12T U2200 ( .A(n1420), .B(n1419), .CI(n1418), .CO(n1451), .S(n895)
         );
  TPNR2D1BWP12T U2201 ( .A1(n1450), .A2(n1451), .ZN(n1421) );
  ND2D1BWP12T U2202 ( .A1(n3135), .A2(n317), .ZN(n1783) );
  NR2D1BWP12T U2203 ( .A1(n1424), .A2(n1423), .ZN(n1427) );
  INVD1BWP12T U2204 ( .I(n1422), .ZN(n1426) );
  CKND2D1BWP12T U2205 ( .A1(n1424), .A2(n1423), .ZN(n1425) );
  OAI21D1BWP12T U2206 ( .A1(n1427), .A2(n1426), .B(n1425), .ZN(n1490) );
  FA1D1BWP12T U2207 ( .A(n1430), .B(n1429), .CI(n1428), .CO(n1464), .S(n1443)
         );
  FA1D0BWP12T U2208 ( .A(n1433), .B(n1432), .CI(n1431), .CO(n1463), .S(n1434)
         );
  FA1D1BWP12T U2209 ( .A(n1436), .B(n1435), .CI(n1434), .CO(n1462), .S(n1422)
         );
  XOR3D1BWP12T U2210 ( .A1(n1439), .A2(n1438), .A3(n1437), .Z(n1478) );
  FA1D2BWP12T U2211 ( .A(n1442), .B(n1441), .CI(n1440), .CO(n1474), .S(n1479)
         );
  FA1D2BWP12T U2212 ( .A(n1445), .B(n1444), .CI(n1443), .CO(n1477), .S(n1447)
         );
  XOR3D2BWP12T U2213 ( .A1(n1478), .A2(n1479), .A3(n1477), .Z(n1488) );
  TPNR2D1BWP12T U2214 ( .A1(n1453), .A2(n1452), .ZN(n1786) );
  TPNR2D1BWP12T U2215 ( .A1(n1783), .A2(n1786), .ZN(n1455) );
  INVD1P75BWP12T U2216 ( .I(n1449), .ZN(n3133) );
  TPAOI21D1BWP12T U2217 ( .A1(n3135), .A2(n3133), .B(n3136), .ZN(n1784) );
  ND2D1BWP12T U2218 ( .A1(n1453), .A2(n1452), .ZN(n1787) );
  TPOAI21D1BWP12T U2219 ( .A1(n1784), .A2(n1786), .B(n1787), .ZN(n1454) );
  FA1D2BWP12T U2220 ( .A(n1458), .B(n1457), .CI(n1456), .CO(n1472), .S(n1483)
         );
  FA1D1BWP12T U2221 ( .A(n1461), .B(n1460), .CI(n1459), .CO(n1469), .S(n1484)
         );
  INVD1BWP12T U2222 ( .I(n1484), .ZN(n1466) );
  INVD1BWP12T U2223 ( .I(n1483), .ZN(n1465) );
  FA1D2BWP12T U2224 ( .A(n1464), .B(n1463), .CI(n1462), .CO(n1482), .S(n1489)
         );
  IOA21D2BWP12T U2225 ( .A1(n1466), .A2(n1465), .B(n1482), .ZN(n1467) );
  IOA21D2BWP12T U2226 ( .A1(n1483), .A2(n1484), .B(n1467), .ZN(n1496) );
  XOR3D2BWP12T U2227 ( .A1(n1470), .A2(n1469), .A3(n1468), .Z(n1495) );
  FA1D1BWP12T U2228 ( .A(n1473), .B(n1472), .CI(n1471), .CO(n1493), .S(n1494)
         );
  FA1D1BWP12T U2229 ( .A(n1476), .B(n1475), .CI(n1474), .CO(n1471), .S(n1487)
         );
  ND2D1BWP12T U2230 ( .A1(n1479), .A2(n1478), .ZN(n1480) );
  ND2D1BWP12T U2231 ( .A1(n1481), .A2(n1480), .ZN(n1486) );
  NR2D2BWP12T U2232 ( .A1(n1500), .A2(n1499), .ZN(n3091) );
  FA1D1BWP12T U2233 ( .A(n1487), .B(n1486), .CI(n1485), .CO(n1499), .S(n1498)
         );
  FA1D1BWP12T U2234 ( .A(n1490), .B(n1489), .CI(n1488), .CO(n1497), .S(n1453)
         );
  TPNR2D1BWP12T U2235 ( .A1(n3091), .A2(n3089), .ZN(n3045) );
  FA1D1BWP12T U2236 ( .A(n1493), .B(n1492), .CI(n1491), .CO(n1507), .S(n1502)
         );
  FA1D1BWP12T U2237 ( .A(n1496), .B(n1495), .CI(n1494), .CO(n1501), .S(n1500)
         );
  ND2D1BWP12T U2238 ( .A1(n3045), .A2(n321), .ZN(n1505) );
  TPOAI21D1BWP12T U2239 ( .A1(n3091), .A2(n3261), .B(n3092), .ZN(n3044) );
  INVD1BWP12T U2240 ( .I(n3046), .ZN(n1503) );
  TPOAI21D1BWP12T U2241 ( .A1(n3043), .A2(n1505), .B(n1504), .ZN(n3454) );
  ND2D1BWP12T U2242 ( .A1(n1506), .A2(n3454), .ZN(n1515) );
  ND2D1BWP12T U2243 ( .A1(n1508), .A2(n1507), .ZN(n3452) );
  CKND2D2BWP12T U2244 ( .A1(n1510), .A2(n1509), .ZN(n3455) );
  OA21D1BWP12T U2245 ( .A1(n1511), .A2(n3452), .B(n3455), .Z(n2991) );
  ND2D1BWP12T U2246 ( .A1(n1513), .A2(n1512), .ZN(n2995) );
  OA21D1BWP12T U2247 ( .A1(n2991), .A2(n2994), .B(n2995), .Z(n1514) );
  CKND2D2BWP12T U2248 ( .A1(n1515), .A2(n1514), .ZN(n2847) );
  XNR2D1BWP12T U2249 ( .A1(n3897), .A2(n4076), .ZN(n1516) );
  CKXOR2D1BWP12T U2250 ( .A1(n1979), .A2(n3897), .Z(n1518) );
  CKXOR2D1BWP12T U2251 ( .A1(n1517), .A2(n3897), .Z(n1590) );
  OAI22D1BWP12T U2252 ( .A1(n2005), .A2(n1518), .B1(n2003), .B2(n1590), .ZN(
        n1599) );
  CKXOR2D1BWP12T U2253 ( .A1(n3920), .A2(n2064), .Z(n1541) );
  OAI22D1BWP12T U2254 ( .A1(n2068), .A2(n1519), .B1(n1541), .B2(n2065), .ZN(
        n1598) );
  XNR2XD1BWP12T U2255 ( .A1(n4068), .A2(b[25]), .ZN(n1594) );
  OAI22D1BWP12T U2256 ( .A1(n2072), .A2(n1520), .B1(n2070), .B2(n1594), .ZN(
        n1597) );
  FA1D0BWP12T U2257 ( .A(n1523), .B(n1522), .CI(n1521), .CO(n1552), .S(n1554)
         );
  XNR2XD1BWP12T U2258 ( .A1(n4075), .A2(n3943), .ZN(n1542) );
  OAI22D1BWP12T U2259 ( .A1(n2083), .A2(n1524), .B1(n1542), .B2(n2080), .ZN(
        n1576) );
  XNR2XD1BWP12T U2260 ( .A1(n3922), .A2(n4157), .ZN(n1543) );
  OAI22D1BWP12T U2261 ( .A1(n2023), .A2(n1525), .B1(n1543), .B2(n2021), .ZN(
        n1575) );
  XNR2D0BWP12T U2262 ( .A1(n595), .A2(b[19]), .ZN(n1591) );
  OAI22D1BWP12T U2263 ( .A1(n2027), .A2(n1526), .B1(n2025), .B2(n1591), .ZN(
        n1574) );
  FA1D0BWP12T U2264 ( .A(n1529), .B(n1528), .CI(n1527), .CO(n1547), .S(n1548)
         );
  CKND2D1BWP12T U2265 ( .A1(n1532), .A2(n1531), .ZN(n1533) );
  ND2D1BWP12T U2266 ( .A1(n1534), .A2(n1533), .ZN(n1546) );
  XNR2D1BWP12T U2267 ( .A1(n3173), .A2(n3957), .ZN(n1580) );
  OAI22D1BWP12T U2268 ( .A1(n2127), .A2(n1535), .B1(n2125), .B2(n1580), .ZN(
        n1540) );
  XNR2D1BWP12T U2269 ( .A1(a[21]), .A2(n3929), .ZN(n1581) );
  OAI22D1BWP12T U2270 ( .A1(n2079), .A2(n1536), .B1(n2077), .B2(n1581), .ZN(
        n1539) );
  XNR2D1BWP12T U2271 ( .A1(n2084), .A2(n3949), .ZN(n1544) );
  OAI22D1BWP12T U2272 ( .A1(n2088), .A2(n1537), .B1(n2086), .B2(n1544), .ZN(
        n1538) );
  FA1D0BWP12T U2273 ( .A(n1540), .B(n1539), .CI(n1538), .CO(n1635), .S(n1545)
         );
  CKXOR2D1BWP12T U2274 ( .A1(n3927), .A2(n2064), .Z(n1652) );
  OAI22D1BWP12T U2275 ( .A1(n2068), .A2(n1541), .B1(n1652), .B2(n2065), .ZN(
        n1638) );
  XNR2D1BWP12T U2276 ( .A1(n2058), .A2(n3933), .ZN(n1568) );
  XNR2XD1BWP12T U2277 ( .A1(n2058), .A2(n3950), .ZN(n1649) );
  OAI22D1BWP12T U2278 ( .A1(n2062), .A2(n1568), .B1(n1649), .B2(n1648), .ZN(
        n1637) );
  XNR2D1BWP12T U2279 ( .A1(n4084), .A2(n3939), .ZN(n1565) );
  XNR2D1BWP12T U2280 ( .A1(n4084), .A2(n3941), .ZN(n1651) );
  OAI22D1BWP12T U2281 ( .A1(n2013), .A2(n1565), .B1(n2011), .B2(n1651), .ZN(
        n1636) );
  XNR2XD1BWP12T U2282 ( .A1(n4075), .A2(n3918), .ZN(n1674) );
  OAI22D1BWP12T U2283 ( .A1(n2083), .A2(n1542), .B1(n1674), .B2(n2080), .ZN(
        n1670) );
  XNR2XD1BWP12T U2284 ( .A1(n2098), .A2(n4157), .ZN(n1655) );
  OAI22D1BWP12T U2285 ( .A1(n2023), .A2(n1543), .B1(n2021), .B2(n1655), .ZN(
        n1669) );
  XNR2D0BWP12T U2286 ( .A1(n2084), .A2(n4191), .ZN(n1676) );
  OAI22D1BWP12T U2287 ( .A1(n2088), .A2(n1544), .B1(n2086), .B2(n1676), .ZN(
        n1668) );
  FA1D2BWP12T U2288 ( .A(n1547), .B(n1546), .CI(n1545), .CO(n1662), .S(n1608)
         );
  FA1D1BWP12T U2289 ( .A(n1550), .B(n1549), .CI(n1548), .CO(n1607), .S(n1603)
         );
  FA1D0BWP12T U2290 ( .A(n1553), .B(n1552), .CI(n1551), .CO(n1663), .S(n1606)
         );
  FA1D1BWP12T U2291 ( .A(n1556), .B(n1555), .CI(n1554), .CO(n1602), .S(n1614)
         );
  FA1D0BWP12T U2292 ( .A(n1562), .B(n1561), .CI(n1560), .CO(n1585), .S(n1557)
         );
  XNR2D1BWP12T U2293 ( .A1(n4060), .A2(n3952), .ZN(n1589) );
  OAI22D1BWP12T U2294 ( .A1(n2009), .A2(n1563), .B1(n1589), .B2(n2006), .ZN(
        n1579) );
  OR2XD1BWP12T U2295 ( .A1(n1979), .A2(n3897), .Z(n1564) );
  OAI22D1BWP12T U2296 ( .A1(n2005), .A2(n3897), .B1(n2003), .B2(n1564), .ZN(
        n1578) );
  OAI22D1BWP12T U2297 ( .A1(n2013), .A2(n1566), .B1(n2011), .B2(n1565), .ZN(
        n1577) );
  OAI22D1BWP12T U2298 ( .A1(n2019), .A2(n1567), .B1(n1592), .B2(n2018), .ZN(
        n1596) );
  OAI22D2BWP12T U2299 ( .A1(n1650), .A2(n1569), .B1(n1568), .B2(n1648), .ZN(
        n1595) );
  XNR2D1BWP12T U2300 ( .A1(n4082), .A2(n3931), .ZN(n1582) );
  OAI22D1BWP12T U2301 ( .A1(n2130), .A2(n1570), .B1(n754), .B2(n1582), .ZN(
        n1587) );
  FA1D0BWP12T U2302 ( .A(n1573), .B(n1572), .CI(n1571), .CO(n1586), .S(n1558)
         );
  FA1D0BWP12T U2303 ( .A(n1576), .B(n1575), .CI(n1574), .CO(n1685), .S(n1551)
         );
  FA1D1BWP12T U2304 ( .A(n1579), .B(n1578), .CI(n1577), .CO(n1684), .S(n1584)
         );
  XNR2D1BWP12T U2305 ( .A1(a[19]), .A2(n3932), .ZN(n1643) );
  OAI22D1BWP12T U2306 ( .A1(n2127), .A2(n1580), .B1(n2125), .B2(n1643), .ZN(
        n1682) );
  XNR2XD1BWP12T U2307 ( .A1(a[21]), .A2(n3928), .ZN(n1675) );
  OAI22D1BWP12T U2308 ( .A1(n2079), .A2(n1581), .B1(n2077), .B2(n1675), .ZN(
        n1681) );
  XNR2D1BWP12T U2309 ( .A1(n4082), .A2(n3930), .ZN(n1642) );
  OAI22D1BWP12T U2310 ( .A1(n2130), .A2(n1582), .B1(n754), .B2(n1642), .ZN(
        n1680) );
  FA1D0BWP12T U2311 ( .A(n1585), .B(n1584), .CI(n1583), .CO(n1659), .S(n1600)
         );
  FA1D1BWP12T U2312 ( .A(n1588), .B(n1587), .CI(n1586), .CO(n1667), .S(n1583)
         );
  XNR2XD1BWP12T U2313 ( .A1(n4060), .A2(n3951), .ZN(n1656) );
  OAI22D1BWP12T U2314 ( .A1(n2009), .A2(n1589), .B1(n1656), .B2(n2006), .ZN(
        n1673) );
  CKXOR2D1BWP12T U2315 ( .A1(n3921), .A2(n3897), .Z(n1647) );
  OAI22D1BWP12T U2316 ( .A1(n2005), .A2(n1590), .B1(n1647), .B2(n2003), .ZN(
        n1672) );
  XNR2XD1BWP12T U2317 ( .A1(n517), .A2(n3938), .ZN(n1657) );
  OAI22D1BWP12T U2318 ( .A1(n2027), .A2(n1591), .B1(n1986), .B2(n1657), .ZN(
        n1671) );
  XNR2D1BWP12T U2319 ( .A1(n1977), .A2(n3944), .ZN(n1644) );
  OAI22D1BWP12T U2320 ( .A1(n2019), .A2(n1592), .B1(n1644), .B2(n2018), .ZN(
        n1641) );
  XNR2D2BWP12T U2321 ( .A1(n3897), .A2(n3895), .ZN(n2099) );
  NR2D1BWP12T U2322 ( .A1(n2099), .A2(n1593), .ZN(n1640) );
  XNR2D0BWP12T U2323 ( .A1(n3885), .A2(n3917), .ZN(n1654) );
  OAI22D1BWP12T U2324 ( .A1(n2072), .A2(n1594), .B1(n2070), .B2(n1654), .ZN(
        n1639) );
  HA1D1BWP12T U2325 ( .A(n1596), .B(n1595), .CO(n1678), .S(n1588) );
  FA1D0BWP12T U2326 ( .A(n1599), .B(n1598), .CI(n1597), .CO(n1677), .S(n1553)
         );
  FA1D1BWP12T U2327 ( .A(n1602), .B(n1601), .CI(n1600), .CO(n1631), .S(n1619)
         );
  FA1D1BWP12T U2328 ( .A(n1605), .B(n1604), .CI(n1603), .CO(n1618), .S(n1624)
         );
  FA1D1BWP12T U2329 ( .A(n1608), .B(n1607), .CI(n1606), .CO(n1632), .S(n1617)
         );
  INVD1P75BWP12T U2330 ( .I(n1688), .ZN(n1609) );
  XNR3XD4BWP12T U2331 ( .A1(n1687), .A2(n1686), .A3(n1609), .ZN(n1629) );
  OAI21D1BWP12T U2332 ( .A1(n1612), .A2(n1613), .B(n1610), .ZN(n1611) );
  IOA21D1BWP12T U2333 ( .A1(n1613), .A2(n1612), .B(n1611), .ZN(n1622) );
  FA1D1BWP12T U2334 ( .A(n1616), .B(n1615), .CI(n1614), .CO(n1621), .S(n1610)
         );
  FA1D1BWP12T U2335 ( .A(n1619), .B(n1618), .CI(n1617), .CO(n1688), .S(n1620)
         );
  TPNR2D2BWP12T U2336 ( .A1(n1629), .A2(n1628), .ZN(n2694) );
  FA1D1BWP12T U2337 ( .A(n1622), .B(n1621), .CI(n1620), .CO(n1628), .S(n1627)
         );
  FA1D1BWP12T U2338 ( .A(n1625), .B(n1624), .CI(n1623), .CO(n1626), .S(n1513)
         );
  TPNR2D1BWP12T U2339 ( .A1(n1627), .A2(n1626), .ZN(n2692) );
  NR2D1BWP12T U2340 ( .A1(n2694), .A2(n2692), .ZN(n2737) );
  ND2D1BWP12T U2341 ( .A1(n1627), .A2(n1626), .ZN(n2844) );
  CKND2D2BWP12T U2342 ( .A1(n1629), .A2(n1628), .ZN(n2695) );
  TPAOI21D1BWP12T U2343 ( .A1(n2847), .A2(n2737), .B(n2742), .ZN(n1694) );
  FA1D1BWP12T U2344 ( .A(n1632), .B(n1631), .CI(n1630), .CO(n1861), .S(n1686)
         );
  FA1D1BWP12T U2345 ( .A(n1635), .B(n1634), .CI(n1633), .CO(n1919), .S(n1661)
         );
  FA1D2BWP12T U2346 ( .A(n1641), .B(n1640), .CI(n1639), .CO(n1884), .S(n1679)
         );
  XNR2D1BWP12T U2347 ( .A1(n4082), .A2(n3949), .ZN(n1902) );
  OAI22D1BWP12T U2348 ( .A1(n2130), .A2(n1642), .B1(n754), .B2(n1902), .ZN(
        n1916) );
  XNR2D1BWP12T U2349 ( .A1(a[19]), .A2(n3933), .ZN(n1888) );
  OAI22D1BWP12T U2350 ( .A1(n2127), .A2(n1643), .B1(n2125), .B2(n1888), .ZN(
        n1915) );
  XNR2D1BWP12T U2351 ( .A1(n1977), .A2(b[29]), .ZN(n1889) );
  OAI22D1BWP12T U2352 ( .A1(n2019), .A2(n1644), .B1(n1889), .B2(n2018), .ZN(
        n1887) );
  CKXOR2D1BWP12T U2353 ( .A1(a[29]), .A2(n4065), .Z(n1645) );
  CKND2D2BWP12T U2354 ( .A1(n1645), .A2(n2099), .ZN(n1911) );
  IND2D0BWP12T U2355 ( .A1(n1979), .B1(a[29]), .ZN(n1646) );
  OAI22D1BWP12T U2356 ( .A1(n1911), .A2(n3894), .B1(n1646), .B2(n2099), .ZN(
        n1886) );
  OAI22D1BWP12T U2357 ( .A1(n2005), .A2(n1647), .B1(n1906), .B2(n2003), .ZN(
        n1896) );
  XNR2XD1BWP12T U2358 ( .A1(n2058), .A2(n3931), .ZN(n1907) );
  OAI22D1BWP12T U2359 ( .A1(n1650), .A2(n1649), .B1(n1907), .B2(n1648), .ZN(
        n1895) );
  XNR2D1BWP12T U2360 ( .A1(n4084), .A2(n3943), .ZN(n1913) );
  OAI22D1BWP12T U2361 ( .A1(n2013), .A2(n1651), .B1(n2011), .B2(n1913), .ZN(
        n1894) );
  CKXOR2D1BWP12T U2362 ( .A1(n3929), .A2(n2064), .Z(n1910) );
  OAI22D1BWP12T U2363 ( .A1(n2068), .A2(n1652), .B1(n1910), .B2(n2065), .ZN(
        n1899) );
  XNR2XD1BWP12T U2364 ( .A1(n1979), .A2(a[29]), .ZN(n1653) );
  XNR2D1BWP12T U2365 ( .A1(a[29]), .A2(n1962), .ZN(n1912) );
  OAI22D1BWP12T U2366 ( .A1(n1653), .A2(n1911), .B1(n1912), .B2(n2099), .ZN(
        n1898) );
  XNR2XD1BWP12T U2367 ( .A1(n3885), .A2(n3942), .ZN(n1890) );
  OAI22D1BWP12T U2368 ( .A1(n2072), .A2(n1654), .B1(n2070), .B2(n1890), .ZN(
        n1897) );
  XNR2D1BWP12T U2369 ( .A1(n4157), .A2(n3920), .ZN(n1880) );
  OAI22D1BWP12T U2370 ( .A1(n2023), .A2(n1655), .B1(n2021), .B2(n1880), .ZN(
        n1879) );
  XNR2XD1BWP12T U2371 ( .A1(n4060), .A2(b[19]), .ZN(n1881) );
  OAI22D1BWP12T U2372 ( .A1(n2009), .A2(n1656), .B1(n1881), .B2(n2006), .ZN(
        n1878) );
  XNR2D0BWP12T U2373 ( .A1(n595), .A2(n3939), .ZN(n1908) );
  OAI22D1BWP12T U2374 ( .A1(n2027), .A2(n1657), .B1(n2025), .B2(n1908), .ZN(
        n1877) );
  FA1D1BWP12T U2375 ( .A(n1660), .B(n1659), .CI(n1658), .CO(n1867), .S(n1630)
         );
  FA1D1BWP12T U2376 ( .A(n1663), .B(n1662), .CI(n1661), .CO(n1869), .S(n1687)
         );
  INVD1BWP12T U2377 ( .I(n1869), .ZN(n1664) );
  XNR3XD4BWP12T U2378 ( .A1(n1870), .A2(n1867), .A3(n1664), .ZN(n1863) );
  FA1D0BWP12T U2379 ( .A(n1670), .B(n1669), .CI(n1668), .CO(n1893), .S(n1633)
         );
  FA1D0BWP12T U2380 ( .A(n1673), .B(n1672), .CI(n1671), .CO(n1892), .S(n1666)
         );
  XNR2XD1BWP12T U2381 ( .A1(n4075), .A2(b[25]), .ZN(n1900) );
  OAI22D1BWP12T U2382 ( .A1(n2083), .A2(n1674), .B1(n1900), .B2(n2080), .ZN(
        n1876) );
  XNR2XD1BWP12T U2383 ( .A1(a[21]), .A2(n3957), .ZN(n1901) );
  OAI22D1BWP12T U2384 ( .A1(n2079), .A2(n1675), .B1(n2077), .B2(n1901), .ZN(
        n1875) );
  XNR2D0BWP12T U2385 ( .A1(n2084), .A2(n3952), .ZN(n1882) );
  OAI22D1BWP12T U2386 ( .A1(n2088), .A2(n1676), .B1(n2086), .B2(n1882), .ZN(
        n1874) );
  FA1D1BWP12T U2387 ( .A(n1679), .B(n1678), .CI(n1677), .CO(n1873), .S(n1665)
         );
  FA1D0BWP12T U2388 ( .A(n1682), .B(n1681), .CI(n1680), .CO(n1872), .S(n1683)
         );
  FA1D0BWP12T U2389 ( .A(n1685), .B(n1684), .CI(n1683), .CO(n1871), .S(n1660)
         );
  XOR3XD4BWP12T U2390 ( .A1(n1861), .A2(n1863), .A3(n1862), .Z(n1692) );
  CKND2D1BWP12T U2391 ( .A1(n1688), .A2(n1687), .ZN(n1689) );
  ND2D1BWP12T U2392 ( .A1(n1690), .A2(n1689), .ZN(n1691) );
  TPNR2D2BWP12T U2393 ( .A1(n1692), .A2(n1691), .ZN(n2738) );
  INVD1BWP12T U2394 ( .I(n2738), .ZN(n2741) );
  ND2D1BWP12T U2395 ( .A1(n2741), .A2(n2739), .ZN(n1693) );
  XOR2D2BWP12T U2396 ( .A1(n1694), .A2(n1693), .Z(n3450) );
  INVD1BWP12T U2397 ( .I(n3944), .ZN(n3849) );
  INVD1BWP12T U2398 ( .I(n3917), .ZN(n3850) );
  OR2XD1BWP12T U2399 ( .A1(n3197), .A2(n1696), .Z(n1698) );
  NR2D1BWP12T U2400 ( .A1(n1698), .A2(n3193), .ZN(n3147) );
  CKBD1BWP12T U2401 ( .I(a[19]), .Z(n1699) );
  NR2D1BWP12T U2402 ( .A1(n1714), .A2(n1699), .ZN(n3148) );
  NR2D1BWP12T U2403 ( .A1(n3817), .A2(n4069), .ZN(n1806) );
  NR2D1BWP12T U2404 ( .A1(n3148), .A2(n1806), .ZN(n3268) );
  INVD1BWP12T U2405 ( .I(n3939), .ZN(n3818) );
  OR2XD1BWP12T U2406 ( .A1(n3818), .A2(a[21]), .Z(n3278) );
  AN2XD1BWP12T U2407 ( .A1(n3268), .A2(n3278), .Z(n1702) );
  AN2XD1BWP12T U2408 ( .A1(n3147), .A2(n1702), .Z(n1704) );
  OA21D1BWP12T U2409 ( .A1(n1696), .A2(n3198), .B(n1695), .Z(n1697) );
  OAI21D1BWP12T U2410 ( .A1(n1698), .A2(n3194), .B(n1697), .ZN(n3146) );
  ND2D1BWP12T U2411 ( .A1(n1714), .A2(n1699), .ZN(n3149) );
  CKND2D1BWP12T U2412 ( .A1(n3817), .A2(n4069), .ZN(n1807) );
  OAI21D1BWP12T U2413 ( .A1(n1806), .A2(n3149), .B(n1807), .ZN(n3270) );
  CKND2D1BWP12T U2414 ( .A1(n3818), .A2(a[21]), .ZN(n3277) );
  INVD1BWP12T U2415 ( .I(n3277), .ZN(n1700) );
  AO21D1BWP12T U2416 ( .A1(n3270), .A2(n3278), .B(n1700), .Z(n1701) );
  AO21D1BWP12T U2417 ( .A1(n3146), .A2(n1702), .B(n1701), .Z(n1703) );
  AOI21D1BWP12T U2418 ( .A1(n3276), .A2(n1704), .B(n1703), .ZN(n3127) );
  INVD1BWP12T U2419 ( .I(n3941), .ZN(n3815) );
  NR2D1BWP12T U2420 ( .A1(n3815), .A2(n4070), .ZN(n3125) );
  ND2D1BWP12T U2421 ( .A1(n3815), .A2(n4070), .ZN(n3126) );
  TPOAI21D1BWP12T U2422 ( .A1(n3127), .A2(n3125), .B(n3126), .ZN(n3055) );
  INVD1BWP12T U2423 ( .I(n3943), .ZN(n3816) );
  OR2XD1BWP12T U2424 ( .A1(n3816), .A2(a[23]), .Z(n3054) );
  ND2D1BWP12T U2425 ( .A1(n3816), .A2(a[23]), .ZN(n3053) );
  INVD1BWP12T U2426 ( .I(n3053), .ZN(n1705) );
  AOI21D1BWP12T U2427 ( .A1(n3055), .A2(n3054), .B(n1705), .ZN(n2231) );
  INVD1BWP12T U2428 ( .I(n3918), .ZN(n3852) );
  NR2D1BWP12T U2429 ( .A1(n3852), .A2(n4064), .ZN(n2228) );
  ND2D1BWP12T U2430 ( .A1(n3852), .A2(n4064), .ZN(n2229) );
  OAI21D1BWP12T U2431 ( .A1(n2231), .A2(n2228), .B(n2229), .ZN(n3496) );
  INVD1BWP12T U2432 ( .I(b[25]), .ZN(n1706) );
  OR2XD1BWP12T U2433 ( .A1(n1706), .A2(n4157), .Z(n3495) );
  ND2D1BWP12T U2434 ( .A1(n1706), .A2(n4157), .ZN(n3494) );
  INVD1BWP12T U2435 ( .I(n3494), .ZN(n1707) );
  AO21D1BWP12T U2436 ( .A1(n3496), .A2(n3495), .B(n1707), .Z(n3038) );
  INVD1BWP12T U2437 ( .I(b[29]), .ZN(n2169) );
  INVD1BWP12T U2438 ( .I(n1708), .ZN(n3190) );
  ND2D1BWP12T U2439 ( .A1(n3190), .A2(n1712), .ZN(n3142) );
  INVD1BWP12T U2440 ( .I(b[19]), .ZN(n1714) );
  CKBD1BWP12T U2441 ( .I(a[19]), .Z(n1713) );
  ND2D1BWP12T U2442 ( .A1(n3145), .A2(n1801), .ZN(n1717) );
  NR2D1BWP12T U2443 ( .A1(n3142), .A2(n1717), .ZN(n1719) );
  CKND2D1BWP12T U2444 ( .A1(n3186), .A2(n1719), .ZN(n1721) );
  NR2XD0BWP12T U2445 ( .A1(n1721), .A2(n2930), .ZN(n1723) );
  CKND0BWP12T U2446 ( .I(n3189), .ZN(n1711) );
  INVD1BWP12T U2447 ( .I(n1709), .ZN(n1710) );
  AOI21D1BWP12T U2448 ( .A1(n1712), .A2(n1711), .B(n1710), .ZN(n3141) );
  ND2D1BWP12T U2449 ( .A1(n1714), .A2(n1713), .ZN(n3144) );
  INVD1BWP12T U2450 ( .I(n3144), .ZN(n1792) );
  CKND2D1BWP12T U2451 ( .A1(n3817), .A2(n4069), .ZN(n1800) );
  INVD1BWP12T U2452 ( .I(n1800), .ZN(n1715) );
  AOI21D1BWP12T U2453 ( .A1(n1801), .A2(n1792), .B(n1715), .ZN(n1716) );
  TPOAI21D0BWP12T U2454 ( .A1(n3141), .A2(n1717), .B(n1716), .ZN(n1718) );
  TPAOI21D0BWP12T U2455 ( .A1(n3185), .A2(n1719), .B(n1718), .ZN(n1720) );
  TPOAI21D0BWP12T U2456 ( .A1(n2929), .A2(n1721), .B(n1720), .ZN(n1722) );
  NR2XD0BWP12T U2457 ( .A1(n3818), .A2(a[21]), .ZN(n3264) );
  ND2D1BWP12T U2458 ( .A1(n3818), .A2(a[21]), .ZN(n3265) );
  OR2XD1BWP12T U2459 ( .A1(n3815), .A2(n4070), .Z(n3097) );
  CKND2D1BWP12T U2460 ( .A1(n3815), .A2(n4070), .ZN(n3096) );
  INVD1BWP12T U2461 ( .I(n3096), .ZN(n1725) );
  NR2XD0BWP12T U2462 ( .A1(n3816), .A2(a[23]), .ZN(n3049) );
  ND2D1BWP12T U2463 ( .A1(n3816), .A2(a[23]), .ZN(n3050) );
  TPOAI21D1BWP12T U2464 ( .A1(n3052), .A2(n3049), .B(n3050), .ZN(n2227) );
  OR2XD1BWP12T U2465 ( .A1(n3852), .A2(n4064), .Z(n2225) );
  ND2D1BWP12T U2466 ( .A1(n3852), .A2(n4064), .ZN(n2224) );
  INVD1BWP12T U2467 ( .I(n2224), .ZN(n1726) );
  NR2D1BWP12T U2468 ( .A1(n1706), .A2(n4157), .ZN(n3506) );
  ND2D1BWP12T U2469 ( .A1(n1706), .A2(n4157), .ZN(n3507) );
  OR2XD1BWP12T U2470 ( .A1(n3850), .A2(n4076), .Z(n3000) );
  ND2D1BWP12T U2471 ( .A1(n3850), .A2(n4076), .ZN(n2999) );
  INVD1BWP12T U2472 ( .I(n2999), .ZN(n1727) );
  AO21D1BWP12T U2473 ( .A1(n3001), .A2(n3000), .B(n1727), .Z(n2848) );
  OR2XD1BWP12T U2474 ( .A1(n3210), .A2(n1737), .Z(n1729) );
  NR2D1BWP12T U2475 ( .A1(n1729), .A2(n3206), .ZN(n3151) );
  CKBD1BWP12T U2476 ( .I(a[19]), .Z(n1730) );
  NR2D1BWP12T U2477 ( .A1(n1730), .A2(b[19]), .ZN(n3152) );
  NR2D1BWP12T U2478 ( .A1(n3938), .A2(n4069), .ZN(n1812) );
  NR2D1BWP12T U2479 ( .A1(n3152), .A2(n1812), .ZN(n3313) );
  OR2XD1BWP12T U2480 ( .A1(a[21]), .A2(n3939), .Z(n3323) );
  AN2XD1BWP12T U2481 ( .A1(n3313), .A2(n3323), .Z(n1732) );
  AN2XD1BWP12T U2482 ( .A1(n3151), .A2(n1732), .Z(n1734) );
  OA21D1BWP12T U2483 ( .A1(n1737), .A2(n3211), .B(n3159), .Z(n1728) );
  OAI21D1BWP12T U2484 ( .A1(n1729), .A2(n3207), .B(n1728), .ZN(n3150) );
  CKND2D1BWP12T U2485 ( .A1(n1730), .A2(b[19]), .ZN(n3153) );
  ND2D1BWP12T U2486 ( .A1(n3938), .A2(n4069), .ZN(n3303) );
  OAI21D1BWP12T U2487 ( .A1(n1812), .A2(n3153), .B(n3303), .ZN(n3315) );
  CKND2D1BWP12T U2488 ( .A1(a[21]), .A2(n3939), .ZN(n3322) );
  AO21D1BWP12T U2489 ( .A1(n3150), .A2(n1732), .B(n1731), .Z(n1733) );
  AOI21D1BWP12T U2490 ( .A1(n3321), .A2(n1734), .B(n1733), .ZN(n3120) );
  TPNR2D0BWP12T U2491 ( .A1(n3941), .A2(n4070), .ZN(n3118) );
  ND2D1BWP12T U2492 ( .A1(n3941), .A2(n4070), .ZN(n3123) );
  OR2XD1BWP12T U2493 ( .A1(a[23]), .A2(n3943), .Z(n3056) );
  NR2D1BWP12T U2494 ( .A1(n3918), .A2(n4064), .ZN(n2232) );
  ND2D1BWP12T U2495 ( .A1(n3918), .A2(n4064), .ZN(n2241) );
  OAI21D1BWP12T U2496 ( .A1(n2233), .A2(n2232), .B(n2241), .ZN(n4131) );
  INVD1BWP12T U2497 ( .I(n4140), .ZN(n1779) );
  BUFFD1BWP12T U2498 ( .I(a[21]), .Z(n1735) );
  NR2D1BWP12T U2499 ( .A1(n1735), .A2(n3939), .ZN(n3309) );
  CKND2D1BWP12T U2500 ( .A1(n1735), .A2(n3939), .ZN(n3310) );
  OAI21D1BWP12T U2501 ( .A1(n3309), .A2(n3303), .B(n3310), .ZN(n3121) );
  OR2XD1BWP12T U2502 ( .A1(n3941), .A2(n4070), .Z(n3124) );
  CKND0BWP12T U2503 ( .I(n3123), .ZN(n1736) );
  AOI21D1BWP12T U2504 ( .A1(n3121), .A2(n3124), .B(n1736), .ZN(n2234) );
  CKND2D1BWP12T U2505 ( .A1(a[23]), .A2(n3943), .ZN(n3060) );
  INVD1BWP12T U2506 ( .I(n3060), .ZN(n2238) );
  TPND2D0BWP12T U2507 ( .A1(n2234), .A2(n1742), .ZN(n1744) );
  NR2D1BWP12T U2508 ( .A1(n3309), .A2(n1812), .ZN(n3122) );
  ND2D1BWP12T U2509 ( .A1(n3122), .A2(n3124), .ZN(n1740) );
  NR2D1BWP12T U2510 ( .A1(a[19]), .A2(b[19]), .ZN(n3161) );
  OR2XD1BWP12T U2511 ( .A1(n3161), .A2(n1737), .Z(n1739) );
  CKND2D0BWP12T U2512 ( .A1(a[19]), .A2(b[19]), .ZN(n3162) );
  OA21D0BWP12T U2513 ( .A1(n3161), .A2(n3159), .B(n3162), .Z(n1738) );
  OAI21D1BWP12T U2514 ( .A1(n3158), .A2(n1739), .B(n1738), .ZN(n3306) );
  INVD1BWP12T U2515 ( .I(n3306), .ZN(n1817) );
  NR2D1BWP12T U2516 ( .A1(n1739), .A2(n3157), .ZN(n3302) );
  INVD1BWP12T U2517 ( .I(n3302), .ZN(n1818) );
  NR2D1BWP12T U2518 ( .A1(n1818), .A2(n1740), .ZN(n1741) );
  NR2D1BWP12T U2519 ( .A1(a[23]), .A2(n3943), .ZN(n2237) );
  OR2XD1BWP12T U2520 ( .A1(n3918), .A2(n4064), .Z(n2242) );
  AOI21D0BWP12T U2521 ( .A1(n2237), .A2(n1742), .B(n2232), .ZN(n1743) );
  OA31D1BWP12T U2522 ( .A1(n1744), .A2(n3058), .A3(n2236), .B(n1743), .Z(n3565) );
  CKND2D1BWP12T U2523 ( .A1(n3607), .A2(n4206), .ZN(n1778) );
  INVD1BWP12T U2524 ( .I(n4157), .ZN(n3618) );
  ND2D1BWP12T U2525 ( .A1(n3866), .A2(n3867), .ZN(n1745) );
  NR2D1BWP12T U2526 ( .A1(n3172), .A2(n1745), .ZN(n3106) );
  CKND0BWP12T U2527 ( .I(a[21]), .ZN(n1746) );
  ND2D1BWP12T U2528 ( .A1(n1746), .A2(n3865), .ZN(n3107) );
  CKMUX2D1BWP12T U2529 ( .I0(n4157), .I1(n4064), .S(b[0]), .Z(n3781) );
  INVD1BWP12T U2530 ( .I(n3781), .ZN(n3706) );
  CKMUX2D1BWP12T U2531 ( .I0(n4077), .I1(n4076), .S(b[0]), .Z(n2191) );
  MUX2D0BWP12T U2532 ( .I0(a[23]), .I1(n4070), .S(b[0]), .Z(n3783) );
  AOI22D0BWP12T U2533 ( .A1(n3227), .A2(n2191), .B1(n3231), .B2(n3783), .ZN(
        n1748) );
  MUX2XD0BWP12T U2534 ( .I0(a[29]), .I1(n4065), .S(b[0]), .Z(n2190) );
  CKND2D0BWP12T U2535 ( .A1(n3707), .A2(n2190), .ZN(n1747) );
  OAI211D0BWP12T U2536 ( .A1(n3706), .A2(n3703), .B(n1748), .C(n1747), .ZN(
        n1759) );
  MUX2XD0BWP12T U2537 ( .I0(n3868), .I1(n4187), .S(b[0]), .Z(n3240) );
  INVD1BWP12T U2538 ( .I(n3240), .ZN(n3232) );
  MUX2XD0BWP12T U2539 ( .I0(a[19]), .I1(a[18]), .S(b[0]), .Z(n3787) );
  INVD1BWP12T U2540 ( .I(n3787), .ZN(n2859) );
  CKMUX2D1BWP12T U2541 ( .I0(n4082), .I1(a[14]), .S(b[0]), .Z(n3226) );
  INVD1BWP12T U2542 ( .I(n3226), .ZN(n3239) );
  AOI22D0BWP12T U2543 ( .A1(n3227), .A2(n2859), .B1(n3231), .B2(n3239), .ZN(
        n1750) );
  MUX2XD0BWP12T U2544 ( .I0(a[21]), .I1(n4069), .S(b[0]), .Z(n3785) );
  INVD1BWP12T U2545 ( .I(n3785), .ZN(n2864) );
  TPND2D0BWP12T U2546 ( .A1(n3707), .A2(n2864), .ZN(n1749) );
  OAI211D1BWP12T U2547 ( .A1(n3232), .A2(n3703), .B(n1750), .C(n1749), .ZN(
        n3296) );
  INVD1BWP12T U2548 ( .I(n4175), .ZN(n3006) );
  OAI22D1BWP12T U2549 ( .A1(n3703), .A2(n2595), .B1(n2808), .B2(n3704), .ZN(
        n1752) );
  INVD1BWP12T U2550 ( .I(n2823), .ZN(n2809) );
  NR2D1BWP12T U2551 ( .A1(n3005), .A2(n2809), .ZN(n1751) );
  TPNR2D1BWP12T U2552 ( .A1(n1752), .A2(n1751), .ZN(n3295) );
  OAI22D0BWP12T U2553 ( .A1(n3296), .A2(n3006), .B1(n3295), .B2(n2760), .ZN(
        n1758) );
  MUX2XD1BWP12T U2554 ( .I0(n3875), .I1(n3876), .S(b[0]), .Z(n3243) );
  TPNR2D0BWP12T U2555 ( .A1(n3005), .A2(n3243), .ZN(n1755) );
  NR2XD0BWP12T U2556 ( .A1(n3703), .A2(n2807), .ZN(n1754) );
  OAI22D1BWP12T U2557 ( .A1(n3705), .A2(n2805), .B1(n3704), .B2(n3244), .ZN(
        n1753) );
  NR3D1BWP12T U2558 ( .A1(n1755), .A2(n1754), .A3(n1753), .ZN(n3301) );
  INVD1BWP12T U2559 ( .I(n3170), .ZN(n3701) );
  NR2D0BWP12T U2560 ( .A1(n3701), .A2(n2771), .ZN(n1756) );
  ND2D1BWP12T U2561 ( .A1(n1756), .A2(n2547), .ZN(n3234) );
  NR2D0BWP12T U2562 ( .A1(n3301), .A2(n3234), .ZN(n1757) );
  AOI211D1BWP12T U2563 ( .A1(n4179), .A2(n1759), .B(n1758), .C(n1757), .ZN(
        n3667) );
  OAI21D0BWP12T U2564 ( .A1(a[29]), .A2(n4182), .B(n4181), .ZN(n1764) );
  OR2XD1BWP12T U2565 ( .A1(n3019), .A2(n3360), .Z(n3289) );
  CKND2D1BWP12T U2566 ( .A1(n3289), .A2(n3353), .ZN(n2781) );
  AOI22D1BWP12T U2567 ( .A1(n2463), .A2(a[30]), .B1(n2462), .B2(a[29]), .ZN(
        n2621) );
  NR2XD0BWP12T U2568 ( .A1(n2781), .A2(n3682), .ZN(n1763) );
  MUX2ND0BWP12T U2569 ( .I0(n4184), .I1(n2664), .S(b[29]), .ZN(n1760) );
  NR2D0BWP12T U2570 ( .A1(n1760), .A2(n4185), .ZN(n1761) );
  MUX2ND0BWP12T U2571 ( .I0(n1761), .I1(n2205), .S(n3894), .ZN(n1762) );
  AOI211XD0BWP12T U2572 ( .A1(b[29]), .A2(n1764), .B(n1763), .C(n1762), .ZN(
        n1775) );
  NR2D1BWP12T U2573 ( .A1(n3841), .A2(n3922), .ZN(n2778) );
  AOI22D0BWP12T U2574 ( .A1(n3241), .A2(n3243), .B1(n3244), .B2(n3238), .ZN(
        n1766) );
  TPND2D0BWP12T U2575 ( .A1(n2807), .A2(n3242), .ZN(n1765) );
  OAI211D1BWP12T U2576 ( .A1(n2822), .A2(n3786), .B(n1766), .C(n1765), .ZN(
        n3282) );
  INVD1BWP12T U2577 ( .I(n3249), .ZN(n3792) );
  OAI22D0BWP12T U2578 ( .A1(n3787), .A2(n3782), .B1(n3785), .B2(n3780), .ZN(
        n1768) );
  NR2D0BWP12T U2579 ( .A1(n3226), .A2(n3786), .ZN(n1767) );
  RCAOI211D0BWP12T U2580 ( .A1(n3242), .A2(n3240), .B(n1768), .C(n1767), .ZN(
        n3283) );
  OAI22D0BWP12T U2581 ( .A1(n2190), .A2(n3780), .B1(n2191), .B2(n3782), .ZN(
        n1770) );
  OAI22D0BWP12T U2582 ( .A1(n3783), .A2(n3786), .B1(n3781), .B2(n3784), .ZN(
        n1769) );
  INVD1BWP12T U2583 ( .I(n3767), .ZN(n3788) );
  OAI21D0BWP12T U2584 ( .A1(n1770), .A2(n1769), .B(n3788), .ZN(n1771) );
  OAI211D0BWP12T U2585 ( .A1(n3792), .A2(n3283), .B(n3986), .C(n1771), .ZN(
        n1773) );
  NR2D0BWP12T U2586 ( .A1(n2478), .A2(n2780), .ZN(n1772) );
  AOI211D1BWP12T U2587 ( .A1(n2778), .A2(n3282), .B(n1773), .C(n1772), .ZN(
        n3762) );
  OAI22D1BWP12T U2588 ( .A1(n2621), .A2(n3921), .B1(n3241), .B2(n3911), .ZN(
        n2461) );
  CKND2D0BWP12T U2589 ( .A1(n2461), .A2(n4044), .ZN(n2971) );
  CKND2D1BWP12T U2590 ( .A1(n2920), .A2(n2970), .ZN(n4043) );
  INVD1BWP12T U2591 ( .I(n4043), .ZN(n3065) );
  NR2D1BWP12T U2592 ( .A1(n2423), .A2(n4036), .ZN(n4046) );
  AOI21D0BWP12T U2593 ( .A1(n2971), .A2(n3065), .B(n4046), .ZN(n4050) );
  AOI22D1BWP12T U2594 ( .A1(n3762), .A2(n4195), .B1(n4050), .B2(n4011), .ZN(
        n1774) );
  OAI211D1BWP12T U2595 ( .A1(n3667), .A2(n4201), .B(n1775), .C(n1774), .ZN(
        n1776) );
  AOI21D1BWP12T U2596 ( .A1(n3644), .A2(n4203), .B(n1776), .ZN(n1777) );
  OAI211D1BWP12T U2597 ( .A1(n1779), .A2(n4164), .B(n1778), .C(n1777), .ZN(
        n1780) );
  AOI21D1BWP12T U2598 ( .A1(n4215), .A2(n3561), .B(n1780), .ZN(n1781) );
  IOA21D1BWP12T U2599 ( .A1(n4173), .A2(n3503), .B(n1781), .ZN(n1782) );
  ND2D1BWP12T U2600 ( .A1(n1785), .A2(n1784), .ZN(n1790) );
  INVD1BWP12T U2601 ( .I(n1786), .ZN(n1788) );
  CKND2D1BWP12T U2602 ( .A1(n1788), .A2(n1787), .ZN(n1789) );
  XNR2XD1BWP12T U2603 ( .A1(n1790), .A2(n1789), .ZN(n3437) );
  ND2D1BWP12T U2604 ( .A1(n3437), .A2(n4171), .ZN(n1844) );
  CKND0BWP12T U2605 ( .I(n3142), .ZN(n1791) );
  CKND2D1BWP12T U2606 ( .A1(n1791), .A2(n3145), .ZN(n1795) );
  NR2D1BWP12T U2607 ( .A1(n3140), .A2(n1795), .ZN(n1797) );
  ND2XD0BWP12T U2608 ( .A1(n1797), .A2(n3510), .ZN(n1799) );
  CKND0BWP12T U2609 ( .I(n3141), .ZN(n1793) );
  TPAOI21D0BWP12T U2610 ( .A1(n1793), .A2(n3145), .B(n1792), .ZN(n1794) );
  OAI21D1BWP12T U2611 ( .A1(n3143), .A2(n1795), .B(n1794), .ZN(n1796) );
  AOI21D1BWP12T U2612 ( .A1(n3516), .A2(n1797), .B(n1796), .ZN(n1798) );
  OAI21D1BWP12T U2613 ( .A1(n3519), .A2(n1799), .B(n1798), .ZN(n1803) );
  ND2D1BWP12T U2614 ( .A1(n1801), .A2(n1800), .ZN(n1802) );
  XNR2D1BWP12T U2615 ( .A1(n1803), .A2(n1802), .ZN(n3554) );
  INVD1BWP12T U2616 ( .I(n3147), .ZN(n3269) );
  NR2D0BWP12T U2617 ( .A1(n3269), .A2(n3148), .ZN(n1805) );
  INVD0BWP12T U2618 ( .I(n3146), .ZN(n3273) );
  TPOAI21D0BWP12T U2619 ( .A1(n3273), .A2(n3148), .B(n3149), .ZN(n1804) );
  AOI21D1BWP12T U2620 ( .A1(n3276), .A2(n1805), .B(n1804), .ZN(n1809) );
  CKND2D1BWP12T U2621 ( .A1(n1801), .A2(n1807), .ZN(n1808) );
  XOR2XD1BWP12T U2622 ( .A1(n1809), .A2(n1808), .Z(n3475) );
  INVD1BWP12T U2623 ( .I(n3151), .ZN(n3314) );
  NR2D0BWP12T U2624 ( .A1(n3314), .A2(n3152), .ZN(n1811) );
  INVD1BWP12T U2625 ( .I(n3150), .ZN(n3318) );
  OAI21D0BWP12T U2626 ( .A1(n3318), .A2(n3152), .B(n3153), .ZN(n1810) );
  AOI21D1BWP12T U2627 ( .A1(n3321), .A2(n1811), .B(n1810), .ZN(n1814) );
  INVD1BWP12T U2628 ( .I(n1812), .ZN(n3305) );
  CKND2D0BWP12T U2629 ( .A1(n3305), .A2(n3303), .ZN(n1813) );
  XOR2XD1BWP12T U2630 ( .A1(n1814), .A2(n1813), .Z(n4099) );
  CKND0BWP12T U2631 ( .I(n2920), .ZN(n3030) );
  MUX2D1BWP12T U2632 ( .I0(n1815), .I1(n1852), .S(n3921), .Z(n2388) );
  NR2D1BWP12T U2633 ( .A1(n3681), .A2(n2949), .ZN(n1816) );
  AOI21D1BWP12T U2634 ( .A1(n2388), .A2(n4044), .B(n1816), .ZN(n2427) );
  TPOAI21D0BWP12T U2635 ( .A1(n3579), .A2(n1818), .B(n1817), .ZN(n1820) );
  ND2XD0BWP12T U2636 ( .A1(n3305), .A2(n3303), .ZN(n1819) );
  XNR2XD1BWP12T U2637 ( .A1(n1820), .A2(n1819), .ZN(n3572) );
  INVD1BWP12T U2638 ( .I(n2427), .ZN(n3724) );
  MUX2XD0BWP12T U2639 ( .I0(n4069), .I1(a[19]), .S(b[0]), .Z(n3015) );
  NR2D0BWP12T U2640 ( .A1(n3703), .A2(n2775), .ZN(n1822) );
  TPOAI22D0BWP12T U2641 ( .A1(n3705), .A2(n2331), .B1(n3704), .B2(n2772), .ZN(
        n1821) );
  RCAOI211D0BWP12T U2642 ( .A1(n3015), .A2(n3707), .B(n1822), .C(n1821), .ZN(
        n2704) );
  INVD1BWP12T U2643 ( .I(n2704), .ZN(n1830) );
  AOI22D0BWP12T U2644 ( .A1(n3227), .A2(n2255), .B1(n3231), .B2(n1838), .ZN(
        n1824) );
  TPND2D0BWP12T U2645 ( .A1(n3707), .A2(n2295), .ZN(n1823) );
  OAI211D1BWP12T U2646 ( .A1(n2333), .A2(n3703), .B(n1824), .C(n1823), .ZN(
        n2702) );
  CKND2D1BWP12T U2647 ( .A1(n3227), .A2(n1832), .ZN(n1826) );
  CKND2D0BWP12T U2648 ( .A1(n1831), .A2(n2629), .ZN(n1825) );
  CKND2D1BWP12T U2649 ( .A1(n1826), .A2(n1825), .ZN(n1829) );
  NR2D1BWP12T U2650 ( .A1(n3005), .A2(n1827), .ZN(n1828) );
  NR2D1BWP12T U2651 ( .A1(n1829), .A2(n1828), .ZN(n2426) );
  INVD1BWP12T U2652 ( .I(n2426), .ZN(n2710) );
  INVD1BWP12T U2653 ( .I(n3234), .ZN(n4177) );
  AOI222D1BWP12T U2654 ( .A1(n1830), .A2(n4179), .B1(n2702), .B2(n4175), .C1(
        n2710), .C2(n4177), .ZN(n3669) );
  TPND2D0BWP12T U2655 ( .A1(n3293), .A2(n3106), .ZN(n3067) );
  CKXOR2D0BWP12T U2656 ( .A1(n3067), .A2(n4069), .Z(n3628) );
  OAI22D0BWP12T U2657 ( .A1(n3015), .A2(n3780), .B1(n2258), .B2(n3782), .ZN(
        n1835) );
  NR2D0BWP12T U2658 ( .A1(n2296), .A2(n3786), .ZN(n1834) );
  RCAOI211D0BWP12T U2659 ( .A1(n3242), .A2(n2775), .B(n1835), .C(n1834), .ZN(
        n2717) );
  INVD0BWP12T U2660 ( .I(n2717), .ZN(n1839) );
  AOI22D0BWP12T U2661 ( .A1(n3238), .A2(n2330), .B1(n2333), .B2(n3242), .ZN(
        n1837) );
  CKND2D0BWP12T U2662 ( .A1(n2332), .A2(n3241), .ZN(n1836) );
  OAI211D1BWP12T U2663 ( .A1(n1838), .A2(n3786), .B(n1837), .C(n1836), .ZN(
        n2720) );
  AOI22D0BWP12T U2664 ( .A1(n3788), .A2(n1839), .B1(n2720), .B2(n3922), .ZN(
        n1840) );
  ND2D1BWP12T U2665 ( .A1(n3986), .A2(n2780), .ZN(n3770) );
  INVD1BWP12T U2666 ( .I(n3770), .ZN(n3285) );
  OAI211D0BWP12T U2667 ( .A1(n3752), .A2(n3841), .B(n1840), .C(n3285), .ZN(
        n3799) );
  MUX2ND0BWP12T U2668 ( .I0(n4184), .I1(n2664), .S(n3938), .ZN(n1841) );
  AOI21D1BWP12T U2669 ( .A1(n3554), .A2(n4215), .B(n1842), .ZN(n1843) );
  CKND2D2BWP12T U2670 ( .A1(n1844), .A2(n1843), .ZN(result[20]) );
  INR2D1BWP12T U2671 ( .A1(b[0]), .B1(n3782), .ZN(n2633) );
  NR2D1BWP12T U2672 ( .A1(n3782), .A2(b[0]), .ZN(n2630) );
  AOI22D1BWP12T U2673 ( .A1(n1845), .A2(n4083), .B1(n2463), .B2(n4075), .ZN(
        n1847) );
  AOI22D1BWP12T U2674 ( .A1(n2454), .A2(n4084), .B1(n2462), .B2(n4081), .ZN(
        n1846) );
  ND2D1BWP12T U2675 ( .A1(n1847), .A2(n1846), .ZN(n2418) );
  NR2D1BWP12T U2676 ( .A1(n1848), .A2(n2955), .ZN(n3748) );
  OAI22D0BWP12T U2677 ( .A1(n3681), .A2(n2948), .B1(n2420), .B2(n2955), .ZN(
        n1851) );
  NR2D0BWP12T U2678 ( .A1(n1849), .A2(n3356), .ZN(n1850) );
  AO211D1BWP12T U2679 ( .A1(n2641), .A2(n1852), .B(n1851), .C(n1850), .Z(n3717) );
  ND2D1BWP12T U2680 ( .A1(n3717), .A2(n3919), .ZN(n1853) );
  OAI22D1BWP12T U2681 ( .A1(n3674), .A2(n3765), .B1(n1853), .B2(n3655), .ZN(
        n4018) );
  INVD1BWP12T U2682 ( .I(n4018), .ZN(n3974) );
  INVD1BWP12T U2683 ( .I(n1853), .ZN(n3677) );
  CKND0BWP12T U2684 ( .I(n3360), .ZN(n2592) );
  INR2D0BWP12T U2685 ( .A1(n1979), .B1(n2018), .ZN(n3408) );
  XNR2D0BWP12T U2686 ( .A1(n1854), .A2(n4066), .ZN(n3533) );
  INVD1BWP12T U2687 ( .I(n1855), .ZN(n1857) );
  TPNR2D1BWP12T U2688 ( .A1(n2694), .A2(n2738), .ZN(n1924) );
  CKND2D1BWP12T U2689 ( .A1(n1861), .A2(n1863), .ZN(n1866) );
  CKND2D1BWP12T U2690 ( .A1(n1861), .A2(n1862), .ZN(n1865) );
  CKND2D1BWP12T U2691 ( .A1(n1863), .A2(n1862), .ZN(n1864) );
  ND3D1BWP12T U2692 ( .A1(n1866), .A2(n1865), .A3(n1864), .ZN(n1926) );
  OAI21D1BWP12T U2693 ( .A1(n1869), .A2(n1870), .B(n1867), .ZN(n1868) );
  IOA21D1BWP12T U2694 ( .A1(n1870), .A2(n1869), .B(n1868), .ZN(n1934) );
  FA1D1BWP12T U2695 ( .A(n1873), .B(n1872), .CI(n1871), .CO(n1996), .S(n1920)
         );
  FA1D0BWP12T U2696 ( .A(n1876), .B(n1875), .CI(n1874), .CO(n1958), .S(n1891)
         );
  FA1D0BWP12T U2697 ( .A(n1879), .B(n1878), .CI(n1877), .CO(n1957), .S(n1903)
         );
  XNR2XD1BWP12T U2698 ( .A1(n4157), .A2(n3927), .ZN(n1969) );
  OAI22D1BWP12T U2699 ( .A1(n2023), .A2(n1880), .B1(n2021), .B2(n1969), .ZN(
        n1943) );
  XNR2D1BWP12T U2700 ( .A1(n4060), .A2(n3938), .ZN(n1984) );
  OAI22D1BWP12T U2701 ( .A1(n2009), .A2(n1881), .B1(n1984), .B2(n2006), .ZN(
        n1942) );
  XNR2D0BWP12T U2702 ( .A1(n2084), .A2(n3951), .ZN(n1970) );
  OAI22D1BWP12T U2703 ( .A1(n2088), .A2(n1882), .B1(n2086), .B2(n1970), .ZN(
        n1941) );
  FA1D1BWP12T U2704 ( .A(n1885), .B(n1884), .CI(n1883), .CO(n1940), .S(n1918)
         );
  XNR2D1BWP12T U2705 ( .A1(a[19]), .A2(n3950), .ZN(n1947) );
  OAI22D1BWP12T U2706 ( .A1(n2127), .A2(n1888), .B1(n2125), .B2(n1947), .ZN(
        n1992) );
  XNR2D1BWP12T U2707 ( .A1(n1977), .A2(n3940), .ZN(n1978) );
  OAI22D1BWP12T U2708 ( .A1(n2019), .A2(n1889), .B1(n1978), .B2(n2018), .ZN(
        n1976) );
  XNR2D2BWP12T U2709 ( .A1(a[29]), .A2(a[30]), .ZN(n2102) );
  INR2D1BWP12T U2710 ( .A1(n1979), .B1(n2102), .ZN(n1975) );
  XNR2XD1BWP12T U2711 ( .A1(n3885), .A2(n3944), .ZN(n1964) );
  OAI22D1BWP12T U2712 ( .A1(n2072), .A2(n1890), .B1(n2070), .B2(n1964), .ZN(
        n1974) );
  FA1D0BWP12T U2713 ( .A(n1893), .B(n1892), .CI(n1891), .CO(n1938), .S(n1921)
         );
  FA1D2BWP12T U2714 ( .A(n1896), .B(n1895), .CI(n1894), .CO(n1973), .S(n1905)
         );
  XNR2XD1BWP12T U2715 ( .A1(n4075), .A2(n3917), .ZN(n1968) );
  OAI22D0BWP12T U2716 ( .A1(n2083), .A2(n1900), .B1(n1968), .B2(n2080), .ZN(
        n1967) );
  XNR2D1BWP12T U2717 ( .A1(a[21]), .A2(n3932), .ZN(n1948) );
  OAI22D1BWP12T U2718 ( .A1(n2079), .A2(n1901), .B1(n2077), .B2(n1948), .ZN(
        n1966) );
  XNR2D1BWP12T U2719 ( .A1(n4082), .A2(n4191), .ZN(n1949) );
  OAI22D1BWP12T U2720 ( .A1(n2130), .A2(n1902), .B1(n754), .B2(n1949), .ZN(
        n1965) );
  FA1D0BWP12T U2721 ( .A(n1905), .B(n1904), .CI(n1903), .CO(n1951), .S(n1917)
         );
  XOR2D1BWP12T U2722 ( .A1(n3897), .A2(n2098), .Z(n1985) );
  OAI22D1BWP12T U2723 ( .A1(n2005), .A2(n1906), .B1(n1985), .B2(n2003), .ZN(
        n1946) );
  XNR2XD1BWP12T U2724 ( .A1(n2058), .A2(n3930), .ZN(n1988) );
  OAI22D1BWP12T U2725 ( .A1(n2062), .A2(n1907), .B1(n1988), .B2(n2059), .ZN(
        n1945) );
  XNR2D0BWP12T U2726 ( .A1(n506), .A2(n3941), .ZN(n1987) );
  OAI22D1BWP12T U2727 ( .A1(n2027), .A2(n1908), .B1(n2025), .B2(n1987), .ZN(
        n1944) );
  XNR2D1BWP12T U2728 ( .A1(n2064), .A2(n1909), .ZN(n1960) );
  OAI22D1BWP12T U2729 ( .A1(n2068), .A2(n1910), .B1(n1960), .B2(n2065), .ZN(
        n1983) );
  XNR2XD1BWP12T U2730 ( .A1(n3921), .A2(a[29]), .ZN(n1989) );
  OAI22D1BWP12T U2731 ( .A1(n1989), .A2(n2099), .B1(n1912), .B2(n2100), .ZN(
        n1982) );
  XNR2XD1BWP12T U2732 ( .A1(n4084), .A2(n3918), .ZN(n1990) );
  OAI22D1BWP12T U2733 ( .A1(n2013), .A2(n1913), .B1(n2011), .B2(n1990), .ZN(
        n1981) );
  FA1D0BWP12T U2734 ( .A(n1916), .B(n1915), .CI(n1914), .CO(n1953), .S(n1883)
         );
  FA1D2BWP12T U2735 ( .A(n1919), .B(n1918), .CI(n1917), .CO(n1936), .S(n1870)
         );
  TPNR2D2BWP12T U2736 ( .A1(n1926), .A2(n1927), .ZN(n2745) );
  TPNR2D1BWP12T U2737 ( .A1(n2745), .A2(n2692), .ZN(n1923) );
  AN2XD2BWP12T U2738 ( .A1(n1924), .A2(n1923), .Z(n1925) );
  ND2D1BWP12T U2739 ( .A1(n1925), .A2(n2847), .ZN(n1931) );
  NR2D1BWP12T U2740 ( .A1(n2738), .A2(n2745), .ZN(n1929) );
  TPOAI21D1BWP12T U2741 ( .A1(n2745), .A2(n2739), .B(n2746), .ZN(n1928) );
  TPAOI21D1BWP12T U2742 ( .A1(n1929), .A2(n2742), .B(n1928), .ZN(n1930) );
  FA1D2BWP12T U2743 ( .A(n1934), .B(n1933), .CI(n1932), .CO(n1999), .S(n1927)
         );
  INVD1BWP12T U2744 ( .I(n1999), .ZN(n1997) );
  FA1D2BWP12T U2745 ( .A(n1937), .B(n1936), .CI(n1935), .CO(n2153), .S(n1932)
         );
  FA1D0BWP12T U2746 ( .A(n1940), .B(n1939), .CI(n1938), .CO(n2144), .S(n1994)
         );
  FA1D0BWP12T U2747 ( .A(n1943), .B(n1942), .CI(n1941), .CO(n2051), .S(n1956)
         );
  FA1D0BWP12T U2748 ( .A(n1946), .B(n1945), .CI(n1944), .CO(n2050), .S(n1955)
         );
  XNR2D1BWP12T U2749 ( .A1(a[19]), .A2(n3931), .ZN(n2126) );
  OAI22D1BWP12T U2750 ( .A1(n2127), .A2(n1947), .B1(n2125), .B2(n2126), .ZN(
        n2057) );
  XNR2XD1BWP12T U2751 ( .A1(a[21]), .A2(n3933), .ZN(n2078) );
  OAI22D1BWP12T U2752 ( .A1(n2079), .A2(n1948), .B1(n2077), .B2(n2078), .ZN(
        n2056) );
  XNR2XD1BWP12T U2753 ( .A1(n4082), .A2(n3952), .ZN(n2129) );
  TPOAI22D0BWP12T U2754 ( .A1(n2130), .A2(n1949), .B1(n754), .B2(n2129), .ZN(
        n2055) );
  FA1D2BWP12T U2755 ( .A(n1952), .B(n1951), .CI(n1950), .CO(n2142), .S(n1937)
         );
  FA1D0BWP12T U2756 ( .A(n1955), .B(n1954), .CI(n1953), .CO(n2042), .S(n1950)
         );
  FA1D0BWP12T U2757 ( .A(n1958), .B(n1957), .CI(n1956), .CO(n2041), .S(n1995)
         );
  XNR2XD1BWP12T U2758 ( .A1(n2064), .A2(n1959), .ZN(n2067) );
  OAI22D1BWP12T U2759 ( .A1(n2068), .A2(n1960), .B1(n2067), .B2(n2065), .ZN(
        n2121) );
  XNR2XD1BWP12T U2760 ( .A1(n1979), .A2(n4089), .ZN(n1963) );
  XOR2XD1BWP12T U2761 ( .A1(n4089), .A2(a[30]), .Z(n1961) );
  ND2D1BWP12T U2762 ( .A1(n1961), .A2(n2102), .ZN(n2103) );
  XNR2XD1BWP12T U2763 ( .A1(n4089), .A2(n1962), .ZN(n2104) );
  OAI22D1BWP12T U2764 ( .A1(n1963), .A2(n2103), .B1(n2104), .B2(n2102), .ZN(
        n2120) );
  XNR2XD1BWP12T U2765 ( .A1(n4068), .A2(b[29]), .ZN(n2071) );
  OAI22D1BWP12T U2766 ( .A1(n2072), .A2(n1964), .B1(n2070), .B2(n2071), .ZN(
        n2119) );
  FA1D0BWP12T U2767 ( .A(n1967), .B(n1966), .CI(n1965), .CO(n2053), .S(n1971)
         );
  XNR2XD0BWP12T U2768 ( .A1(n4075), .A2(n3942), .ZN(n2082) );
  OAI22D0BWP12T U2769 ( .A1(n2083), .A2(n1968), .B1(n2082), .B2(n2080), .ZN(
        n2124) );
  XNR2D1BWP12T U2770 ( .A1(n4157), .A2(n3929), .ZN(n2022) );
  OAI22D1BWP12T U2771 ( .A1(n2023), .A2(n1969), .B1(n2021), .B2(n2022), .ZN(
        n2123) );
  XNR2D0BWP12T U2772 ( .A1(n2084), .A2(b[19]), .ZN(n2087) );
  OAI22D0BWP12T U2773 ( .A1(n2088), .A2(n1970), .B1(n2086), .B2(n2087), .ZN(
        n2122) );
  FA1D0BWP12T U2774 ( .A(n1973), .B(n1972), .CI(n1971), .CO(n2039), .S(n1952)
         );
  FA1D0BWP12T U2775 ( .A(n1976), .B(n1975), .CI(n1974), .CO(n2033), .S(n1991)
         );
  XNR2D1BWP12T U2776 ( .A1(n1977), .A2(b[31]), .ZN(n2017) );
  OAI22D1BWP12T U2777 ( .A1(n2019), .A2(n1978), .B1(n2017), .B2(n2018), .ZN(
        n2132) );
  IND2D0BWP12T U2778 ( .A1(n1979), .B1(n4089), .ZN(n1980) );
  OAI22D1BWP12T U2779 ( .A1(n2103), .A2(n3395), .B1(n1980), .B2(n2102), .ZN(
        n2131) );
  FA1D2BWP12T U2780 ( .A(n1983), .B(n1982), .CI(n1981), .CO(n2031), .S(n1954)
         );
  XNR2D1BWP12T U2781 ( .A1(n4060), .A2(n3939), .ZN(n2008) );
  OAI22D1BWP12T U2782 ( .A1(n2009), .A2(n1984), .B1(n2008), .B2(n2006), .ZN(
        n2112) );
  XOR2XD1BWP12T U2783 ( .A1(n3897), .A2(n3920), .Z(n2004) );
  OAI22D1BWP12T U2784 ( .A1(n2005), .A2(n1985), .B1(n2003), .B2(n2004), .ZN(
        n2111) );
  XNR2D0BWP12T U2785 ( .A1(n506), .A2(n3943), .ZN(n2026) );
  OAI22D1BWP12T U2786 ( .A1(n2027), .A2(n1987), .B1(n1986), .B2(n2026), .ZN(
        n2110) );
  XNR2D0BWP12T U2787 ( .A1(n2058), .A2(n3949), .ZN(n2061) );
  OAI22D0BWP12T U2788 ( .A1(n2062), .A2(n1988), .B1(n2061), .B2(n2059), .ZN(
        n2109) );
  XNR2XD1BWP12T U2789 ( .A1(n3922), .A2(a[29]), .ZN(n2101) );
  OAI22D1BWP12T U2790 ( .A1(n2101), .A2(n2099), .B1(n1989), .B2(n2100), .ZN(
        n2108) );
  XNR2XD1BWP12T U2791 ( .A1(n4084), .A2(b[25]), .ZN(n2012) );
  OAI22D1BWP12T U2792 ( .A1(n2013), .A2(n1990), .B1(n2011), .B2(n2012), .ZN(
        n2107) );
  FA1D0BWP12T U2793 ( .A(n1993), .B(n1992), .CI(n1991), .CO(n2116), .S(n1939)
         );
  FA1D1BWP12T U2794 ( .A(n1996), .B(n1995), .CI(n1994), .CO(n2046), .S(n1933)
         );
  INR2D1BWP12T U2795 ( .A1(n1997), .B1(n2000), .ZN(n1998) );
  INVD1BWP12T U2796 ( .I(n1998), .ZN(n2161) );
  ND2D1BWP12T U2797 ( .A1(n2000), .A2(n1999), .ZN(n2160) );
  CKND1BWP12T U2798 ( .I(n2160), .ZN(n2001) );
  TPAOI21D1BWP12T U2799 ( .A1(n2163), .A2(n2161), .B(n2001), .ZN(n2159) );
  XOR2D1BWP12T U2800 ( .A1(n3897), .A2(n3927), .Z(n2002) );
  TPOAI22D0BWP12T U2801 ( .A1(n2005), .A2(n2004), .B1(n2003), .B2(n2002), .ZN(
        n2016) );
  XNR2XD0BWP12T U2802 ( .A1(n4060), .A2(n3941), .ZN(n2007) );
  OAI22D1BWP12T U2803 ( .A1(n2009), .A2(n2008), .B1(n2007), .B2(n2006), .ZN(
        n2015) );
  XNR2XD1BWP12T U2804 ( .A1(n4084), .A2(n3917), .ZN(n2010) );
  OAI22D0BWP12T U2805 ( .A1(n2013), .A2(n2012), .B1(n2011), .B2(n2010), .ZN(
        n2014) );
  XOR3D1BWP12T U2806 ( .A1(n2016), .A2(n2015), .A3(n2014), .Z(n2036) );
  AO21D0BWP12T U2807 ( .A1(n2019), .A2(n2018), .B(n2017), .Z(n2030) );
  XNR2D0BWP12T U2808 ( .A1(n4157), .A2(n3928), .ZN(n2020) );
  OAI22D1BWP12T U2809 ( .A1(n2023), .A2(n2022), .B1(n2021), .B2(n2020), .ZN(
        n2029) );
  XNR2XD0BWP12T U2810 ( .A1(n595), .A2(n3918), .ZN(n2024) );
  OAI22D0BWP12T U2811 ( .A1(n2027), .A2(n2026), .B1(n2025), .B2(n2024), .ZN(
        n2028) );
  XOR3D1BWP12T U2812 ( .A1(n2030), .A2(n2029), .A3(n2028), .Z(n2035) );
  FA1D0BWP12T U2813 ( .A(n2033), .B(n2032), .CI(n2031), .CO(n2034), .S(n2038)
         );
  XOR3D1BWP12T U2814 ( .A1(n2036), .A2(n2035), .A3(n2034), .Z(n2045) );
  FA1D0BWP12T U2815 ( .A(n2039), .B(n2038), .CI(n2037), .CO(n2044), .S(n2047)
         );
  FA1D1BWP12T U2816 ( .A(n2042), .B(n2041), .CI(n2040), .CO(n2043), .S(n2048)
         );
  XOR3D1BWP12T U2817 ( .A1(n2045), .A2(n2044), .A3(n2043), .Z(n2150) );
  FA1D0BWP12T U2818 ( .A(n2051), .B(n2050), .CI(n2049), .CO(n2097), .S(n2143)
         );
  FA1D0BWP12T U2819 ( .A(n2057), .B(n2056), .CI(n2055), .CO(n2094), .S(n2049)
         );
  XNR2XD0BWP12T U2820 ( .A1(n2058), .A2(n4191), .ZN(n2060) );
  OAI22D0BWP12T U2821 ( .A1(n2062), .A2(n2061), .B1(n2060), .B2(n2059), .ZN(
        n2075) );
  XNR2D0BWP12T U2822 ( .A1(n2064), .A2(n2063), .ZN(n2066) );
  OAI22D1BWP12T U2823 ( .A1(n2068), .A2(n2067), .B1(n2066), .B2(n2065), .ZN(
        n2074) );
  XNR2D0BWP12T U2824 ( .A1(n3885), .A2(n3940), .ZN(n2069) );
  OAI22D1BWP12T U2825 ( .A1(n2072), .A2(n2071), .B1(n2070), .B2(n2069), .ZN(
        n2073) );
  XOR3D1BWP12T U2826 ( .A1(n2075), .A2(n2074), .A3(n2073), .Z(n2093) );
  XNR2D0BWP12T U2827 ( .A1(a[21]), .A2(n3950), .ZN(n2076) );
  OAI22D1BWP12T U2828 ( .A1(n2079), .A2(n2078), .B1(n2077), .B2(n2076), .ZN(
        n2091) );
  XNR2XD0BWP12T U2829 ( .A1(n4075), .A2(n3944), .ZN(n2081) );
  OAI22D0BWP12T U2830 ( .A1(n2083), .A2(n2082), .B1(n2081), .B2(n2080), .ZN(
        n2090) );
  XNR2D0BWP12T U2831 ( .A1(n2084), .A2(n3938), .ZN(n2085) );
  OAI22D0BWP12T U2832 ( .A1(n2088), .A2(n2087), .B1(n2086), .B2(n2085), .ZN(
        n2089) );
  XOR3D1BWP12T U2833 ( .A1(n2091), .A2(n2090), .A3(n2089), .Z(n2092) );
  XOR3D1BWP12T U2834 ( .A1(n2094), .A2(n2093), .A3(n2092), .Z(n2095) );
  XOR3D1BWP12T U2835 ( .A1(n2097), .A2(n2096), .A3(n2095), .Z(n2147) );
  XNR2D1BWP12T U2836 ( .A1(n2106), .A2(n2105), .ZN(n2115) );
  FA1D0BWP12T U2837 ( .A(n2109), .B(n2108), .CI(n2107), .CO(n2114), .S(n2117)
         );
  FA1D0BWP12T U2838 ( .A(n2112), .B(n2111), .CI(n2110), .CO(n2113), .S(n2118)
         );
  XOR3D1BWP12T U2839 ( .A1(n2115), .A2(n2114), .A3(n2113), .Z(n2141) );
  FA1D0BWP12T U2840 ( .A(n2118), .B(n2117), .CI(n2116), .CO(n2140), .S(n2037)
         );
  FA1D0BWP12T U2841 ( .A(n2121), .B(n2120), .CI(n2119), .CO(n2138), .S(n2054)
         );
  FA1D0BWP12T U2842 ( .A(n2124), .B(n2123), .CI(n2122), .CO(n2137), .S(n2052)
         );
  XNR2D0BWP12T U2843 ( .A1(n4082), .A2(n3951), .ZN(n2128) );
  OAI22D1BWP12T U2844 ( .A1(n2130), .A2(n2129), .B1(n754), .B2(n2128), .ZN(
        n2134) );
  HA1D0BWP12T U2845 ( .A(n2132), .B(n2131), .CO(n2133), .S(n2032) );
  XOR3D1BWP12T U2846 ( .A1(n2135), .A2(n2134), .A3(n2133), .Z(n2136) );
  XOR3D1BWP12T U2847 ( .A1(n2138), .A2(n2137), .A3(n2136), .Z(n2139) );
  XOR3D1BWP12T U2848 ( .A1(n2141), .A2(n2140), .A3(n2139), .Z(n2146) );
  FA1D0BWP12T U2849 ( .A(n2144), .B(n2143), .CI(n2142), .CO(n2145), .S(n2152)
         );
  XOR3D1BWP12T U2850 ( .A1(n2147), .A2(n2146), .A3(n2145), .Z(n2148) );
  XOR3D1BWP12T U2851 ( .A1(n2150), .A2(n2149), .A3(n2148), .Z(n2155) );
  FA1D1BWP12T U2852 ( .A(n2153), .B(n2152), .CI(n2151), .CO(n2154), .S(n2000)
         );
  CKND2D1BWP12T U2853 ( .A1(n2155), .A2(n2154), .ZN(n2157) );
  NR2D1BWP12T U2854 ( .A1(n2155), .A2(n2154), .ZN(n2156) );
  INR2D1BWP12T U2855 ( .A1(n2157), .B1(n2156), .ZN(n2158) );
  XNR2D2BWP12T U2856 ( .A1(n2159), .A2(n2158), .ZN(n3393) );
  ND2D1BWP12T U2857 ( .A1(n2161), .A2(n2160), .ZN(n2162) );
  XNR2D2BWP12T U2858 ( .A1(n2163), .A2(n2162), .ZN(n3451) );
  XNR2D1BWP12T U2859 ( .A1(n3393), .A2(n3451), .ZN(n2178) );
  HA1D1BWP12T U2860 ( .A(n3894), .B(n2164), .CO(n2752), .S(n3644) );
  NR2XD0BWP12T U2861 ( .A1(n2165), .A2(n4089), .ZN(n3399) );
  XNR2D1BWP12T U2862 ( .A1(n2165), .A2(n4089), .ZN(n3660) );
  INVD1BWP12T U2863 ( .I(n3940), .ZN(n3848) );
  INVD1BWP12T U2864 ( .I(n2167), .ZN(n2172) );
  FA1D0BWP12T U2865 ( .A(a[29]), .B(n2169), .CI(n2168), .CO(n2750), .S(n3561)
         );
  INVD1BWP12T U2866 ( .I(n2170), .ZN(n2171) );
  AOI22D1BWP12T U2867 ( .A1(n4173), .A2(n2172), .B1(n2171), .B2(n4215), .ZN(
        n3401) );
  CKND2D0BWP12T U2868 ( .A1(n3395), .A2(n3479), .ZN(n2173) );
  XOR2XD1BWP12T U2869 ( .A1(b[31]), .A2(n4089), .Z(n3905) );
  OAI21D1BWP12T U2870 ( .A1(n4215), .A2(n2173), .B(n3905), .ZN(n2174) );
  AOI21D0BWP12T U2871 ( .A1(n3401), .A2(n4089), .B(n2174), .ZN(n2175) );
  NR2D1BWP12T U2872 ( .A1(n2176), .A2(n2175), .ZN(n2177) );
  CKND2D1BWP12T U2873 ( .A1(n3562), .A2(n4215), .ZN(n2220) );
  FA1D1BWP12T U2874 ( .A(a[29]), .B(b[29]), .CI(n2180), .CO(n2751), .S(n4140)
         );
  FA1D1BWP12T U2875 ( .A(a[29]), .B(b[29]), .CI(n2181), .CO(n2753), .S(n3607)
         );
  INVD1BWP12T U2876 ( .I(n2191), .ZN(n2862) );
  AOI22D0BWP12T U2877 ( .A1(n3227), .A2(n2190), .B1(n3231), .B2(n3781), .ZN(
        n2183) );
  CKND2D0BWP12T U2878 ( .A1(n3707), .A2(a[30]), .ZN(n2182) );
  OAI211D0BWP12T U2879 ( .A1(n2862), .A2(n3703), .B(n2183), .C(n2182), .ZN(
        n2187) );
  TPNR2D0BWP12T U2880 ( .A1(n3005), .A2(n3783), .ZN(n2186) );
  TPNR2D0BWP12T U2881 ( .A1(n3703), .A2(n3787), .ZN(n2185) );
  OAI22D1BWP12T U2882 ( .A1(n3705), .A2(n3232), .B1(n3704), .B2(n3785), .ZN(
        n2184) );
  NR3D1BWP12T U2883 ( .A1(n2186), .A2(n2185), .A3(n2184), .ZN(n3061) );
  INVD1BWP12T U2884 ( .I(n3243), .ZN(n3228) );
  AOI222D1BWP12T U2885 ( .A1(n2187), .A2(n4179), .B1(n3061), .B2(n4175), .C1(
        n3062), .C2(n4177), .ZN(n3741) );
  TPOAI21D0BWP12T U2886 ( .A1(n3064), .A2(n2760), .B(n3741), .ZN(n2213) );
  INVD1BWP12T U2887 ( .I(n3783), .ZN(n2863) );
  AOI22D0BWP12T U2888 ( .A1(n3241), .A2(n2863), .B1(n2864), .B2(n3238), .ZN(
        n2189) );
  AOI22D0BWP12T U2889 ( .A1(n3245), .A2(n3240), .B1(n2859), .B2(n3242), .ZN(
        n2188) );
  ND2D1BWP12T U2890 ( .A1(n2189), .A2(n2188), .ZN(n3072) );
  OAI22D0BWP12T U2891 ( .A1(n3781), .A2(n3786), .B1(n2190), .B2(n3782), .ZN(
        n2193) );
  CKND0BWP12T U2892 ( .I(n2632), .ZN(n2770) );
  OAI22D0BWP12T U2893 ( .A1(n2191), .A2(n3784), .B1(n2770), .B2(a[30]), .ZN(
        n2192) );
  OAI21D0BWP12T U2894 ( .A1(n2193), .A2(n2192), .B(n3788), .ZN(n2194) );
  OAI211D0BWP12T U2895 ( .A1(n4089), .A2(n3710), .B(n2194), .C(n3986), .ZN(
        n2199) );
  OAI22D0BWP12T U2896 ( .A1(n3226), .A2(n3780), .B1(n3228), .B2(n3782), .ZN(
        n2196) );
  OAI22D0BWP12T U2897 ( .A1(n3230), .A2(n3784), .B1(n2821), .B2(n3786), .ZN(
        n2195) );
  NR2D1BWP12T U2898 ( .A1(n2196), .A2(n2195), .ZN(n3074) );
  CKND0BWP12T U2899 ( .I(n2778), .ZN(n2197) );
  OAI22D0BWP12T U2900 ( .A1(n3753), .A2(n2780), .B1(n3074), .B2(n2197), .ZN(
        n2198) );
  AO211D1BWP12T U2901 ( .A1(n3249), .A2(n3072), .B(n2199), .C(n2198), .Z(n3776) );
  INVD1BWP12T U2902 ( .I(n3289), .ZN(n3079) );
  NR2D0BWP12T U2903 ( .A1(n3922), .A2(n3911), .ZN(n2200) );
  ND2D1BWP12T U2904 ( .A1(n2582), .A2(n2200), .ZN(n3680) );
  NR2D1BWP12T U2905 ( .A1(n3079), .A2(n3680), .ZN(n2210) );
  CKND0BWP12T U2906 ( .I(b[31]), .ZN(n2207) );
  CKND2D0BWP12T U2907 ( .A1(n2207), .A2(n2201), .ZN(n2203) );
  AOI22D0BWP12T U2908 ( .A1(n2203), .A2(n2202), .B1(n3910), .B2(n2207), .ZN(
        n2204) );
  MUX2NXD0BWP12T U2909 ( .I0(n2205), .I1(n2204), .S(n4089), .ZN(n2209) );
  CKND2D1BWP12T U2910 ( .A1(n3905), .A2(n2667), .ZN(n2206) );
  OAI21D0BWP12T U2911 ( .A1(n4181), .A2(n2207), .B(n2206), .ZN(n2208) );
  NR3D1BWP12T U2912 ( .A1(n2210), .A2(n2209), .A3(n2208), .ZN(n2211) );
  OAI21D1BWP12T U2913 ( .A1(n3776), .A2(n3773), .B(n2211), .ZN(n2212) );
  AO21D1BWP12T U2914 ( .A1(n4163), .A2(n2213), .B(n2212), .Z(n2214) );
  AOI21D1BWP12T U2915 ( .A1(n3660), .A2(n4203), .B(n2214), .ZN(n2215) );
  IOA21D1BWP12T U2916 ( .A1(n3609), .A2(n4206), .B(n2215), .ZN(n2216) );
  AOI21D1BWP12T U2917 ( .A1(n4210), .A2(n4142), .B(n2216), .ZN(n2219) );
  FA1D1BWP12T U2918 ( .A(n3395), .B(b[31]), .CI(n2217), .CO(n2167), .S(n3505)
         );
  AN3XD2BWP12T U2919 ( .A1(n2220), .A2(n2219), .A3(n2218), .Z(n2221) );
  XNR2XD4BWP12T U2920 ( .A1(n2993), .A2(n2223), .ZN(n3443) );
  ND2XD0BWP12T U2921 ( .A1(n2225), .A2(n2224), .ZN(n2226) );
  XNR2D1BWP12T U2922 ( .A1(n2227), .A2(n2226), .ZN(n3557) );
  CKND2D0BWP12T U2923 ( .A1(n2225), .A2(n2229), .ZN(n2230) );
  XOR2XD1BWP12T U2924 ( .A1(n2231), .A2(n2230), .Z(n3497) );
  INVD0BWP12T U2925 ( .I(n2234), .ZN(n2235) );
  OR2D1BWP12T U2926 ( .A1(n2236), .A2(n2235), .Z(n3059) );
  ND2D1BWP12T U2927 ( .A1(n3059), .A2(n3056), .ZN(n2240) );
  TPAOI21D0BWP12T U2928 ( .A1(n3058), .A2(n3056), .B(n2238), .ZN(n2239) );
  ND2D1BWP12T U2929 ( .A1(n2240), .A2(n2239), .ZN(n2244) );
  CKND2D0BWP12T U2930 ( .A1(n2242), .A2(n2241), .ZN(n2243) );
  XNR2D1BWP12T U2931 ( .A1(n2244), .A2(n2243), .ZN(n3597) );
  INVD1BWP12T U2932 ( .I(n3293), .ZN(n3619) );
  MUX2XD0BWP12T U2933 ( .I0(n4070), .I1(a[21]), .S(b[0]), .Z(n3014) );
  INVD1BWP12T U2934 ( .I(n3014), .ZN(n2774) );
  AOI22D0BWP12T U2935 ( .A1(n3227), .A2(n2774), .B1(n3231), .B2(n2772), .ZN(
        n2247) );
  CKMUX2D1BWP12T U2936 ( .I0(n4064), .I1(a[23]), .S(b[0]), .Z(n3017) );
  INVD1BWP12T U2937 ( .I(n3017), .ZN(n2768) );
  TPND2D0BWP12T U2938 ( .A1(n3707), .A2(n2768), .ZN(n2246) );
  OAI211D1BWP12T U2939 ( .A1(n3015), .A2(n3703), .B(n2247), .C(n2246), .ZN(
        n2253) );
  CKND2D0BWP12T U2940 ( .A1(n2547), .A2(n3170), .ZN(n2250) );
  AOI22D0BWP12T U2941 ( .A1(n3231), .A2(n2255), .B1(n3227), .B2(n2296), .ZN(
        n2249) );
  TPND2D0BWP12T U2942 ( .A1(n3707), .A2(n2756), .ZN(n2248) );
  OAI211D1BWP12T U2943 ( .A1(n3703), .A2(n2332), .B(n2249), .C(n2248), .ZN(
        n4180) );
  OAI22D1BWP12T U2944 ( .A1(n4176), .A2(n2250), .B1(n4180), .B2(n3006), .ZN(
        n2252) );
  TPOAI21D0BWP12T U2945 ( .A1(n2760), .A2(n4178), .B(n3710), .ZN(n2251) );
  AOI211D1BWP12T U2946 ( .A1(n4179), .A2(n2253), .B(n2252), .C(n2251), .ZN(
        n3670) );
  ND2D1BWP12T U2947 ( .A1(n4036), .A2(n4011), .ZN(n3290) );
  INVD1BWP12T U2948 ( .I(n3290), .ZN(n2254) );
  NR2D1BWP12T U2949 ( .A1(n3289), .A2(n2254), .ZN(n4198) );
  OAI22D0BWP12T U2950 ( .A1(n2756), .A2(n3780), .B1(n2296), .B2(n3782), .ZN(
        n2257) );
  NR2D0BWP12T U2951 ( .A1(n2255), .A2(n3786), .ZN(n2256) );
  AOI211D1BWP12T U2952 ( .A1(n3242), .A2(n2332), .B(n2257), .C(n2256), .ZN(
        n3768) );
  NR2D1BWP12T U2953 ( .A1(n3768), .A2(n3792), .ZN(n2263) );
  OAI22D0BWP12T U2954 ( .A1(n3015), .A2(n3784), .B1(n2258), .B2(n3786), .ZN(
        n2260) );
  OAI22D0BWP12T U2955 ( .A1(n3017), .A2(n3780), .B1(n3014), .B2(n3782), .ZN(
        n2259) );
  OAI21D0BWP12T U2956 ( .A1(n2260), .A2(n2259), .B(n3788), .ZN(n2261) );
  OAI211D0BWP12T U2957 ( .A1(n4178), .A2(n2780), .B(n2261), .C(n3986), .ZN(
        n2262) );
  AOI211D1BWP12T U2958 ( .A1(n2778), .A2(n2264), .B(n2263), .C(n2262), .ZN(
        n3808) );
  OAI21D0BWP12T U2959 ( .A1(n4064), .A2(n4182), .B(n4181), .ZN(n2268) );
  MUX2ND0BWP12T U2960 ( .I0(n4184), .I1(n2664), .S(n3918), .ZN(n2265) );
  NR2XD0BWP12T U2961 ( .A1(n2265), .A2(n4185), .ZN(n2266) );
  MUX2ND0BWP12T U2962 ( .I0(n2266), .I1(n2205), .S(n3898), .ZN(n2267) );
  RCAOI21D0BWP12T U2963 ( .A1(n3918), .A2(n2268), .B(n2267), .ZN(n2269) );
  OAI21D1BWP12T U2964 ( .A1(n3065), .A2(n3029), .B(n2269), .ZN(n2270) );
  AOI21D1BWP12T U2965 ( .A1(n3808), .A2(n4195), .B(n2270), .ZN(n2271) );
  OAI21D1BWP12T U2966 ( .A1(n4014), .A2(n4198), .B(n2271), .ZN(n2272) );
  AO21D1BWP12T U2967 ( .A1(n4163), .A2(n3670), .B(n2272), .Z(n2273) );
  AOI21D1BWP12T U2968 ( .A1(n4203), .A2(n3641), .B(n2273), .ZN(n2274) );
  IOA21D1BWP12T U2969 ( .A1(n3597), .A2(n4206), .B(n2274), .ZN(n2275) );
  AOI21D1BWP12T U2970 ( .A1(n4210), .A2(n4133), .B(n2275), .ZN(n2276) );
  IOA21D1BWP12T U2971 ( .A1(n3497), .A2(n4173), .B(n2276), .ZN(n2277) );
  AOI21D1BWP12T U2972 ( .A1(n3557), .A2(n4215), .B(n2277), .ZN(n2278) );
  INVD1BWP12T U2973 ( .I(n2890), .ZN(n2928) );
  OAI21D1BWP12T U2974 ( .A1(n2928), .A2(n2280), .B(n2926), .ZN(n2286) );
  CKND2D1BWP12T U2975 ( .A1(n2282), .A2(n2281), .ZN(n2283) );
  ND2D1BWP12T U2976 ( .A1(n2284), .A2(n2283), .ZN(n2285) );
  XNR2XD2BWP12T U2977 ( .A1(n2286), .A2(n2285), .ZN(n3431) );
  CKND2D1BWP12T U2978 ( .A1(n3431), .A2(n4171), .ZN(n2362) );
  TPND2D0BWP12T U2979 ( .A1(n3510), .A2(n2932), .ZN(n2289) );
  AOI21D1BWP12T U2980 ( .A1(n3516), .A2(n2932), .B(n2287), .ZN(n2288) );
  OAI21D1BWP12T U2981 ( .A1(n3519), .A2(n2289), .B(n2288), .ZN(n2293) );
  CKND2D1BWP12T U2982 ( .A1(n2291), .A2(n2290), .ZN(n2292) );
  XNR2D1BWP12T U2983 ( .A1(n2293), .A2(n2292), .ZN(n3550) );
  AOI22D0BWP12T U2984 ( .A1(n3227), .A2(n2295), .B1(n3231), .B2(n2294), .ZN(
        n2298) );
  TPND2D0BWP12T U2985 ( .A1(n3707), .A2(n2296), .ZN(n2297) );
  OAI211D1BWP12T U2986 ( .A1(n2330), .A2(n3703), .B(n2298), .C(n2297), .ZN(
        n3099) );
  MUX2ND0BWP12T U2987 ( .I0(n3100), .I1(n3099), .S(n2547), .ZN(n2306) );
  MUX2ND0BWP12T U2988 ( .I0(n2299), .I1(n3026), .S(n3921), .ZN(n2300) );
  CKND2D0BWP12T U2989 ( .A1(n2300), .A2(n3841), .ZN(n2303) );
  OAI22D0BWP12T U2990 ( .A1(n3357), .A2(n2955), .B1(n2301), .B2(n3356), .ZN(
        n2302) );
  TPAOI21D0BWP12T U2991 ( .A1(n2303), .A2(n3767), .B(n2302), .ZN(n2315) );
  AOI21D0BWP12T U2992 ( .A1(n2304), .A2(n3353), .B(n3841), .ZN(n2305) );
  NR2D1BWP12T U2993 ( .A1(n2315), .A2(n2305), .ZN(n3989) );
  INVD1BWP12T U2994 ( .I(n3989), .ZN(n2312) );
  OAI21D0BWP12T U2995 ( .A1(n2306), .A2(n3170), .B(n2312), .ZN(n3732) );
  INVD1BWP12T U2996 ( .I(n2401), .ZN(n2958) );
  ND2XD0BWP12T U2997 ( .A1(n2958), .A2(n2907), .ZN(n2308) );
  INVD1BWP12T U2998 ( .I(n2400), .ZN(n2962) );
  AOI21D1BWP12T U2999 ( .A1(n2962), .A2(n2907), .B(n2908), .ZN(n2307) );
  OAI21D1BWP12T U3000 ( .A1(n3388), .A2(n2308), .B(n2307), .ZN(n2310) );
  INVD1BWP12T U3001 ( .I(n2910), .ZN(n2325) );
  CKND2D1BWP12T U3002 ( .A1(n2325), .A2(n2909), .ZN(n2309) );
  XNR2XD1BWP12T U3003 ( .A1(n2310), .A2(n2309), .ZN(n3574) );
  CKND2D1BWP12T U3004 ( .A1(n3574), .A2(n4206), .ZN(n2311) );
  OAI21D1BWP12T U3005 ( .A1(n2978), .A2(n2312), .B(n2311), .ZN(n2313) );
  TPAOI21D0BWP12T U3006 ( .A1(n4163), .A2(n3732), .B(n2313), .ZN(n2359) );
  OAI21D0BWP12T U3007 ( .A1(n2314), .A2(b[3]), .B(n2970), .ZN(n4039) );
  NR2D0BWP12T U3008 ( .A1(n4039), .A2(n3841), .ZN(n2316) );
  OAI31D0BWP12T U3009 ( .A1(n3655), .A2(n2316), .A3(n2315), .B(n3384), .ZN(
        n4030) );
  CKND0BWP12T U3010 ( .I(n2943), .ZN(n2317) );
  NR2D0BWP12T U3011 ( .A1(n2317), .A2(n2945), .ZN(n2322) );
  INVD1BWP12T U3012 ( .I(n2318), .ZN(n2941) );
  ND2XD0BWP12T U3013 ( .A1(n2322), .A2(n2941), .ZN(n2324) );
  INVD1BWP12T U3014 ( .I(n2319), .ZN(n2944) );
  CKND0BWP12T U3015 ( .I(n2942), .ZN(n2320) );
  OAI21D0BWP12T U3016 ( .A1(n2320), .A2(n2945), .B(n2946), .ZN(n2321) );
  AOI21D1BWP12T U3017 ( .A1(n2944), .A2(n2322), .B(n2321), .ZN(n2323) );
  OAI21D1BWP12T U3018 ( .A1(n3379), .A2(n2324), .B(n2323), .ZN(n2327) );
  ND2XD0BWP12T U3019 ( .A1(n2325), .A2(n2909), .ZN(n2326) );
  XNR2D1BWP12T U3020 ( .A1(n2327), .A2(n2326), .ZN(n4095) );
  INVD0BWP12T U3021 ( .I(n2391), .ZN(n2977) );
  NR2D0BWP12T U3022 ( .A1(n2977), .A2(n2917), .ZN(n2328) );
  ND2XD0BWP12T U3023 ( .A1(n2328), .A2(n3351), .ZN(n2329) );
  CKXOR2D0BWP12T U3024 ( .A1(n2329), .A2(a[14]), .Z(n3632) );
  AOI22D0BWP12T U3025 ( .A1(n3241), .A2(n2331), .B1(n2330), .B2(n3242), .ZN(
        n2335) );
  AOI22D0BWP12T U3026 ( .A1(n3245), .A2(n2333), .B1(n2332), .B2(n3238), .ZN(
        n2334) );
  ND2D1BWP12T U3027 ( .A1(n2335), .A2(n2334), .ZN(n2779) );
  INVD1BWP12T U3028 ( .I(n2779), .ZN(n3105) );
  MUX2NXD0BWP12T U3029 ( .I0(n3105), .I1(n3754), .S(n3922), .ZN(n2336) );
  NR2XD0BWP12T U3030 ( .A1(n2336), .A2(n3765), .ZN(n3810) );
  OAI21D0BWP12T U3031 ( .A1(a[14]), .A2(n4182), .B(n4181), .ZN(n2340) );
  MUX2ND0BWP12T U3032 ( .I0(n4184), .I1(n2664), .S(n3930), .ZN(n2337) );
  NR2D0BWP12T U3033 ( .A1(n2337), .A2(n4185), .ZN(n2338) );
  MUX2ND0BWP12T U3034 ( .I0(n2338), .I1(n2205), .S(n3873), .ZN(n2339) );
  RCAOI21D0BWP12T U3035 ( .A1(n3930), .A2(n2340), .B(n2339), .ZN(n2341) );
  IOA21D1BWP12T U3036 ( .A1(n3810), .A2(n4195), .B(n2341), .ZN(n2342) );
  AOI21D1BWP12T U3037 ( .A1(n4203), .A2(n3632), .B(n2342), .ZN(n2343) );
  IOA21D1BWP12T U3038 ( .A1(n4095), .A2(n4210), .B(n2343), .ZN(n2344) );
  AOI21D1BWP12T U3039 ( .A1(n4011), .A2(n4030), .B(n2344), .ZN(n2358) );
  CKND0BWP12T U3040 ( .I(n2937), .ZN(n2345) );
  NR2XD0BWP12T U3041 ( .A1(n2345), .A2(n2939), .ZN(n2350) );
  INVD1BWP12T U3042 ( .I(n2346), .ZN(n2935) );
  CKND2D1BWP12T U3043 ( .A1(n2350), .A2(n2935), .ZN(n2352) );
  INVD1BWP12T U3044 ( .I(n2347), .ZN(n2938) );
  CKND0BWP12T U3045 ( .I(n2936), .ZN(n2348) );
  OAI21D0BWP12T U3046 ( .A1(n2348), .A2(n2939), .B(n2940), .ZN(n2349) );
  AOI21D1BWP12T U3047 ( .A1(n2938), .A2(n2350), .B(n2349), .ZN(n2351) );
  OAI21D1BWP12T U3048 ( .A1(n3345), .A2(n2352), .B(n2351), .ZN(n2356) );
  CKND2D1BWP12T U3049 ( .A1(n2291), .A2(n2354), .ZN(n2355) );
  XNR2XD1BWP12T U3050 ( .A1(n2356), .A2(n2355), .ZN(n3471) );
  CKND2D1BWP12T U3051 ( .A1(n3471), .A2(n4173), .ZN(n2357) );
  ND3D1BWP12T U3052 ( .A1(n2359), .A2(n2358), .A3(n2357), .ZN(n2360) );
  AOI21D1BWP12T U3053 ( .A1(n3550), .A2(n4215), .B(n2360), .ZN(n2361) );
  INVD1BWP12T U3054 ( .I(n2363), .ZN(n2364) );
  AOI21D1BWP12T U3055 ( .A1(n2366), .A2(n2365), .B(n2364), .ZN(n2371) );
  INVD1BWP12T U3056 ( .I(n2367), .ZN(n2369) );
  CKND2D1BWP12T U3057 ( .A1(n2369), .A2(n2368), .ZN(n2370) );
  XOR2XD1BWP12T U3058 ( .A1(n2371), .A2(n2370), .Z(n3421) );
  AOI22D1BWP12T U3059 ( .A1(n4215), .A2(n3527), .B1(n3465), .B2(n4173), .ZN(
        n2408) );
  CKND2D1BWP12T U3060 ( .A1(n2941), .A2(n2382), .ZN(n2384) );
  INVD1BWP12T U3061 ( .I(n2380), .ZN(n2381) );
  AOI21D1BWP12T U3062 ( .A1(n2944), .A2(n2382), .B(n2381), .ZN(n2383) );
  OAI21D1BWP12T U3063 ( .A1(n3379), .A2(n2384), .B(n2383), .ZN(n2387) );
  INVD1BWP12T U3064 ( .I(n2385), .ZN(n2961) );
  CKND2D1BWP12T U3065 ( .A1(n2961), .A2(n2959), .ZN(n2386) );
  XNR2D1BWP12T U3066 ( .A1(n2387), .A2(n2386), .ZN(n4097) );
  MUX2NXD0BWP12T U3067 ( .I0(n2710), .I1(n2702), .S(n2547), .ZN(n2390) );
  OAI21D0BWP12T U3068 ( .A1(n3681), .A2(n2955), .B(n3919), .ZN(n2389) );
  ND2D1BWP12T U3069 ( .A1(n2404), .A2(n2389), .ZN(n3967) );
  OA21D1BWP12T U3070 ( .A1(n2390), .A2(n3170), .B(n3967), .Z(n3739) );
  MAOI22D0BWP12T U3071 ( .A1(n4210), .A2(n4097), .B1(n3739), .B2(n4201), .ZN(
        n2407) );
  INVD1BWP12T U3072 ( .I(n3752), .ZN(n2428) );
  MUX2ND0BWP12T U3073 ( .I0(n2720), .I1(n2428), .S(n3922), .ZN(n2392) );
  CKND2D1BWP12T U3074 ( .A1(n2392), .A2(n3997), .ZN(n3804) );
  MUX2ND0BWP12T U3075 ( .I0(n3364), .I1(n3363), .S(n3950), .ZN(n2393) );
  CKND2D0BWP12T U3076 ( .A1(n2393), .A2(n4181), .ZN(n2394) );
  MUX2NXD0BWP12T U3077 ( .I0(n2394), .I1(n3366), .S(n3876), .ZN(n2397) );
  OAI21D0BWP12T U3078 ( .A1(n4078), .A2(n4182), .B(n4181), .ZN(n2395) );
  TPND2D0BWP12T U3079 ( .A1(n3950), .A2(n2395), .ZN(n2396) );
  OAI211D1BWP12T U3080 ( .A1(n3773), .A2(n3804), .B(n2397), .C(n2396), .ZN(
        n2399) );
  NR2XD0BWP12T U3081 ( .A1(n3967), .A2(n2978), .ZN(n2398) );
  AOI211D1BWP12T U3082 ( .A1(n3626), .A2(n4203), .B(n2399), .C(n2398), .ZN(
        n2406) );
  MUX2NXD0BWP12T U3083 ( .I0(n4089), .I1(n2402), .S(n3353), .ZN(n2713) );
  CKND2D0BWP12T U3084 ( .A1(n2713), .A2(n3919), .ZN(n2403) );
  TPAOI31D0BWP12T U3085 ( .A1(n2404), .A2(n2403), .A3(n3986), .B(n2423), .ZN(
        n4053) );
  MAOI22D0BWP12T U3086 ( .A1(n3576), .A2(n4206), .B1(n4053), .B2(n3029), .ZN(
        n2405) );
  ND4D1BWP12T U3087 ( .A1(n2408), .A2(n2407), .A3(n2406), .A4(n2405), .ZN(
        n2409) );
  AO21D2BWP12T U3088 ( .A1(n3421), .A2(n4171), .B(n2409), .Z(result[12]) );
  OAI211D0BWP12T U3089 ( .A1(n3886), .A2(n2970), .B(n2427), .C(n3919), .ZN(
        n2424) );
  TPAOI21D0BWP12T U3090 ( .A1(n2413), .A2(n2579), .B(n3919), .ZN(n2417) );
  INVD0BWP12T U3091 ( .I(n2414), .ZN(n2415) );
  ND2D0BWP12T U3092 ( .A1(n2415), .A2(n2641), .ZN(n2416) );
  AN2XD1BWP12T U3093 ( .A1(n2417), .A2(n2416), .Z(n2422) );
  TPND2D0BWP12T U3094 ( .A1(n2418), .A2(n3353), .ZN(n2419) );
  OA21D0BWP12T U3095 ( .A1(n2420), .A2(n2948), .B(n2419), .Z(n2421) );
  ND2D1BWP12T U3096 ( .A1(n2422), .A2(n2421), .ZN(n2435) );
  TPAOI31D0BWP12T U3097 ( .A1(n2424), .A2(n3986), .A3(n2435), .B(n2423), .ZN(
        n4054) );
  ND2D0BWP12T U3098 ( .A1(n3724), .A2(n3986), .ZN(n2425) );
  INVD1BWP12T U3099 ( .I(n2435), .ZN(n3720) );
  TPAOI21D0BWP12T U3100 ( .A1(n2425), .A2(n3765), .B(n3720), .ZN(n3968) );
  TPOAI22D1BWP12T U3101 ( .A1(n3720), .A2(n2427), .B1(n2426), .B2(n3711), .ZN(
        n3731) );
  INVD1BWP12T U3102 ( .I(n3731), .ZN(n2442) );
  OAI22D1BWP12T U3103 ( .A1(n320), .A2(n3613), .B1(n2428), .B2(n2675), .ZN(
        n2434) );
  AOI21D1BWP12T U3104 ( .A1(n3893), .A2(n2667), .B(n4185), .ZN(n2432) );
  MUX2ND0BWP12T U3105 ( .I0(n3364), .I1(n3363), .S(n3919), .ZN(n2429) );
  CKND2D0BWP12T U3106 ( .A1(n2429), .A2(n4181), .ZN(n2430) );
  MUX2NXD0BWP12T U3107 ( .I0(n2430), .I1(n3366), .S(n3893), .ZN(n2431) );
  OAI21D0BWP12T U3108 ( .A1(n2432), .A2(n3841), .B(n2431), .ZN(n2433) );
  AOI211D1BWP12T U3109 ( .A1(n3360), .A2(n2435), .B(n2434), .C(n2433), .ZN(
        n2441) );
  INVD1BWP12T U3110 ( .I(n2436), .ZN(n2534) );
  INVD0BWP12T U3111 ( .I(n2437), .ZN(n2439) );
  AOI22D0BWP12T U3112 ( .A1(n4109), .A2(n4210), .B1(n3588), .B2(n4206), .ZN(
        n2440) );
  OAI211D1BWP12T U3113 ( .A1(n2442), .A2(n4201), .B(n2441), .C(n2440), .ZN(
        n2443) );
  AOI21D1BWP12T U3114 ( .A1(n3973), .A2(n3968), .B(n2443), .ZN(n2449) );
  INVD1BWP12T U3115 ( .I(n2444), .ZN(n2537) );
  INVD1BWP12T U3116 ( .I(n2447), .ZN(n2503) );
  RCAOI22D0BWP12T U3117 ( .A1(n4173), .A2(n3483), .B1(n3542), .B2(n4215), .ZN(
        n2448) );
  OAI211D1BWP12T U3118 ( .A1(n4054), .A2(n3029), .B(n2449), .C(n2448), .ZN(
        n2450) );
  AO21D2BWP12T U3119 ( .A1(n3414), .A2(n4171), .B(n2450), .Z(result[4]) );
  ND2D1BWP12T U3120 ( .A1(n318), .A2(n2451), .ZN(n2453) );
  XNR2D1BWP12T U3121 ( .A1(n2453), .A2(n2452), .ZN(n3412) );
  AOI22D0BWP12T U3122 ( .A1(n2454), .A2(n4064), .B1(n2462), .B2(a[21]), .ZN(
        n2458) );
  TPNR2D0BWP12T U3123 ( .A1(n2471), .A2(n3863), .ZN(n2456) );
  NR2XD0BWP12T U3124 ( .A1(n2470), .A2(n3862), .ZN(n2455) );
  NR2D1BWP12T U3125 ( .A1(n2456), .A2(n2455), .ZN(n2457) );
  ND2D1BWP12T U3126 ( .A1(n2458), .A2(n2457), .ZN(n2578) );
  INVD1BWP12T U3127 ( .I(n2578), .ZN(n2950) );
  TPOAI22D0BWP12T U3128 ( .A1(n2469), .A2(n4160), .B1(n2470), .B2(n3896), .ZN(
        n2460) );
  OAI22D1BWP12T U3129 ( .A1(n2471), .A2(n3897), .B1(n2468), .B2(n3895), .ZN(
        n2459) );
  NR2D1BWP12T U3130 ( .A1(n2460), .A2(n2459), .ZN(n3712) );
  INVD1BWP12T U3131 ( .I(n2577), .ZN(n2947) );
  OAI22D1BWP12T U3132 ( .A1(n2469), .A2(n3879), .B1(n2468), .B2(n3876), .ZN(
        n2465) );
  TPOAI22D0BWP12T U3133 ( .A1(n2471), .A2(n3878), .B1(n2470), .B2(n3877), .ZN(
        n2464) );
  NR2D1BWP12T U3134 ( .A1(n2465), .A2(n2464), .ZN(n2812) );
  TPOAI22D0BWP12T U3135 ( .A1(n2947), .A2(n2948), .B1(n2812), .B2(n3356), .ZN(
        n2476) );
  OAI22D1BWP12T U3136 ( .A1(n2469), .A2(n3875), .B1(n2468), .B2(n4187), .ZN(
        n2467) );
  OAI22D1BWP12T U3137 ( .A1(n2471), .A2(n3874), .B1(n2470), .B2(n3873), .ZN(
        n2466) );
  NR2D1BWP12T U3138 ( .A1(n2467), .A2(n2466), .ZN(n2951) );
  OAI21D0BWP12T U3139 ( .A1(n2951), .A2(n2949), .B(n3841), .ZN(n2475) );
  TPOAI22D0BWP12T U3140 ( .A1(n2469), .A2(n3892), .B1(n2468), .B2(n3880), .ZN(
        n2473) );
  OAI22D1BWP12T U3141 ( .A1(n2471), .A2(n3891), .B1(n2470), .B2(n3890), .ZN(
        n2472) );
  NR2D1BWP12T U3142 ( .A1(n2473), .A2(n2472), .ZN(n2585) );
  NR2D0BWP12T U3143 ( .A1(n2585), .A2(n2955), .ZN(n2474) );
  NR3D1BWP12T U3144 ( .A1(n2476), .A2(n2475), .A3(n2474), .ZN(n2494) );
  NR2D1BWP12T U3145 ( .A1(n2494), .A2(n3655), .ZN(n3975) );
  OAI21D0BWP12T U3146 ( .A1(n3288), .A2(n3841), .B(n3975), .ZN(n2477) );
  CKND2D0BWP12T U3147 ( .A1(n2477), .A2(n3384), .ZN(n4023) );
  INVD1BWP12T U3148 ( .I(n2478), .ZN(n3757) );
  CKND2D1BWP12T U3149 ( .A1(n3621), .A2(n4203), .ZN(n2487) );
  OAI21D0BWP12T U3150 ( .A1(n4075), .A2(n4182), .B(n4181), .ZN(n2485) );
  NR2D1BWP12T U3151 ( .A1(n3295), .A2(n2480), .ZN(n2484) );
  MUX2ND0BWP12T U3152 ( .I0(n4184), .I1(n2664), .S(n3920), .ZN(n2481) );
  NR2XD0BWP12T U3153 ( .A1(n2481), .A2(n4185), .ZN(n2482) );
  MUX2ND0BWP12T U3154 ( .I0(n2482), .I1(n2205), .S(n3892), .ZN(n2483) );
  AOI211D1BWP12T U3155 ( .A1(n3920), .A2(n2485), .B(n2484), .C(n2483), .ZN(
        n2486) );
  OAI211D1BWP12T U3156 ( .A1(n3757), .A2(n2675), .B(n2487), .C(n2486), .ZN(
        n2488) );
  AOI21D1BWP12T U3157 ( .A1(n4011), .A2(n4023), .B(n2488), .ZN(n2514) );
  INVD0BWP12T U3158 ( .I(n2491), .ZN(n2493) );
  INVD1BWP12T U3159 ( .I(n2494), .ZN(n3692) );
  INVD1BWP12T U3160 ( .I(n3682), .ZN(n3713) );
  AO21D0BWP12T U3161 ( .A1(n3723), .A2(n4163), .B(n3360), .Z(n2496) );
  AOI22D1BWP12T U3162 ( .A1(n3581), .A2(n4206), .B1(n3692), .B2(n2496), .ZN(
        n2513) );
  NR2D1BWP12T U3163 ( .A1(n3723), .A2(n3841), .ZN(n3981) );
  NR2D1BWP12T U3164 ( .A1(n3981), .A2(n2834), .ZN(n2501) );
  AOI22D1BWP12T U3165 ( .A1(n4107), .A2(n4210), .B1(n3975), .B2(n2501), .ZN(
        n2512) );
  INVD0BWP12T U3166 ( .I(n2509), .ZN(n2511) );
  CKND2D1BWP12T U3167 ( .A1(n2516), .A2(n2515), .ZN(n2518) );
  XNR2D1BWP12T U3168 ( .A1(n2518), .A2(n2517), .ZN(n3409) );
  MUX2NXD0BWP12T U3169 ( .I0(n2520), .I1(n2519), .S(n3921), .ZN(n2521) );
  NR2D1BWP12T U3170 ( .A1(n2521), .A2(b[3]), .ZN(n2572) );
  INVD1BWP12T U3171 ( .I(n2572), .ZN(n2522) );
  OA21D1BWP12T U3172 ( .A1(n2523), .A2(n4044), .B(n2522), .Z(n3725) );
  AOI22D0BWP12T U3173 ( .A1(n4075), .A2(n2630), .B1(n2633), .B2(n4083), .ZN(
        n2527) );
  INVD1BWP12T U3174 ( .I(n2573), .ZN(n2528) );
  OAI21D1BWP12T U3175 ( .A1(n3725), .A2(n3841), .B(n2528), .ZN(n3736) );
  NR2D1BWP12T U3176 ( .A1(n3736), .A2(n2529), .ZN(n2569) );
  INVD1BWP12T U3177 ( .I(n2530), .ZN(n2663) );
  INVD1BWP12T U3178 ( .I(n4206), .ZN(n3582) );
  MOAI22D0BWP12T U3179 ( .A1(n322), .A2(n3582), .B1(n4108), .B2(n4210), .ZN(
        n2567) );
  CKND2D0BWP12T U3180 ( .A1(n2537), .A2(n2536), .ZN(n2538) );
  XNR2XD1BWP12T U3181 ( .A1(n2539), .A2(n2538), .ZN(n3484) );
  INR2D1BWP12T U3182 ( .A1(n3756), .B1(n2675), .ZN(n2540) );
  AOI21D0BWP12T U3183 ( .A1(n3484), .A2(n4173), .B(n2540), .ZN(n2558) );
  CKND0BWP12T U3184 ( .I(n2541), .ZN(n2672) );
  CKND2D0BWP12T U3185 ( .A1(n2586), .A2(n4163), .ZN(n2543) );
  NR2D1BWP12T U3186 ( .A1(n3170), .A2(n2543), .ZN(n2544) );
  IND3D1BWP12T U3187 ( .A1(n3300), .B1(n2544), .B2(n2806), .ZN(n2549) );
  CKND2D0BWP12T U3188 ( .A1(n2824), .A2(n4163), .ZN(n2545) );
  TPNR2D0BWP12T U3189 ( .A1(n3170), .A2(n2545), .ZN(n2546) );
  ND3D0BWP12T U3190 ( .A1(n2547), .A2(n3707), .A3(n2546), .ZN(n2548) );
  CKND2D1BWP12T U3191 ( .A1(n2549), .A2(n2548), .ZN(n2556) );
  CKND0BWP12T U3192 ( .I(n4068), .ZN(n2550) );
  AOI21D0BWP12T U3193 ( .A1(n2667), .A2(n2550), .B(n4185), .ZN(n2554) );
  MUX2ND0BWP12T U3194 ( .I0(n3364), .I1(n3363), .S(b[3]), .ZN(n2551) );
  CKND2D0BWP12T U3195 ( .A1(n2551), .A2(n4181), .ZN(n2552) );
  MUX2NXD0BWP12T U3196 ( .I0(n3366), .I1(n2552), .S(n3885), .ZN(n2553) );
  OAI21D0BWP12T U3197 ( .A1(n2554), .A2(n4044), .B(n2553), .ZN(n2555) );
  AO211D1BWP12T U3198 ( .A1(n3615), .A2(n4203), .B(n2556), .C(n2555), .Z(n2557) );
  INR2D1BWP12T U3199 ( .A1(n2558), .B1(n2557), .ZN(n2566) );
  INVD1BWP12T U3200 ( .I(n2559), .ZN(n2681) );
  OAI21D1BWP12T U3201 ( .A1(n2681), .A2(n2677), .B(n2678), .ZN(n2564) );
  INVD0BWP12T U3202 ( .I(n2560), .ZN(n2562) );
  TPND2D0BWP12T U3203 ( .A1(n2562), .A2(n2561), .ZN(n2563) );
  XNR2XD1BWP12T U3204 ( .A1(n2564), .A2(n2563), .ZN(n3538) );
  ND2D0BWP12T U3205 ( .A1(n3538), .A2(n4215), .ZN(n2565) );
  IND3D1BWP12T U3206 ( .A1(n2567), .B1(n2566), .B2(n2565), .ZN(n2568) );
  AOI211D1BWP12T U3207 ( .A1(n3409), .A2(n4171), .B(n2569), .C(n2568), .ZN(
        n2576) );
  OAI22D0BWP12T U3208 ( .A1(n2570), .A2(n2949), .B1(n4089), .B2(n2948), .ZN(
        n2571) );
  NR2D1BWP12T U3209 ( .A1(n2572), .A2(n2571), .ZN(n3171) );
  AOI21D1BWP12T U3210 ( .A1(n3171), .A2(n3986), .B(n3997), .ZN(n2574) );
  OAI21D1BWP12T U3211 ( .A1(n2574), .A2(n2573), .B(n3384), .ZN(n4019) );
  ND2D1BWP12T U3212 ( .A1(n4019), .A2(n4011), .ZN(n2575) );
  CKND2D2BWP12T U3213 ( .A1(n2576), .A2(n2575), .ZN(result[3]) );
  AOI22D1BWP12T U3214 ( .A1(n2579), .A2(n2578), .B1(n2577), .B2(n3353), .ZN(
        n2623) );
  INVD1BWP12T U3215 ( .I(n2623), .ZN(n2581) );
  AOI21D0BWP12T U3216 ( .A1(n3712), .A2(n3886), .B(n4044), .ZN(n2580) );
  OAI22D1BWP12T U3217 ( .A1(n2581), .A2(n2580), .B1(n2948), .B2(n3713), .ZN(
        n3990) );
  CKND2D1BWP12T U3218 ( .A1(n3990), .A2(n3919), .ZN(n3976) );
  AOI22D1BWP12T U3219 ( .A1(n2630), .A2(n4068), .B1(n2633), .B2(n4081), .ZN(
        n2584) );
  CKND2D0BWP12T U3220 ( .A1(n2582), .A2(n496), .ZN(n2583) );
  AOI21D1BWP12T U3221 ( .A1(n3719), .A2(n3841), .B(n3655), .ZN(n3977) );
  AN3XD1BWP12T U3222 ( .A1(n3976), .A2(n3977), .A3(n3973), .Z(n2627) );
  ND2D1BWP12T U3223 ( .A1(n3707), .A2(n2586), .ZN(n3233) );
  OAI22D1BWP12T U3224 ( .A1(n3990), .A2(n3841), .B1(n3711), .B2(n3233), .ZN(
        n3678) );
  INVD0BWP12T U3225 ( .I(n2587), .ZN(n2589) );
  CKND2D1BWP12T U3226 ( .A1(n2589), .A2(n2588), .ZN(n2591) );
  XOR2XD1BWP12T U3227 ( .A1(n2591), .A2(n2590), .Z(n3534) );
  MOAI22D0BWP12T U3228 ( .A1(n3719), .A2(n2592), .B1(n3534), .B2(n4215), .ZN(
        n2620) );
  INVD1BWP12T U3229 ( .I(n2593), .ZN(n2657) );
  TPND2D0BWP12T U3230 ( .A1(n2589), .A2(n2655), .ZN(n2594) );
  XOR2XD1BWP12T U3231 ( .A1(n2657), .A2(n2594), .Z(n3481) );
  NR2D1BWP12T U3232 ( .A1(n2595), .A2(n3780), .ZN(n3755) );
  TPAOI22D0BWP12T U3233 ( .A1(n3481), .A2(n4173), .B1(n2596), .B2(n3755), .ZN(
        n2618) );
  INVD1BWP12T U3234 ( .I(n3406), .ZN(n2616) );
  INVD1BWP12T U3235 ( .I(n2600), .ZN(n2684) );
  ND2XD0BWP12T U3236 ( .A1(n2604), .A2(n2682), .ZN(n2601) );
  XOR2XD1BWP12T U3237 ( .A1(n2684), .A2(n2601), .Z(n4104) );
  CKND2D0BWP12T U3238 ( .A1(n4104), .A2(n4210), .ZN(n2614) );
  CKND0BWP12T U3239 ( .I(n2602), .ZN(n2604) );
  CKND2D1BWP12T U3240 ( .A1(n2604), .A2(n2603), .ZN(n2606) );
  XOR2XD1BWP12T U3241 ( .A1(n2606), .A2(n2605), .Z(n3584) );
  XNR2XD0BWP12T U3242 ( .A1(n496), .A2(n2018), .ZN(n3614) );
  MUX2ND0BWP12T U3243 ( .I0(n4184), .I1(n2664), .S(n3916), .ZN(n2607) );
  NR2D0BWP12T U3244 ( .A1(n2607), .A2(n4185), .ZN(n2608) );
  MUX2ND0BWP12T U3245 ( .I0(n2608), .I1(n2205), .S(n484), .ZN(n2611) );
  AOI21D0BWP12T U3246 ( .A1(n484), .A2(n2667), .B(n4185), .ZN(n2609) );
  NR2D0BWP12T U3247 ( .A1(n3853), .A2(n2609), .ZN(n2610) );
  RCAOI211D0BWP12T U3248 ( .A1(n3614), .A2(n4203), .B(n2611), .C(n2610), .ZN(
        n2612) );
  IOA21D1BWP12T U3249 ( .A1(n4206), .A2(n3584), .B(n2612), .ZN(n2613) );
  INR2D1BWP12T U3250 ( .A1(n2614), .B1(n2613), .ZN(n2615) );
  OA21D0BWP12T U3251 ( .A1(n2616), .A2(n3407), .B(n2615), .Z(n2617) );
  CKND2D1BWP12T U3252 ( .A1(n2618), .A2(n2617), .ZN(n2619) );
  AOI211D1BWP12T U3253 ( .A1(n4163), .A2(n3678), .B(n2620), .C(n2619), .ZN(
        n2626) );
  MUX2NXD0BWP12T U3254 ( .I0(n3712), .I1(n2621), .S(n3921), .ZN(n2622) );
  AOI21D1BWP12T U3255 ( .A1(n4089), .A2(n3245), .B(n2622), .ZN(n4042) );
  OAI21D1BWP12T U3256 ( .A1(n4042), .A2(n4044), .B(n2623), .ZN(n3215) );
  TPOAI21D0BWP12T U3257 ( .A1(n3215), .A2(n3841), .B(n3977), .ZN(n2624) );
  CKND2D1BWP12T U3258 ( .A1(n2624), .A2(n3384), .ZN(n4020) );
  CKND2D1BWP12T U3259 ( .A1(n4020), .A2(n4011), .ZN(n2625) );
  IND3D1BWP12T U3260 ( .A1(n2627), .B1(n2626), .B2(n2625), .ZN(result[1]) );
  ND2XD0BWP12T U3261 ( .A1(n3992), .A2(n3986), .ZN(n2645) );
  NR2D0BWP12T U3262 ( .A1(n2628), .A2(n3886), .ZN(n2640) );
  OAI21D0BWP12T U3263 ( .A1(n2629), .A2(n4067), .B(n4044), .ZN(n2638) );
  INVD1BWP12T U3264 ( .I(n2630), .ZN(n2631) );
  CKND0BWP12T U3265 ( .I(n4075), .ZN(n2634) );
  INVD1BWP12T U3266 ( .I(n2635), .ZN(n2636) );
  IND3D1BWP12T U3267 ( .A1(n2638), .B1(n2637), .B2(n2636), .ZN(n2639) );
  NR2XD0BWP12T U3268 ( .A1(n2640), .A2(n2639), .ZN(n2644) );
  TPAOI21D0BWP12T U3269 ( .A1(n3354), .A2(n2641), .B(n3919), .ZN(n2642) );
  OAI21D1BWP12T U3270 ( .A1(n3357), .A2(n2948), .B(n2642), .ZN(n2643) );
  TPNR2D1BWP12T U3271 ( .A1(n2644), .A2(n2643), .ZN(n2652) );
  AOI21D1BWP12T U3272 ( .A1(n2645), .A2(n3765), .B(n2652), .ZN(n3969) );
  INVD1BWP12T U3273 ( .I(n3969), .ZN(n2691) );
  AOI21D1BWP12T U3274 ( .A1(n2649), .A2(n3986), .B(n3997), .ZN(n2650) );
  RCOAI21D1BWP12T U3275 ( .A1(n2650), .A2(n2652), .B(n3384), .ZN(n4032) );
  AOI22D1BWP12T U3276 ( .A1(n3411), .A2(n4171), .B1(n4011), .B2(n4032), .ZN(
        n2690) );
  INVD1BWP12T U3277 ( .I(n3018), .ZN(n3676) );
  NR2D1BWP12T U3278 ( .A1(n3676), .A2(n2780), .ZN(n2651) );
  RCAOI211D1BWP12T U3279 ( .A1(n3352), .A2(n2778), .B(n2652), .C(n2651), .ZN(
        n2653) );
  AOI21D1BWP12T U3280 ( .A1(n2654), .A2(n4179), .B(n2653), .ZN(n3729) );
  CKND0BWP12T U3281 ( .I(n2660), .ZN(n2662) );
  MUX2ND0BWP12T U3282 ( .I0(n4184), .I1(n2664), .S(n3921), .ZN(n2665) );
  NR2D0BWP12T U3283 ( .A1(n2665), .A2(n4185), .ZN(n2666) );
  MUX2NXD0BWP12T U3284 ( .I0(n2205), .I1(n2666), .S(n4067), .ZN(n2671) );
  AOI21D0BWP12T U3285 ( .A1(n2668), .A2(n2667), .B(n4185), .ZN(n2669) );
  TPNR2D0BWP12T U3286 ( .A1(n3886), .A2(n2669), .ZN(n2670) );
  AOI211D1BWP12T U3287 ( .A1(n3585), .A2(n4206), .B(n2671), .C(n2670), .ZN(
        n2674) );
  XNR2D0BWP12T U3288 ( .A1(n2672), .A2(n4067), .ZN(n3616) );
  ND2D0BWP12T U3289 ( .A1(n3616), .A2(n4203), .ZN(n2673) );
  OAI211D1BWP12T U3290 ( .A1(n2675), .A2(n3010), .B(n2674), .C(n2673), .ZN(
        n2676) );
  AOI21D1BWP12T U3291 ( .A1(n4173), .A2(n3482), .B(n2676), .ZN(n2688) );
  INVD0BWP12T U3292 ( .I(n2677), .ZN(n2679) );
  CKND2D1BWP12T U3293 ( .A1(n2679), .A2(n2678), .ZN(n2680) );
  XOR2XD1BWP12T U3294 ( .A1(n2681), .A2(n2680), .Z(n3531) );
  AOI22D0BWP12T U3295 ( .A1(n4215), .A2(n3531), .B1(n4105), .B2(n4210), .ZN(
        n2687) );
  OA211D1BWP12T U3296 ( .A1(n3729), .A2(n4201), .B(n2688), .C(n2687), .Z(n2689) );
  OAI211D2BWP12T U3297 ( .A1(n2834), .A2(n2691), .B(n2690), .C(n2689), .ZN(
        result[2]) );
  INVD1BWP12T U3298 ( .I(n2692), .ZN(n2845) );
  INVD1BWP12T U3299 ( .I(n2844), .ZN(n2693) );
  INVD1BWP12T U3300 ( .I(n2694), .ZN(n2696) );
  ND2D1BWP12T U3301 ( .A1(n2696), .A2(n2695), .ZN(n2697) );
  XOR2XD1BWP12T U3302 ( .A1(n2698), .A2(n2697), .Z(n3460) );
  INVD1P75BWP12T U3303 ( .I(n3460), .ZN(n2736) );
  FA1D0BWP12T U3304 ( .A(n3849), .B(n4065), .CI(n2699), .CO(n2166), .S(n3499)
         );
  CKND2D1BWP12T U3305 ( .A1(n3499), .A2(n4173), .ZN(n2734) );
  FA1D0BWP12T U3306 ( .A(n3849), .B(n4065), .CI(n2700), .CO(n2168), .S(n3560)
         );
  CKND2D1BWP12T U3307 ( .A1(n3560), .A2(n4215), .ZN(n2733) );
  FA1D0BWP12T U3308 ( .A(n3944), .B(n4065), .CI(n2701), .CO(n2181), .S(n3602)
         );
  CKND0BWP12T U3309 ( .I(n2760), .ZN(n2711) );
  CKND0BWP12T U3310 ( .I(n2702), .ZN(n2703) );
  OAI22D0BWP12T U3311 ( .A1(n2704), .A2(n3006), .B1(n2703), .B2(n3234), .ZN(
        n2709) );
  CKND2D0BWP12T U3312 ( .A1(n3229), .A2(n3017), .ZN(n2707) );
  CKMUX2D1BWP12T U3313 ( .I0(n4076), .I1(n4157), .S(b[0]), .Z(n3016) );
  AOI22D0BWP12T U3314 ( .A1(n3227), .A2(n3016), .B1(n3231), .B2(n3014), .ZN(
        n2706) );
  MUX2D0BWP12T U3315 ( .I0(n4065), .I1(n4077), .S(b[0]), .Z(n2769) );
  CKND2D0BWP12T U3316 ( .A1(n3707), .A2(n2769), .ZN(n2705) );
  AOI31D1BWP12T U3317 ( .A1(n2707), .A2(n2706), .A3(n2705), .B(n3711), .ZN(
        n2708) );
  AOI211D1BWP12T U3318 ( .A1(n2711), .A2(n2710), .B(n2709), .C(n2708), .ZN(
        n3742) );
  HA1D1BWP12T U3319 ( .A(n3895), .B(n2712), .CO(n2164), .S(n3646) );
  ND2D1BWP12T U3320 ( .A1(n3646), .A2(n4203), .ZN(n2728) );
  AOI21D0BWP12T U3321 ( .A1(n2713), .A2(n2920), .B(n4046), .ZN(n4017) );
  OAI22D0BWP12T U3322 ( .A1(n3014), .A2(n3786), .B1(n2769), .B2(n3780), .ZN(
        n2715) );
  OAI22D0BWP12T U3323 ( .A1(n3017), .A2(n3784), .B1(n3016), .B2(n3782), .ZN(
        n2714) );
  OAI21D0BWP12T U3324 ( .A1(n2715), .A2(n2714), .B(n3788), .ZN(n2716) );
  OAI211D0BWP12T U3325 ( .A1(n2717), .A2(n3792), .B(n2716), .C(n3986), .ZN(
        n2719) );
  NR2D0BWP12T U3326 ( .A1(n3752), .A2(n2780), .ZN(n2718) );
  AOI211XD0BWP12T U3327 ( .A1(n2720), .A2(n2778), .B(n2719), .C(n2718), .ZN(
        n3763) );
  MOAI22D0BWP12T U3328 ( .A1(n2781), .A2(n3681), .B1(n4195), .B2(n3763), .ZN(
        n2726) );
  OAI21D0BWP12T U3329 ( .A1(n4065), .A2(n4182), .B(n4181), .ZN(n2724) );
  MUX2ND0BWP12T U3330 ( .I0(n4184), .I1(n2664), .S(n3944), .ZN(n2721) );
  NR2D0BWP12T U3331 ( .A1(n2721), .A2(n4185), .ZN(n2722) );
  MUX2ND0BWP12T U3332 ( .I0(n2722), .I1(n2205), .S(n3895), .ZN(n2723) );
  AO21D0BWP12T U3333 ( .A1(n3944), .A2(n2724), .B(n2723), .Z(n2725) );
  RCAOI211D0BWP12T U3334 ( .A1(n4017), .A2(n4011), .B(n2726), .C(n2725), .ZN(
        n2727) );
  OAI211D1BWP12T U3335 ( .A1(n3742), .A2(n4201), .B(n2728), .C(n2727), .ZN(
        n2729) );
  AOI21D1BWP12T U3336 ( .A1(n3602), .A2(n4206), .B(n2729), .ZN(n2732) );
  FA1D1BWP12T U3337 ( .A(n3944), .B(n4065), .CI(n2730), .CO(n2180), .S(n4135)
         );
  CKND2D1BWP12T U3338 ( .A1(n4135), .A2(n4210), .ZN(n2731) );
  AN4XD1BWP12T U3339 ( .A1(n2734), .A2(n2733), .A3(n2732), .A4(n2731), .Z(
        n2735) );
  TPOAI21D2BWP12T U3340 ( .A1(n2736), .A2(n3407), .B(n2735), .ZN(result[28])
         );
  IND3D1BWP12T U3341 ( .A1(n2738), .B1(n2737), .B2(n2847), .ZN(n2744) );
  INVD1BWP12T U3342 ( .I(n2739), .ZN(n2740) );
  AOI21D1BWP12T U3343 ( .A1(n2742), .A2(n2741), .B(n2740), .ZN(n2743) );
  ND2D1BWP12T U3344 ( .A1(n2744), .A2(n2743), .ZN(n2749) );
  INVD1BWP12T U3345 ( .I(n2745), .ZN(n2747) );
  ND2D1BWP12T U3346 ( .A1(n2747), .A2(n2746), .ZN(n2748) );
  XNR2XD4BWP12T U3347 ( .A1(n2749), .A2(n2748), .ZN(n3403) );
  FA1D1BWP12T U3348 ( .A(n3848), .B(a[30]), .CI(n2750), .CO(n2179), .S(n3563)
         );
  FA1D1BWP12T U3349 ( .A(n3940), .B(a[30]), .CI(n2751), .CO(n3397), .S(n4141)
         );
  INVD1BWP12T U3350 ( .I(n3662), .ZN(n2787) );
  FA1D1BWP12T U3351 ( .A(n3940), .B(a[30]), .CI(n2753), .CO(n3394), .S(n3608)
         );
  CKND2D1BWP12T U3352 ( .A1(n3608), .A2(n4206), .ZN(n2786) );
  INVD1BWP12T U3353 ( .I(n3016), .ZN(n2767) );
  AOI22D0BWP12T U3354 ( .A1(n3227), .A2(n2769), .B1(n3231), .B2(n3017), .ZN(
        n2755) );
  CKND2D0BWP12T U3355 ( .A1(n3707), .A2(a[29]), .ZN(n2754) );
  OAI211D0BWP12T U3356 ( .A1(n2767), .A2(n3703), .B(n2755), .C(n2754), .ZN(
        n2759) );
  AOI22D0BWP12T U3357 ( .A1(n3227), .A2(n3015), .B1(n3231), .B2(n2756), .ZN(
        n2758) );
  TPND2D0BWP12T U3358 ( .A1(n3707), .A2(n3014), .ZN(n2757) );
  OAI211D1BWP12T U3359 ( .A1(n2772), .A2(n3703), .B(n2758), .C(n2757), .ZN(
        n3101) );
  AOI222D0BWP12T U3360 ( .A1(n2759), .A2(n4179), .B1(n3101), .B2(n4175), .C1(
        n3099), .C2(n4177), .ZN(n3666) );
  OAI21D0BWP12T U3361 ( .A1(n3688), .A2(n2760), .B(n3666), .ZN(n2784) );
  INVD1BWP12T U3362 ( .I(n4039), .ZN(n2766) );
  OAI21D0BWP12T U3363 ( .A1(a[30]), .A2(n4182), .B(n4181), .ZN(n2764) );
  NR2D1BWP12T U3364 ( .A1(n2920), .A2(n3029), .ZN(n3216) );
  MUX2ND0BWP12T U3365 ( .I0(n4184), .I1(n2664), .S(n3940), .ZN(n2761) );
  NR2D0BWP12T U3366 ( .A1(n2761), .A2(n4185), .ZN(n2762) );
  MUX2NXD0BWP12T U3367 ( .I0(n2762), .I1(n2205), .S(n3899), .ZN(n2763) );
  AOI211XD0BWP12T U3368 ( .A1(n3940), .A2(n2764), .B(n3216), .C(n2763), .ZN(
        n2765) );
  OAI21D1BWP12T U3369 ( .A1(n2766), .A2(n3290), .B(n2765), .ZN(n2783) );
  CKND2D0BWP12T U3370 ( .A1(n2771), .A2(n3899), .ZN(n3658) );
  INVD0BWP12T U3371 ( .I(n3015), .ZN(n2773) );
  AOI22D0BWP12T U3372 ( .A1(n3238), .A2(n2773), .B1(n2772), .B2(n3242), .ZN(
        n2777) );
  AOI22D0BWP12T U3373 ( .A1(n3245), .A2(n2775), .B1(n2774), .B2(n3241), .ZN(
        n2776) );
  CKND2D1BWP12T U3374 ( .A1(n2777), .A2(n2776), .ZN(n3102) );
  OAI22D1BWP12T U3375 ( .A1(n2781), .A2(n3679), .B1(n3775), .B2(n3773), .ZN(
        n2782) );
  AOI211D1BWP12T U3376 ( .A1(n2784), .A2(n4163), .B(n2783), .C(n2782), .ZN(
        n2785) );
  OAI211D1BWP12T U3377 ( .A1(n2787), .A2(n3613), .B(n2786), .C(n2785), .ZN(
        n2788) );
  AOI21D1BWP12T U3378 ( .A1(n4210), .A2(n4141), .B(n2788), .ZN(n2790) );
  TPAOI21D1BWP12T U3379 ( .A1(n2794), .A2(n2793), .B(n2792), .ZN(n2798) );
  ND2D1BWP12T U3380 ( .A1(n2796), .A2(n2795), .ZN(n2797) );
  XOR2XD1BWP12T U3381 ( .A1(n2798), .A2(n2797), .Z(n3420) );
  INVD1BWP12T U3382 ( .I(n2803), .ZN(n3341) );
  AOI22D1BWP12T U3383 ( .A1(n4215), .A2(n3530), .B1(n3492), .B2(n4173), .ZN(
        n2842) );
  INVD1BWP12T U3384 ( .I(n2804), .ZN(n3377) );
  AOI22D1BWP12T U3385 ( .A1(n3707), .A2(n2807), .B1(n2806), .B2(n2805), .ZN(
        n2811) );
  AOI22D0BWP12T U3386 ( .A1(n3229), .A2(n2809), .B1(n3231), .B2(n2808), .ZN(
        n2810) );
  ND2D1BWP12T U3387 ( .A1(n2811), .A2(n2810), .ZN(n3225) );
  MUX2NXD0BWP12T U3388 ( .I0(n3233), .I1(n3225), .S(n2547), .ZN(n3702) );
  INVD0BWP12T U3389 ( .I(n2812), .ZN(n2815) );
  OAI22D0BWP12T U3390 ( .A1(n2950), .A2(n2948), .B1(n2951), .B2(n3356), .ZN(
        n2814) );
  OAI21D0BWP12T U3391 ( .A1(n2947), .A2(n2949), .B(n3841), .ZN(n2813) );
  AOI211D1BWP12T U3392 ( .A1(n3353), .A2(n2815), .B(n2814), .C(n2813), .ZN(
        n2837) );
  OAI22D1BWP12T U3393 ( .A1(n3682), .A2(n3356), .B1(n3712), .B2(n2955), .ZN(
        n4158) );
  MAOI22D0BWP12T U3394 ( .A1(n4210), .A2(n4125), .B1(n3743), .B2(n4201), .ZN(
        n2841) );
  CKND2D0BWP12T U3395 ( .A1(n4158), .A2(n3986), .ZN(n2820) );
  AO21D0BWP12T U3396 ( .A1(n3765), .A2(n2820), .B(n2837), .Z(n3971) );
  CKND2D1BWP12T U3397 ( .A1(n3624), .A2(n4203), .ZN(n2833) );
  OAI21D0BWP12T U3398 ( .A1(n4063), .A2(n4182), .B(n4181), .ZN(n2831) );
  OAI22D0BWP12T U3399 ( .A1(n2822), .A2(n3782), .B1(n2821), .B2(n3780), .ZN(
        n2826) );
  OAI22D0BWP12T U3400 ( .A1(n2824), .A2(n3786), .B1(n2823), .B2(n3784), .ZN(
        n2825) );
  NR2D1BWP12T U3401 ( .A1(n2826), .A2(n2825), .ZN(n3248) );
  MUX2D1BWP12T U3402 ( .I0(n3755), .I1(n3248), .S(n4044), .Z(n3749) );
  INVD1BWP12T U3403 ( .I(n3749), .ZN(n3795) );
  NR2D1BWP12T U3404 ( .A1(n3795), .A2(n3372), .ZN(n2830) );
  MUX2ND0BWP12T U3405 ( .I0(n4184), .I1(n2664), .S(n3957), .ZN(n2827) );
  NR2D0BWP12T U3406 ( .A1(n2827), .A2(n4185), .ZN(n2828) );
  MUX2NXD0BWP12T U3407 ( .I0(n2828), .I1(n2205), .S(n3879), .ZN(n2829) );
  RCAOI211D0BWP12T U3408 ( .A1(n3957), .A2(n2831), .B(n2830), .C(n2829), .ZN(
        n2832) );
  OAI211D1BWP12T U3409 ( .A1(n3971), .A2(n2834), .B(n2833), .C(n2832), .ZN(
        n2835) );
  AOI21D1BWP12T U3410 ( .A1(n4206), .A2(n3592), .B(n2835), .ZN(n2840) );
  AOI21D0BWP12T U3411 ( .A1(n3919), .A2(n4042), .B(n3770), .ZN(n2836) );
  NR2D1BWP12T U3412 ( .A1(n2836), .A2(n3027), .ZN(n2838) );
  OAI21D1BWP12T U3413 ( .A1(n2838), .A2(n2837), .B(n3384), .ZN(n4051) );
  CKND2D1BWP12T U3414 ( .A1(n4051), .A2(n4011), .ZN(n2839) );
  ND4D1BWP12T U3415 ( .A1(n2842), .A2(n2841), .A3(n2840), .A4(n2839), .ZN(
        n2843) );
  ND2D1BWP12T U3416 ( .A1(n2845), .A2(n2844), .ZN(n2846) );
  XNR2XD4BWP12T U3417 ( .A1(n2847), .A2(n2846), .ZN(n3445) );
  ND2XD3BWP12T U3418 ( .A1(n3445), .A2(n4171), .ZN(n2888) );
  FA1D0BWP12T U3419 ( .A(n3851), .B(n4077), .CI(n2848), .CO(n2700), .S(n3559)
         );
  INVD1BWP12T U3420 ( .I(n3559), .ZN(n2886) );
  FA1D0BWP12T U3421 ( .A(n4077), .B(n3942), .CI(n2849), .CO(n2730), .S(n4138)
         );
  FA1D0BWP12T U3422 ( .A(n4077), .B(n3942), .CI(n2850), .CO(n2701), .S(n3605)
         );
  INVD1BWP12T U3423 ( .I(n3605), .ZN(n2881) );
  TPNR2D0BWP12T U3424 ( .A1(n3703), .A2(n3226), .ZN(n2852) );
  TPOAI22D0BWP12T U3425 ( .A1(n3705), .A2(n3228), .B1(n3704), .B2(n3232), .ZN(
        n2851) );
  RCAOI211D0BWP12T U3426 ( .A1(n3707), .A2(n2859), .B(n2852), .C(n2851), .ZN(
        n3168) );
  CKND0BWP12T U3427 ( .I(n3168), .ZN(n2858) );
  NR2D0BWP12T U3428 ( .A1(n3693), .A2(n3701), .ZN(n2857) );
  NR2D0BWP12T U3429 ( .A1(n3703), .A2(n3783), .ZN(n2854) );
  OAI22D0BWP12T U3430 ( .A1(n3705), .A2(n3785), .B1(n3704), .B2(n3781), .ZN(
        n2853) );
  AOI211D0BWP12T U3431 ( .A1(n3707), .A2(n2862), .B(n2854), .C(n2853), .ZN(
        n2855) );
  OAI21D0BWP12T U3432 ( .A1(n2855), .A2(n3711), .B(n3710), .ZN(n2856) );
  RCAOI211D0BWP12T U3433 ( .A1(n4175), .A2(n2858), .B(n2857), .C(n2856), .ZN(
        n3714) );
  AOI22D0BWP12T U3434 ( .A1(n3241), .A2(n2859), .B1(n3240), .B2(n3238), .ZN(
        n2861) );
  AOI22D0BWP12T U3435 ( .A1(n3245), .A2(n3243), .B1(n3239), .B2(n3242), .ZN(
        n2860) );
  CKND2D1BWP12T U3436 ( .A1(n2861), .A2(n2860), .ZN(n3164) );
  AOI22D0BWP12T U3437 ( .A1(n3241), .A2(n2862), .B1(n3706), .B2(n3238), .ZN(
        n2866) );
  AOI22D0BWP12T U3438 ( .A1(n3245), .A2(n2864), .B1(n2863), .B2(n3242), .ZN(
        n2865) );
  AOI21D0BWP12T U3439 ( .A1(n2866), .A2(n2865), .B(n3767), .ZN(n2867) );
  AOI211D0BWP12T U3440 ( .A1(n3249), .A2(n3164), .B(n2867), .C(n3655), .ZN(
        n2868) );
  OAI21D0BWP12T U3441 ( .A1(n3751), .A2(n3841), .B(n2868), .ZN(n3811) );
  NR2D0BWP12T U3442 ( .A1(n3811), .A2(n3773), .ZN(n2877) );
  CKND2D0BWP12T U3443 ( .A1(n2869), .A2(n4036), .ZN(n4012) );
  INVD1BWP12T U3444 ( .I(n3994), .ZN(n3722) );
  CKND2D0BWP12T U3445 ( .A1(n3722), .A2(n3289), .ZN(n2875) );
  OAI21D0BWP12T U3446 ( .A1(n4077), .A2(n4182), .B(n4181), .ZN(n2873) );
  MUX2ND0BWP12T U3447 ( .I0(n4184), .I1(n2664), .S(n3942), .ZN(n2870) );
  NR2D0BWP12T U3448 ( .A1(n2870), .A2(n4185), .ZN(n2871) );
  MUX2NXD0BWP12T U3449 ( .I0(n2871), .I1(n2205), .S(n3897), .ZN(n2872) );
  AOI211XD0BWP12T U3450 ( .A1(n3942), .A2(n2873), .B(n3216), .C(n2872), .ZN(
        n2874) );
  OAI211D0BWP12T U3451 ( .A1(n4012), .A2(n3029), .B(n2875), .C(n2874), .ZN(
        n2876) );
  RCAOI211D0BWP12T U3452 ( .A1(n3714), .A2(n4163), .B(n2877), .C(n2876), .ZN(
        n2880) );
  HA1D1BWP12T U3453 ( .A(n3897), .B(n2878), .CO(n2712), .S(n3645) );
  ND2D1BWP12T U3454 ( .A1(n3645), .A2(n4203), .ZN(n2879) );
  OAI211D1BWP12T U3455 ( .A1(n3582), .A2(n2881), .B(n2880), .C(n2879), .ZN(
        n2882) );
  AOI21D1BWP12T U3456 ( .A1(n4210), .A2(n4138), .B(n2882), .ZN(n2885) );
  FA1D0BWP12T U3457 ( .A(n3851), .B(n4077), .CI(n2883), .CO(n2699), .S(n3501)
         );
  CKND2D1BWP12T U3458 ( .A1(n3501), .A2(n4173), .ZN(n2884) );
  OA211D1BWP12T U3459 ( .A1(n2886), .A2(n3532), .B(n2885), .C(n2884), .Z(n2887) );
  ND2D8BWP12T U3460 ( .A1(n2888), .A2(n2887), .ZN(result[27]) );
  ND2D1BWP12T U3461 ( .A1(n2892), .A2(n2891), .ZN(n2897) );
  INVD1BWP12T U3462 ( .I(n2893), .ZN(n2895) );
  CKND2D1BWP12T U3463 ( .A1(n2895), .A2(n2894), .ZN(n2896) );
  XNR2XD1BWP12T U3464 ( .A1(n2897), .A2(n2896), .ZN(n3434) );
  INVD0BWP12T U3465 ( .I(n3509), .ZN(n2899) );
  TPND2D0BWP12T U3466 ( .A1(n3510), .A2(n2899), .ZN(n2901) );
  INVD1BWP12T U3467 ( .I(n3513), .ZN(n2898) );
  AOI21D1BWP12T U3468 ( .A1(n3516), .A2(n2899), .B(n2898), .ZN(n2900) );
  OAI21D1BWP12T U3469 ( .A1(n3519), .A2(n2901), .B(n2900), .ZN(n2904) );
  CKND2D1BWP12T U3470 ( .A1(n2902), .A2(n3511), .ZN(n2903) );
  XNR2D1BWP12T U3471 ( .A1(n2904), .A2(n2903), .ZN(n3549) );
  INVD1BWP12T U3472 ( .I(n3549), .ZN(n2924) );
  CKND2D1BWP12T U3473 ( .A1(n2905), .A2(n4117), .ZN(n2906) );
  XNR2D1BWP12T U3474 ( .A1(n3321), .A2(n2906), .ZN(n4116) );
  MUX2NXD0BWP12T U3475 ( .I0(n3074), .I1(n3753), .S(b[3]), .ZN(n2913) );
  NR2D0BWP12T U3476 ( .A1(n2913), .A2(n3765), .ZN(n3760) );
  MUX2ND0BWP12T U3477 ( .I0(n4184), .I1(n2664), .S(n3949), .ZN(n2914) );
  NR2D0BWP12T U3478 ( .A1(n2914), .A2(n4185), .ZN(n2915) );
  NR2D0BWP12T U3479 ( .A1(n4082), .A2(n4182), .ZN(n2916) );
  AOI22D0BWP12T U3480 ( .A1(n4179), .A2(n3062), .B1(n3686), .B2(n4175), .ZN(
        n3728) );
  AOI22D1BWP12T U3481 ( .A1(n3788), .A2(n2919), .B1(n2918), .B2(n3249), .ZN(
        n3735) );
  OAI21D0BWP12T U3482 ( .A1(n3735), .A2(n3655), .B(n2920), .ZN(n4024) );
  NR2D0BWP12T U3483 ( .A1(n3680), .A2(n3841), .ZN(n3988) );
  CKND2D1BWP12T U3484 ( .A1(n3474), .A2(n4173), .ZN(n2922) );
  OAI211D1BWP12T U3485 ( .A1(n3532), .A2(n2924), .B(n2923), .C(n2922), .ZN(
        n2925) );
  AO21D4BWP12T U3486 ( .A1(n3434), .A2(n4171), .B(n2925), .Z(result[15]) );
  OAI21D1BWP12T U3487 ( .A1(n3519), .A2(n2930), .B(n2929), .ZN(n2934) );
  ND2D1BWP12T U3488 ( .A1(n2932), .A2(n2931), .ZN(n2933) );
  XNR2XD1BWP12T U3489 ( .A1(n2934), .A2(n2933), .ZN(n3545) );
  AOI22D1BWP12T U3490 ( .A1(n4215), .A2(n3545), .B1(n3464), .B2(n4173), .ZN(
        n2989) );
  MUX2NXD0BWP12T U3491 ( .I0(n3295), .I1(n3301), .S(n2547), .ZN(n2957) );
  OAI22D0BWP12T U3492 ( .A1(n3712), .A2(n2948), .B1(n2947), .B2(n3356), .ZN(
        n2954) );
  OAI21D0BWP12T U3493 ( .A1(n2950), .A2(n2949), .B(n3841), .ZN(n2953) );
  NR2D0BWP12T U3494 ( .A1(n2951), .A2(n2955), .ZN(n2952) );
  NR3D1BWP12T U3495 ( .A1(n2954), .A2(n2953), .A3(n2952), .ZN(n2973) );
  INVD1BWP12T U3496 ( .I(n3966), .ZN(n2956) );
  AOI21D1BWP12T U3497 ( .A1(n2957), .A2(n3701), .B(n2956), .ZN(n3737) );
  ND2XD0BWP12T U3498 ( .A1(n2958), .A2(n2961), .ZN(n2964) );
  INVD0BWP12T U3499 ( .I(n2959), .ZN(n2960) );
  AOI21D1BWP12T U3500 ( .A1(n2962), .A2(n2961), .B(n2960), .ZN(n2963) );
  OAI21D1BWP12T U3501 ( .A1(n3388), .A2(n2964), .B(n2963), .ZN(n2969) );
  INVD0BWP12T U3502 ( .I(n2965), .ZN(n2967) );
  CKND2D1BWP12T U3503 ( .A1(n2967), .A2(n2966), .ZN(n2968) );
  XNR2XD1BWP12T U3504 ( .A1(n2969), .A2(n2968), .ZN(n3575) );
  CKND2D0BWP12T U3505 ( .A1(n2971), .A2(n2970), .ZN(n2972) );
  AOI21D0BWP12T U3506 ( .A1(n2972), .A2(n3986), .B(n3997), .ZN(n2974) );
  OAI21D0BWP12T U3507 ( .A1(n2974), .A2(n2973), .B(n3384), .ZN(n4021) );
  AOI22D0BWP12T U3508 ( .A1(n3575), .A2(n4206), .B1(n4011), .B2(n4021), .ZN(
        n2975) );
  OAI21D1BWP12T U3509 ( .A1(n3737), .A2(n4201), .B(n2975), .ZN(n2987) );
  MUX2ND0BWP12T U3510 ( .I0(n3282), .I1(n3757), .S(b[3]), .ZN(n2976) );
  CKND2D1BWP12T U3511 ( .A1(n2976), .A2(n3997), .ZN(n3805) );
  CKND2D1BWP12T U3512 ( .A1(n3633), .A2(n4203), .ZN(n2985) );
  OAI21D1BWP12T U3513 ( .A1(a[13]), .A2(n4182), .B(n4181), .ZN(n2983) );
  NR2XD0BWP12T U3514 ( .A1(n3966), .A2(n2978), .ZN(n2982) );
  MUX2ND0BWP12T U3515 ( .I0(n4184), .I1(n2664), .S(n3931), .ZN(n2979) );
  NR2D0BWP12T U3516 ( .A1(n2979), .A2(n4185), .ZN(n2980) );
  MUX2ND0BWP12T U3517 ( .I0(n2980), .I1(n2205), .S(n3875), .ZN(n2981) );
  AOI211XD0BWP12T U3518 ( .A1(n3931), .A2(n2983), .B(n2982), .C(n2981), .ZN(
        n2984) );
  OAI211D1BWP12T U3519 ( .A1(n3773), .A2(n3805), .B(n2985), .C(n2984), .ZN(
        n2986) );
  RCAOI211D0BWP12T U3520 ( .A1(n4210), .A2(n4096), .B(n2987), .C(n2986), .ZN(
        n2988) );
  ND2D1BWP12T U3521 ( .A1(n2989), .A2(n2988), .ZN(n2990) );
  AO21D4BWP12T U3522 ( .A1(n3426), .A2(n4171), .B(n2990), .Z(result[13]) );
  OAI21D1BWP12T U3523 ( .A1(n2993), .A2(n2992), .B(n2991), .ZN(n2998) );
  INVD1BWP12T U3524 ( .I(n2994), .ZN(n2996) );
  ND2D1BWP12T U3525 ( .A1(n2996), .A2(n2995), .ZN(n2997) );
  XNR2XD2BWP12T U3526 ( .A1(n2998), .A2(n2997), .ZN(n3459) );
  INVD1BWP12T U3527 ( .I(n3555), .ZN(n3041) );
  FA1D0BWP12T U3528 ( .A(n3917), .B(n4076), .CI(n3002), .CO(n2849), .S(n4137)
         );
  AOI21D1BWP12T U3529 ( .A1(n3676), .A2(n3788), .B(n3715), .ZN(n3036) );
  FA1D0BWP12T U3530 ( .A(n3917), .B(n4076), .CI(n3008), .CO(n2850), .S(n3604)
         );
  CKND2D1BWP12T U3531 ( .A1(n3604), .A2(n4206), .ZN(n3035) );
  HA1D1BWP12T U3532 ( .A(n3896), .B(n3009), .CO(n2878), .S(n3642) );
  MUX2ND0BWP12T U3533 ( .I0(n3011), .I1(n3010), .S(b[3]), .ZN(n3750) );
  INVD1BWP12T U3534 ( .I(n3750), .ZN(n3371) );
  OAI21D0BWP12T U3535 ( .A1(n4076), .A2(n4182), .B(n4181), .ZN(n3024) );
  INR2D1BWP12T U3536 ( .A1(n4044), .B1(n3018), .ZN(n3391) );
  INVD1BWP12T U3537 ( .I(n3391), .ZN(n3993) );
  INVD0BWP12T U3538 ( .I(n3019), .ZN(n4159) );
  NR2D1BWP12T U3539 ( .A1(n3993), .A2(n4159), .ZN(n3023) );
  MUX2ND0BWP12T U3540 ( .I0(n4184), .I1(n2664), .S(n3917), .ZN(n3020) );
  NR2D0BWP12T U3541 ( .A1(n3020), .A2(n4185), .ZN(n3021) );
  MUX2ND0BWP12T U3542 ( .I0(n3021), .I1(n2205), .S(n3896), .ZN(n3022) );
  RCAOI211D0BWP12T U3543 ( .A1(n3917), .A2(n3024), .B(n3023), .C(n3022), .ZN(
        n3032) );
  MUX2D0BWP12T U3544 ( .I0(n3026), .I1(n3025), .S(n3921), .Z(n3028) );
  TPAOI21D0BWP12T U3545 ( .A1(n3028), .A2(n4044), .B(n3027), .ZN(n4047) );
  INVD1BWP12T U3546 ( .I(n4047), .ZN(n3383) );
  NR2D1BWP12T U3547 ( .A1(n4046), .A2(n3029), .ZN(n4154) );
  TPOAI21D0BWP12T U3548 ( .A1(n3383), .A2(n3030), .B(n4154), .ZN(n3031) );
  OAI211D1BWP12T U3549 ( .A1(n3773), .A2(n3812), .B(n3032), .C(n3031), .ZN(
        n3033) );
  AOI21D1BWP12T U3550 ( .A1(n3642), .A2(n4203), .B(n3033), .ZN(n3034) );
  OAI211D1BWP12T U3551 ( .A1(n3036), .A2(n4201), .B(n3035), .C(n3034), .ZN(
        n3037) );
  AOI21D1BWP12T U3552 ( .A1(n4210), .A2(n4137), .B(n3037), .ZN(n3040) );
  FA1D1BWP12T U3553 ( .A(n3850), .B(n4076), .CI(n3038), .CO(n2883), .S(n3500)
         );
  CKND2D1BWP12T U3554 ( .A1(n3500), .A2(n4173), .ZN(n3039) );
  OAI211D1BWP12T U3555 ( .A1(n3041), .A2(n3532), .B(n3040), .C(n3039), .ZN(
        n3042) );
  AO21D4BWP12T U3556 ( .A1(n3459), .A2(n4171), .B(n3042), .Z(result[26]) );
  INVD1BWP12T U3557 ( .I(n3043), .ZN(n3263) );
  AOI21D1BWP12T U3558 ( .A1(n3263), .A2(n3045), .B(n3044), .ZN(n3048) );
  ND2D1BWP12T U3559 ( .A1(n321), .A2(n3046), .ZN(n3047) );
  XOR2XD2BWP12T U3560 ( .A1(n3048), .A2(n3047), .Z(n3404) );
  ND2XD0BWP12T U3561 ( .A1(n3054), .A2(n3050), .ZN(n3051) );
  XOR2XD1BWP12T U3562 ( .A1(n3052), .A2(n3051), .Z(n3547) );
  INVD1BWP12T U3563 ( .I(n3547), .ZN(n3087) );
  CKND2D1BWP12T U3564 ( .A1(n3498), .A2(n4173), .ZN(n3086) );
  INVD1BWP12T U3565 ( .I(n3571), .ZN(n3083) );
  OAI22D1BWP12T U3566 ( .A1(n3062), .A2(n2547), .B1(n3061), .B2(n3711), .ZN(
        n3063) );
  RCAOI211D0BWP12T U3567 ( .A1(n3170), .A2(n3064), .B(n3063), .C(n3298), .ZN(
        n3695) );
  OAI21D1BWP12T U3568 ( .A1(n3066), .A2(n4013), .B(n3065), .ZN(n4048) );
  AOI22D1BWP12T U3569 ( .A1(n3695), .A2(n4163), .B1(n4011), .B2(n4048), .ZN(
        n3082) );
  OAI21D0BWP12T U3570 ( .A1(a[23]), .A2(n4182), .B(n4181), .ZN(n3071) );
  MUX2ND0BWP12T U3571 ( .I0(n4184), .I1(n2664), .S(n3943), .ZN(n3068) );
  NR2D0BWP12T U3572 ( .A1(n3068), .A2(n4185), .ZN(n3069) );
  MUX2ND0BWP12T U3573 ( .I0(n3069), .I1(n2205), .S(n3863), .ZN(n3070) );
  RCAOI21D0BWP12T U3574 ( .A1(n3943), .A2(n3071), .B(n3070), .ZN(n3078) );
  INVD1BWP12T U3575 ( .I(n3072), .ZN(n3073) );
  OAI22D0BWP12T U3576 ( .A1(n3074), .A2(n4044), .B1(n3073), .B2(n3767), .ZN(
        n3075) );
  AOI211XD0BWP12T U3577 ( .A1(n3919), .A2(n3076), .B(n3075), .C(n3770), .ZN(
        n3807) );
  CKND2D1BWP12T U3578 ( .A1(n3807), .A2(n4195), .ZN(n3077) );
  OAI211D1BWP12T U3579 ( .A1(n3079), .A2(n3684), .B(n3078), .C(n3077), .ZN(
        n3080) );
  AOI21D1BWP12T U3580 ( .A1(n3623), .A2(n4203), .B(n3080), .ZN(n3081) );
  OAI211D1BWP12T U3581 ( .A1(n3582), .A2(n3083), .B(n3082), .C(n3081), .ZN(
        n3084) );
  AOI21D1BWP12T U3582 ( .A1(n4134), .A2(n4210), .B(n3084), .ZN(n3085) );
  OAI211D1BWP12T U3583 ( .A1(n3087), .A2(n3532), .B(n3086), .C(n3085), .ZN(
        n3088) );
  AO21D4BWP12T U3584 ( .A1(n3404), .A2(n4171), .B(n3088), .Z(result[23]) );
  INVD1BWP12T U3585 ( .I(n3089), .ZN(n3262) );
  INVD1BWP12T U3586 ( .I(n3261), .ZN(n3090) );
  TPAOI21D1BWP12T U3587 ( .A1(n3263), .A2(n3262), .B(n3090), .ZN(n3095) );
  CKND0BWP12T U3588 ( .I(n3091), .ZN(n3093) );
  ND2D1BWP12T U3589 ( .A1(n3093), .A2(n3092), .ZN(n3094) );
  XOR2XD1BWP12T U3590 ( .A1(n3095), .A2(n3094), .Z(n3405) );
  CKND2D1BWP12T U3591 ( .A1(n3548), .A2(n4215), .ZN(n3131) );
  AOI222D1BWP12T U3592 ( .A1(n3101), .A2(n4179), .B1(n3100), .B2(n4177), .C1(
        n3099), .C2(n4175), .ZN(n3668) );
  INVD1BWP12T U3593 ( .I(n3668), .ZN(n3117) );
  CKND0BWP12T U3594 ( .I(n3754), .ZN(n3103) );
  AOI22D0BWP12T U3595 ( .A1(n3919), .A2(n3103), .B1(n3102), .B2(n3788), .ZN(
        n3104) );
  OAI211D1BWP12T U3596 ( .A1(n3105), .A2(n4044), .B(n3104), .C(n3285), .ZN(
        n3777) );
  INVD1BWP12T U3597 ( .I(n3106), .ZN(n3291) );
  MOAI22D0BWP12T U3598 ( .A1(n3777), .A2(n3773), .B1(n3612), .B2(n4203), .ZN(
        n3116) );
  INVD1BWP12T U3599 ( .I(n4038), .ZN(n3114) );
  TPND2D0BWP12T U3600 ( .A1(n3289), .A2(n3683), .ZN(n3113) );
  OAI21D0BWP12T U3601 ( .A1(n4070), .A2(n4182), .B(n4181), .ZN(n3111) );
  MUX2ND0BWP12T U3602 ( .I0(n4184), .I1(n2664), .S(n3941), .ZN(n3108) );
  NR2D0BWP12T U3603 ( .A1(n3108), .A2(n4185), .ZN(n3109) );
  MUX2ND0BWP12T U3604 ( .I0(n3109), .I1(n2205), .S(n3862), .ZN(n3110) );
  AOI211XD0BWP12T U3605 ( .A1(n3941), .A2(n3111), .B(n3216), .C(n3110), .ZN(
        n3112) );
  OAI211D1BWP12T U3606 ( .A1(n3114), .A2(n3290), .B(n3113), .C(n3112), .ZN(
        n3115) );
  RCAOI211D0BWP12T U3607 ( .A1(n4163), .A2(n3117), .B(n3116), .C(n3115), .ZN(
        n3130) );
  ND2XD0BWP12T U3608 ( .A1(n3124), .A2(n3123), .ZN(n3119) );
  XOR2XD1BWP12T U3609 ( .A1(n3120), .A2(n3119), .Z(n4114) );
  AOI22D1BWP12T U3610 ( .A1(n4114), .A2(n4210), .B1(n4206), .B2(n3570), .ZN(
        n3129) );
  CKND2D1BWP12T U3611 ( .A1(n3473), .A2(n4173), .ZN(n3128) );
  ND4D1BWP12T U3612 ( .A1(n3131), .A2(n3130), .A3(n3129), .A4(n3128), .ZN(
        n3132) );
  AO21D4BWP12T U3613 ( .A1(n3405), .A2(n4171), .B(n3132), .Z(result[22]) );
  IND2XD1BWP12T U3614 ( .A1(n3136), .B1(n3135), .ZN(n3137) );
  INVD1BWP12T U3615 ( .I(n3137), .ZN(n3138) );
  XNR2XD1BWP12T U3616 ( .A1(n3139), .A2(n3138), .ZN(n3436) );
  AOI21D1BWP12T U3617 ( .A1(n3321), .A2(n3151), .B(n3150), .ZN(n3156) );
  INVD0BWP12T U3618 ( .I(n3152), .ZN(n3154) );
  CKND2D1BWP12T U3619 ( .A1(n3154), .A2(n3153), .ZN(n3155) );
  XOR2XD1BWP12T U3620 ( .A1(n3156), .A2(n3155), .Z(n4100) );
  ND3D0BWP12T U3621 ( .A1(n3986), .A2(n4044), .A3(n3756), .ZN(n3163) );
  AO222D1BWP12T U3622 ( .A1(n3165), .A2(n3249), .B1(n3164), .B2(n3788), .C1(
        n3163), .C2(n3765), .Z(n3798) );
  MUX2ND0BWP12T U3623 ( .I0(n4184), .I1(n2664), .S(b[19]), .ZN(n3166) );
  OAI22D0BWP12T U3624 ( .A1(n3168), .A2(n3711), .B1(n3167), .B2(n2547), .ZN(
        n3169) );
  AOI211XD0BWP12T U3625 ( .A1(n3170), .A2(n3687), .B(n3169), .C(n3298), .ZN(
        n3696) );
  INVD1BWP12T U3626 ( .I(n3171), .ZN(n4033) );
  AOI21D1BWP12T U3627 ( .A1(n4173), .A2(n3468), .B(n3174), .ZN(n3175) );
  IOA21D1BWP12T U3628 ( .A1(n3525), .A2(n4215), .B(n3175), .ZN(n3176) );
  AO21D4BWP12T U3629 ( .A1(n3436), .A2(n4171), .B(n3176), .Z(result[19]) );
  INVD0BWP12T U3630 ( .I(n3430), .ZN(n3178) );
  AOI21D1BWP12T U3631 ( .A1(n3178), .A2(n3428), .B(n3177), .ZN(n3184) );
  CKND2D1BWP12T U3632 ( .A1(n3180), .A2(n3179), .ZN(n3181) );
  ND2D1BWP12T U3633 ( .A1(n3182), .A2(n3181), .ZN(n3183) );
  XOR2XD1BWP12T U3634 ( .A1(n3184), .A2(n3183), .Z(n3433) );
  INVD1BWP12T U3635 ( .I(n3433), .ZN(n3260) );
  ND2XD0BWP12T U3636 ( .A1(n3510), .A2(n3186), .ZN(n3188) );
  AOI21D1BWP12T U3637 ( .A1(n3516), .A2(n3186), .B(n3185), .ZN(n3187) );
  OAI21D1BWP12T U3638 ( .A1(n3519), .A2(n3188), .B(n3187), .ZN(n3192) );
  ND2D1BWP12T U3639 ( .A1(n3190), .A2(n3189), .ZN(n3191) );
  XNR2D1BWP12T U3640 ( .A1(n3192), .A2(n3191), .ZN(n3524) );
  INVD0BWP12T U3641 ( .I(n3193), .ZN(n3196) );
  INVD1BWP12T U3642 ( .I(n3194), .ZN(n3195) );
  AOI21D1BWP12T U3643 ( .A1(n3276), .A2(n3196), .B(n3195), .ZN(n3200) );
  CKND2D1BWP12T U3644 ( .A1(n3190), .A2(n3198), .ZN(n3199) );
  XOR2XD1BWP12T U3645 ( .A1(n3200), .A2(n3199), .Z(n3470) );
  TPOAI21D0BWP12T U3646 ( .A1(n3579), .A2(n3201), .B(n4120), .ZN(n3205) );
  CKND2D1BWP12T U3647 ( .A1(n3203), .A2(n3202), .ZN(n3204) );
  XNR2XD1BWP12T U3648 ( .A1(n3205), .A2(n3204), .ZN(n3569) );
  INVD0BWP12T U3649 ( .I(n3206), .ZN(n3209) );
  INVD1BWP12T U3650 ( .I(n3207), .ZN(n3208) );
  AOI21D1BWP12T U3651 ( .A1(n3321), .A2(n3209), .B(n3208), .ZN(n3213) );
  CKND2D1BWP12T U3652 ( .A1(n3203), .A2(n3211), .ZN(n3212) );
  XOR2XD1BWP12T U3653 ( .A1(n3213), .A2(n3212), .Z(n4102) );
  CKND2D1BWP12T U3654 ( .A1(n4102), .A2(n4210), .ZN(n3214) );
  IOA21D1BWP12T U3655 ( .A1(n3569), .A2(n4206), .B(n3214), .ZN(n3256) );
  INVD1BWP12T U3656 ( .I(n3215), .ZN(n4035) );
  INVD0BWP12T U3657 ( .I(n3990), .ZN(n3223) );
  INVD1BWP12T U3658 ( .I(n3216), .ZN(n4193) );
  OAI21D0BWP12T U3659 ( .A1(a[17]), .A2(n4182), .B(n4181), .ZN(n3220) );
  MUX2ND0BWP12T U3660 ( .I0(n4184), .I1(n2664), .S(n3952), .ZN(n3217) );
  NR2XD0BWP12T U3661 ( .A1(n3217), .A2(n4185), .ZN(n3218) );
  MUX2NXD0BWP12T U3662 ( .I0(n3218), .I1(n2205), .S(n3868), .ZN(n3219) );
  RCAOI21D0BWP12T U3663 ( .A1(n3952), .A2(n3220), .B(n3219), .ZN(n3221) );
  CKND2D1BWP12T U3664 ( .A1(n4193), .A2(n3221), .ZN(n3222) );
  TPAOI21D0BWP12T U3665 ( .A1(n3223), .A2(n3289), .B(n3222), .ZN(n3224) );
  OAI21D1BWP12T U3666 ( .A1(n4035), .A2(n3290), .B(n3224), .ZN(n3255) );
  INVD0BWP12T U3667 ( .I(n3225), .ZN(n3237) );
  AOI22D0BWP12T U3668 ( .A1(n3229), .A2(n3228), .B1(n3227), .B2(n3226), .ZN(
        n3709) );
  AOI22D0BWP12T U3669 ( .A1(n3707), .A2(n3232), .B1(n3231), .B2(n3230), .ZN(
        n3708) );
  AOI21D1BWP12T U3670 ( .A1(n3709), .A2(n3708), .B(n3711), .ZN(n3236) );
  TPNR2D0BWP12T U3671 ( .A1(n3234), .A2(n3233), .ZN(n3235) );
  RCAOI211D0BWP12T U3672 ( .A1(n3237), .A2(n4175), .B(n3236), .C(n3235), .ZN(
        n3664) );
  AOI22D0BWP12T U3673 ( .A1(n3241), .A2(n3240), .B1(n3239), .B2(n3238), .ZN(
        n3247) );
  AOI22D0BWP12T U3674 ( .A1(n3245), .A2(n3244), .B1(n3243), .B2(n3242), .ZN(
        n3246) );
  ND2D1BWP12T U3675 ( .A1(n3247), .A2(n3246), .ZN(n3779) );
  INVD1BWP12T U3676 ( .I(n3248), .ZN(n3250) );
  AOI22D1BWP12T U3677 ( .A1(n3788), .A2(n3779), .B1(n3250), .B2(n3249), .ZN(
        n3251) );
  OAI211D1BWP12T U3678 ( .A1(n3755), .A2(n3841), .B(n3251), .C(n3285), .ZN(
        n3797) );
  NR2D1BWP12T U3679 ( .A1(n3797), .A2(n3773), .ZN(n3252) );
  AOI21D1BWP12T U3680 ( .A1(n3611), .A2(n4203), .B(n3252), .ZN(n3253) );
  OAI21D1BWP12T U3681 ( .A1(n3664), .A2(n4201), .B(n3253), .ZN(n3254) );
  NR3D1BWP12T U3682 ( .A1(n3256), .A2(n3255), .A3(n3254), .ZN(n3257) );
  IOA21D1BWP12T U3683 ( .A1(n3470), .A2(n4173), .B(n3257), .ZN(n3258) );
  AOI21D1BWP12T U3684 ( .A1(n3524), .A2(n4215), .B(n3258), .ZN(n3259) );
  RCOAI21D1BWP12T U3685 ( .A1(n3260), .A2(n3407), .B(n3259), .ZN(result[17])
         );
  ND2XD0BWP12T U3686 ( .A1(n3278), .A2(n3265), .ZN(n3266) );
  XOR2XD1BWP12T U3687 ( .A1(n3267), .A2(n3266), .Z(n3543) );
  INVD1BWP12T U3688 ( .I(n3268), .ZN(n3272) );
  NR2D1BWP12T U3689 ( .A1(n3269), .A2(n3272), .ZN(n3275) );
  INVD1BWP12T U3690 ( .I(n3270), .ZN(n3271) );
  OAI21D1BWP12T U3691 ( .A1(n3273), .A2(n3272), .B(n3271), .ZN(n3274) );
  AOI21D1BWP12T U3692 ( .A1(n3276), .A2(n3275), .B(n3274), .ZN(n3280) );
  CKND2D1BWP12T U3693 ( .A1(n3278), .A2(n3277), .ZN(n3279) );
  XOR2XD1BWP12T U3694 ( .A1(n3280), .A2(n3279), .Z(n3472) );
  CKND2D1BWP12T U3695 ( .A1(n3472), .A2(n4173), .ZN(n3281) );
  IOA21D1BWP12T U3696 ( .A1(n3543), .A2(n4215), .B(n3281), .ZN(n3328) );
  INVD1BWP12T U3697 ( .I(n3282), .ZN(n3287) );
  INVD0BWP12T U3698 ( .I(n3283), .ZN(n3284) );
  AOI22D0BWP12T U3699 ( .A1(n3284), .A2(n3788), .B1(n3919), .B2(n3757), .ZN(
        n3286) );
  OAI211D1BWP12T U3700 ( .A1(n3287), .A2(n4044), .B(n3286), .C(n3285), .ZN(
        n3796) );
  INVD1BWP12T U3701 ( .I(n3288), .ZN(n4034) );
  NR2XD0BWP12T U3702 ( .A1(n3291), .A2(n4069), .ZN(n3292) );
  TPND2D0BWP12T U3703 ( .A1(n3293), .A2(n3292), .ZN(n3294) );
  XOR2D1BWP12T U3704 ( .A1(n3294), .A2(a[21]), .Z(n3617) );
  INVD1BWP12T U3705 ( .I(n3295), .ZN(n3685) );
  INVD1BWP12T U3706 ( .I(n3296), .ZN(n3297) );
  OAI22D1BWP12T U3707 ( .A1(n3685), .A2(n3701), .B1(n3297), .B2(n3711), .ZN(
        n3299) );
  AOI211D1BWP12T U3708 ( .A1(n3301), .A2(n3300), .B(n3299), .C(n3298), .ZN(
        n3671) );
  TPND2D0BWP12T U3709 ( .A1(n3302), .A2(n3305), .ZN(n3308) );
  INVD0BWP12T U3710 ( .I(n3303), .ZN(n3304) );
  TPAOI21D0BWP12T U3711 ( .A1(n3306), .A2(n3305), .B(n3304), .ZN(n3307) );
  OAI21D1BWP12T U3712 ( .A1(n3579), .A2(n3308), .B(n3307), .ZN(n3312) );
  CKND2D1BWP12T U3713 ( .A1(n3323), .A2(n3310), .ZN(n3311) );
  XNR2XD1BWP12T U3714 ( .A1(n3312), .A2(n3311), .ZN(n3573) );
  INVD1BWP12T U3715 ( .I(n3313), .ZN(n3317) );
  NR2D1BWP12T U3716 ( .A1(n3314), .A2(n3317), .ZN(n3320) );
  INVD1BWP12T U3717 ( .I(n3315), .ZN(n3316) );
  OAI21D1BWP12T U3718 ( .A1(n3318), .A2(n3317), .B(n3316), .ZN(n3319) );
  AOI21D1BWP12T U3719 ( .A1(n3321), .A2(n3320), .B(n3319), .ZN(n3325) );
  ND2D1BWP12T U3720 ( .A1(n3323), .A2(n3322), .ZN(n3324) );
  XOR2XD1BWP12T U3721 ( .A1(n3325), .A2(n3324), .Z(n4113) );
  NR3D1BWP12T U3722 ( .A1(n3328), .A2(n3327), .A3(n3326), .ZN(n3329) );
  INVD0BWP12T U3723 ( .I(n3335), .ZN(n3337) );
  CKND2D0BWP12T U3724 ( .A1(n3338), .A2(n3341), .ZN(n3344) );
  INVD0BWP12T U3725 ( .I(n3339), .ZN(n3340) );
  TPAOI21D0BWP12T U3726 ( .A1(n3342), .A2(n3341), .B(n3340), .ZN(n3343) );
  OAI21D1BWP12T U3727 ( .A1(n3345), .A2(n3344), .B(n3343), .ZN(n3349) );
  TPND2D0BWP12T U3728 ( .A1(n3337), .A2(n3347), .ZN(n3348) );
  XNR2XD1BWP12T U3729 ( .A1(n3349), .A2(n3348), .ZN(n3467) );
  INVD1BWP12T U3730 ( .I(n3467), .ZN(n3382) );
  INVD1BWP12T U3731 ( .I(n3352), .ZN(n3359) );
  AOI21D0BWP12T U3732 ( .A1(n3354), .A2(n3353), .B(n3919), .ZN(n3355) );
  OAI21D0BWP12T U3733 ( .A1(n3357), .A2(n3356), .B(n3355), .ZN(n3358) );
  AOI21D1BWP12T U3734 ( .A1(b[3]), .A2(n3359), .B(n3358), .ZN(n3730) );
  AOI21D0BWP12T U3735 ( .A1(n3391), .A2(n4163), .B(n3360), .ZN(n3362) );
  MOAI22D0BWP12T U3736 ( .A1(n3730), .A2(n3362), .B1(n3694), .B2(n3361), .ZN(
        n3374) );
  MUX2ND0BWP12T U3737 ( .I0(n3364), .I1(n3363), .S(n3932), .ZN(n3365) );
  CKND2D0BWP12T U3738 ( .A1(n3365), .A2(n4181), .ZN(n3367) );
  MUX2NXD0BWP12T U3739 ( .I0(n3367), .I1(n3366), .S(n3877), .ZN(n3370) );
  OAI21D0BWP12T U3740 ( .A1(n4061), .A2(n4182), .B(n4181), .ZN(n3368) );
  TPND2D0BWP12T U3741 ( .A1(n3932), .A2(n3368), .ZN(n3369) );
  OAI211D1BWP12T U3742 ( .A1(n3372), .A2(n3371), .B(n3370), .C(n3369), .ZN(
        n3373) );
  AOI211D1BWP12T U3743 ( .A1(n4203), .A2(n3622), .B(n3374), .C(n3373), .ZN(
        n3381) );
  CKND2D1BWP12T U3744 ( .A1(n4124), .A2(n4210), .ZN(n3380) );
  AOI21D0BWP12T U3745 ( .A1(n3383), .A2(n3986), .B(n3997), .ZN(n3385) );
  OAI21D0BWP12T U3746 ( .A1(n3385), .A2(n3730), .B(n3384), .ZN(n4058) );
  CKND2D0BWP12T U3747 ( .A1(n3391), .A2(n3986), .ZN(n3392) );
  AOI21D1BWP12T U3748 ( .A1(n3392), .A2(n3765), .B(n3730), .ZN(n3982) );
  INVD1BWP12T U3749 ( .I(n3393), .ZN(n3402) );
  FA1D1BWP12T U3750 ( .A(n4089), .B(b[31]), .CI(n3397), .CO(n3398), .S(n4142)
         );
  OAI211D1BWP12T U3751 ( .A1(n3407), .A2(n3402), .B(n3401), .C(n3400), .ZN(
        c_out) );
  CKND2BWP12T U3752 ( .I(n3403), .ZN(n3449) );
  NR2D0BWP12T U3753 ( .A1(n3405), .A2(n3404), .ZN(n3442) );
  OR3D0BWP12T U3754 ( .A1(n3408), .A2(n3407), .A3(n3406), .Z(n3410) );
  OR3D0BWP12T U3755 ( .A1(n3411), .A2(n3410), .A3(n3409), .Z(n3413) );
  OR3D0BWP12T U3756 ( .A1(n3414), .A2(n3413), .A3(n3412), .Z(n3416) );
  OR3D0BWP12T U3757 ( .A1(n3417), .A2(n3416), .A3(n3415), .Z(n3419) );
  OR3D2BWP12T U3758 ( .A1(n3420), .A2(n3419), .A3(n3418), .Z(n3422) );
  OR3XD4BWP12T U3759 ( .A1(n3423), .A2(n3422), .A3(n3421), .Z(n3424) );
  TPNR3D2BWP12T U3760 ( .A1(n3426), .A2(n3425), .A3(n3424), .ZN(n3432) );
  ND2D1BWP12T U3761 ( .A1(n3428), .A2(n3427), .ZN(n3429) );
  XOR2D1BWP12T U3762 ( .A1(n3430), .A2(n3429), .Z(n4172) );
  INR3XD0BWP12T U3763 ( .A1(n3432), .B1(n3431), .B2(n4172), .ZN(n3440) );
  NR3D0BWP12T U3764 ( .A1(n3435), .A2(n3434), .A3(n3433), .ZN(n3439) );
  NR2D0BWP12T U3765 ( .A1(n3437), .A2(n3436), .ZN(n3438) );
  AN3D2BWP12T U3766 ( .A1(n3440), .A2(n3439), .A3(n3438), .Z(n3441) );
  CKND2D1BWP12T U3767 ( .A1(n3442), .A2(n3441), .ZN(n3447) );
  OR2XD1BWP12T U3768 ( .A1(n3444), .A2(n3443), .Z(n3446) );
  TPNR3D2BWP12T U3769 ( .A1(n3447), .A2(n3446), .A3(n3445), .ZN(n3448) );
  IND3D1BWP12T U3770 ( .A1(n3450), .B1(n3449), .B2(n3448), .ZN(n4151) );
  CKND1BWP12T U3771 ( .I(n3451), .ZN(n3463) );
  INVD1BWP12T U3772 ( .I(n3452), .ZN(n3453) );
  TPAOI21D1BWP12T U3773 ( .A1(n3454), .A2(n319), .B(n3453), .ZN(n3458) );
  AN2XD2BWP12T U3774 ( .A1(n3456), .A2(n3455), .Z(n3457) );
  XNR2XD1BWP12T U3775 ( .A1(n3458), .A2(n3457), .ZN(n4170) );
  OR2XD1BWP12T U3776 ( .A1(n4170), .A2(n3459), .Z(n3461) );
  TPNR2D0BWP12T U3777 ( .A1(n3461), .A2(n3460), .ZN(n3462) );
  CKND2D1BWP12T U3778 ( .A1(n3463), .A2(n3462), .ZN(n4150) );
  TPOAI21D0BWP12T U3779 ( .A1(n3487), .A2(n3486), .B(n3485), .ZN(n3491) );
  CKND2D1BWP12T U3780 ( .A1(n3489), .A2(n3488), .ZN(n3490) );
  XNR2XD1BWP12T U3781 ( .A1(n3491), .A2(n3490), .ZN(n4174) );
  NR4D0BWP12T U3782 ( .A1(n3505), .A2(n3504), .A3(n3503), .A4(n3502), .ZN(
        n4148) );
  NR2D0BWP12T U3783 ( .A1(n3509), .A2(n3512), .ZN(n3515) );
  TPND2D0BWP12T U3784 ( .A1(n3510), .A2(n3515), .ZN(n3518) );
  OAI21D0BWP12T U3785 ( .A1(n3513), .A2(n3512), .B(n3511), .ZN(n3514) );
  AOI21D1BWP12T U3786 ( .A1(n3516), .A2(n3515), .B(n3514), .ZN(n3517) );
  OAI21D1BWP12T U3787 ( .A1(n3519), .A2(n3518), .B(n3517), .ZN(n3523) );
  CKND2D1BWP12T U3788 ( .A1(n3521), .A2(n3520), .ZN(n3522) );
  XNR2D1BWP12T U3789 ( .A1(n3523), .A2(n3522), .ZN(n4216) );
  NR4D0BWP12T U3790 ( .A1(n3526), .A2(n3525), .A3(n4216), .A4(n3524), .ZN(
        n3553) );
  OR4D1BWP12T U3791 ( .A1(n3530), .A2(n3529), .A3(n3528), .A4(n3527), .Z(n3546) );
  OR4D1BWP12T U3792 ( .A1(n3534), .A2(n3533), .A3(n3532), .A4(n3531), .Z(n3535) );
  OR4D1BWP12T U3793 ( .A1(n3538), .A2(n3537), .A3(n3536), .A4(n3535), .Z(n3539) );
  OR4D1BWP12T U3794 ( .A1(n3542), .A2(n3541), .A3(n3540), .A4(n3539), .Z(n3544) );
  NR4D0BWP12T U3795 ( .A1(n3546), .A2(n3545), .A3(n3544), .A4(n3543), .ZN(
        n3552) );
  NR4D0BWP12T U3796 ( .A1(n3550), .A2(n3549), .A3(n3548), .A4(n3547), .ZN(
        n3551) );
  IND4D1BWP12T U3797 ( .A1(n3554), .B1(n3553), .B2(n3552), .B3(n3551), .ZN(
        n3556) );
  OR4D1BWP12T U3798 ( .A1(n3557), .A2(n4166), .A3(n3556), .A4(n3555), .Z(n3558) );
  NR4D0BWP12T U3799 ( .A1(n3561), .A2(n3560), .A3(n3559), .A4(n3558), .ZN(
        n3564) );
  INR3XD0BWP12T U3800 ( .A1(n3564), .B1(n3563), .B2(n3562), .ZN(n4147) );
  FA1D0BWP12T U3801 ( .A(n4157), .B(b[25]), .CI(n3565), .CO(n3008), .S(n4153)
         );
  NR4D0BWP12T U3802 ( .A1(n3569), .A2(n3568), .A3(n3567), .A4(n3566), .ZN(
        n3601) );
  NR4D0BWP12T U3803 ( .A1(n3573), .A2(n3572), .A3(n3571), .A4(n3570), .ZN(
        n3600) );
  NR4D0BWP12T U3804 ( .A1(n3577), .A2(n3576), .A3(n3575), .A4(n3574), .ZN(
        n3596) );
  CKND2D0BWP12T U3805 ( .A1(n4121), .A2(n4120), .ZN(n3578) );
  XOR2XD1BWP12T U3806 ( .A1(n3579), .A2(n3578), .Z(n4207) );
  NR3D0BWP12T U3807 ( .A1(n4207), .A2(n3581), .A3(n3580), .ZN(n3595) );
  NR4D0BWP12T U3808 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(
        n3586) );
  CKND2D0BWP12T U3809 ( .A1(n322), .A2(n3586), .ZN(n3590) );
  NR4D0BWP12T U3810 ( .A1(n3590), .A2(n3589), .A3(n3588), .A4(n3587), .ZN(
        n3594) );
  NR2D0BWP12T U3811 ( .A1(n3592), .A2(n3591), .ZN(n3593) );
  ND4D1BWP12T U3812 ( .A1(n3596), .A2(n3595), .A3(n3594), .A4(n3593), .ZN(
        n3598) );
  NR2D0BWP12T U3813 ( .A1(n3598), .A2(n3597), .ZN(n3599) );
  IND4D1BWP12T U3814 ( .A1(n4153), .B1(n3601), .B2(n3600), .B3(n3599), .ZN(
        n3603) );
  OR4D1BWP12T U3815 ( .A1(n3605), .A2(n3604), .A3(n3603), .A4(n3602), .Z(n3606) );
  NR4D0BWP12T U3816 ( .A1(n3609), .A2(n3608), .A3(n3607), .A4(n3606), .ZN(
        n4145) );
  XOR2D1BWP12T U3817 ( .A1(n3619), .A2(n4183), .Z(n4204) );
  OR4D1BWP12T U3818 ( .A1(n3621), .A2(n3620), .A3(n4156), .A4(n4204), .Z(n3625) );
  NR4D0BWP12T U3819 ( .A1(n3625), .A2(n3624), .A3(n3623), .A4(n3622), .ZN(
        n3638) );
  NR2D0BWP12T U3820 ( .A1(n3627), .A2(n3626), .ZN(n3637) );
  NR3D0BWP12T U3821 ( .A1(n3630), .A2(n3629), .A3(n3628), .ZN(n3636) );
  NR4D0BWP12T U3822 ( .A1(n3634), .A2(n3633), .A3(n3632), .A4(n3631), .ZN(
        n3635) );
  ND4D1BWP12T U3823 ( .A1(n3638), .A2(n3637), .A3(n3636), .A4(n3635), .ZN(
        n3639) );
  OR4D1BWP12T U3824 ( .A1(n3642), .A2(n3641), .A3(n3640), .A4(n3639), .Z(n3643) );
  OR4D1BWP12T U3825 ( .A1(n3646), .A2(n3645), .A3(n3644), .A4(n3643), .Z(n3661) );
  NR4D0BWP12T U3826 ( .A1(n4089), .A2(n4076), .A3(n4077), .A4(n4064), .ZN(
        n3650) );
  NR4D0BWP12T U3827 ( .A1(a[29]), .A2(n4065), .A3(n4157), .A4(n4061), .ZN(
        n3649) );
  NR4D0BWP12T U3828 ( .A1(a[14]), .A2(n4063), .A3(n4062), .A4(n4060), .ZN(
        n3648) );
  NR4D0BWP12T U3829 ( .A1(a[18]), .A2(n4082), .A3(a[13]), .A4(n4078), .ZN(
        n3647) );
  ND4D1BWP12T U3830 ( .A1(n3650), .A2(n3649), .A3(n3648), .A4(n3647), .ZN(
        n3657) );
  NR4D0BWP12T U3831 ( .A1(a[21]), .A2(n4069), .A3(a[19]), .A4(n4070), .ZN(
        n3654) );
  NR4D0BWP12T U3832 ( .A1(a[17]), .A2(n4183), .A3(n4083), .A4(n4084), .ZN(
        n3653) );
  NR4D0BWP12T U3833 ( .A1(n4075), .A2(n4081), .A3(n4068), .A4(n581), .ZN(n3651) );
  INR3XD0BWP12T U3834 ( .A1(n3651), .B1(n4181), .B2(n4067), .ZN(n3652) );
  ND4D0BWP12T U3835 ( .A1(n3654), .A2(n3653), .A3(n3652), .A4(n3863), .ZN(
        n3656) );
  OR4D0BWP12T U3836 ( .A1(n3658), .A2(n3657), .A3(n3656), .A4(n3655), .Z(n3659) );
  TPOAI31D0BWP12T U3837 ( .A1(n3662), .A2(n3661), .A3(n3660), .B(n3659), .ZN(
        n3663) );
  CKND2D0BWP12T U3838 ( .A1(n3663), .A2(n2018), .ZN(n4094) );
  CKND2D0BWP12T U3839 ( .A1(n3665), .A2(n3664), .ZN(n3673) );
  ND4D0BWP12T U3840 ( .A1(n3669), .A2(n3668), .A3(n3667), .A4(n3666), .ZN(
        n3672) );
  NR4D0BWP12T U3841 ( .A1(n3673), .A2(n3672), .A3(n3671), .A4(n3670), .ZN(
        n3700) );
  CKND0BWP12T U3842 ( .I(n3674), .ZN(n3675) );
  NR4D0BWP12T U3843 ( .A1(n3678), .A2(n3677), .A3(n3676), .A4(n3675), .ZN(
        n3699) );
  CKND0BWP12T U3844 ( .I(n3981), .ZN(n3691) );
  NR2D0BWP12T U3845 ( .A1(n3686), .A2(n3685), .ZN(n3689) );
  ND4D0BWP12T U3846 ( .A1(n3689), .A2(n3688), .A3(n4163), .A4(n3687), .ZN(
        n3690) );
  AOI211D0BWP12T U3847 ( .A1(n3692), .A2(n3691), .B(n3999), .C(n3690), .ZN(
        n3698) );
  NR4D0BWP12T U3848 ( .A1(n3696), .A2(n3695), .A3(n3694), .A4(n3693), .ZN(
        n3697) );
  ND4D1BWP12T U3849 ( .A1(n3700), .A2(n3699), .A3(n3698), .A4(n3697), .ZN(
        n3716) );
  NR4D0BWP12T U3850 ( .A1(n3716), .A2(n3715), .A3(n3714), .A4(n4162), .ZN(
        n4010) );
  INVD1BWP12T U3851 ( .I(n3717), .ZN(n4199) );
  ND4D0BWP12T U3852 ( .A1(n3720), .A2(n4199), .A3(n3719), .A4(n3718), .ZN(
        n3721) );
  INR3XD0BWP12T U3853 ( .A1(n3990), .B1(n3722), .B2(n3721), .ZN(n3727) );
  NR2D0BWP12T U3854 ( .A1(n3724), .A2(n3723), .ZN(n3995) );
  CKND0BWP12T U3855 ( .I(n3725), .ZN(n3991) );
  ND4D0BWP12T U3856 ( .A1(n3727), .A2(n3995), .A3(n3726), .A4(n3991), .ZN(
        n3747) );
  OAI211D0BWP12T U3857 ( .A1(n3919), .A2(n3730), .B(n3729), .C(n3728), .ZN(
        n3733) );
  NR3D0BWP12T U3858 ( .A1(n3733), .A2(n3732), .A3(n3731), .ZN(n3740) );
  ND3D0BWP12T U3859 ( .A1(n3736), .A2(n3735), .A3(n3734), .ZN(n3987) );
  INVD0BWP12T U3860 ( .I(n3987), .ZN(n3738) );
  ND4D0BWP12T U3861 ( .A1(n3740), .A2(n3739), .A3(n3738), .A4(n3737), .ZN(
        n3746) );
  ND4D0BWP12T U3862 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(
        n3745) );
  AOI211D0BWP12T U3863 ( .A1(n3841), .A2(n3747), .B(n3746), .C(n3745), .ZN(
        n4009) );
  NR4D0BWP12T U3864 ( .A1(n3751), .A2(n3750), .A3(n3749), .A4(n3748), .ZN(
        n3766) );
  NR3D0BWP12T U3865 ( .A1(n3754), .A2(n3753), .A3(n3752), .ZN(n3759) );
  NR2D0BWP12T U3866 ( .A1(n3756), .A2(n3755), .ZN(n3758) );
  AOI31D0BWP12T U3867 ( .A1(n3759), .A2(n3758), .A3(n3757), .B(n3765), .ZN(
        n3761) );
  NR4D0BWP12T U3868 ( .A1(n3763), .A2(n3762), .A3(n3761), .A4(n3760), .ZN(
        n3764) );
  OAI21D0BWP12T U3869 ( .A1(n3766), .A2(n3765), .B(n3764), .ZN(n3802) );
  OAI22D0BWP12T U3870 ( .A1(n3769), .A2(n4044), .B1(n3768), .B2(n3767), .ZN(
        n3771) );
  RCAOI211D0BWP12T U3871 ( .A1(n3919), .A2(n3772), .B(n3771), .C(n3770), .ZN(
        n4196) );
  AOI211D0BWP12T U3872 ( .A1(n3774), .A2(n3997), .B(n4196), .C(n3773), .ZN(
        n3778) );
  ND4D0BWP12T U3873 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(
        n3801) );
  INVD0BWP12T U3874 ( .I(n3779), .ZN(n3793) );
  OAI22D0BWP12T U3875 ( .A1(n3783), .A2(n3782), .B1(n3781), .B2(n3780), .ZN(
        n3790) );
  OAI22D0BWP12T U3876 ( .A1(n3787), .A2(n3786), .B1(n3785), .B2(n3784), .ZN(
        n3789) );
  TPOAI21D0BWP12T U3877 ( .A1(n3790), .A2(n3789), .B(n3788), .ZN(n3791) );
  OAI211D1BWP12T U3878 ( .A1(n3793), .A2(n3792), .B(n3791), .C(n3986), .ZN(
        n3794) );
  AOI21D1BWP12T U3879 ( .A1(n3795), .A2(n3919), .B(n3794), .ZN(n4155) );
  ND4D0BWP12T U3880 ( .A1(n3799), .A2(n3798), .A3(n3797), .A4(n3796), .ZN(
        n3800) );
  NR4D0BWP12T U3881 ( .A1(n3802), .A2(n3801), .A3(n4155), .A4(n3800), .ZN(
        n3814) );
  ND4D0BWP12T U3882 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(
        n3809) );
  NR4D0BWP12T U3883 ( .A1(n3810), .A2(n3809), .A3(n3808), .A4(n3807), .ZN(
        n3813) );
  ND4D0BWP12T U3884 ( .A1(n3814), .A2(n3813), .A3(n3812), .A4(n3811), .ZN(
        n4007) );
  AOI22D1BWP12T U3885 ( .A1(n4070), .A2(n3815), .B1(n1706), .B2(n4157), .ZN(
        n3825) );
  AOI22D0BWP12T U3886 ( .A1(n4069), .A2(n3817), .B1(n3816), .B2(a[23]), .ZN(
        n3824) );
  AOI22D0BWP12T U3887 ( .A1(n3820), .A2(n3819), .B1(n3818), .B2(a[21]), .ZN(
        n3823) );
  AOI22D0BWP12T U3888 ( .A1(n4183), .A2(n3821), .B1(n1714), .B2(a[19]), .ZN(
        n3822) );
  ND4D1BWP12T U3889 ( .A1(n3825), .A2(n3824), .A3(n3823), .A4(n3822), .ZN(
        n3861) );
  AOI22D1BWP12T U3890 ( .A1(a[14]), .A2(n3827), .B1(n3826), .B2(a[17]), .ZN(
        n3837) );
  AOI22D1BWP12T U3891 ( .A1(n4078), .A2(n3829), .B1(n3828), .B2(n4082), .ZN(
        n3836) );
  AOI22D0BWP12T U3892 ( .A1(n4061), .A2(n3831), .B1(n3830), .B2(a[13]), .ZN(
        n3835) );
  AOI22D0BWP12T U3893 ( .A1(n4060), .A2(n3833), .B1(n3832), .B2(n4062), .ZN(
        n3834) );
  ND4D1BWP12T U3894 ( .A1(n3837), .A2(n3836), .A3(n3835), .A4(n3834), .ZN(
        n3860) );
  AOI22D0BWP12T U3895 ( .A1(n4083), .A2(n3839), .B1(n3838), .B2(n4063), .ZN(
        n3847) );
  AOI22D0BWP12T U3896 ( .A1(n4081), .A2(n3841), .B1(n3840), .B2(n4084), .ZN(
        n3846) );
  AOI22D0BWP12T U3897 ( .A1(n4067), .A2(n3886), .B1(n3842), .B2(n4075), .ZN(
        n3845) );
  CKND0BWP12T U3898 ( .I(b[0]), .ZN(n3843) );
  AOI22D0BWP12T U3899 ( .A1(n3885), .A2(n4044), .B1(n3843), .B2(n4066), .ZN(
        n3844) );
  ND4D1BWP12T U3900 ( .A1(n3847), .A2(n3846), .A3(n3845), .A4(n3844), .ZN(
        n3859) );
  AOI22D1BWP12T U3901 ( .A1(n4065), .A2(n3849), .B1(n3848), .B2(a[30]), .ZN(
        n3857) );
  AOI22D1BWP12T U3902 ( .A1(n4076), .A2(n3850), .B1(n2169), .B2(a[29]), .ZN(
        n3856) );
  AOI22D1BWP12T U3903 ( .A1(n4064), .A2(n3852), .B1(n3851), .B2(n4077), .ZN(
        n3855) );
  CKND2D0BWP12T U3904 ( .A1(n3853), .A2(n581), .ZN(n3854) );
  ND4D1BWP12T U3905 ( .A1(n3857), .A2(n3856), .A3(n3855), .A4(n3854), .ZN(
        n3858) );
  NR4D0BWP12T U3906 ( .A1(n3861), .A2(n3860), .A3(n3859), .A4(n3858), .ZN(
        n3965) );
  AOI22D0BWP12T U3907 ( .A1(n3943), .A2(n3863), .B1(n3941), .B2(n3862), .ZN(
        n3872) );
  AOI22D0BWP12T U3908 ( .A1(n3938), .A2(n3865), .B1(n3939), .B2(n3864), .ZN(
        n3871) );
  AOI22D0BWP12T U3909 ( .A1(n3951), .A2(n3867), .B1(b[19]), .B2(n3866), .ZN(
        n3870) );
  AOI22D1BWP12T U3910 ( .A1(n4191), .A2(n4187), .B1(n3952), .B2(n3868), .ZN(
        n3869) );
  ND4D1BWP12T U3911 ( .A1(n3872), .A2(n3871), .A3(n3870), .A4(n3869), .ZN(
        n3915) );
  AOI22D0BWP12T U3912 ( .A1(n3949), .A2(n3874), .B1(n3930), .B2(n3873), .ZN(
        n3884) );
  AOI22D0BWP12T U3913 ( .A1(n3950), .A2(n3876), .B1(n3931), .B2(n3875), .ZN(
        n3883) );
  AOI22D0BWP12T U3914 ( .A1(n3933), .A2(n3878), .B1(n3932), .B2(n3877), .ZN(
        n3882) );
  AOI22D1BWP12T U3915 ( .A1(n3928), .A2(n3880), .B1(n3957), .B2(n3879), .ZN(
        n3881) );
  ND4D1BWP12T U3916 ( .A1(n3884), .A2(n3883), .A3(n3882), .A4(n3881), .ZN(
        n3914) );
  OAI22D0BWP12T U3917 ( .A1(n4067), .A2(n3886), .B1(n4044), .B2(n3885), .ZN(
        n3889) );
  CKND0BWP12T U3918 ( .I(n3887), .ZN(n3888) );
  AOI211D0BWP12T U3919 ( .A1(n3916), .A2(n484), .B(n3889), .C(n3888), .ZN(
        n3909) );
  AOI22D0BWP12T U3920 ( .A1(n3929), .A2(n3891), .B1(n3927), .B2(n3890), .ZN(
        n3908) );
  AOI22D0BWP12T U3921 ( .A1(n3919), .A2(n3893), .B1(n3920), .B2(n3892), .ZN(
        n3907) );
  AOI22D1BWP12T U3922 ( .A1(n3944), .A2(n3895), .B1(b[29]), .B2(n3894), .ZN(
        n3903) );
  AOI22D0BWP12T U3923 ( .A1(n3942), .A2(n3897), .B1(n3917), .B2(n3896), .ZN(
        n3902) );
  AOI22D1BWP12T U3924 ( .A1(n3918), .A2(n3898), .B1(b[25]), .B2(n4160), .ZN(
        n3901) );
  AOI21D0BWP12T U3925 ( .A1(n3899), .A2(n3940), .B(n4182), .ZN(n3900) );
  ND4D1BWP12T U3926 ( .A1(n3903), .A2(n3902), .A3(n3901), .A4(n3900), .ZN(
        n3904) );
  NR2D0BWP12T U3927 ( .A1(n3905), .A2(n3904), .ZN(n3906) );
  ND4D1BWP12T U3928 ( .A1(n3909), .A2(n3908), .A3(n3907), .A4(n3906), .ZN(
        n3913) );
  OAI21D0BWP12T U3929 ( .A1(b[31]), .A2(n3911), .B(n3910), .ZN(n3912) );
  OAI31D1BWP12T U3930 ( .A1(n3915), .A2(n3914), .A3(n3913), .B(n3912), .ZN(
        n3964) );
  AOI22D0BWP12T U3931 ( .A1(n3917), .A2(n4076), .B1(n3916), .B2(n496), .ZN(
        n3926) );
  AOI22D0BWP12T U3932 ( .A1(n3918), .A2(n4064), .B1(b[25]), .B2(n4157), .ZN(
        n3925) );
  AOI22D0BWP12T U3933 ( .A1(n3920), .A2(n4075), .B1(n3919), .B2(n4081), .ZN(
        n3924) );
  AOI22D0BWP12T U3934 ( .A1(n3922), .A2(n4068), .B1(n3921), .B2(n4067), .ZN(
        n3923) );
  ND4D1BWP12T U3935 ( .A1(n3926), .A2(n3925), .A3(n3924), .A4(n3923), .ZN(
        n3962) );
  AOI22D0BWP12T U3936 ( .A1(n3928), .A2(n4062), .B1(n3927), .B2(n4083), .ZN(
        n3937) );
  AOI22D0BWP12T U3937 ( .A1(n4089), .A2(b[31]), .B1(n3929), .B2(n4084), .ZN(
        n3936) );
  AOI22D0BWP12T U3938 ( .A1(n3931), .A2(a[13]), .B1(n3930), .B2(a[14]), .ZN(
        n3935) );
  AOI22D0BWP12T U3939 ( .A1(n3933), .A2(n4060), .B1(n3932), .B2(n4061), .ZN(
        n3934) );
  ND4D1BWP12T U3940 ( .A1(n3937), .A2(n3936), .A3(n3935), .A4(n3934), .ZN(
        n3961) );
  AOI22D0BWP12T U3941 ( .A1(n3939), .A2(a[21]), .B1(n3938), .B2(n4069), .ZN(
        n3948) );
  AOI22D0BWP12T U3942 ( .A1(n3941), .A2(n4070), .B1(n3940), .B2(a[30]), .ZN(
        n3947) );
  AOI22D0BWP12T U3943 ( .A1(n3942), .A2(n4077), .B1(b[29]), .B2(a[29]), .ZN(
        n3946) );
  AOI22D0BWP12T U3944 ( .A1(n3944), .A2(n4065), .B1(n3943), .B2(a[23]), .ZN(
        n3945) );
  ND4D1BWP12T U3945 ( .A1(n3948), .A2(n3947), .A3(n3946), .A4(n3945), .ZN(
        n3960) );
  AOI22D0BWP12T U3946 ( .A1(n3950), .A2(n4078), .B1(n3949), .B2(n4082), .ZN(
        n3955) );
  AOI22D0BWP12T U3947 ( .A1(n3951), .A2(a[18]), .B1(n4191), .B2(n4183), .ZN(
        n3954) );
  AOI22D0BWP12T U3948 ( .A1(b[19]), .A2(a[19]), .B1(n3952), .B2(a[17]), .ZN(
        n3953) );
  ND3D1BWP12T U3949 ( .A1(n3955), .A2(n3954), .A3(n3953), .ZN(n3956) );
  AOI211D0BWP12T U3950 ( .A1(n3957), .A2(n4063), .B(n2664), .C(n3956), .ZN(
        n3958) );
  IOA21D0BWP12T U3951 ( .A1(b[0]), .A2(n4066), .B(n3958), .ZN(n3959) );
  NR4D0BWP12T U3952 ( .A1(n3962), .A2(n3961), .A3(n3960), .A4(n3959), .ZN(
        n3963) );
  AOI21D1BWP12T U3953 ( .A1(n3965), .A2(n3964), .B(n3963), .ZN(n4006) );
  CKND2D0BWP12T U3954 ( .A1(n3967), .A2(n3966), .ZN(n3970) );
  AOI211D0BWP12T U3955 ( .A1(n3986), .A2(n3970), .B(n3969), .C(n3968), .ZN(
        n4004) );
  ND4D0BWP12T U3956 ( .A1(n3974), .A2(n3973), .A3(n3972), .A4(n3971), .ZN(
        n3984) );
  CKND0BWP12T U3957 ( .I(n3975), .ZN(n3980) );
  CKND2D0BWP12T U3958 ( .A1(n3977), .A2(n3976), .ZN(n3979) );
  OAI211D0BWP12T U3959 ( .A1(n3981), .A2(n3980), .B(n3979), .C(n3978), .ZN(
        n3983) );
  NR4D0BWP12T U3960 ( .A1(n3985), .A2(n3984), .A3(n3983), .A4(n3982), .ZN(
        n4003) );
  OAI31D0BWP12T U3961 ( .A1(n3989), .A2(n3988), .A3(n3987), .B(n3986), .ZN(
        n4002) );
  IND4D0BWP12T U3962 ( .A1(n4158), .B1(n3991), .B2(n4199), .B3(n3990), .ZN(
        n4000) );
  CKND0BWP12T U3963 ( .I(n3992), .ZN(n3996) );
  ND4D0BWP12T U3964 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(
        n3998) );
  OAI31D0BWP12T U3965 ( .A1(n4000), .A2(n3999), .A3(n3998), .B(n3997), .ZN(
        n4001) );
  ND4D1BWP12T U3966 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(
        n4005) );
  ND3D1BWP12T U3967 ( .A1(n4007), .A2(n4006), .A3(n4005), .ZN(n4008) );
  AOI21D1BWP12T U3968 ( .A1(n4010), .A2(n4009), .B(n4008), .ZN(n4093) );
  OAI211D0BWP12T U3969 ( .A1(n4014), .A2(n4013), .B(n4012), .C(n4011), .ZN(
        n4015) );
  NR4D0BWP12T U3970 ( .A1(n4018), .A2(n4017), .A3(n4016), .A4(n4015), .ZN(
        n4028) );
  NR2D0BWP12T U3971 ( .A1(n4020), .A2(n4019), .ZN(n4027) );
  NR4D0BWP12T U3972 ( .A1(n4024), .A2(n4023), .A3(n4022), .A4(n4021), .ZN(
        n4025) );
  ND4D0BWP12T U3973 ( .A1(n4028), .A2(n4027), .A3(n4026), .A4(n4025), .ZN(
        n4029) );
  OR4D0BWP12T U3974 ( .A1(n4032), .A2(n4031), .A3(n4030), .A4(n4029), .Z(n4059) );
  ND4D0BWP12T U3975 ( .A1(n4035), .A2(n4199), .A3(n4034), .A4(n4033), .ZN(
        n4037) );
  OAI31D0BWP12T U3976 ( .A1(n4039), .A2(n4038), .A3(n4037), .B(n4036), .ZN(
        n4040) );
  CKND2D0BWP12T U3977 ( .A1(n4041), .A2(n4040), .ZN(n4057) );
  INVD0BWP12T U3978 ( .I(n4042), .ZN(n4045) );
  AOI21D0BWP12T U3979 ( .A1(n4045), .A2(n4044), .B(n4043), .ZN(n4161) );
  AOI21D0BWP12T U3980 ( .A1(n4047), .A2(n4161), .B(n4046), .ZN(n4049) );
  NR4D0BWP12T U3981 ( .A1(n4051), .A2(n4050), .A3(n4049), .A4(n4048), .ZN(
        n4055) );
  ND4D0BWP12T U3982 ( .A1(n4055), .A2(n4054), .A3(n4053), .A4(n4052), .ZN(
        n4056) );
  NR4D0BWP12T U3983 ( .A1(n4059), .A2(n4058), .A3(n4057), .A4(n4056), .ZN(
        n4091) );
  ND4D0BWP12T U3984 ( .A1(n4063), .A2(n4062), .A3(n4061), .A4(n4060), .ZN(
        n4074) );
  ND4D0BWP12T U3985 ( .A1(a[29]), .A2(n4065), .A3(n4157), .A4(n4064), .ZN(
        n4073) );
  ND4D0BWP12T U3986 ( .A1(n4068), .A2(n4067), .A3(n496), .A4(n4066), .ZN(n4072) );
  ND4D0BWP12T U3987 ( .A1(a[23]), .A2(n4070), .A3(a[21]), .A4(n4069), .ZN(
        n4071) );
  NR4D0BWP12T U3988 ( .A1(n4074), .A2(n4073), .A3(n4072), .A4(n4071), .ZN(
        n4088) );
  ND4D0BWP12T U3989 ( .A1(a[19]), .A2(n4077), .A3(n4076), .A4(n4075), .ZN(
        n4087) );
  ND4D0BWP12T U3990 ( .A1(a[17]), .A2(n4183), .A3(a[13]), .A4(n4078), .ZN(
        n4079) );
  NR2D0BWP12T U3991 ( .A1(n2205), .A2(n4079), .ZN(n4080) );
  ND4D0BWP12T U3992 ( .A1(a[14]), .A2(n4082), .A3(n4081), .A4(n4080), .ZN(
        n4086) );
  ND4D0BWP12T U3993 ( .A1(a[18]), .A2(a[30]), .A3(n4084), .A4(n4083), .ZN(
        n4085) );
  INR4D0BWP12T U3994 ( .A1(n4088), .B1(n4087), .B2(n4086), .B3(n4085), .ZN(
        n4090) );
  MUX2ND0BWP12T U3995 ( .I0(n4091), .I1(n4090), .S(n4089), .ZN(n4092) );
  ND3D1BWP12T U3996 ( .A1(n4094), .A2(n4093), .A3(n4092), .ZN(n4144) );
  NR4D0BWP12T U3997 ( .A1(n4098), .A2(n4097), .A3(n4096), .A4(n4095), .ZN(
        n4130) );
  NR4D0BWP12T U3998 ( .A1(n4102), .A2(n4101), .A3(n4100), .A4(n4099), .ZN(
        n4129) );
  NR4D0BWP12T U3999 ( .A1(n4105), .A2(n4104), .A3(n4103), .A4(n4164), .ZN(
        n4111) );
  NR4D0BWP12T U4000 ( .A1(n4109), .A2(n4108), .A3(n4107), .A4(n4106), .ZN(
        n4110) );
  IND3D1BWP12T U4001 ( .A1(n4112), .B1(n4111), .B2(n4110), .ZN(n4115) );
  NR4D0BWP12T U4002 ( .A1(n4116), .A2(n4115), .A3(n4114), .A4(n4113), .ZN(
        n4128) );
  TPOAI21D0BWP12T U4003 ( .A1(n4119), .A2(n4118), .B(n4117), .ZN(n4123) );
  CKND2D0BWP12T U4004 ( .A1(n4121), .A2(n4120), .ZN(n4122) );
  XNR2D1BWP12T U4005 ( .A1(n4123), .A2(n4122), .ZN(n4209) );
  NR4D0BWP12T U4006 ( .A1(n4126), .A2(n4125), .A3(n4124), .A4(n4209), .ZN(
        n4127) );
  ND4D1BWP12T U4007 ( .A1(n4130), .A2(n4129), .A3(n4128), .A4(n4127), .ZN(
        n4132) );
  FA1D0BWP12T U4008 ( .A(n4157), .B(b[25]), .CI(n4131), .CO(n3002), .S(n4152)
         );
  OR4D1BWP12T U4009 ( .A1(n4134), .A2(n4133), .A3(n4132), .A4(n4152), .Z(n4136) );
  OR4D1BWP12T U4010 ( .A1(n4138), .A2(n4137), .A3(n4136), .A4(n4135), .Z(n4139) );
  NR4D0BWP12T U4011 ( .A1(n4142), .A2(n4141), .A3(n4140), .A4(n4139), .ZN(
        n4143) );
  OR3XD2BWP12T U4012 ( .A1(n4145), .A2(n4144), .A3(n4143), .Z(n4146) );
  NR3D1BWP12T U4013 ( .A1(n4148), .A2(n4147), .A3(n4146), .ZN(n4149) );
  OAI21D1BWP12T U4014 ( .A1(n4151), .A2(n4150), .B(n4149), .ZN(z) );
  AOI21D1BWP12T U4015 ( .A1(n4215), .A2(n4166), .B(n4165), .ZN(n4167) );
  IOA21D1BWP12T U4016 ( .A1(n4173), .A2(n4168), .B(n4167), .ZN(n4169) );
  ND2D1BWP12T U4017 ( .A1(n4172), .A2(n4171), .ZN(n4218) );
  CKND2D1BWP12T U4018 ( .A1(n4174), .A2(n4173), .ZN(n4213) );
  AOI222D0BWP12T U4019 ( .A1(n4180), .A2(n4179), .B1(n4178), .B2(n4177), .C1(
        n4176), .C2(n4175), .ZN(n4202) );
  OAI21D0BWP12T U4020 ( .A1(n4183), .A2(n4182), .B(n4181), .ZN(n4190) );
  MUX2ND0BWP12T U4021 ( .I0(n4184), .I1(n2664), .S(n4191), .ZN(n4186) );
  NR2D0BWP12T U4022 ( .A1(n4186), .A2(n4185), .ZN(n4188) );
  MUX2ND0BWP12T U4023 ( .I0(n4188), .I1(n2205), .S(n4187), .ZN(n4189) );
  RCAOI21D0BWP12T U4024 ( .A1(n4191), .A2(n4190), .B(n4189), .ZN(n4192) );
  CKND2D1BWP12T U4025 ( .A1(n4193), .A2(n4192), .ZN(n4194) );
  AOI21D1BWP12T U4026 ( .A1(n4196), .A2(n4195), .B(n4194), .ZN(n4197) );
  OAI21D1BWP12T U4027 ( .A1(n4199), .A2(n4198), .B(n4197), .ZN(n4200) );
  IAO21D1BWP12T U4028 ( .A1(n4202), .A2(n4201), .B(n4200), .ZN(n4212) );
  CKND2D1BWP12T U4029 ( .A1(n4204), .A2(n4203), .ZN(n4205) );
  IOA21D1BWP12T U4030 ( .A1(n4207), .A2(n4206), .B(n4205), .ZN(n4208) );
  AOI21D1BWP12T U4031 ( .A1(n4210), .A2(n4209), .B(n4208), .ZN(n4211) );
  ND3D1BWP12T U4032 ( .A1(n4213), .A2(n4212), .A3(n4211), .ZN(n4214) );
  AOI21D1BWP12T U4033 ( .A1(n4216), .A2(n4215), .B(n4214), .ZN(n4217) );
  ND2D1BWP12T U4034 ( .A1(n4218), .A2(n4217), .ZN(result[16]) );
endmodule


module top7 ( clk, reset, MEM_MEMCTRL_from_mem_data, 
        MEMCTRL_MEM_to_mem_read_enable, MEMCTRL_MEM_to_mem_write_enable, 
        MEMCTRL_MEM_to_mem_mem_enable, MEMCTRL_MEM_to_mem_address, 
        MEMCTRL_MEM_to_mem_data );
  input [15:0] MEM_MEMCTRL_from_mem_data;
  output [11:0] MEMCTRL_MEM_to_mem_address;
  output [15:0] MEMCTRL_MEM_to_mem_data;
  input clk, reset;
  output MEMCTRL_MEM_to_mem_read_enable, MEMCTRL_MEM_to_mem_write_enable,
         MEMCTRL_MEM_to_mem_mem_enable;
  wire   DEC_CPSR_update_flag_n, new_n, ALU_OUT_n, RF_OUT_n,
         DEC_CPSR_update_flag_c, new_c, ALU_OUT_c, RF_OUT_c,
         DEC_CPSR_update_flag_z, new_z, ALU_OUT_z, RF_OUT_z,
         DEC_CPSR_update_flag_v, new_v, ALU_OUT_v, RF_OUT_v,
         DEC_RF_alu_write_to_reg_enable, DEC_RF_memory_write_to_reg_enable,
         DEC_MISC_OUT_memory_address_source_is_reg,
         DEC_MEMCTRL_memorycontroller_sign_extend,
         DEC_MEMCTRL_memory_load_request, DEC_MEMCTRL_memory_store_request,
         DEC_IF_stall_to_instructionfetch, ALU_IN_c, irdecode_inst1_N912,
         irdecode_inst1_N911, irdecode_inst1_N907, irdecode_inst1_N906,
         irdecode_inst1_N707, irdecode_inst1_N706, irdecode_inst1_N705,
         irdecode_inst1_N704, irdecode_inst1_N703, irdecode_inst1_N702,
         irdecode_inst1_N701, irdecode_inst1_N546, irdecode_inst1_N545,
         irdecode_inst1_N544, irdecode_inst1_N543, irdecode_inst1_N542,
         irdecode_inst1_N541, irdecode_inst1_N540, irdecode_inst1_N539,
         irdecode_inst1_split_instruction, irdecode_inst1_next_step_0_,
         irdecode_inst1_next_step_1_, irdecode_inst1_next_step_2_,
         irdecode_inst1_next_step_3_, irdecode_inst1_next_step_4_,
         irdecode_inst1_next_step_5_, irdecode_inst1_next_step_6_,
         irdecode_inst1_next_step_7_, irdecode_inst1_itstate_0_,
         irdecode_inst1_itstate_1_, irdecode_inst1_itstate_2_,
         irdecode_inst1_itstate_3_, irdecode_inst1_itstate_4_,
         irdecode_inst1_itstate_5_, irdecode_inst1_itstate_6_,
         irdecode_inst1_itstate_7_,
         irdecode_inst1_next_alu_write_to_reg_enable,
         irdecode_inst1_next_update_flag_v, irdecode_inst1_next_update_flag_c,
         irdecode_inst1_next_update_flag_n,
         memory_interface_inst1_delayed_is_signed, Instruction_Fetch_inst1_N98,
         Instruction_Fetch_inst1_N97, Instruction_Fetch_inst1_N96,
         Instruction_Fetch_inst1_N95, Instruction_Fetch_inst1_N94,
         Instruction_Fetch_inst1_N93, Instruction_Fetch_inst1_N92,
         Instruction_Fetch_inst1_N91, Instruction_Fetch_inst1_N90,
         Instruction_Fetch_inst1_N89, Instruction_Fetch_inst1_N88,
         Instruction_Fetch_inst1_N87, Instruction_Fetch_inst1_N86,
         Instruction_Fetch_inst1_N85, Instruction_Fetch_inst1_N84,
         Instruction_Fetch_inst1_N83, Instruction_Fetch_inst1_N80,
         Instruction_Fetch_inst1_N79,
         Instruction_Fetch_inst1_first_instruction_fetched,
         Instruction_Fetch_inst1_fetched_instruction_reg_0_,
         Instruction_Fetch_inst1_fetched_instruction_reg_1_,
         Instruction_Fetch_inst1_fetched_instruction_reg_2_,
         Instruction_Fetch_inst1_fetched_instruction_reg_3_,
         Instruction_Fetch_inst1_fetched_instruction_reg_4_,
         Instruction_Fetch_inst1_fetched_instruction_reg_5_,
         Instruction_Fetch_inst1_fetched_instruction_reg_6_,
         Instruction_Fetch_inst1_fetched_instruction_reg_7_,
         Instruction_Fetch_inst1_fetched_instruction_reg_8_,
         Instruction_Fetch_inst1_fetched_instruction_reg_9_,
         Instruction_Fetch_inst1_fetched_instruction_reg_10_,
         Instruction_Fetch_inst1_fetched_instruction_reg_11_,
         Instruction_Fetch_inst1_fetched_instruction_reg_12_,
         Instruction_Fetch_inst1_fetched_instruction_reg_13_,
         Instruction_Fetch_inst1_fetched_instruction_reg_14_,
         Instruction_Fetch_inst1_fetched_instruction_reg_15_,
         Instruction_Fetch_inst1_currentState_0_,
         Instruction_Fetch_inst1_currentState_1_,
         memory_interface_inst1_fsm_N35, memory_interface_inst1_fsm_N34,
         memory_interface_inst1_fsm_N33, memory_interface_inst1_fsm_N32,
         memory_interface_inst1_fsm_state_0_,
         memory_interface_inst1_fsm_state_1_,
         memory_interface_inst1_fsm_state_2_,
         memory_interface_inst1_fsm_state_3_, n754, n777, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n822, n823, n824, n825, n826,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53;
  wire   [7:0] IF_DEC_instruction;
  wire   [4:0] DEC_RF_operand_a;
  wire   [4:0] DEC_RF_operand_b;
  wire   [31:0] DEC_RF_offset_b;
  wire   [4:0] DEC_ALU_alu_opcode;
  wire   [4:0] DEC_RF_alu_write_to_reg;
  wire   [4:0] DEC_RF_memory_write_to_reg;
  wire   [4:0] DEC_RF_memory_store_data_reg;
  wire   [4:0] DEC_RF_memory_store_address_reg;
  wire   [1:0] DEC_MEMCTRL_load_store_width;
  wire   [31:0] ALU_MISC_OUT_result;
  wire   [31:0] MEMCTRL_RF_IF_data_in;
  wire   [31:0] IF_RF_incremented_pc_out;
  wire   [31:0] RF_ALU_operand_a;
  wire   [31:0] RF_ALU_operand_b;
  wire   [31:0] RF_MEMCTRL_data_reg;
  wire   [12:2] RF_MEMCTRL_address_reg;
  wire   [31:0] RF_pc_out;
  wire   [11:0] MEMCTRL_IN_address;
  wire   [7:0] irdecode_inst1_step;
  wire   [15:0] memory_interface_inst1_delay_first_two_bytes_out;
  wire   [31:0] memory_interface_inst1_delay_data_in32;
  wire   [11:0] memory_interface_inst1_delay_addr_for_adder;

  register_file register_file_inst1 ( .readA_sel(DEC_RF_operand_a), 
        .readB_sel(DEC_RF_operand_b), .readC_sel(DEC_RF_memory_store_data_reg), 
        .readD_sel(DEC_RF_memory_store_address_reg), .write1_sel(
        DEC_RF_alu_write_to_reg), .write2_sel(DEC_RF_memory_write_to_reg), 
        .write1_en(DEC_RF_alu_write_to_reg_enable), .write2_en(
        DEC_RF_memory_write_to_reg_enable), .write1_in(ALU_MISC_OUT_result), 
        .write2_in(MEMCTRL_RF_IF_data_in), .immediate1_in({n864, n864, n864, 
        n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, 
        n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, 
        n864, n864, n864, n864, n864}), .immediate2_in(DEC_RF_offset_b), 
        .next_pc_in({IF_RF_incremented_pc_out[31], n1745, n1754, n1747, n1751, 
        n1746, n1753, n1752, n1749, n1748, IF_RF_incremented_pc_out[21], n1750, 
        IF_RF_incremented_pc_out[19], n1757, IF_RF_incremented_pc_out[17], 
        n1756, IF_RF_incremented_pc_out[15], n1755, 
        IF_RF_incremented_pc_out[13:2], MEMCTRL_IN_address[0], 
        IF_RF_incremented_pc_out[0]}), .next_cpsr_in({new_n, new_c, new_z, 
        new_v}), .next_sp_in({n864, n864, n864, n864, n864, n864, n864, n864, 
        n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, 
        n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864, n864}), .clk(clk), .reset(reset), .regA_out(RF_ALU_operand_a), .regB_out(
        RF_ALU_operand_b), .regC_out(RF_MEMCTRL_data_reg), .regD_out({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        RF_MEMCTRL_address_reg, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21}), .pc_out(RF_pc_out), .cpsr_out({RF_OUT_n, 
        RF_OUT_c, RF_OUT_z, RF_OUT_v}), .sp_out({SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53}), .next_pc_en_BAR(n754) );
  ALU_VARIABLE ALU_VARIABLE_inst1 ( .a({RF_ALU_operand_a[31:30], n1767, 
        RF_ALU_operand_a[28:24], n1766, RF_ALU_operand_a[22], n1765, 
        RF_ALU_operand_a[20], n1764, RF_ALU_operand_a[18:4], n1763, 
        RF_ALU_operand_a[2:0]}), .b({RF_ALU_operand_b[31:4], n1762, 
        RF_ALU_operand_b[2:1], n1761}), .op(DEC_ALU_alu_opcode[3:0]), .c_in(
        ALU_IN_c), .result(ALU_MISC_OUT_result), .c_out(ALU_OUT_c), .z(
        ALU_OUT_z), .n(ALU_OUT_n), .v(ALU_OUT_v) );
  CKAN2D2BWP12T irdecode_inst1_C5193 ( .A1(irdecode_inst1_next_step_7_), .A2(
        IF_DEC_instruction[7]), .Z(irdecode_inst1_N539) );
  CKAN2D2BWP12T irdecode_inst1_C5194 ( .A1(irdecode_inst1_next_step_6_), .A2(
        IF_DEC_instruction[6]), .Z(irdecode_inst1_N540) );
  CKAN2D2BWP12T irdecode_inst1_C5195 ( .A1(irdecode_inst1_next_step_5_), .A2(
        IF_DEC_instruction[5]), .Z(irdecode_inst1_N541) );
  CKAN2D2BWP12T irdecode_inst1_C5196 ( .A1(irdecode_inst1_next_step_4_), .A2(
        IF_DEC_instruction[4]), .Z(irdecode_inst1_N542) );
  CKAN2D2BWP12T irdecode_inst1_C5197 ( .A1(irdecode_inst1_next_step_3_), .A2(
        IF_DEC_instruction[3]), .Z(irdecode_inst1_N543) );
  CKAN2D2BWP12T irdecode_inst1_C5198 ( .A1(irdecode_inst1_next_step_2_), .A2(
        IF_DEC_instruction[2]), .Z(irdecode_inst1_N544) );
  CKAN2D2BWP12T irdecode_inst1_C5199 ( .A1(irdecode_inst1_next_step_1_), .A2(
        IF_DEC_instruction[1]), .Z(irdecode_inst1_N545) );
  CKAN2D2BWP12T irdecode_inst1_C5200 ( .A1(irdecode_inst1_next_step_0_), .A2(
        IF_DEC_instruction[0]), .Z(irdecode_inst1_N546) );
  CKAN2D2BWP12T irdecode_inst1_C5280 ( .A1(irdecode_inst1_next_step_6_), .A2(
        IF_DEC_instruction[6]), .Z(irdecode_inst1_N701) );
  CKAN2D2BWP12T irdecode_inst1_C5281 ( .A1(irdecode_inst1_next_step_5_), .A2(
        IF_DEC_instruction[5]), .Z(irdecode_inst1_N702) );
  CKAN2D2BWP12T irdecode_inst1_C5282 ( .A1(irdecode_inst1_next_step_4_), .A2(
        IF_DEC_instruction[4]), .Z(irdecode_inst1_N703) );
  CKAN2D2BWP12T irdecode_inst1_C5283 ( .A1(irdecode_inst1_next_step_3_), .A2(
        IF_DEC_instruction[3]), .Z(irdecode_inst1_N704) );
  CKAN2D2BWP12T irdecode_inst1_C5284 ( .A1(irdecode_inst1_next_step_2_), .A2(
        IF_DEC_instruction[2]), .Z(irdecode_inst1_N705) );
  CKAN2D2BWP12T irdecode_inst1_C5285 ( .A1(irdecode_inst1_next_step_1_), .A2(
        IF_DEC_instruction[1]), .Z(irdecode_inst1_N706) );
  CKAN2D2BWP12T irdecode_inst1_C5286 ( .A1(irdecode_inst1_next_step_0_), .A2(
        IF_DEC_instruction[0]), .Z(irdecode_inst1_N707) );
  CKAN2D2BWP12T irdecode_inst1_C2476 ( .A1(irdecode_inst1_next_step_1_), .A2(
        irdecode_inst1_next_step_0_), .Z(irdecode_inst1_N906) );
  CKAN2D2BWP12T irdecode_inst1_C2482 ( .A1(irdecode_inst1_N907), .A2(n1768), 
        .Z(irdecode_inst1_N911) );
  OR2XD4BWP12T irdecode_inst1_C2484 ( .A1(irdecode_inst1_next_step_1_), .A2(
        n1768), .Z(irdecode_inst1_N912) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_0_ ( .D(
        MEM_MEMCTRL_from_mem_data[8]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[0]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_1_ ( .D(
        MEM_MEMCTRL_from_mem_data[9]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[1]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_2_ ( .D(
        MEM_MEMCTRL_from_mem_data[10]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_3_ ( .D(
        MEM_MEMCTRL_from_mem_data[11]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_4_ ( .D(
        MEM_MEMCTRL_from_mem_data[12]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[4]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_5_ ( .D(
        MEM_MEMCTRL_from_mem_data[13]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[5]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_6_ ( .D(
        MEM_MEMCTRL_from_mem_data[14]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_7_ ( .D(
        MEM_MEMCTRL_from_mem_data[15]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_8_ ( .D(
        MEM_MEMCTRL_from_mem_data[0]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_9_ ( .D(
        MEM_MEMCTRL_from_mem_data[1]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_10_ ( .D(
        MEM_MEMCTRL_from_mem_data[2]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_11_ ( .D(
        MEM_MEMCTRL_from_mem_data[3]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[11]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_12_ ( .D(
        MEM_MEMCTRL_from_mem_data[4]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[12]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_13_ ( .D(
        MEM_MEMCTRL_from_mem_data[5]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[13]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_14_ ( .D(
        MEM_MEMCTRL_from_mem_data[6]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[14]) );
  DFQD1BWP12T memory_interface_inst1_delay_first_two_bytes_out_reg_15_ ( .D(
        MEM_MEMCTRL_from_mem_data[7]), .CP(clk), .Q(
        memory_interface_inst1_delay_first_two_bytes_out[15]) );
  DFQD1BWP12T irdecode_inst1_load_store_width_reg_0_ ( .D(n838), .CP(clk), .Q(
        DEC_MEMCTRL_load_store_width[0]) );
  DFQD1BWP12T irdecode_inst1_load_store_width_reg_1_ ( .D(n837), .CP(clk), .Q(
        DEC_MEMCTRL_load_store_width[1]) );
  DFQD1BWP12T irdecode_inst1_memory_load_request_reg ( .D(n861), .CP(clk), .Q(
        DEC_MEMCTRL_memory_load_request) );
  DFQD1BWP12T irdecode_inst1_stall_to_instructionfetch_reg ( .D(n845), .CP(clk), .Q(DEC_IF_stall_to_instructionfetch) );
  DFQD1BWP12T irdecode_inst1_step_reg_1_ ( .D(irdecode_inst1_next_step_1_), 
        .CP(clk), .Q(irdecode_inst1_step[1]) );
  DFQD1BWP12T irdecode_inst1_split_instruction_reg ( .D(n847), .CP(clk), .Q(
        irdecode_inst1_split_instruction) );
  DFQD1BWP12T irdecode_inst1_step_reg_6_ ( .D(irdecode_inst1_next_step_6_), 
        .CP(clk), .Q(irdecode_inst1_step[6]) );
  DFQD1BWP12T irdecode_inst1_step_reg_5_ ( .D(irdecode_inst1_next_step_5_), 
        .CP(clk), .Q(irdecode_inst1_step[5]) );
  DFQD1BWP12T irdecode_inst1_step_reg_0_ ( .D(irdecode_inst1_next_step_0_), 
        .CP(clk), .Q(irdecode_inst1_step[0]) );
  DFQD1BWP12T irdecode_inst1_step_reg_2_ ( .D(irdecode_inst1_next_step_2_), 
        .CP(clk), .Q(irdecode_inst1_step[2]) );
  DFQD1BWP12T irdecode_inst1_step_reg_3_ ( .D(irdecode_inst1_next_step_3_), 
        .CP(clk), .Q(irdecode_inst1_step[3]) );
  DFQD1BWP12T irdecode_inst1_step_reg_4_ ( .D(irdecode_inst1_next_step_4_), 
        .CP(clk), .Q(irdecode_inst1_step[4]) );
  DFQD1BWP12T irdecode_inst1_step_reg_7_ ( .D(irdecode_inst1_next_step_7_), 
        .CP(clk), .Q(irdecode_inst1_step[7]) );
  DFQD1BWP12T irdecode_inst1_memory_store_request_reg ( .D(n852), .CP(clk), 
        .Q(DEC_MEMCTRL_memory_store_request) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_0_ ( .D(n860), .CP(clk), .Q(
        irdecode_inst1_itstate_0_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_1_ ( .D(n859), .CP(clk), .Q(
        irdecode_inst1_itstate_1_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_2_ ( .D(n858), .CP(clk), .Q(
        irdecode_inst1_itstate_2_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_3_ ( .D(n857), .CP(clk), .Q(
        irdecode_inst1_itstate_3_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_4_ ( .D(n856), .CP(clk), .Q(
        irdecode_inst1_itstate_4_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_5_ ( .D(n855), .CP(clk), .Q(
        irdecode_inst1_itstate_5_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_6_ ( .D(n854), .CP(clk), .Q(
        irdecode_inst1_itstate_6_) );
  DFQD1BWP12T irdecode_inst1_itstate_reg_7_ ( .D(n853), .CP(clk), .Q(
        irdecode_inst1_itstate_7_) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_0_ ( .D(n835), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[0]) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_2_ ( .D(n833), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[2]) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_3_ ( .D(n832), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[3]) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_4_ ( .D(n831), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[4]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_0_ ( .D(n830), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[0]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_2_ ( .D(n828), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[2]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_3_ ( .D(n1759), .CP(clk), .Q(DEC_RF_memory_store_data_reg[3]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_4_ ( .D(n826), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[4]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_0_ ( .D(n824), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[0]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_2_ ( .D(n822), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[2]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_4_ ( .D(n848), .CP(clk), .Q(
        DEC_ALU_alu_opcode[4]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_3_ ( .D(n1758), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[3]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_4_ ( .D(n820), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[4]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_1_ ( .D(n850), .CP(clk), .Q(
        DEC_ALU_alu_opcode[1]) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_2_ ( .D(n846), .CP(clk), .Q(
        DEC_ALU_alu_opcode[2]) );
  DFQD1BWP12T irdecode_inst1_update_flag_v_reg ( .D(
        irdecode_inst1_next_update_flag_v), .CP(clk), .Q(
        DEC_CPSR_update_flag_v) );
  DFQD1BWP12T irdecode_inst1_update_flag_c_reg ( .D(
        irdecode_inst1_next_update_flag_c), .CP(clk), .Q(
        DEC_CPSR_update_flag_c) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_0_ ( .D(n851), .CP(clk), .Q(
        DEC_ALU_alu_opcode[0]) );
  DFQD1BWP12T irdecode_inst1_update_flag_n_reg ( .D(
        irdecode_inst1_next_update_flag_n), .CP(clk), .Q(
        DEC_CPSR_update_flag_n) );
  DFQD1BWP12T irdecode_inst1_update_flag_z_reg ( .D(
        irdecode_inst1_next_update_flag_n), .CP(clk), .Q(
        DEC_CPSR_update_flag_z) );
  DFQD1BWP12T irdecode_inst1_alu_opcode_reg_3_ ( .D(n849), .CP(clk), .Q(
        DEC_ALU_alu_opcode[3]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_2_ ( .D(n818), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[2]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_3_ ( .D(n817), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[3]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_4_ ( .D(n815), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[4]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_0_ ( .D(n816), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[0]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_enable_reg ( .D(
        irdecode_inst1_next_alu_write_to_reg_enable), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg_enable) );
  DFQD1BWP12T irdecode_inst1_memory_address_source_is_reg_reg ( .D(n836), .CP(
        clk), .Q(DEC_MISC_OUT_memory_address_source_is_reg) );
  DFQD1BWP12T irdecode_inst1_memory_store_address_reg_reg_1_ ( .D(n834), .CP(
        clk), .Q(DEC_RF_memory_store_address_reg[1]) );
  DFQD1BWP12T irdecode_inst1_memory_store_data_reg_reg_1_ ( .D(n829), .CP(clk), 
        .Q(DEC_RF_memory_store_data_reg[1]) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_enable_reg ( .D(n825), .CP(
        clk), .Q(DEC_RF_memory_write_to_reg_enable) );
  DFQD1BWP12T irdecode_inst1_memory_write_to_reg_reg_1_ ( .D(n823), .CP(clk), 
        .Q(DEC_RF_memory_write_to_reg[1]) );
  DFQD1BWP12T irdecode_inst1_alu_write_to_reg_reg_1_ ( .D(n819), .CP(clk), .Q(
        DEC_RF_alu_write_to_reg[1]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_0_ ( .D(n809), .CP(clk), .Q(
        DEC_RF_offset_b[0]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_1_ ( .D(n808), .CP(clk), .Q(
        DEC_RF_offset_b[1]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_2_ ( .D(n807), .CP(clk), .Q(
        DEC_RF_offset_b[2]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_3_ ( .D(n806), .CP(clk), .Q(
        DEC_RF_offset_b[3]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_4_ ( .D(n805), .CP(clk), .Q(
        DEC_RF_offset_b[4]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_5_ ( .D(n804), .CP(clk), .Q(
        DEC_RF_offset_b[5]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_6_ ( .D(n803), .CP(clk), .Q(
        DEC_RF_offset_b[6]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_7_ ( .D(n802), .CP(clk), .Q(
        DEC_RF_offset_b[7]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_8_ ( .D(n801), .CP(clk), .Q(
        DEC_RF_offset_b[8]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_9_ ( .D(n800), .CP(clk), .Q(
        DEC_RF_offset_b[9]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_10_ ( .D(n799), .CP(clk), .Q(
        DEC_RF_offset_b[10]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_11_ ( .D(n798), .CP(clk), .Q(
        DEC_RF_offset_b[11]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_12_ ( .D(n797), .CP(clk), .Q(
        DEC_RF_offset_b[12]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_13_ ( .D(n796), .CP(clk), .Q(
        DEC_RF_offset_b[13]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_14_ ( .D(n795), .CP(clk), .Q(
        DEC_RF_offset_b[14]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_15_ ( .D(n794), .CP(clk), .Q(
        DEC_RF_offset_b[15]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_16_ ( .D(n793), .CP(clk), .Q(
        DEC_RF_offset_b[16]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_17_ ( .D(n792), .CP(clk), .Q(
        DEC_RF_offset_b[17]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_18_ ( .D(n791), .CP(clk), .Q(
        DEC_RF_offset_b[18]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_19_ ( .D(n790), .CP(clk), .Q(
        DEC_RF_offset_b[19]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_20_ ( .D(n789), .CP(clk), .Q(
        DEC_RF_offset_b[20]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_21_ ( .D(n788), .CP(clk), .Q(
        DEC_RF_offset_b[21]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_22_ ( .D(n787), .CP(clk), .Q(
        DEC_RF_offset_b[22]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_23_ ( .D(n786), .CP(clk), .Q(
        DEC_RF_offset_b[23]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_24_ ( .D(n785), .CP(clk), .Q(
        DEC_RF_offset_b[24]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_25_ ( .D(n784), .CP(clk), .Q(
        DEC_RF_offset_b[25]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_1_ ( .D(
        MEMCTRL_IN_address[1]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[1]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_2_ ( .D(
        MEMCTRL_IN_address[2]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_3_ ( .D(
        MEMCTRL_IN_address[3]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_4_ ( .D(
        MEMCTRL_IN_address[4]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[4]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_5_ ( .D(
        MEMCTRL_IN_address[5]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[5]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_6_ ( .D(
        MEMCTRL_IN_address[6]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_7_ ( .D(
        MEMCTRL_IN_address[7]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_8_ ( .D(
        MEMCTRL_IN_address[8]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_9_ ( .D(
        MEMCTRL_IN_address[9]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_10_ ( .D(
        MEMCTRL_IN_address[10]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_11_ ( .D(
        MEMCTRL_IN_address[11]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[11]) );
  DFQD4BWP12T irdecode_inst1_operand_a_reg_4_ ( .D(n810), .CP(clk), .Q(
        DEC_RF_operand_a[4]) );
  DFQD4BWP12T irdecode_inst1_operand_a_reg_0_ ( .D(n811), .CP(clk), .Q(
        DEC_RF_operand_a[0]) );
  DFQD4BWP12T irdecode_inst1_operand_a_reg_3_ ( .D(n812), .CP(clk), .Q(
        DEC_RF_operand_a[3]) );
  DFQD4BWP12T irdecode_inst1_operand_a_reg_1_ ( .D(n814), .CP(clk), .Q(
        DEC_RF_operand_a[1]) );
  DFQD4BWP12T irdecode_inst1_operand_a_reg_2_ ( .D(n813), .CP(clk), .Q(
        DEC_RF_operand_a[2]) );
  DFQD4BWP12T irdecode_inst1_operand_b_reg_0_ ( .D(n844), .CP(clk), .Q(
        DEC_RF_operand_b[0]) );
  DFQD4BWP12T irdecode_inst1_operand_b_reg_2_ ( .D(n842), .CP(clk), .Q(
        DEC_RF_operand_b[2]) );
  DFQD4BWP12T irdecode_inst1_operand_b_reg_3_ ( .D(n841), .CP(clk), .Q(
        DEC_RF_operand_b[3]) );
  DFQD4BWP12T irdecode_inst1_operand_b_reg_1_ ( .D(n843), .CP(clk), .Q(
        DEC_RF_operand_b[1]) );
  DFQD4BWP12T irdecode_inst1_operand_b_reg_4_ ( .D(n840), .CP(clk), .Q(
        DEC_RF_operand_b[4]) );
  DFQD1BWP12T memory_interface_inst1_delayed_is_signed_reg ( .D(
        DEC_MEMCTRL_memorycontroller_sign_extend), .CP(clk), .Q(
        memory_interface_inst1_delayed_is_signed) );
  DFQD1BWP12T memory_interface_inst1_delay_addr_for_adder_reg_0_ ( .D(
        MEMCTRL_IN_address[0]), .CP(clk), .Q(
        memory_interface_inst1_delay_addr_for_adder[0]) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_1_ ( .D(
        memory_interface_inst1_fsm_N33), .CP(clk), .Q(
        memory_interface_inst1_fsm_state_1_) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_3_ ( .D(
        memory_interface_inst1_fsm_N35), .CP(clk), .Q(
        memory_interface_inst1_fsm_state_3_) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_2_ ( .D(
        memory_interface_inst1_fsm_N34), .CP(clk), .Q(
        memory_interface_inst1_fsm_state_2_) );
  DFQD1BWP12T memory_interface_inst1_fsm_state_reg_0_ ( .D(
        memory_interface_inst1_fsm_N32), .CP(clk), .Q(
        memory_interface_inst1_fsm_state_0_) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_31_ ( .D(
        RF_MEMCTRL_data_reg[31]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[31]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_3_ ( .D(
        RF_MEMCTRL_data_reg[3]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[3]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_2_ ( .D(
        RF_MEMCTRL_data_reg[2]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[2]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_21_ ( .D(
        RF_MEMCTRL_data_reg[21]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[21]) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_7_ ( .D(
        Instruction_Fetch_inst1_N90), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_7_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_6_ ( .D(
        Instruction_Fetch_inst1_N89), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_6_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_5_ ( .D(
        Instruction_Fetch_inst1_N88), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_5_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_4_ ( .D(
        Instruction_Fetch_inst1_N87), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_4_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_3_ ( .D(
        Instruction_Fetch_inst1_N86), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_3_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_2_ ( .D(
        Instruction_Fetch_inst1_N85), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_2_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_1_ ( .D(
        Instruction_Fetch_inst1_N84), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_1_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_0_ ( .D(
        Instruction_Fetch_inst1_N83), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_0_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_8_ ( .D(
        Instruction_Fetch_inst1_N91), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_8_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_12_ ( .D(
        Instruction_Fetch_inst1_N95), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_12_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_10_ ( .D(
        Instruction_Fetch_inst1_N93), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_10_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_9_ ( .D(
        Instruction_Fetch_inst1_N92), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_9_) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_11_ ( .D(
        Instruction_Fetch_inst1_N94), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_11_) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_13_ ( .D(
        RF_MEMCTRL_data_reg[13]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[13]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_23_ ( .D(
        RF_MEMCTRL_data_reg[23]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[23]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_0_ ( .D(
        RF_MEMCTRL_data_reg[0]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[0]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_5_ ( .D(
        RF_MEMCTRL_data_reg[5]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[5]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_9_ ( .D(
        RF_MEMCTRL_data_reg[9]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[9]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_19_ ( .D(
        RF_MEMCTRL_data_reg[19]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[19]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_16_ ( .D(
        RF_MEMCTRL_data_reg[16]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[16]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_30_ ( .D(
        RF_MEMCTRL_data_reg[30]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[30]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_27_ ( .D(
        RF_MEMCTRL_data_reg[27]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[27]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_29_ ( .D(
        RF_MEMCTRL_data_reg[29]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[29]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_28_ ( .D(
        RF_MEMCTRL_data_reg[28]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[28]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_25_ ( .D(
        RF_MEMCTRL_data_reg[25]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[25]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_20_ ( .D(
        RF_MEMCTRL_data_reg[20]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[20]) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_13_ ( .D(
        Instruction_Fetch_inst1_N96), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_13_) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_24_ ( .D(
        RF_MEMCTRL_data_reg[24]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[24]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_17_ ( .D(
        RF_MEMCTRL_data_reg[17]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[17]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_4_ ( .D(
        RF_MEMCTRL_data_reg[4]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[4]) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_15_ ( .D(
        Instruction_Fetch_inst1_N98), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_15_) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_14_ ( .D(
        RF_MEMCTRL_data_reg[14]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[14]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_22_ ( .D(
        RF_MEMCTRL_data_reg[22]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[22]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_26_ ( .D(
        RF_MEMCTRL_data_reg[26]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[26]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_6_ ( .D(
        RF_MEMCTRL_data_reg[6]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[6]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_11_ ( .D(
        RF_MEMCTRL_data_reg[11]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[11]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_10_ ( .D(
        RF_MEMCTRL_data_reg[10]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[10]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_12_ ( .D(
        RF_MEMCTRL_data_reg[12]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[12]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_7_ ( .D(
        RF_MEMCTRL_data_reg[7]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[7]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_18_ ( .D(
        RF_MEMCTRL_data_reg[18]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[18]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_8_ ( .D(
        RF_MEMCTRL_data_reg[8]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[8]) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_15_ ( .D(
        RF_MEMCTRL_data_reg[15]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[15]) );
  DFQD1BWP12T Instruction_Fetch_inst1_fetched_instruction_reg_reg_14_ ( .D(
        Instruction_Fetch_inst1_N97), .CP(clk), .Q(
        Instruction_Fetch_inst1_fetched_instruction_reg_14_) );
  DFQD1BWP12T memory_interface_inst1_delay_data_in32_reg_1_ ( .D(
        RF_MEMCTRL_data_reg[1]), .CP(clk), .Q(
        memory_interface_inst1_delay_data_in32[1]) );
  DFQD1BWP12T Instruction_Fetch_inst1_first_instruction_fetched_reg ( .D(n862), 
        .CP(clk), .Q(Instruction_Fetch_inst1_first_instruction_fetched) );
  DFQD1BWP12T irdecode_inst1_memorycontroller_sign_extend_reg ( .D(n839), .CP(
        clk), .Q(DEC_MEMCTRL_memorycontroller_sign_extend) );
  DFQD1BWP12T Instruction_Fetch_inst1_currentState_reg_1_ ( .D(
        Instruction_Fetch_inst1_N80), .CP(clk), .Q(
        Instruction_Fetch_inst1_currentState_1_) );
  DFQD1BWP12T Instruction_Fetch_inst1_currentState_reg_0_ ( .D(
        Instruction_Fetch_inst1_N79), .CP(clk), .Q(
        Instruction_Fetch_inst1_currentState_0_) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_31_ ( .D(n777), .CP(clk), .Q(
        DEC_RF_offset_b[31]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_30_ ( .D(n779), .CP(clk), .Q(
        DEC_RF_offset_b[30]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_29_ ( .D(n780), .CP(clk), .Q(
        DEC_RF_offset_b[29]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_28_ ( .D(n781), .CP(clk), .Q(
        DEC_RF_offset_b[28]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_27_ ( .D(n782), .CP(clk), .Q(
        DEC_RF_offset_b[27]) );
  DFQD1BWP12T irdecode_inst1_offset_b_reg_26_ ( .D(n783), .CP(clk), .Q(
        DEC_RF_offset_b[26]) );
  TIELBWP12T U1022 ( .ZN(n864) );
  INVD1BWP12T U1023 ( .I(n864), .ZN(MEMCTRL_MEM_to_mem_mem_enable) );
  NR2D1BWP12T U1024 ( .A1(memory_interface_inst1_fsm_state_0_), .A2(
        memory_interface_inst1_fsm_state_3_), .ZN(n1010) );
  OAI22D1BWP12T U1025 ( .A1(n1551), .A2(n1574), .B1(n1542), .B2(n1567), .ZN(
        n1122) );
  INR2D1BWP12T U1026 ( .A1(n1299), .B1(n1602), .ZN(n1584) );
  INVD1BWP12T U1027 ( .I(n1687), .ZN(n1711) );
  INVD1BWP12T U1028 ( .I(n1696), .ZN(n1738) );
  ND2D1BWP12T U1029 ( .A1(n1232), .A2(n1308), .ZN(n1743) );
  IND2D1BWP12T U1030 ( .A1(Instruction_Fetch_inst1_currentState_1_), .B1(
        Instruction_Fetch_inst1_currentState_0_), .ZN(n1132) );
  AN2D1BWP12T U1031 ( .A1(n1304), .A2(n1308), .Z(n1570) );
  INR4D0BWP12T U1032 ( .A1(n1205), .B1(n1095), .B2(IF_DEC_instruction[7]), 
        .B3(irdecode_inst1_N706), .ZN(n1099) );
  MAOI22D0BWP12T U1033 ( .A1(n1410), .A2(DEC_MEMCTRL_memory_load_request), 
        .B1(n1449), .B2(n1511), .ZN(n1087) );
  ND3D0BWP12T U1034 ( .A1(IF_DEC_instruction[7]), .A2(n1220), .A3(n1102), .ZN(
        n1530) );
  CKND0BWP12T U1035 ( .I(n1226), .ZN(n865) );
  OA211D0BWP12T U1036 ( .A1(n1088), .A2(n865), .B(n1552), .C(n1553), .Z(n1643)
         );
  IOA21D0BWP12T U1037 ( .A1(n1731), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[11]), .B(n1034), .ZN(
        n866) );
  AO21D0BWP12T U1038 ( .A1(MEM_MEMCTRL_from_mem_data[3]), .A2(n1033), .B(n866), 
        .Z(MEMCTRL_RF_IF_data_in[11]) );
  IIND4D1BWP12T U1039 ( .A1(irdecode_inst1_N706), .A2(n1096), .B1(
        irdecode_inst1_N704), .B2(n1102), .ZN(n1209) );
  IND2D0BWP12T U1040 ( .A1(n1417), .B1(n1415), .ZN(n1418) );
  NR4D0BWP12T U1041 ( .A1(n1277), .A2(n1606), .A3(n1699), .A4(n1671), .ZN(
        n1547) );
  IOA21D0BWP12T U1042 ( .A1(n1710), .A2(n1739), .B(n1713), .ZN(n1635) );
  IAO21D0BWP12T U1043 ( .A1(n1551), .A2(n1640), .B(n1732), .ZN(n1697) );
  CKND0BWP12T U1044 ( .I(n1554), .ZN(n867) );
  OAI32D0BWP12T U1045 ( .A1(n1071), .A2(irdecode_inst1_N541), .A3(n867), .B1(
        n1527), .B2(n1071), .ZN(n868) );
  INR2D0BWP12T U1046 ( .A1(n1641), .B1(n868), .ZN(n1067) );
  CKND0BWP12T U1047 ( .I(n1413), .ZN(n869) );
  OA21D0BWP12T U1048 ( .A1(n1008), .A2(n869), .B(n1728), .Z(n1015) );
  AN3D0BWP12T U1049 ( .A1(n1534), .A2(n1223), .A3(n1545), .Z(n1252) );
  IIND4D1BWP12T U1050 ( .A1(n1096), .A2(irdecode_inst1_N704), .B1(
        irdecode_inst1_N706), .B2(n1102), .ZN(n1218) );
  IND3D0BWP12T U1051 ( .A1(n1236), .B1(n1523), .B2(n870), .ZN(n1690) );
  CKND0BWP12T U1052 ( .I(n1110), .ZN(n870) );
  NR2D1BWP12T U1053 ( .A1(n1603), .A2(irdecode_inst1_N539), .ZN(n871) );
  ND2D1BWP12T U1054 ( .A1(n871), .A2(n1075), .ZN(n1405) );
  ND3D1BWP12T U1055 ( .A1(irdecode_inst1_N703), .A2(n1220), .A3(n1533), .ZN(
        n1545) );
  IOA21D0BWP12T U1056 ( .A1(n1479), .A2(n1485), .B(n1486), .ZN(n1483) );
  AOI21D0BWP12T U1057 ( .A1(n1361), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_12_), .B(n1031), .ZN(
        n872) );
  IOA21D0BWP12T U1058 ( .A1(n1016), .A2(MEMCTRL_RF_IF_data_in[12]), .B(n872), 
        .ZN(n1111) );
  IND2D0BWP12T U1059 ( .A1(n1083), .B1(n1551), .ZN(n1552) );
  IOA21D0BWP12T U1060 ( .A1(n1479), .A2(n1475), .B(n1486), .ZN(n1473) );
  IND2D0BWP12T U1061 ( .A1(n1405), .B1(n1570), .ZN(n1538) );
  INR3D0BWP12T U1062 ( .A1(n1112), .B1(n1114), .B2(n1111), .ZN(n1735) );
  INR2D0BWP12T U1063 ( .A1(n1544), .B1(n1562), .ZN(n1568) );
  IOA21D1BWP12T U1064 ( .A1(n1731), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[8]), .B(n1034), .ZN(
        n873) );
  AO21D1BWP12T U1065 ( .A1(MEM_MEMCTRL_from_mem_data[0]), .A2(n1033), .B(n873), 
        .Z(MEMCTRL_RF_IF_data_in[8]) );
  AOI31D0BWP12T U1066 ( .A1(n1256), .A2(n1255), .A3(n1240), .B(n1668), .ZN(
        n874) );
  CKND2D0BWP12T U1067 ( .A1(n1567), .A2(n1574), .ZN(n875) );
  AOI21D0BWP12T U1068 ( .A1(n875), .A2(n1696), .B(n874), .ZN(n1539) );
  CKND0BWP12T U1069 ( .I(n1550), .ZN(n876) );
  MAOI22D0BWP12T U1070 ( .A1(n1551), .A2(n876), .B1(n1084), .B2(n1564), .ZN(
        n877) );
  AOI21D0BWP12T U1071 ( .A1(n1643), .A2(n877), .B(n1640), .ZN(n1732) );
  CKND0BWP12T U1072 ( .I(n1509), .ZN(n878) );
  AOI222D0BWP12T U1073 ( .A1(n878), .A2(RF_MEMCTRL_data_reg[16]), .B1(n1506), 
        .B2(memory_interface_inst1_delay_data_in32[0]), .C1(n1507), .C2(
        memory_interface_inst1_delay_data_in32[16]), .ZN(n879) );
  IOA21D0BWP12T U1074 ( .A1(n1508), .A2(RF_MEMCTRL_data_reg[0]), .B(n879), 
        .ZN(MEMCTRL_MEM_to_mem_data[8]) );
  CKND2D0BWP12T U1075 ( .A1(n1530), .A2(n1531), .ZN(n880) );
  AOI211D1BWP12T U1076 ( .A1(n1533), .A2(irdecode_inst1_N706), .B(n1532), .C(
        n880), .ZN(n881) );
  AOI31D1BWP12T U1077 ( .A1(n1543), .A2(n881), .A3(n1534), .B(n1567), .ZN(n882) );
  AN4D0BWP12T U1078 ( .A1(n1528), .A2(n1529), .A3(n1553), .A4(n1549), .Z(n883)
         );
  ND2D1BWP12T U1079 ( .A1(n1526), .A2(irdecode_inst1_N545), .ZN(n884) );
  AOI31D1BWP12T U1080 ( .A1(n1527), .A2(n883), .A3(n884), .B(n1574), .ZN(n885)
         );
  OAI21D0BWP12T U1081 ( .A1(n1536), .A2(n1634), .B(n1535), .ZN(n886) );
  NR4D0BWP12T U1082 ( .A1(n882), .A2(n1572), .A3(n885), .A4(n886), .ZN(n1580)
         );
  AOI21D0BWP12T U1083 ( .A1(n1361), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_10_), .B(n1031), .ZN(
        n887) );
  IOA21D0BWP12T U1084 ( .A1(n1016), .A2(MEMCTRL_RF_IF_data_in[10]), .B(n887), 
        .ZN(n1701) );
  CKND0BWP12T U1085 ( .I(n1509), .ZN(n888) );
  AOI222D0BWP12T U1086 ( .A1(n888), .A2(RF_MEMCTRL_data_reg[17]), .B1(n1506), 
        .B2(memory_interface_inst1_delay_data_in32[1]), .C1(n1507), .C2(
        memory_interface_inst1_delay_data_in32[17]), .ZN(n889) );
  IOA21D0BWP12T U1087 ( .A1(RF_MEMCTRL_data_reg[1]), .A2(n1508), .B(n889), 
        .ZN(MEMCTRL_MEM_to_mem_data[9]) );
  NR2D1BWP12T U1088 ( .A1(irdecode_inst1_N543), .A2(irdecode_inst1_N545), .ZN(
        n890) );
  ND2D1BWP12T U1089 ( .A1(n890), .A2(n1076), .ZN(n1063) );
  CKND0BWP12T U1090 ( .I(n1144), .ZN(n891) );
  AOI21D0BWP12T U1091 ( .A1(memory_interface_inst1_delayed_is_signed), .A2(
        n891), .B(n1145), .ZN(n892) );
  ND3D0BWP12T U1092 ( .A1(n1143), .A2(memory_interface_inst1_delayed_is_signed), .A3(MEM_MEMCTRL_from_mem_data[7]), .ZN(n893) );
  MOAI22D0BWP12T U1093 ( .A1(n892), .A2(MEM_MEMCTRL_from_mem_data[15]), .B1(
        n892), .B2(n893), .ZN(n1730) );
  AN3XD2BWP12T U1094 ( .A1(n1207), .A2(n1099), .A3(irdecode_inst1_N707), .Z(
        n1219) );
  INR2D0BWP12T U1095 ( .A1(n1527), .B1(n1554), .ZN(n1564) );
  IOA21D1BWP12T U1096 ( .A1(n1731), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[14]), .B(n1034), .ZN(
        n894) );
  AO21D1BWP12T U1097 ( .A1(MEM_MEMCTRL_from_mem_data[6]), .A2(n1033), .B(n894), 
        .Z(MEMCTRL_RF_IF_data_in[14]) );
  CKND0BWP12T U1098 ( .I(n1522), .ZN(n895) );
  OAI32D0BWP12T U1099 ( .A1(n1713), .A2(n1295), .A3(n895), .B1(n1264), .B2(
        n1713), .ZN(n1611) );
  INR4D0BWP12T U1100 ( .A1(n1640), .B1(n1606), .B2(n1735), .B3(n1275), .ZN(
        n1283) );
  CKND0BWP12T U1101 ( .I(n1509), .ZN(n896) );
  AOI222D0BWP12T U1102 ( .A1(n896), .A2(RF_MEMCTRL_data_reg[18]), .B1(n1506), 
        .B2(memory_interface_inst1_delay_data_in32[2]), .C1(n1507), .C2(
        memory_interface_inst1_delay_data_in32[18]), .ZN(n897) );
  IOA21D0BWP12T U1103 ( .A1(RF_MEMCTRL_data_reg[2]), .A2(n1508), .B(n897), 
        .ZN(MEMCTRL_MEM_to_mem_data[10]) );
  NR2D1BWP12T U1104 ( .A1(n1207), .A2(irdecode_inst1_N706), .ZN(n898) );
  ND2D1BWP12T U1105 ( .A1(n898), .A2(n1533), .ZN(n1544) );
  IOA21D0BWP12T U1106 ( .A1(
        Instruction_Fetch_inst1_fetched_instruction_reg_11_), .A2(n1361), .B(
        n1363), .ZN(n899) );
  AOI21D1BWP12T U1107 ( .A1(n1016), .A2(MEMCTRL_RF_IF_data_in[11]), .B(n899), 
        .ZN(n1696) );
  CKND0BWP12T U1108 ( .I(n1570), .ZN(n900) );
  AOI32D0BWP12T U1109 ( .A1(n1564), .A2(n1656), .A3(n1575), .B1(n900), .B2(
        n1656), .ZN(n1665) );
  CKND0BWP12T U1110 ( .I(n1509), .ZN(n901) );
  AOI222D0BWP12T U1111 ( .A1(n901), .A2(RF_MEMCTRL_data_reg[19]), .B1(n1506), 
        .B2(memory_interface_inst1_delay_data_in32[3]), .C1(n1507), .C2(
        memory_interface_inst1_delay_data_in32[19]), .ZN(n902) );
  IOA21D0BWP12T U1112 ( .A1(RF_MEMCTRL_data_reg[3]), .A2(n1508), .B(n902), 
        .ZN(MEMCTRL_MEM_to_mem_data[11]) );
  OAI21D0BWP12T U1113 ( .A1(n1378), .A2(n1377), .B(n1016), .ZN(n903) );
  AOI21D0BWP12T U1114 ( .A1(n1378), .A2(n1377), .B(n903), .ZN(
        IF_RF_incremented_pc_out[13]) );
  AN2D0BWP12T U1115 ( .A1(n1016), .A2(n1288), .Z(n1752) );
  IIND4D0BWP12T U1116 ( .A1(n1540), .A2(n1541), .B1(n1543), .B2(n1542), .ZN(
        n1562) );
  INR2D0BWP12T U1117 ( .A1(n1553), .B1(n1569), .ZN(n1575) );
  CKND0BWP12T U1118 ( .I(n1509), .ZN(n904) );
  AOI222D0BWP12T U1119 ( .A1(n904), .A2(RF_MEMCTRL_data_reg[20]), .B1(n1506), 
        .B2(memory_interface_inst1_delay_data_in32[4]), .C1(n1507), .C2(
        memory_interface_inst1_delay_data_in32[20]), .ZN(n905) );
  IOA21D0BWP12T U1120 ( .A1(RF_MEMCTRL_data_reg[4]), .A2(n1508), .B(n905), 
        .ZN(MEMCTRL_MEM_to_mem_data[12]) );
  AN2D0BWP12T U1121 ( .A1(n1016), .A2(n1374), .Z(n1755) );
  ND4D0BWP12T U1122 ( .A1(n1302), .A2(n1303), .A3(n1611), .A4(n1612), .ZN(n906) );
  NR3D0BWP12T U1123 ( .A1(n1693), .A2(n1304), .A3(n906), .ZN(n907) );
  CKND0BWP12T U1124 ( .I(n1687), .ZN(n908) );
  AOI22D0BWP12T U1125 ( .A1(n1687), .A2(RF_OUT_n), .B1(RF_OUT_v), .B2(n908), 
        .ZN(n909) );
  MOAI22D0BWP12T U1126 ( .A1(n1707), .A2(n909), .B1(n1707), .B2(n909), .ZN(
        n910) );
  CKND0BWP12T U1127 ( .I(n1696), .ZN(n911) );
  AOI22D0BWP12T U1128 ( .A1(n1687), .A2(n1291), .B1(n1292), .B2(n908), .ZN(
        n912) );
  MAOI22D0BWP12T U1129 ( .A1(n1707), .A2(n912), .B1(n1707), .B2(n912), .ZN(
        n913) );
  AOI22D0BWP12T U1130 ( .A1(n1294), .A2(n1521), .B1(n1678), .B2(n1293), .ZN(
        n914) );
  MOAI22D0BWP12T U1131 ( .A1(n1701), .A2(n913), .B1(n1701), .B2(n914), .ZN(
        n915) );
  AOI32D0BWP12T U1132 ( .A1(n1701), .A2(n1696), .A3(n910), .B1(n911), .B2(n915), .ZN(n916) );
  OAI22D0BWP12T U1133 ( .A1(RF_OUT_z), .A2(n1521), .B1(n1625), .B2(n1295), 
        .ZN(n917) );
  OAI22D0BWP12T U1134 ( .A1(RF_OUT_c), .A2(n1297), .B1(n1296), .B2(n1678), 
        .ZN(n918) );
  OAI21D0BWP12T U1135 ( .A1(n917), .A2(n918), .B(n1298), .ZN(n919) );
  IOA21D0BWP12T U1136 ( .A1(n916), .A2(n919), .B(n1299), .ZN(n920) );
  AOI31D0BWP12T U1137 ( .A1(n1300), .A2(n907), .A3(n920), .B(n1743), .ZN(
        irdecode_inst1_next_alu_write_to_reg_enable) );
  CKND0BWP12T U1138 ( .I(n1538), .ZN(n921) );
  AO211D0BWP12T U1139 ( .A1(n1742), .A2(DEC_RF_memory_write_to_reg[3]), .B(
        n1406), .C(n921), .Z(n1758) );
  NR2D1BWP12T U1140 ( .A1(n1207), .A2(irdecode_inst1_N707), .ZN(n922) );
  ND2D1BWP12T U1141 ( .A1(n922), .A2(n1099), .ZN(n1210) );
  IND2D0BWP12T U1142 ( .A1(n1221), .B1(n1312), .ZN(n1320) );
  INR3D0BWP12T U1143 ( .A1(n1510), .B1(n1514), .B2(n1449), .ZN(n1479) );
  AN2D0BWP12T U1144 ( .A1(n1016), .A2(n996), .Z(n1753) );
  IOA21D0BWP12T U1145 ( .A1(n1731), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[9]), .B(n1034), .ZN(
        n923) );
  AO21D0BWP12T U1146 ( .A1(MEM_MEMCTRL_from_mem_data[1]), .A2(n1033), .B(n923), 
        .Z(MEMCTRL_RF_IF_data_in[9]) );
  INR2D0BWP12T U1147 ( .A1(irdecode_inst1_N911), .B1(n1323), .ZN(n1637) );
  AN3D0BWP12T U1148 ( .A1(n1551), .A2(n1549), .A3(n1550), .Z(n1563) );
  ND3D0BWP12T U1149 ( .A1(n1545), .A2(n1546), .A3(n1568), .ZN(n1664) );
  CKND0BWP12T U1150 ( .I(n1509), .ZN(n924) );
  AOI222D0BWP12T U1151 ( .A1(n924), .A2(RF_MEMCTRL_data_reg[21]), .B1(n1506), 
        .B2(memory_interface_inst1_delay_data_in32[5]), .C1(n1507), .C2(
        memory_interface_inst1_delay_data_in32[21]), .ZN(n925) );
  IOA21D0BWP12T U1152 ( .A1(RF_MEMCTRL_data_reg[5]), .A2(n1508), .B(n925), 
        .ZN(MEMCTRL_MEM_to_mem_data[13]) );
  OAI21D0BWP12T U1153 ( .A1(n1402), .A2(n1401), .B(n1016), .ZN(n926) );
  AOI21D0BWP12T U1154 ( .A1(n1402), .A2(n1401), .B(n926), .ZN(
        IF_RF_incremented_pc_out[3]) );
  AN2D0BWP12T U1155 ( .A1(n1016), .A2(n1366), .Z(IF_RF_incremented_pc_out[15])
         );
  AOI222D0BWP12T U1156 ( .A1(n1577), .A2(n1652), .B1(
        DEC_RF_memory_write_to_reg[0]), .B2(n1742), .C1(n1576), .C2(n1537), 
        .ZN(n927) );
  ND4D0BWP12T U1157 ( .A1(n1538), .A2(n1539), .A3(n927), .A4(n1580), .ZN(n824)
         );
  AN2D0BWP12T U1158 ( .A1(n1006), .A2(n1413), .Z(n1143) );
  INR2D0BWP12T U1159 ( .A1(memory_interface_inst1_delay_addr_for_adder[6]), 
        .B1(n1478), .ZN(n1462) );
  AN2D0BWP12T U1160 ( .A1(n1016), .A2(n1261), .Z(n1746) );
  IOA21D1BWP12T U1161 ( .A1(n1731), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[13]), .B(n1034), .ZN(
        n928) );
  AO21D1BWP12T U1162 ( .A1(MEM_MEMCTRL_from_mem_data[5]), .A2(n1033), .B(n928), 
        .Z(MEMCTRL_RF_IF_data_in[13]) );
  IND3D0BWP12T U1163 ( .A1(n1219), .B1(n1218), .B2(n1531), .ZN(n929) );
  NR4D0BWP12T U1164 ( .A1(n1217), .A2(n1663), .A3(n1540), .A4(n929), .ZN(n930)
         );
  AOI31D0BWP12T U1165 ( .A1(n1649), .A2(n1545), .A3(n930), .B(n1648), .ZN(n931) );
  OAI31D0BWP12T U1166 ( .A1(n1231), .A2(n931), .A3(n1683), .B(n1738), .ZN(n932) );
  AOI21D0BWP12T U1167 ( .A1(n1241), .A2(n932), .B(n1743), .ZN(n1222) );
  INR2D1BWP12T U1168 ( .A1(irdecode_inst1_N540), .B1(n1069), .ZN(n1566) );
  CKND0BWP12T U1169 ( .I(n1509), .ZN(n933) );
  AOI222D0BWP12T U1170 ( .A1(n933), .A2(RF_MEMCTRL_data_reg[22]), .B1(n1506), 
        .B2(memory_interface_inst1_delay_data_in32[6]), .C1(n1507), .C2(
        memory_interface_inst1_delay_data_in32[22]), .ZN(n934) );
  IOA21D0BWP12T U1171 ( .A1(RF_MEMCTRL_data_reg[6]), .A2(n1508), .B(n934), 
        .ZN(MEMCTRL_MEM_to_mem_data[14]) );
  INR2D0BWP12T U1172 ( .A1(n1400), .B1(n1401), .ZN(n935) );
  OAI21D0BWP12T U1173 ( .A1(RF_pc_out[4]), .A2(n935), .B(n1016), .ZN(n936) );
  AOI21D0BWP12T U1174 ( .A1(RF_pc_out[4]), .A2(n935), .B(n936), .ZN(
        IF_RF_incremented_pc_out[4]) );
  AN2D0BWP12T U1175 ( .A1(n1016), .A2(n1359), .Z(n1756) );
  OAI211D0BWP12T U1176 ( .A1(n1690), .A2(n1603), .B(n1523), .C(n1312), .ZN(
        n937) );
  NR2D0BWP12T U1177 ( .A1(n1301), .A2(n937), .ZN(n938) );
  AOI31D0BWP12T U1178 ( .A1(n1283), .A2(n1300), .A3(n938), .B(n1668), .ZN(n939) );
  AO211D0BWP12T U1179 ( .A1(DEC_ALU_alu_opcode[2]), .A2(n1742), .B(n939), .C(
        n1671), .Z(n846) );
  CKND2D0BWP12T U1180 ( .A1(irdecode_inst1_step[2]), .A2(n1742), .ZN(n940) );
  OAI211D0BWP12T U1181 ( .A1(n1574), .A2(n1563), .B(n1656), .C(n940), .ZN(n941) );
  AO21D0BWP12T U1182 ( .A1(n1662), .A2(n1562), .B(n941), .Z(
        irdecode_inst1_next_step_2_) );
  CKND0BWP12T U1183 ( .I(RF_pc_out[31]), .ZN(n942) );
  OAI21D0BWP12T U1184 ( .A1(n1409), .A2(n942), .B(n1016), .ZN(n943) );
  AOI21D0BWP12T U1185 ( .A1(n1409), .A2(n942), .B(n943), .ZN(
        IF_RF_incremented_pc_out[31]) );
  ND3D1BWP12T U1186 ( .A1(n1550), .A2(irdecode_inst1_N543), .A3(n1076), .ZN(
        n1529) );
  IOA21D0BWP12T U1187 ( .A1(n1731), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[10]), .B(n1034), .ZN(
        n944) );
  AO21D0BWP12T U1188 ( .A1(MEM_MEMCTRL_from_mem_data[2]), .A2(n1033), .B(n944), 
        .Z(MEMCTRL_RF_IF_data_in[10]) );
  CKND2D0BWP12T U1189 ( .A1(memory_interface_inst1_fsm_state_2_), .A2(
        memory_interface_inst1_fsm_state_3_), .ZN(n945) );
  TPNR2D1BWP12T U1190 ( .A1(n1008), .A2(n945), .ZN(n1507) );
  INR2D1BWP12T U1191 ( .A1(n1151), .B1(n1323), .ZN(n1733) );
  CKND0BWP12T U1192 ( .I(MEMCTRL_IN_address[10]), .ZN(n946) );
  CKND2D0BWP12T U1193 ( .A1(memory_interface_inst1_delay_addr_for_adder[9]), 
        .A2(n1459), .ZN(n947) );
  OAI22D0BWP12T U1194 ( .A1(n1479), .A2(n946), .B1(
        memory_interface_inst1_delay_addr_for_adder[10]), .B2(n947), .ZN(n948)
         );
  AO21D0BWP12T U1195 ( .A1(memory_interface_inst1_delay_addr_for_adder[10]), 
        .A2(n1457), .B(n948), .Z(MEMCTRL_MEM_to_mem_address[10]) );
  CKND0BWP12T U1196 ( .I(n1629), .ZN(n949) );
  CKND0BWP12T U1197 ( .I(n1630), .ZN(n950) );
  AOI32D0BWP12T U1198 ( .A1(n1628), .A2(n1630), .A3(n949), .B1(n1631), .B2(
        n950), .ZN(MEMCTRL_MEM_to_mem_read_enable) );
  AN2D0BWP12T U1199 ( .A1(RF_pc_out[0]), .A2(n1016), .Z(
        IF_RF_incremented_pc_out[0]) );
  NR3D0BWP12T U1200 ( .A1(n1395), .A2(n1401), .A3(n1396), .ZN(n951) );
  OAI21D0BWP12T U1201 ( .A1(n951), .A2(RF_pc_out[6]), .B(n1016), .ZN(n952) );
  AOI21D0BWP12T U1202 ( .A1(n951), .A2(RF_pc_out[6]), .B(n952), .ZN(
        IF_RF_incremented_pc_out[6]) );
  AN2D0BWP12T U1203 ( .A1(n1016), .A2(n1330), .Z(n1757) );
  CKND0BWP12T U1204 ( .I(n1521), .ZN(n953) );
  OAI22D0BWP12T U1205 ( .A1(n1694), .A2(n1678), .B1(n1707), .B2(n1522), .ZN(
        n954) );
  OAI21D0BWP12T U1206 ( .A1(n953), .A2(n954), .B(n1264), .ZN(n955) );
  OAI211D0BWP12T U1207 ( .A1(n1523), .A2(n1721), .B(n1688), .C(n955), .ZN(n956) );
  IOA21D0BWP12T U1208 ( .A1(n1524), .A2(n956), .B(n1525), .ZN(
        irdecode_inst1_next_update_flag_c) );
  CKND0BWP12T U1209 ( .I(n1600), .ZN(n957) );
  AOI21D0BWP12T U1210 ( .A1(irdecode_inst1_step[4]), .A2(n957), .B(n1572), 
        .ZN(n958) );
  OAI211D0BWP12T U1211 ( .A1(n1575), .A2(n1574), .B(n1573), .C(n958), .ZN(
        irdecode_inst1_next_step_4_) );
  INR2D0BWP12T U1212 ( .A1(n1631), .B1(n1449), .ZN(n1417) );
  IND4D0BWP12T U1213 ( .A1(n1541), .B1(n1210), .B2(n1209), .B3(n1223), .ZN(
        n959) );
  NR2D0BWP12T U1214 ( .A1(n1253), .A2(n959), .ZN(n1649) );
  IND2XD2BWP12T U1215 ( .A1(irdecode_inst1_N906), .B1(irdecode_inst1_N912), 
        .ZN(n1151) );
  IND2D0BWP12T U1216 ( .A1(n1485), .B1(
        memory_interface_inst1_delay_addr_for_adder[5]), .ZN(n1478) );
  AN2D0BWP12T U1217 ( .A1(n1016), .A2(n1202), .Z(n1754) );
  IOA21D0BWP12T U1218 ( .A1(n1731), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[12]), .B(n1034), .ZN(
        n960) );
  AO21D0BWP12T U1219 ( .A1(MEM_MEMCTRL_from_mem_data[4]), .A2(n1033), .B(n960), 
        .Z(MEMCTRL_RF_IF_data_in[12]) );
  MAOI22D0BWP12T U1220 ( .A1(memory_interface_inst1_delay_addr_for_adder[9]), 
        .A2(n1460), .B1(memory_interface_inst1_delay_addr_for_adder[9]), .B2(
        n1459), .ZN(n961) );
  AO21D0BWP12T U1221 ( .A1(MEMCTRL_IN_address[9]), .A2(n1501), .B(n961), .Z(
        MEMCTRL_MEM_to_mem_address[9]) );
  OAI21D0BWP12T U1222 ( .A1(RF_pc_out[2]), .A2(RF_pc_out[1]), .B(n1016), .ZN(
        n962) );
  AOI21D0BWP12T U1223 ( .A1(RF_pc_out[2]), .A2(RF_pc_out[1]), .B(n962), .ZN(
        IF_RF_incremented_pc_out[2]) );
  OR2D0BWP12T U1224 ( .A1(n1395), .A2(n1401), .Z(n963) );
  OAI21D0BWP12T U1225 ( .A1(n1396), .A2(n963), .B(n1016), .ZN(n964) );
  AOI21D0BWP12T U1226 ( .A1(n1396), .A2(n963), .B(n964), .ZN(
        IF_RF_incremented_pc_out[5]) );
  OAI21D0BWP12T U1227 ( .A1(RF_pc_out[8]), .A2(n1394), .B(n1016), .ZN(n965) );
  AOI21D0BWP12T U1228 ( .A1(RF_pc_out[8]), .A2(n1394), .B(n965), .ZN(
        IF_RF_incremented_pc_out[8]) );
  OAI21D0BWP12T U1229 ( .A1(n1381), .A2(n1380), .B(n1016), .ZN(n966) );
  AOI21D0BWP12T U1230 ( .A1(n1381), .A2(n1380), .B(n966), .ZN(
        IF_RF_incremented_pc_out[11]) );
  AN2D0BWP12T U1231 ( .A1(n1016), .A2(n1142), .Z(n1750) );
  CKND0BWP12T U1232 ( .I(n1628), .ZN(n967) );
  OA21D0BWP12T U1233 ( .A1(n1511), .A2(DEC_MEMCTRL_load_store_width[1]), .B(
        n1628), .Z(n968) );
  AO211D0BWP12T U1234 ( .A1(DEC_MEMCTRL_load_store_width[0]), .A2(n967), .B(
        n1510), .C(n968), .Z(n969) );
  AOI21D0BWP12T U1235 ( .A1(n1512), .A2(n969), .B(reset), .ZN(
        memory_interface_inst1_fsm_N33) );
  CKND0BWP12T U1236 ( .I(n1522), .ZN(n970) );
  CKND2D0BWP12T U1237 ( .A1(IF_DEC_instruction[7]), .A2(n1722), .ZN(n971) );
  AOI211D0BWP12T U1238 ( .A1(n1522), .A2(n971), .B(n1690), .C(n1521), .ZN(n972) );
  AOI211D0BWP12T U1239 ( .A1(n1520), .A2(n970), .B(n1673), .C(n972), .ZN(n973)
         );
  CKND0BWP12T U1240 ( .I(n1524), .ZN(n974) );
  AOI32D0BWP12T U1241 ( .A1(n973), .A2(n1525), .A3(n1679), .B1(n974), .B2(
        n1525), .ZN(irdecode_inst1_next_update_flag_v) );
  CKND0BWP12T U1242 ( .I(n1664), .ZN(n975) );
  IND2D0BWP12T U1243 ( .A1(n1554), .B1(n1575), .ZN(n976) );
  AOI22D0BWP12T U1244 ( .A1(irdecode_inst1_step[5]), .A2(n1742), .B1(n1570), 
        .B2(n976), .ZN(n977) );
  OAI211D0BWP12T U1245 ( .A1(n1567), .A2(n975), .B(n1656), .C(n977), .ZN(
        irdecode_inst1_next_step_5_) );
  NR2D0BWP12T U1246 ( .A1(irdecode_inst1_N705), .A2(irdecode_inst1_N707), .ZN(
        n978) );
  CKND2D0BWP12T U1247 ( .A1(n978), .A2(n1694), .ZN(n1096) );
  ND3D0BWP12T U1248 ( .A1(n1082), .A2(irdecode_inst1_N543), .A3(n1551), .ZN(
        n1553) );
  IND2D0BWP12T U1249 ( .A1(memory_interface_inst1_fsm_state_0_), .B1(n1143), 
        .ZN(n1510) );
  MUX2ND0BWP12T U1250 ( .I0(RF_OUT_n), .I1(n1043), .S(RF_OUT_v), .ZN(n1292) );
  IND2D0BWP12T U1251 ( .A1(n1087), .B1(n1375), .ZN(n1600) );
  CKND0BWP12T U1252 ( .I(n1509), .ZN(n979) );
  AOI222D0BWP12T U1253 ( .A1(n979), .A2(RF_MEMCTRL_data_reg[23]), .B1(n1506), 
        .B2(memory_interface_inst1_delay_data_in32[7]), .C1(n1507), .C2(
        memory_interface_inst1_delay_data_in32[23]), .ZN(n980) );
  IOA21D0BWP12T U1254 ( .A1(RF_MEMCTRL_data_reg[7]), .A2(n1508), .B(n980), 
        .ZN(MEMCTRL_MEM_to_mem_data[15]) );
  OAI21D0BWP12T U1255 ( .A1(n1390), .A2(n1389), .B(n1016), .ZN(n981) );
  AOI21D0BWP12T U1256 ( .A1(n1390), .A2(n1389), .B(n981), .ZN(
        IF_RF_incremented_pc_out[9]) );
  OAI21D0BWP12T U1257 ( .A1(RF_pc_out[12]), .A2(n1379), .B(n1016), .ZN(n982)
         );
  AOI21D0BWP12T U1258 ( .A1(RF_pc_out[12]), .A2(n1379), .B(n982), .ZN(
        IF_RF_incremented_pc_out[12]) );
  OAI21D0BWP12T U1259 ( .A1(n1140), .A2(n1139), .B(n1016), .ZN(n983) );
  AOI21D0BWP12T U1260 ( .A1(n1140), .A2(n1139), .B(n983), .ZN(
        IF_RF_incremented_pc_out[21]) );
  INR2D0BWP12T U1261 ( .A1(n1016), .B1(RF_pc_out[1]), .ZN(
        MEMCTRL_IN_address[0]) );
  AO222D0BWP12T U1262 ( .A1(ALU_MISC_OUT_result[7]), .A2(n1498), .B1(n1016), 
        .B2(n1477), .C1(n1499), .C2(RF_MEMCTRL_address_reg[7]), .Z(
        MEMCTRL_IN_address[6]) );
  CKND0BWP12T U1263 ( .I(n1710), .ZN(n984) );
  OAI22D0BWP12T U1264 ( .A1(n1721), .A2(n984), .B1(n1111), .B2(n1688), .ZN(
        n985) );
  NR3D0BWP12T U1265 ( .A1(n1733), .A2(n1263), .A3(n985), .ZN(n986) );
  OAI32D0BWP12T U1266 ( .A1(n1743), .A2(n1679), .A3(n1687), .B1(n986), .B2(
        n1743), .ZN(n987) );
  AOI211D0BWP12T U1267 ( .A1(n1742), .A2(DEC_ALU_alu_opcode[1]), .B(n1259), 
        .C(n987), .ZN(n988) );
  CKND0BWP12T U1268 ( .I(n1609), .ZN(n989) );
  AOI32D0BWP12T U1269 ( .A1(n1680), .A2(n988), .A3(n1690), .B1(n989), .B2(n988), .ZN(n850) );
  CKND0BWP12T U1270 ( .I(n1538), .ZN(n990) );
  AO211D0BWP12T U1271 ( .A1(n1742), .A2(DEC_RF_memory_store_data_reg[3]), .B(
        n1407), .C(n990), .Z(n1759) );
  OAI32D0BWP12T U1272 ( .A1(n1665), .A2(n1664), .A3(n1663), .B1(n1662), .B2(
        n1665), .ZN(n991) );
  IOA21D0BWP12T U1273 ( .A1(irdecode_inst1_step[6]), .A2(n1742), .B(n991), 
        .ZN(irdecode_inst1_next_step_6_) );
  NR2D1BWP12T U1274 ( .A1(n1266), .A2(n1101), .ZN(n1248) );
  TPND2D1BWP12T U1275 ( .A1(n1542), .A2(n1103), .ZN(n1215) );
  TPOAI21D1BWP12T U1276 ( .A1(n1543), .A2(n1567), .B(n1535), .ZN(n1101) );
  TPND2D1BWP12T U1277 ( .A1(n1533), .A2(n1099), .ZN(n1543) );
  NR3D1BWP12T U1278 ( .A1(n1097), .A2(n1219), .A3(n1532), .ZN(n1542) );
  HICOND2BWP12T U1279 ( .A(RF_pc_out[18]), .CI(n1329), .CON(n1178), .S(n1330)
         );
  TPND2D2BWP12T U1280 ( .A1(RF_pc_out[2]), .A2(RF_pc_out[1]), .ZN(n1402) );
  TPND2D2BWP12T U1281 ( .A1(n1248), .A2(n1104), .ZN(n1230) );
  TPNR2D2BWP12T U1282 ( .A1(irdecode_inst1_N907), .A2(n1323), .ZN(n1183) );
  TPNR2D2BWP12T U1283 ( .A1(n1549), .A2(n1574), .ZN(n1266) );
  ND2D3BWP12T U1284 ( .A1(n1699), .A2(n1151), .ZN(n1681) );
  IND4D4BWP12T U1285 ( .A1(n1078), .B1(n1077), .B2(n1405), .B3(n1529), .ZN(
        n1639) );
  NR2D2BWP12T U1286 ( .A1(n1528), .A2(n1707), .ZN(n1078) );
  OAI211D2BWP12T U1287 ( .A1(n1668), .A2(n1681), .B(n1153), .C(n1152), .ZN(
        n1154) );
  BUFFD2BWP12T U1288 ( .I(RF_ALU_operand_a[23]), .Z(n1766) );
  BUFFD6BWP12T U1289 ( .I(RF_ALU_operand_b[3]), .Z(n1762) );
  INR2D2BWP12T U1290 ( .A1(Instruction_Fetch_inst1_currentState_1_), .B1(
        Instruction_Fetch_inst1_currentState_0_), .ZN(n1016) );
  BUFFD2BWP12T U1291 ( .I(RF_ALU_operand_a[29]), .Z(n1767) );
  INVD1BWP12T U1292 ( .I(n1668), .ZN(n1308) );
  ND2D1BWP12T U1293 ( .A1(n1087), .A2(n1057), .ZN(n1668) );
  BUFFXD3BWP12T U1294 ( .I(RF_ALU_operand_a[3]), .Z(n1763) );
  CKND1BWP12T U1295 ( .I(RF_pc_out[3]), .ZN(n1401) );
  INVD1BWP12T U1296 ( .I(n1402), .ZN(n1400) );
  CKND1BWP12T U1297 ( .I(RF_pc_out[5]), .ZN(n1396) );
  ND2XD0BWP12T U1298 ( .A1(RF_pc_out[6]), .A2(RF_pc_out[4]), .ZN(n992) );
  INR3XD1BWP12T U1299 ( .A1(n1400), .B1(n1396), .B2(n992), .ZN(n993) );
  ND2D1BWP12T U1300 ( .A1(RF_pc_out[3]), .A2(n993), .ZN(n1398) );
  INVD0BWP12T U1301 ( .I(RF_pc_out[7]), .ZN(n1397) );
  TPNR2D1BWP12T U1302 ( .A1(n1398), .A2(n1397), .ZN(n1394) );
  CKND2D1BWP12T U1303 ( .A1(n1394), .A2(RF_pc_out[8]), .ZN(n1390) );
  INVD1BWP12T U1304 ( .I(RF_pc_out[9]), .ZN(n1389) );
  TPNR2D1BWP12T U1305 ( .A1(n1390), .A2(n1389), .ZN(n1383) );
  CKND2D1BWP12T U1306 ( .A1(n1383), .A2(RF_pc_out[10]), .ZN(n1381) );
  INVD1BWP12T U1307 ( .I(RF_pc_out[11]), .ZN(n1380) );
  TPNR2D1BWP12T U1308 ( .A1(n1381), .A2(n1380), .ZN(n1379) );
  TPND2D1BWP12T U1309 ( .A1(n1379), .A2(RF_pc_out[12]), .ZN(n1378) );
  INVD1BWP12T U1310 ( .I(RF_pc_out[13]), .ZN(n1377) );
  NR2XD1BWP12T U1311 ( .A1(n1378), .A2(n1377), .ZN(n1373) );
  INVD1BWP12T U1312 ( .I(RF_pc_out[21]), .ZN(n1139) );
  NR2XD1BWP12T U1313 ( .A1(n1140), .A2(n1139), .ZN(n997) );
  AN2D0BWP12T U1314 ( .A1(n994), .A2(n1016), .Z(n1747) );
  NR4D0BWP12T U1315 ( .A1(RF_pc_out[4]), .A2(RF_pc_out[3]), .A3(RF_pc_out[2]), 
        .A4(RF_pc_out[1]), .ZN(n1339) );
  IND2D1BWP12T U1316 ( .A1(RF_pc_out[5]), .B1(n1339), .ZN(n1335) );
  MOAI22D0BWP12T U1317 ( .A1(RF_pc_out[6]), .A2(n1335), .B1(RF_pc_out[6]), 
        .B2(n1335), .ZN(n1346) );
  INR2D1BWP12T U1318 ( .A1(DEC_MISC_OUT_memory_address_source_is_reg), .B1(
        Instruction_Fetch_inst1_currentState_1_), .ZN(n1499) );
  NR2D1BWP12T U1319 ( .A1(DEC_MISC_OUT_memory_address_source_is_reg), .A2(
        Instruction_Fetch_inst1_currentState_1_), .ZN(n1498) );
  AO222D0BWP12T U1320 ( .A1(n1016), .A2(n1346), .B1(n1499), .B2(
        RF_MEMCTRL_address_reg[6]), .C1(n1498), .C2(ALU_MISC_OUT_result[6]), 
        .Z(MEMCTRL_IN_address[5]) );
  HICIND1BWP12T U1321 ( .A(RF_pc_out[25]), .CIN(n995), .CO(n1260), .S(n996) );
  HICOND1BWP12T U1322 ( .A(RF_pc_out[22]), .CI(n997), .CON(n1318), .S(n998) );
  AN2D0BWP12T U1323 ( .A1(n998), .A2(n1016), .Z(n1748) );
  INVD1BWP12T U1324 ( .I(memory_interface_inst1_fsm_state_1_), .ZN(n1006) );
  ND2D1BWP12T U1325 ( .A1(n1006), .A2(memory_interface_inst1_fsm_state_0_), 
        .ZN(n1008) );
  INVD0BWP12T U1326 ( .I(n1008), .ZN(n999) );
  INR2D1BWP12T U1327 ( .A1(memory_interface_inst1_fsm_state_3_), .B1(n999), 
        .ZN(n1004) );
  INR2D1BWP12T U1328 ( .A1(memory_interface_inst1_fsm_state_1_), .B1(
        memory_interface_inst1_fsm_state_2_), .ZN(n1011) );
  CKND0BWP12T U1329 ( .I(n1011), .ZN(n1001) );
  INR2D1BWP12T U1330 ( .A1(memory_interface_inst1_fsm_state_2_), .B1(
        memory_interface_inst1_fsm_state_1_), .ZN(n1007) );
  CKND0BWP12T U1331 ( .I(n1007), .ZN(n1000) );
  CKND2D1BWP12T U1332 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  MUX2NXD0BWP12T U1333 ( .I0(n1002), .I1(memory_interface_inst1_fsm_state_2_), 
        .S(memory_interface_inst1_fsm_state_0_), .ZN(n1003) );
  INR2D1BWP12T U1334 ( .A1(n1004), .B1(n1003), .ZN(n1449) );
  INVD1BWP12T U1335 ( .I(n1507), .ZN(n1416) );
  CKND2D1BWP12T U1336 ( .A1(n1011), .A2(memory_interface_inst1_fsm_state_0_), 
        .ZN(n1150) );
  ND2D1BWP12T U1337 ( .A1(n1416), .A2(n1150), .ZN(n1005) );
  NR2XD0BWP12T U1338 ( .A1(n1449), .A2(n1005), .ZN(n1411) );
  NR2D1BWP12T U1339 ( .A1(memory_interface_inst1_fsm_state_2_), .A2(
        memory_interface_inst1_fsm_state_3_), .ZN(n1413) );
  ND2D1BWP12T U1340 ( .A1(n1411), .A2(n1510), .ZN(n1145) );
  ND2D2BWP12T U1341 ( .A1(n1007), .A2(n1010), .ZN(n1728) );
  INVD0BWP12T U1342 ( .I(n1015), .ZN(n1009) );
  NR2D1BWP12T U1343 ( .A1(n1145), .A2(n1009), .ZN(n1014) );
  INVD3BWP12T U1344 ( .I(n1728), .ZN(n1731) );
  TPNR2D1BWP12T U1345 ( .A1(n1014), .A2(n1731), .ZN(n1033) );
  ND2D1BWP12T U1346 ( .A1(n1011), .A2(n1010), .ZN(n1144) );
  TPNR2D0BWP12T U1347 ( .A1(n1144), .A2(
        memory_interface_inst1_delayed_is_signed), .ZN(n1012) );
  NR2D1BWP12T U1348 ( .A1(n1012), .A2(MEM_MEMCTRL_from_mem_data[15]), .ZN(
        n1013) );
  CKND2D2BWP12T U1349 ( .A1(n1014), .A2(n1013), .ZN(n1034) );
  ND2D1BWP12T U1350 ( .A1(n1015), .A2(n1144), .ZN(n1514) );
  TPND2D2BWP12T U1351 ( .A1(n1514), .A2(n1016), .ZN(n754) );
  INR2D1BWP12T U1352 ( .A1(n754), .B1(reset), .ZN(n1180) );
  INVD1BWP12T U1353 ( .I(n1180), .ZN(n1388) );
  INVD1BWP12T U1354 ( .I(Instruction_Fetch_inst1_fetched_instruction_reg_5_), 
        .ZN(n1017) );
  INVD1BWP12T U1355 ( .I(reset), .ZN(n1375) );
  INR2D1BWP12T U1356 ( .A1(n1375), .B1(n754), .ZN(n1356) );
  CKND0BWP12T U1357 ( .I(n1356), .ZN(n1386) );
  MUX2D1BWP12T U1358 ( .I0(MEM_MEMCTRL_from_mem_data[13]), .I1(
        memory_interface_inst1_delay_first_two_bytes_out[5]), .S(n1731), .Z(
        MEMCTRL_RF_IF_data_in[5]) );
  INVD1BWP12T U1359 ( .I(MEMCTRL_RF_IF_data_in[5]), .ZN(n1018) );
  OAI22D0BWP12T U1360 ( .A1(n1388), .A2(n1017), .B1(n1386), .B2(n1018), .ZN(
        Instruction_Fetch_inst1_N88) );
  INVD1BWP12T U1361 ( .I(Instruction_Fetch_inst1_fetched_instruction_reg_4_), 
        .ZN(n1021) );
  MUX2D1BWP12T U1362 ( .I0(MEM_MEMCTRL_from_mem_data[12]), .I1(
        memory_interface_inst1_delay_first_two_bytes_out[4]), .S(n1731), .Z(
        MEMCTRL_RF_IF_data_in[4]) );
  INVD1BWP12T U1363 ( .I(MEMCTRL_RF_IF_data_in[4]), .ZN(n1022) );
  OAI22D0BWP12T U1364 ( .A1(n1388), .A2(n1021), .B1(n1386), .B2(n1022), .ZN(
        Instruction_Fetch_inst1_N87) );
  INVD1BWP12T U1365 ( .I(Instruction_Fetch_inst1_fetched_instruction_reg_1_), 
        .ZN(n1131) );
  MUX2D1BWP12T U1366 ( .I0(MEM_MEMCTRL_from_mem_data[9]), .I1(
        memory_interface_inst1_delay_first_two_bytes_out[1]), .S(n1731), .Z(
        MEMCTRL_RF_IF_data_in[1]) );
  INVD1BWP12T U1367 ( .I(MEMCTRL_RF_IF_data_in[1]), .ZN(n1133) );
  OAI22D0BWP12T U1368 ( .A1(n1388), .A2(n1131), .B1(n1386), .B2(n1133), .ZN(
        Instruction_Fetch_inst1_N84) );
  INVD1BWP12T U1369 ( .I(Instruction_Fetch_inst1_fetched_instruction_reg_2_), 
        .ZN(n1019) );
  MUX2D1BWP12T U1370 ( .I0(MEM_MEMCTRL_from_mem_data[10]), .I1(
        memory_interface_inst1_delay_first_two_bytes_out[2]), .S(n1731), .Z(
        MEMCTRL_RF_IF_data_in[2]) );
  INVD1BWP12T U1371 ( .I(MEMCTRL_RF_IF_data_in[2]), .ZN(n1020) );
  OAI22D0BWP12T U1372 ( .A1(n1388), .A2(n1019), .B1(n1386), .B2(n1020), .ZN(
        Instruction_Fetch_inst1_N85) );
  MUX2D1BWP12T U1373 ( .I0(MEM_MEMCTRL_from_mem_data[8]), .I1(
        memory_interface_inst1_delay_first_two_bytes_out[0]), .S(n1731), .Z(
        MEMCTRL_RF_IF_data_in[0]) );
  INVD1BWP12T U1374 ( .I(MEMCTRL_RF_IF_data_in[0]), .ZN(n1181) );
  INVD1BWP12T U1375 ( .I(Instruction_Fetch_inst1_fetched_instruction_reg_0_), 
        .ZN(n1182) );
  OAI22D1BWP12T U1376 ( .A1(n1181), .A2(n754), .B1(n1132), .B2(n1182), .ZN(
        IF_DEC_instruction[0]) );
  OAI22D1BWP12T U1377 ( .A1(n1018), .A2(n754), .B1(n1132), .B2(n1017), .ZN(
        IF_DEC_instruction[5]) );
  OAI22D1BWP12T U1378 ( .A1(n1020), .A2(n754), .B1(n1132), .B2(n1019), .ZN(
        IF_DEC_instruction[2]) );
  OAI22D1BWP12T U1379 ( .A1(n1022), .A2(n754), .B1(n1132), .B2(n1021), .ZN(
        IF_DEC_instruction[4]) );
  AOI211D0BWP12T U1380 ( .A1(DEC_MEMCTRL_load_store_width[0]), .A2(
        DEC_MEMCTRL_load_store_width[1]), .B(n1510), .C(reset), .ZN(n1391) );
  NR2D0BWP12T U1381 ( .A1(DEC_MEMCTRL_memory_load_request), .A2(
        Instruction_Fetch_inst1_currentState_1_), .ZN(n1628) );
  ND3XD0BWP12T U1382 ( .A1(n1391), .A2(DEC_MEMCTRL_memory_store_request), .A3(
        n1628), .ZN(n1392) );
  NR2D1BWP12T U1383 ( .A1(DEC_MEMCTRL_load_store_width[1]), .A2(
        DEC_MEMCTRL_load_store_width[0]), .ZN(n1629) );
  IAO21D0BWP12T U1384 ( .A1(n1150), .A2(memory_interface_inst1_fsm_state_3_), 
        .B(n1507), .ZN(n1023) );
  TPOAI22D0BWP12T U1385 ( .A1(n1392), .A2(n1629), .B1(reset), .B2(n1023), .ZN(
        memory_interface_inst1_fsm_N34) );
  INVD1BWP12T U1386 ( .I(n1132), .ZN(n1361) );
  ND2D2BWP12T U1387 ( .A1(n754), .A2(n1132), .ZN(n1363) );
  IOA21D1BWP12T U1388 ( .A1(n1361), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_13_), .B(n1363), .ZN(
        n1024) );
  AOI21D1BWP12T U1389 ( .A1(MEMCTRL_RF_IF_data_in[13]), .A2(n1016), .B(n1024), 
        .ZN(n1100) );
  INVD1BWP12T U1390 ( .I(n1100), .ZN(n1036) );
  INVD0BWP12T U1391 ( .I(n754), .ZN(n1025) );
  ND2D1BWP12T U1392 ( .A1(MEMCTRL_RF_IF_data_in[14]), .A2(n1025), .ZN(n1027)
         );
  ND2D1BWP12T U1393 ( .A1(n1361), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_14_), .ZN(n1026) );
  CKND2D1BWP12T U1394 ( .A1(n1027), .A2(n1026), .ZN(n1112) );
  CKND2D1BWP12T U1395 ( .A1(n1036), .A2(n1112), .ZN(n1109) );
  CKND2D1BWP12T U1396 ( .A1(n1033), .A2(MEM_MEMCTRL_from_mem_data[7]), .ZN(
        n1029) );
  CKND2D1BWP12T U1397 ( .A1(n1731), .A2(
        memory_interface_inst1_delay_first_two_bytes_out[15]), .ZN(n1028) );
  ND3D2BWP12T U1398 ( .A1(n1029), .A2(n1034), .A3(n1028), .ZN(
        MEMCTRL_RF_IF_data_in[15]) );
  IOA21D1BWP12T U1399 ( .A1(n1361), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_15_), .B(n1363), .ZN(
        n1030) );
  AOI21D1BWP12T U1400 ( .A1(MEMCTRL_RF_IF_data_in[15]), .A2(n1016), .B(n1030), 
        .ZN(n1085) );
  NR2D1BWP12T U1401 ( .A1(n1109), .A2(n1085), .ZN(n1119) );
  INVD1BWP12T U1402 ( .I(n1363), .ZN(n1031) );
  INVD1BWP12T U1403 ( .I(n1111), .ZN(n1523) );
  INR2D1BWP12T U1404 ( .A1(n1119), .B1(n1523), .ZN(n1699) );
  ND2D1BWP12T U1405 ( .A1(n1699), .A2(n1738), .ZN(n1323) );
  NR2D1BWP12T U1406 ( .A1(n1738), .A2(n1111), .ZN(n1162) );
  ND3D1BWP12T U1407 ( .A1(n1112), .A2(n1085), .A3(n1100), .ZN(n1110) );
  INR2D1BWP12T U1408 ( .A1(n1162), .B1(n1110), .ZN(n1557) );
  ND2D1BWP12T U1409 ( .A1(n1557), .A2(n1701), .ZN(n1677) );
  IOA21D1BWP12T U1410 ( .A1(n1361), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_8_), .B(n1363), .ZN(
        n1032) );
  TPAOI21D1BWP12T U1411 ( .A1(MEMCTRL_RF_IF_data_in[8]), .A2(n1016), .B(n1032), 
        .ZN(n1603) );
  INVD1BWP12T U1412 ( .I(n1603), .ZN(n1707) );
  IOA21D0BWP12T U1413 ( .A1(n1361), .A2(
        Instruction_Fetch_inst1_fetched_instruction_reg_9_), .B(n1363), .ZN(
        n1035) );
  AOI21D1BWP12T U1414 ( .A1(MEMCTRL_RF_IF_data_in[9]), .A2(n1016), .B(n1035), 
        .ZN(n1687) );
  ND2XD0BWP12T U1415 ( .A1(n1707), .A2(n1687), .ZN(n1521) );
  NR2D1BWP12T U1416 ( .A1(n1111), .A2(n1696), .ZN(n1686) );
  CKND0BWP12T U1417 ( .I(n1686), .ZN(n1037) );
  INVD1BWP12T U1418 ( .I(n1085), .ZN(n1108) );
  NR2D1BWP12T U1419 ( .A1(n1108), .A2(n1112), .ZN(n1107) );
  ND2D1BWP12T U1420 ( .A1(n1107), .A2(n1036), .ZN(n1721) );
  OAI22D1BWP12T U1421 ( .A1(n1677), .A2(n1521), .B1(n1037), .B2(n1721), .ZN(
        n1263) );
  INR2XD0BWP12T U1422 ( .A1(n1111), .B1(n1696), .ZN(n1710) );
  CKND2D0BWP12T U1423 ( .A1(n1710), .A2(n1107), .ZN(n1679) );
  CKND2D1BWP12T U1424 ( .A1(n1107), .A2(n1100), .ZN(n1688) );
  INVD0BWP12T U1425 ( .I(irdecode_inst1_itstate_6_), .ZN(n1517) );
  AOI22D0BWP12T U1426 ( .A1(irdecode_inst1_itstate_6_), .A2(RF_OUT_n), .B1(
        RF_OUT_z), .B2(n1517), .ZN(n1039) );
  INVD1BWP12T U1427 ( .I(RF_OUT_n), .ZN(n1043) );
  INVD1BWP12T U1428 ( .I(RF_OUT_z), .ZN(n1296) );
  ND2D1BWP12T U1429 ( .A1(n1292), .A2(n1296), .ZN(n1294) );
  INVD1BWP12T U1430 ( .I(n1294), .ZN(n1293) );
  INR2D1BWP12T U1431 ( .A1(RF_OUT_c), .B1(RF_OUT_z), .ZN(n1291) );
  OR2XD1BWP12T U1432 ( .A1(n1291), .A2(irdecode_inst1_itstate_6_), .Z(n1045)
         );
  INVD1BWP12T U1433 ( .I(irdecode_inst1_itstate_5_), .ZN(n1516) );
  OAI211D1BWP12T U1434 ( .A1(n1293), .A2(n1517), .B(n1045), .C(n1516), .ZN(
        n1038) );
  INVD1BWP12T U1435 ( .I(irdecode_inst1_itstate_7_), .ZN(n1325) );
  OAI32D1BWP12T U1436 ( .A1(irdecode_inst1_itstate_7_), .A2(
        irdecode_inst1_itstate_5_), .A3(n1039), .B1(n1038), .B2(n1325), .ZN(
        n1052) );
  NR2D1BWP12T U1437 ( .A1(irdecode_inst1_itstate_6_), .A2(
        irdecode_inst1_itstate_7_), .ZN(n1054) );
  AOI22D0BWP12T U1438 ( .A1(irdecode_inst1_itstate_6_), .A2(RF_OUT_v), .B1(
        RF_OUT_c), .B2(n1054), .ZN(n1041) );
  TPOAI21D0BWP12T U1439 ( .A1(irdecode_inst1_itstate_6_), .A2(n1292), .B(
        irdecode_inst1_itstate_7_), .ZN(n1040) );
  AOI21D1BWP12T U1440 ( .A1(n1041), .A2(n1040), .B(n1516), .ZN(n1049) );
  INVD0BWP12T U1441 ( .I(irdecode_inst1_itstate_4_), .ZN(n1042) );
  IND2XD1BWP12T U1442 ( .A1(n1049), .B1(n1042), .ZN(n1051) );
  TPND2D0BWP12T U1443 ( .A1(irdecode_inst1_itstate_6_), .A2(n1294), .ZN(n1046)
         );
  TPND2D0BWP12T U1444 ( .A1(irdecode_inst1_itstate_6_), .A2(n1043), .ZN(n1044)
         );
  AOI32D1BWP12T U1445 ( .A1(n1046), .A2(irdecode_inst1_itstate_7_), .A3(n1045), 
        .B1(n1044), .B2(n1325), .ZN(n1047) );
  RCAOI211D0BWP12T U1446 ( .A1(n1054), .A2(n1296), .B(
        irdecode_inst1_itstate_5_), .C(n1047), .ZN(n1048) );
  OAI21D1BWP12T U1447 ( .A1(n1049), .A2(n1048), .B(irdecode_inst1_itstate_4_), 
        .ZN(n1050) );
  OAI21D1BWP12T U1448 ( .A1(n1052), .A2(n1051), .B(n1050), .ZN(n1055) );
  NR2D1BWP12T U1449 ( .A1(irdecode_inst1_itstate_1_), .A2(
        irdecode_inst1_itstate_0_), .ZN(n1176) );
  NR4D0BWP12T U1450 ( .A1(irdecode_inst1_itstate_5_), .A2(
        irdecode_inst1_itstate_4_), .A3(irdecode_inst1_itstate_2_), .A4(
        irdecode_inst1_itstate_3_), .ZN(n1053) );
  ND3D1BWP12T U1451 ( .A1(n1054), .A2(n1176), .A3(n1053), .ZN(n1127) );
  ND2D1BWP12T U1452 ( .A1(n1055), .A2(n1127), .ZN(n1232) );
  INVD1BWP12T U1453 ( .I(DEC_MEMCTRL_memory_store_request), .ZN(n1511) );
  INVD1BWP12T U1454 ( .I(n1514), .ZN(n1410) );
  AN3XD1BWP12T U1455 ( .A1(DEC_IF_stall_to_instructionfetch), .A2(
        irdecode_inst1_split_instruction), .A3(n1375), .Z(n1056) );
  OR2XD1BWP12T U1456 ( .A1(n1356), .A2(n1056), .Z(n1057) );
  INVD1BWP12T U1457 ( .I(irdecode_inst1_N543), .ZN(n1062) );
  INVD1BWP12T U1458 ( .I(irdecode_inst1_N545), .ZN(n1058) );
  INVD1BWP12T U1459 ( .I(irdecode_inst1_N546), .ZN(n1526) );
  ND2D1BWP12T U1460 ( .A1(n1058), .A2(n1526), .ZN(n1072) );
  TPNR2D1BWP12T U1461 ( .A1(n1072), .A2(irdecode_inst1_N544), .ZN(n1082) );
  ND2D2BWP12T U1462 ( .A1(n1062), .A2(n1082), .ZN(n1080) );
  TPNR2D1BWP12T U1463 ( .A1(n1080), .A2(irdecode_inst1_N542), .ZN(n1065) );
  ND2D1BWP12T U1464 ( .A1(n1065), .A2(irdecode_inst1_N541), .ZN(n1527) );
  INVD1BWP12T U1465 ( .I(irdecode_inst1_N542), .ZN(n1060) );
  NR2D1BWP12T U1466 ( .A1(n1080), .A2(n1060), .ZN(n1554) );
  NR2XD0BWP12T U1467 ( .A1(irdecode_inst1_N540), .A2(irdecode_inst1_N539), 
        .ZN(n1088) );
  CKND2D1BWP12T U1468 ( .A1(n1088), .A2(n1603), .ZN(n1071) );
  TPNR2D0BWP12T U1469 ( .A1(irdecode_inst1_N541), .A2(irdecode_inst1_N544), 
        .ZN(n1059) );
  CKND2D1BWP12T U1470 ( .A1(n1060), .A2(n1059), .ZN(n1061) );
  NR2D1BWP12T U1471 ( .A1(n1071), .A2(n1061), .ZN(n1076) );
  TPND3D0BWP12T U1472 ( .A1(n1076), .A2(irdecode_inst1_N545), .A3(n1062), .ZN(
        n1064) );
  MUX2D1BWP12T U1473 ( .I0(n1064), .I1(n1063), .S(irdecode_inst1_N546), .Z(
        n1068) );
  INVD1BWP12T U1474 ( .I(n1065), .ZN(n1069) );
  TPNR3D0BWP12T U1475 ( .A1(irdecode_inst1_N541), .A2(n1707), .A3(
        irdecode_inst1_N539), .ZN(n1066) );
  ND2D1BWP12T U1476 ( .A1(n1566), .A2(n1066), .ZN(n1641) );
  ND2D1BWP12T U1477 ( .A1(n1068), .A2(n1067), .ZN(n1079) );
  NR2D1BWP12T U1478 ( .A1(irdecode_inst1_N540), .A2(irdecode_inst1_N541), .ZN(
        n1070) );
  INR2D1BWP12T U1479 ( .A1(n1070), .B1(n1069), .ZN(n1075) );
  CKND2D1BWP12T U1480 ( .A1(n1075), .A2(irdecode_inst1_N539), .ZN(n1528) );
  INVD0BWP12T U1481 ( .I(n1071), .ZN(n1074) );
  INVD1BWP12T U1482 ( .I(n1072), .ZN(n1550) );
  ND2D1BWP12T U1483 ( .A1(n1550), .A2(irdecode_inst1_N544), .ZN(n1083) );
  NR4D0BWP12T U1484 ( .A1(irdecode_inst1_N542), .A2(irdecode_inst1_N543), .A3(
        irdecode_inst1_N541), .A4(n1083), .ZN(n1073) );
  ND2D1BWP12T U1485 ( .A1(n1074), .A2(n1073), .ZN(n1077) );
  TPNR2D1BWP12T U1486 ( .A1(n1079), .A2(n1639), .ZN(n1551) );
  INVD1BWP12T U1487 ( .I(n1080), .ZN(n1081) );
  ND2D1BWP12T U1488 ( .A1(n1551), .A2(n1081), .ZN(n1084) );
  INR2D1BWP12T U1489 ( .A1(n1564), .B1(n1084), .ZN(n1226) );
  NR3D1BWP12T U1490 ( .A1(n1112), .A2(n1100), .A3(n1085), .ZN(n1169) );
  CKND2D1BWP12T U1491 ( .A1(n1169), .A2(n1111), .ZN(n1117) );
  TPND2D0BWP12T U1492 ( .A1(n1701), .A2(n1687), .ZN(n1086) );
  NR2D1BWP12T U1493 ( .A1(n1117), .A2(n1086), .ZN(n1304) );
  INVD1BWP12T U1494 ( .I(n1304), .ZN(n1640) );
  NR3XD0BWP12T U1495 ( .A1(n1697), .A2(n1738), .A3(n1743), .ZN(n1259) );
  CKND2D1BWP12T U1496 ( .A1(n1687), .A2(n1603), .ZN(n1678) );
  INVD1BWP12T U1497 ( .I(n1701), .ZN(n1739) );
  CKND2D1BWP12T U1498 ( .A1(n1739), .A2(n1696), .ZN(n1236) );
  NR3D1BWP12T U1499 ( .A1(n1117), .A2(n1678), .A3(n1236), .ZN(n1693) );
  CKND0BWP12T U1500 ( .I(n1693), .ZN(n1680) );
  MUX2D1BWP12T U1501 ( .I0(MEM_MEMCTRL_from_mem_data[15]), .I1(
        memory_interface_inst1_delay_first_two_bytes_out[7]), .S(n1731), .Z(
        MEMCTRL_RF_IF_data_in[7]) );
  INVD1BWP12T U1502 ( .I(MEMCTRL_RF_IF_data_in[7]), .ZN(n1385) );
  INVD1BWP12T U1503 ( .I(Instruction_Fetch_inst1_fetched_instruction_reg_7_), 
        .ZN(n1387) );
  OAI22D1BWP12T U1504 ( .A1(n1385), .A2(n754), .B1(n1132), .B2(n1387), .ZN(
        IF_DEC_instruction[7]) );
  INVD1BWP12T U1505 ( .I(IF_DEC_instruction[7]), .ZN(n1694) );
  OR2XD1BWP12T U1506 ( .A1(n1743), .A2(n1694), .Z(n1602) );
  INVD0BWP12T U1507 ( .I(n1602), .ZN(n1609) );
  INVD3BWP12T U1508 ( .I(n1600), .ZN(n1742) );
  MUX2D1BWP12T U1509 ( .I0(MEM_MEMCTRL_from_mem_data[11]), .I1(
        memory_interface_inst1_delay_first_two_bytes_out[3]), .S(n1731), .Z(
        MEMCTRL_RF_IF_data_in[3]) );
  INVD1BWP12T U1510 ( .I(MEMCTRL_RF_IF_data_in[3]), .ZN(n1146) );
  INVD1BWP12T U1511 ( .I(Instruction_Fetch_inst1_fetched_instruction_reg_3_), 
        .ZN(n1147) );
  OAI22D1BWP12T U1512 ( .A1(n1146), .A2(n754), .B1(n1132), .B2(n1147), .ZN(
        IF_DEC_instruction[3]) );
  ND2D1BWP12T U1513 ( .A1(n1226), .A2(n1088), .ZN(n1549) );
  INVD1BWP12T U1514 ( .I(n1570), .ZN(n1574) );
  NR2D1BWP12T U1515 ( .A1(irdecode_inst1_N707), .A2(irdecode_inst1_N706), .ZN(
        n1214) );
  INVD1BWP12T U1516 ( .I(irdecode_inst1_N705), .ZN(n1207) );
  ND2D1BWP12T U1517 ( .A1(n1214), .A2(n1207), .ZN(n1204) );
  NR2XD0BWP12T U1518 ( .A1(irdecode_inst1_N704), .A2(n1204), .ZN(n1220) );
  INVD1BWP12T U1519 ( .I(irdecode_inst1_N703), .ZN(n1091) );
  ND2D1BWP12T U1520 ( .A1(n1220), .A2(n1091), .ZN(n1212) );
  CKND2D0BWP12T U1521 ( .A1(irdecode_inst1_N702), .A2(n1694), .ZN(n1089) );
  NR3XD0BWP12T U1522 ( .A1(n1212), .A2(irdecode_inst1_N701), .A3(n1089), .ZN(
        n1216) );
  NR2D0BWP12T U1523 ( .A1(irdecode_inst1_N702), .A2(IF_DEC_instruction[7]), 
        .ZN(n1090) );
  TPND2D0BWP12T U1524 ( .A1(n1220), .A2(n1090), .ZN(n1092) );
  NR3XD0BWP12T U1525 ( .A1(n1092), .A2(irdecode_inst1_N701), .A3(n1091), .ZN(
        n1217) );
  NR2D1BWP12T U1526 ( .A1(n1216), .A2(n1217), .ZN(n1224) );
  INVD1BWP12T U1527 ( .I(irdecode_inst1_N701), .ZN(n1094) );
  NR2D1BWP12T U1528 ( .A1(irdecode_inst1_N703), .A2(irdecode_inst1_N702), .ZN(
        n1093) );
  ND2D1BWP12T U1529 ( .A1(n1094), .A2(n1093), .ZN(n1095) );
  INVD1BWP12T U1530 ( .I(irdecode_inst1_N704), .ZN(n1205) );
  CKND2D1BWP12T U1531 ( .A1(n1224), .A2(n1210), .ZN(n1097) );
  INVD1BWP12T U1532 ( .I(n1095), .ZN(n1102) );
  ND2D1BWP12T U1533 ( .A1(n1209), .A2(n1218), .ZN(n1532) );
  INVD1BWP12T U1534 ( .I(irdecode_inst1_N702), .ZN(n1211) );
  ND2D1BWP12T U1535 ( .A1(n1211), .A2(irdecode_inst1_N701), .ZN(n1098) );
  NR2D1BWP12T U1536 ( .A1(n1212), .A2(n1098), .ZN(n1208) );
  CKND2D1BWP12T U1537 ( .A1(n1208), .A2(n1694), .ZN(n1103) );
  NR2D1BWP12T U1538 ( .A1(n1215), .A2(irdecode_inst1_N707), .ZN(n1533) );
  ND2D1BWP12T U1539 ( .A1(n1108), .A2(n1100), .ZN(n1114) );
  ND2D1BWP12T U1540 ( .A1(n1735), .A2(n1308), .ZN(n1567) );
  INR2D1BWP12T U1541 ( .A1(n1600), .B1(n1308), .ZN(n1671) );
  INVD1BWP12T U1542 ( .I(n1671), .ZN(n1535) );
  ND2D1BWP12T U1543 ( .A1(n1103), .A2(n1530), .ZN(n1541) );
  INVD1BWP12T U1544 ( .I(n1567), .ZN(n1662) );
  ND2D1BWP12T U1545 ( .A1(n1541), .A2(n1662), .ZN(n1104) );
  INVD1BWP12T U1546 ( .I(n1230), .ZN(n1125) );
  CKND2D1BWP12T U1547 ( .A1(n1169), .A2(n1523), .ZN(n1582) );
  INVD1BWP12T U1548 ( .I(n1582), .ZN(n1235) );
  NR2D1BWP12T U1549 ( .A1(n1693), .A2(n1235), .ZN(n1105) );
  INR2D1BWP12T U1550 ( .A1(n1686), .B1(n1110), .ZN(n1653) );
  NR3D1BWP12T U1551 ( .A1(n1114), .A2(n1523), .A3(n1112), .ZN(n1644) );
  NR2D1BWP12T U1552 ( .A1(n1653), .A2(n1644), .ZN(n1583) );
  ND2D1BWP12T U1553 ( .A1(n1105), .A2(n1583), .ZN(n1606) );
  ND2XD0BWP12T U1554 ( .A1(n1699), .A2(n1696), .ZN(n1128) );
  TPND2D0BWP12T U1555 ( .A1(n1699), .A2(irdecode_inst1_N911), .ZN(n1106) );
  TPND2D0BWP12T U1556 ( .A1(n1128), .A2(n1106), .ZN(n1121) );
  NR2D1BWP12T U1557 ( .A1(n1557), .A2(n1107), .ZN(n1282) );
  NR3D1BWP12T U1558 ( .A1(n1114), .A2(n1112), .A3(n1111), .ZN(n1740) );
  NR2D1BWP12T U1559 ( .A1(n1109), .A2(n1108), .ZN(n1708) );
  NR2D1BWP12T U1560 ( .A1(n1740), .A2(n1708), .ZN(n1312) );
  INR2D1BWP12T U1561 ( .A1(n1111), .B1(n1110), .ZN(n1221) );
  INR2XD0BWP12T U1562 ( .A1(n1282), .B1(n1320), .ZN(n1120) );
  ND2D1BWP12T U1563 ( .A1(n1119), .A2(n1162), .ZN(n1302) );
  ND2XD0BWP12T U1564 ( .A1(n1112), .A2(n1111), .ZN(n1113) );
  NR2D1BWP12T U1565 ( .A1(n1114), .A2(n1113), .ZN(n1299) );
  INR2D1BWP12T U1566 ( .A1(n1302), .B1(n1299), .ZN(n1234) );
  CKND2D0BWP12T U1567 ( .A1(n1696), .A2(n1603), .ZN(n1115) );
  TPAOI21D0BWP12T U1568 ( .A1(n1739), .A2(n1115), .B(n1711), .ZN(n1116) );
  TPNR2D0BWP12T U1569 ( .A1(n1117), .A2(n1116), .ZN(n1118) );
  AOI21D1BWP12T U1570 ( .A1(n1119), .A2(n1686), .B(n1118), .ZN(n1233) );
  ND4D1BWP12T U1571 ( .A1(n1120), .A2(n1234), .A3(n1233), .A4(n1232), .ZN(
        n1277) );
  TPOAI31D0BWP12T U1572 ( .A1(n1606), .A2(n1121), .A3(n1277), .B(n1308), .ZN(
        n1123) );
  INR2D1BWP12T U1573 ( .A1(n1123), .B1(n1122), .ZN(n1124) );
  TPND2D1BWP12T U1574 ( .A1(n1125), .A2(n1124), .ZN(n1155) );
  INR2XD0BWP12T U1575 ( .A1(irdecode_inst1_step[0]), .B1(n1600), .ZN(n1126) );
  NR2D2BWP12T U1576 ( .A1(n1155), .A2(n1126), .ZN(n1768) );
  MUX2D1BWP12T U1577 ( .I0(MEM_MEMCTRL_from_mem_data[14]), .I1(
        memory_interface_inst1_delay_first_two_bytes_out[6]), .S(n1731), .Z(
        MEMCTRL_RF_IF_data_in[6]) );
  INVD1BWP12T U1578 ( .I(MEMCTRL_RF_IF_data_in[6]), .ZN(n1148) );
  INVD1BWP12T U1579 ( .I(Instruction_Fetch_inst1_fetched_instruction_reg_6_), 
        .ZN(n1149) );
  OAI22D1BWP12T U1580 ( .A1(n1148), .A2(n754), .B1(n1132), .B2(n1149), .ZN(
        IF_DEC_instruction[6]) );
  CKND2D0BWP12T U1581 ( .A1(n1694), .A2(IF_DEC_instruction[6]), .ZN(n1522) );
  INVD1BWP12T U1582 ( .I(n1690), .ZN(n1264) );
  NR2D0BWP12T U1583 ( .A1(n1668), .A2(n1127), .ZN(n1524) );
  INVD1BWP12T U1584 ( .I(n1743), .ZN(n1682) );
  CKND2D0BWP12T U1585 ( .A1(n1711), .A2(n1603), .ZN(n1295) );
  NR2D1BWP12T U1586 ( .A1(n1690), .A2(n1295), .ZN(n1520) );
  AOI22D1BWP12T U1587 ( .A1(n1263), .A2(n1682), .B1(n1609), .B2(n1520), .ZN(
        n1525) );
  CKND0BWP12T U1588 ( .I(IF_DEC_instruction[0]), .ZN(n1634) );
  INVD1BWP12T U1589 ( .I(n1128), .ZN(n1674) );
  ND2D1BWP12T U1590 ( .A1(n1674), .A2(n1682), .ZN(n1404) );
  TPND2D0BWP12T U1591 ( .A1(n1742), .A2(DEC_RF_offset_b[12]), .ZN(n1129) );
  INVD1BWP12T U1592 ( .I(n1584), .ZN(n1587) );
  OAI211D0BWP12T U1593 ( .A1(n1634), .A2(n1404), .B(n1129), .C(n1587), .ZN(
        n797) );
  INVD0BWP12T U1594 ( .I(IF_DEC_instruction[2]), .ZN(n1716) );
  TPND2D0BWP12T U1595 ( .A1(n1742), .A2(DEC_RF_offset_b[14]), .ZN(n1130) );
  OAI211D0BWP12T U1596 ( .A1(n1716), .A2(n1404), .B(n1130), .C(n1587), .ZN(
        n795) );
  TPOAI22D1BWP12T U1597 ( .A1(n1133), .A2(n754), .B1(n1132), .B2(n1131), .ZN(
        IF_DEC_instruction[1]) );
  INVD1BWP12T U1598 ( .I(IF_DEC_instruction[1]), .ZN(n1608) );
  CKND2D0BWP12T U1599 ( .A1(n1742), .A2(DEC_RF_offset_b[13]), .ZN(n1134) );
  OAI211D0BWP12T U1600 ( .A1(n1608), .A2(n1404), .B(n1134), .C(n1587), .ZN(
        n796) );
  CKND0BWP12T U1601 ( .I(IF_DEC_instruction[3]), .ZN(n1704) );
  CKND2D0BWP12T U1602 ( .A1(n1742), .A2(DEC_RF_offset_b[15]), .ZN(n1135) );
  OAI211D0BWP12T U1603 ( .A1(n1704), .A2(n1404), .B(n1135), .C(n1587), .ZN(
        n794) );
  CKND0BWP12T U1604 ( .I(IF_DEC_instruction[4]), .ZN(n1719) );
  CKND2D0BWP12T U1605 ( .A1(n1742), .A2(DEC_RF_offset_b[16]), .ZN(n1136) );
  OAI211D0BWP12T U1606 ( .A1(n1719), .A2(n1404), .B(n1136), .C(n1587), .ZN(
        n793) );
  CKND0BWP12T U1607 ( .I(IF_DEC_instruction[5]), .ZN(n1555) );
  TPND2D0BWP12T U1608 ( .A1(n1742), .A2(DEC_RF_offset_b[17]), .ZN(n1137) );
  OAI211D0BWP12T U1609 ( .A1(n1555), .A2(n1404), .B(n1137), .C(n1587), .ZN(
        n792) );
  INVD1BWP12T U1610 ( .I(IF_DEC_instruction[6]), .ZN(n1722) );
  CKND2D0BWP12T U1611 ( .A1(n1742), .A2(DEC_RF_offset_b[18]), .ZN(n1138) );
  OAI211D0BWP12T U1612 ( .A1(n1722), .A2(n1404), .B(n1138), .C(n1587), .ZN(
        n791) );
  HICOND2BWP12T U1613 ( .A(RF_pc_out[20]), .CI(n1141), .CON(n1140), .S(n1142)
         );
  INVD1BWP12T U1614 ( .I(MEM_MEMCTRL_from_mem_data[0]), .ZN(n1442) );
  OAI21D1BWP12T U1615 ( .A1(n1442), .A2(n1728), .B(n1730), .ZN(
        MEMCTRL_RF_IF_data_in[24]) );
  OAI22D0BWP12T U1616 ( .A1(n1388), .A2(n1147), .B1(n1386), .B2(n1146), .ZN(
        Instruction_Fetch_inst1_N86) );
  OAI22D0BWP12T U1617 ( .A1(n1388), .A2(n1149), .B1(n1386), .B2(n1148), .ZN(
        Instruction_Fetch_inst1_N89) );
  INR2D0BWP12T U1618 ( .A1(memory_interface_inst1_fsm_state_3_), .B1(n1150), 
        .ZN(n1414) );
  NR2D0BWP12T U1619 ( .A1(n1414), .A2(n1507), .ZN(n1412) );
  OAI21D0BWP12T U1620 ( .A1(reset), .A2(n1412), .B(n1392), .ZN(
        memory_interface_inst1_fsm_N35) );
  ND2D1BWP12T U1621 ( .A1(n1570), .A2(irdecode_inst1_N546), .ZN(n1153) );
  AOI22D1BWP12T U1622 ( .A1(n1662), .A2(irdecode_inst1_N707), .B1(n1742), .B2(
        irdecode_inst1_step[1]), .ZN(n1152) );
  NR2D1BWP12T U1623 ( .A1(n1155), .A2(n1154), .ZN(irdecode_inst1_N907) );
  NR2D0BWP12T U1624 ( .A1(RF_pc_out[2]), .A2(RF_pc_out[1]), .ZN(n1156) );
  MAOI22D0BWP12T U1625 ( .A1(RF_pc_out[3]), .A2(n1156), .B1(RF_pc_out[3]), 
        .B2(n1156), .ZN(n1342) );
  AO222D1BWP12T U1626 ( .A1(n1016), .A2(n1342), .B1(n1499), .B2(
        RF_MEMCTRL_address_reg[3]), .C1(n1498), .C2(ALU_MISC_OUT_result[3]), 
        .Z(MEMCTRL_IN_address[2]) );
  AOI21D1BWP12T U1627 ( .A1(n1520), .A2(n1522), .B(n1263), .ZN(n1196) );
  INVD1BWP12T U1628 ( .I(n1688), .ZN(n1713) );
  INVD1BWP12T U1629 ( .I(n1611), .ZN(n1157) );
  NR2XD0BWP12T U1630 ( .A1(n1721), .A2(n1686), .ZN(n1301) );
  OAI21D1BWP12T U1631 ( .A1(n1157), .A2(n1301), .B(n1524), .ZN(n1158) );
  OAI21D1BWP12T U1632 ( .A1(n1196), .A2(n1743), .B(n1158), .ZN(
        irdecode_inst1_next_update_flag_n) );
  INVD0BWP12T U1633 ( .I(n1234), .ZN(n1322) );
  NR4D0BWP12T U1634 ( .A1(n1304), .A2(n1699), .A3(n1322), .A4(n1606), .ZN(
        n1311) );
  ND4D0BWP12T U1635 ( .A1(n1312), .A2(n1311), .A3(n1232), .A4(n1535), .ZN(
        n1160) );
  INVD1BWP12T U1636 ( .I(n1721), .ZN(n1709) );
  NR2XD0BWP12T U1637 ( .A1(n1709), .A2(n1735), .ZN(n1270) );
  CKND2D1BWP12T U1638 ( .A1(n1635), .A2(n1270), .ZN(n1314) );
  INVD1BWP12T U1639 ( .I(n1233), .ZN(n1194) );
  NR2D1BWP12T U1640 ( .A1(n1671), .A2(n1308), .ZN(n1548) );
  INVD1BWP12T U1641 ( .I(n1548), .ZN(n1159) );
  OAI31D1BWP12T U1642 ( .A1(n1160), .A2(n1314), .A3(n1194), .B(n1159), .ZN(
        n1559) );
  IOA21D0BWP12T U1643 ( .A1(n1742), .A2(DEC_RF_operand_b[4]), .B(n1559), .ZN(
        n840) );
  CKND0BWP12T U1644 ( .I(n1699), .ZN(n1303) );
  ND2XD0BWP12T U1645 ( .A1(n1303), .A2(n1234), .ZN(n1659) );
  OAI22D0BWP12T U1646 ( .A1(n1270), .A2(n1687), .B1(n1738), .B2(n1582), .ZN(
        n1161) );
  AOI211D0BWP12T U1647 ( .A1(n1557), .A2(IF_DEC_instruction[1]), .B(n1161), 
        .C(n1653), .ZN(n1164) );
  INVD1BWP12T U1648 ( .I(n1677), .ZN(n1276) );
  AOI22D0BWP12T U1649 ( .A1(n1276), .A2(n1711), .B1(n1162), .B2(n1709), .ZN(
        n1190) );
  NR2D1BWP12T U1650 ( .A1(n1713), .A2(n1221), .ZN(n1561) );
  CKND2D1BWP12T U1651 ( .A1(n1561), .A2(n1312), .ZN(n1272) );
  CKND2D0BWP12T U1652 ( .A1(n1272), .A2(IF_DEC_instruction[4]), .ZN(n1163) );
  IND4D0BWP12T U1653 ( .A1(n1659), .B1(n1164), .B2(n1190), .B3(n1163), .ZN(
        n1165) );
  AO22XD0BWP12T U1654 ( .A1(n1165), .A2(n1682), .B1(n1742), .B2(
        DEC_RF_operand_a[1]), .Z(n814) );
  CKND2D0BWP12T U1655 ( .A1(n1742), .A2(DEC_RF_offset_b[19]), .ZN(n1166) );
  OAI211D0BWP12T U1656 ( .A1(n1694), .A2(n1404), .B(n1166), .C(n1587), .ZN(
        n790) );
  TPND2D0BWP12T U1657 ( .A1(n1742), .A2(DEC_RF_offset_b[20]), .ZN(n1167) );
  OAI211D0BWP12T U1658 ( .A1(n1603), .A2(n1404), .B(n1167), .C(n1587), .ZN(
        n789) );
  CKND2D0BWP12T U1659 ( .A1(n1742), .A2(DEC_RF_offset_b[22]), .ZN(n1168) );
  OAI211D0BWP12T U1660 ( .A1(n1739), .A2(n1404), .B(n1168), .C(n1587), .ZN(
        n787) );
  ND2XD0BWP12T U1661 ( .A1(n1710), .A2(n1701), .ZN(n1171) );
  CKND0BWP12T U1662 ( .I(n1169), .ZN(n1170) );
  ND2D1BWP12T U1663 ( .A1(n1711), .A2(n1707), .ZN(n1297) );
  NR3D1BWP12T U1664 ( .A1(n1171), .A2(n1170), .A3(n1297), .ZN(n1175) );
  NR4D0BWP12T U1665 ( .A1(IF_DEC_instruction[3]), .A2(IF_DEC_instruction[2]), 
        .A3(IF_DEC_instruction[0]), .A4(IF_DEC_instruction[1]), .ZN(n1173) );
  NR2D0BWP12T U1666 ( .A1(n1173), .A2(n1668), .ZN(n1172) );
  ND2D1BWP12T U1667 ( .A1(n1175), .A2(n1172), .ZN(n1633) );
  INVD1BWP12T U1668 ( .I(n1633), .ZN(n1327) );
  TPND2D0BWP12T U1669 ( .A1(n1175), .A2(n1173), .ZN(n1174) );
  AOI21D1BWP12T U1670 ( .A1(n1174), .A2(n1308), .B(reset), .ZN(n1632) );
  INR2D0BWP12T U1671 ( .A1(irdecode_inst1_itstate_3_), .B1(
        irdecode_inst1_itstate_2_), .ZN(n1177) );
  AOI211XD0BWP12T U1672 ( .A1(n1177), .A2(n1176), .B(n1175), .C(n1668), .ZN(
        n1326) );
  AO222D0BWP12T U1673 ( .A1(IF_DEC_instruction[1]), .A2(n1327), .B1(n1632), 
        .B2(irdecode_inst1_itstate_1_), .C1(irdecode_inst1_itstate_0_), .C2(
        n1326), .Z(n859) );
  HICIND2BWP12T U1674 ( .A(RF_pc_out[19]), .CIN(n1178), .CO(n1141), .S(n1179)
         );
  CKAN2D0BWP12T U1675 ( .A1(n1179), .A2(n1016), .Z(
        IF_RF_incremented_pc_out[19]) );
  AO22XD0BWP12T U1676 ( .A1(MEMCTRL_RF_IF_data_in[14]), .A2(n1356), .B1(
        Instruction_Fetch_inst1_fetched_instruction_reg_14_), .B2(n1180), .Z(
        Instruction_Fetch_inst1_N97) );
  OAI22D0BWP12T U1677 ( .A1(n1388), .A2(n1182), .B1(n1386), .B2(n1181), .ZN(
        Instruction_Fetch_inst1_N83) );
  ND2D1BWP12T U1678 ( .A1(n1183), .A2(n1768), .ZN(n1186) );
  TPND2D1BWP12T U1679 ( .A1(n1186), .A2(n1234), .ZN(n1726) );
  AOI22D0BWP12T U1680 ( .A1(n1726), .A2(IF_DEC_instruction[6]), .B1(n1606), 
        .B2(IF_DEC_instruction[5]), .ZN(n1185) );
  CKND0BWP12T U1681 ( .I(DEC_RF_offset_b[7]), .ZN(n1184) );
  OAI222D0BWP12T U1682 ( .A1(n1602), .A2(n1721), .B1(n1743), .B2(n1185), .C1(
        n1600), .C2(n1184), .ZN(n802) );
  AO21D1BWP12T U1683 ( .A1(n1186), .A2(n1302), .B(n1743), .Z(n1589) );
  CKND2D1BWP12T U1684 ( .A1(n1742), .A2(DEC_RF_offset_b[10]), .ZN(n1187) );
  OAI211D1BWP12T U1685 ( .A1(n1687), .A2(n1589), .B(n1187), .C(n1587), .ZN(
        n799) );
  INVD1BWP12T U1686 ( .I(irdecode_inst1_N907), .ZN(irdecode_inst1_next_step_1_) );
  AOI211D0BWP12T U1687 ( .A1(n1557), .A2(IF_DEC_instruction[0]), .B(n1322), 
        .C(n1674), .ZN(n1188) );
  OAI211D0BWP12T U1688 ( .A1(n1603), .A2(n1270), .B(n1188), .C(n1681), .ZN(
        n1189) );
  AOI211XD0BWP12T U1689 ( .A1(IF_DEC_instruction[3]), .A2(n1272), .B(n1189), 
        .C(n1606), .ZN(n1192) );
  ND3XD0BWP12T U1690 ( .A1(n1190), .A2(n1233), .A3(n1232), .ZN(n1268) );
  CKND0BWP12T U1691 ( .I(n1268), .ZN(n1191) );
  AOI21D0BWP12T U1692 ( .A1(n1192), .A2(n1191), .B(n1668), .ZN(n1193) );
  CKND2D1BWP12T U1693 ( .A1(n1574), .A2(n1535), .ZN(n1616) );
  AO211D1BWP12T U1694 ( .A1(n1742), .A2(DEC_RF_operand_a[0]), .B(n1193), .C(
        n1616), .Z(n811) );
  CKND0BWP12T U1695 ( .I(DEC_RF_alu_write_to_reg[4]), .ZN(n1198) );
  TPNR2D0BWP12T U1696 ( .A1(n1194), .A2(n1320), .ZN(n1195) );
  ND4D0BWP12T U1697 ( .A1(n1196), .A2(n1583), .A3(n1195), .A4(n1232), .ZN(
        n1285) );
  OAI21D0BWP12T U1698 ( .A1(n1285), .A2(n1733), .B(n1308), .ZN(n1197) );
  OAI211D0BWP12T U1699 ( .A1(n1600), .A2(n1198), .B(n1197), .C(n1535), .ZN(
        n815) );
  HICOND1BWP12T U1700 ( .A(RF_pc_out[28]), .CI(n1199), .CON(n1201), .S(n994)
         );
  AN2D0BWP12T U1701 ( .A1(n1200), .A2(n1016), .Z(n1745) );
  HICIND2BWP12T U1702 ( .A(RF_pc_out[29]), .CIN(n1201), .CO(n1408), .S(n1202)
         );
  NR3D0BWP12T U1703 ( .A1(RF_pc_out[3]), .A2(RF_pc_out[2]), .A3(RF_pc_out[1]), 
        .ZN(n1203) );
  MAOI22D0BWP12T U1704 ( .A1(RF_pc_out[4]), .A2(n1203), .B1(RF_pc_out[4]), 
        .B2(n1203), .ZN(n1341) );
  AO222D1BWP12T U1705 ( .A1(n1016), .A2(n1341), .B1(n1499), .B2(
        RF_MEMCTRL_address_reg[4]), .C1(n1498), .C2(ALU_MISC_OUT_result[4]), 
        .Z(MEMCTRL_IN_address[3]) );
  ND2D1BWP12T U1706 ( .A1(n1221), .A2(n1711), .ZN(n1737) );
  INR2D1BWP12T U1707 ( .A1(n1236), .B1(n1737), .ZN(n1652) );
  NR2D1BWP12T U1708 ( .A1(n1653), .A2(n1652), .ZN(n1241) );
  NR2D0BWP12T U1709 ( .A1(n1205), .A2(n1204), .ZN(n1206) );
  CKND2D1BWP12T U1710 ( .A1(n1533), .A2(n1206), .ZN(n1546) );
  ND2D0BWP12T U1711 ( .A1(n1546), .A2(n1544), .ZN(n1253) );
  CKND2D0BWP12T U1712 ( .A1(n1533), .A2(n1208), .ZN(n1223) );
  NR2D0BWP12T U1713 ( .A1(n1212), .A2(n1211), .ZN(n1213) );
  TPND2D0BWP12T U1714 ( .A1(n1533), .A2(n1213), .ZN(n1534) );
  INVD1BWP12T U1715 ( .I(n1534), .ZN(n1663) );
  TPNR2D0BWP12T U1716 ( .A1(n1215), .A2(n1214), .ZN(n1540) );
  CKND0BWP12T U1717 ( .I(n1216), .ZN(n1531) );
  INVD0BWP12T U1718 ( .I(n1735), .ZN(n1648) );
  CKND2D0BWP12T U1719 ( .A1(n1221), .A2(n1687), .ZN(n1280) );
  CKND2D1BWP12T U1720 ( .A1(n1280), .A2(n1312), .ZN(n1645) );
  OR2XD1BWP12T U1721 ( .A1(n1645), .A2(n1644), .Z(n1231) );
  INVD0BWP12T U1722 ( .I(n1697), .ZN(n1683) );
  AO21D0BWP12T U1723 ( .A1(n1742), .A2(DEC_MEMCTRL_memory_load_request), .B(
        n1222), .Z(n861) );
  AO21D0BWP12T U1724 ( .A1(n1742), .A2(DEC_RF_memory_write_to_reg_enable), .B(
        n1222), .Z(n825) );
  AOI21D0BWP12T U1725 ( .A1(n1252), .A2(n1224), .B(n1567), .ZN(n1229) );
  ND4D0BWP12T U1726 ( .A1(n1564), .A2(n1641), .A3(n1528), .A4(n1405), .ZN(
        n1225) );
  TPNR2D0BWP12T U1727 ( .A1(n1226), .A2(n1225), .ZN(n1227) );
  CKND2D0BWP12T U1728 ( .A1(n1645), .A2(n1308), .ZN(n1536) );
  OAI22D0BWP12T U1729 ( .A1(n1227), .A2(n1574), .B1(n1716), .B2(n1536), .ZN(
        n1228) );
  TPNR3D0BWP12T U1730 ( .A1(n1230), .A2(n1229), .A3(n1228), .ZN(n1245) );
  CKND2D0BWP12T U1731 ( .A1(n1231), .A2(n1696), .ZN(n1256) );
  ND4D0BWP12T U1732 ( .A1(n1234), .A2(n1233), .A3(n1232), .A4(n1303), .ZN(
        n1275) );
  INR4D0BWP12T U1733 ( .A1(n1282), .B1(n1235), .B2(n1693), .B3(n1275), .ZN(
        n1240) );
  INVD0BWP12T U1734 ( .I(n1236), .ZN(n1298) );
  INR2D1BWP12T U1735 ( .A1(n1298), .B1(n1737), .ZN(n1650) );
  INVD1BWP12T U1736 ( .I(n1650), .ZN(n1255) );
  CKND0BWP12T U1737 ( .I(n1652), .ZN(n1237) );
  OAI22D0BWP12T U1738 ( .A1(n1237), .A2(n1716), .B1(n1739), .B2(n1583), .ZN(
        n1238) );
  AOI22D0BWP12T U1739 ( .A1(n1238), .A2(n1308), .B1(n1742), .B2(
        DEC_RF_memory_write_to_reg[2]), .ZN(n1239) );
  TPND3D0BWP12T U1740 ( .A1(n1245), .A2(n1539), .A3(n1239), .ZN(n822) );
  CKND2D1BWP12T U1741 ( .A1(n1241), .A2(n1240), .ZN(n1247) );
  CKND0BWP12T U1742 ( .I(n1644), .ZN(n1242) );
  OAI21D0BWP12T U1743 ( .A1(n1242), .A2(n1298), .B(n1696), .ZN(n1243) );
  AOI211D0BWP12T U1744 ( .A1(n1650), .A2(IF_DEC_instruction[2]), .B(n1247), 
        .C(n1243), .ZN(n1246) );
  CKND2D0BWP12T U1745 ( .A1(n1742), .A2(DEC_RF_memory_store_data_reg[2]), .ZN(
        n1244) );
  OAI211D0BWP12T U1746 ( .A1(n1668), .A2(n1246), .B(n1245), .C(n1244), .ZN(
        n828) );
  TPND2D0BWP12T U1747 ( .A1(n1248), .A2(n1539), .ZN(n1406) );
  AO21D0BWP12T U1748 ( .A1(n1742), .A2(DEC_RF_memory_write_to_reg[4]), .B(
        n1406), .Z(n820) );
  NR2D0BWP12T U1749 ( .A1(n1648), .A2(n1743), .ZN(n1328) );
  AO211D0BWP12T U1750 ( .A1(n1742), .A2(
        DEC_MISC_OUT_memory_address_source_is_reg), .B(n1259), .C(n1328), .Z(
        n836) );
  MAOI22D0BWP12T U1751 ( .A1(n1247), .A2(n1308), .B1(n1696), .B2(n1668), .ZN(
        n1581) );
  ND2XD0BWP12T U1752 ( .A1(n1581), .A2(n1248), .ZN(n1407) );
  AO21D0BWP12T U1753 ( .A1(n1742), .A2(DEC_RF_memory_store_data_reg[4]), .B(
        n1407), .Z(n826) );
  HICIND2BWP12T U1754 ( .A(RF_pc_out[27]), .CIN(n1249), .CO(n1199), .S(n1250)
         );
  AN2XD0BWP12T U1755 ( .A1(n1250), .A2(n1016), .Z(n1751) );
  NR2D0BWP12T U1756 ( .A1(n1542), .A2(n1738), .ZN(n1254) );
  INVD0BWP12T U1757 ( .I(n1540), .ZN(n1251) );
  IND3D1BWP12T U1758 ( .A1(n1253), .B1(n1252), .B2(n1251), .ZN(n1734) );
  OAI31D0BWP12T U1759 ( .A1(n1254), .A2(n1541), .A3(n1734), .B(n1735), .ZN(
        n1257) );
  AOI31D0BWP12T U1760 ( .A1(n1257), .A2(n1256), .A3(n1255), .B(n1743), .ZN(
        n1258) );
  AO211D0BWP12T U1761 ( .A1(n1742), .A2(DEC_MEMCTRL_memory_store_request), .B(
        n1259), .C(n1258), .Z(n852) );
  HICOND1BWP12T U1762 ( .A(RF_pc_out[26]), .CI(n1260), .CON(n1249), .S(n1261)
         );
  OAI21D0BWP12T U1763 ( .A1(n1268), .A2(n1637), .B(n1308), .ZN(n1262) );
  CKND2D1BWP12T U1764 ( .A1(n1262), .A2(n1535), .ZN(n1519) );
  AOI21D0BWP12T U1765 ( .A1(n1264), .A2(n1711), .B(n1263), .ZN(n1265) );
  MOAI22D0BWP12T U1766 ( .A1(n1265), .A2(n1668), .B1(n1742), .B2(
        DEC_ALU_alu_opcode[3]), .ZN(n1267) );
  OR3D1BWP12T U1767 ( .A1(n1519), .A2(n1267), .A3(n1266), .Z(n849) );
  IND2XD1BWP12T U1768 ( .A1(n1268), .B1(n1311), .ZN(n1307) );
  AOI21D0BWP12T U1769 ( .A1(n1557), .A2(IF_DEC_instruction[2]), .B(n1307), 
        .ZN(n1269) );
  OAI21D0BWP12T U1770 ( .A1(n1270), .A2(n1739), .B(n1269), .ZN(n1271) );
  AOI21D0BWP12T U1771 ( .A1(IF_DEC_instruction[5]), .A2(n1272), .B(n1271), 
        .ZN(n1274) );
  CKND2D0BWP12T U1772 ( .A1(n1742), .A2(DEC_RF_operand_a[2]), .ZN(n1273) );
  OAI211D0BWP12T U1773 ( .A1(n1668), .A2(n1274), .B(n1535), .C(n1273), .ZN(
        n813) );
  TPND2D0BWP12T U1774 ( .A1(n1276), .A2(n1521), .ZN(n1300) );
  AO21D1BWP12T U1775 ( .A1(n1640), .A2(n1547), .B(n1548), .Z(n1657) );
  AOI22D0BWP12T U1776 ( .A1(n1662), .A2(n1701), .B1(n1742), .B2(
        DEC_RF_memory_store_address_reg[2]), .ZN(n1278) );
  CKND2D1BWP12T U1777 ( .A1(n1657), .A2(n1278), .ZN(n833) );
  AOI22D0BWP12T U1778 ( .A1(n1662), .A2(n1707), .B1(n1742), .B2(
        DEC_RF_memory_store_address_reg[0]), .ZN(n1279) );
  CKND2D1BWP12T U1779 ( .A1(n1657), .A2(n1279), .ZN(n835) );
  MAOI22D0BWP12T U1780 ( .A1(n1523), .A2(n1708), .B1(n1280), .B2(n1701), .ZN(
        n1281) );
  AOI31D0BWP12T U1781 ( .A1(n1283), .A2(n1282), .A3(n1281), .B(n1668), .ZN(
        n1284) );
  AO211D0BWP12T U1782 ( .A1(n1742), .A2(DEC_MEMCTRL_load_store_width[1]), .B(
        n1284), .C(n1671), .Z(n837) );
  NR2XD0BWP12T U1783 ( .A1(n1677), .A2(n1297), .ZN(n1658) );
  NR3XD0BWP12T U1784 ( .A1(n1285), .A2(n1693), .A3(n1658), .ZN(n1614) );
  INR3XD0BWP12T U1785 ( .A1(n1614), .B1(n1304), .B2(n1659), .ZN(n1670) );
  NR2D0BWP12T U1786 ( .A1(n1677), .A2(n1668), .ZN(n1289) );
  AOI21D0BWP12T U1787 ( .A1(n1289), .A2(IF_DEC_instruction[7]), .B(n1671), 
        .ZN(n1310) );
  CKND2D0BWP12T U1788 ( .A1(n1742), .A2(DEC_RF_alu_write_to_reg[3]), .ZN(n1286) );
  OAI211D0BWP12T U1789 ( .A1(n1668), .A2(n1670), .B(n1310), .C(n1286), .ZN(
        n817) );
  HICOND1BWP12T U1790 ( .A(RF_pc_out[24]), .CI(n1287), .CON(n995), .S(n1288)
         );
  AOI22D0BWP12T U1791 ( .A1(n1289), .A2(IF_DEC_instruction[6]), .B1(n1742), 
        .B2(DEC_RF_operand_b[3]), .ZN(n1290) );
  TPND2D0BWP12T U1792 ( .A1(n1559), .A2(n1290), .ZN(n841) );
  INVD1BWP12T U1793 ( .I(RF_OUT_c), .ZN(n1625) );
  ND2XD0BWP12T U1794 ( .A1(n1648), .A2(n1582), .ZN(n1321) );
  NR2D1BWP12T U1795 ( .A1(n1301), .A2(n1321), .ZN(n1612) );
  CKND0BWP12T U1796 ( .I(n1557), .ZN(n1313) );
  OAI22D0BWP12T U1797 ( .A1(n1722), .A2(n1561), .B1(n1313), .B2(n1704), .ZN(
        n1305) );
  AOI22D0BWP12T U1798 ( .A1(n1305), .A2(n1308), .B1(n1742), .B2(
        DEC_RF_operand_b[0]), .ZN(n1306) );
  TPND2D0BWP12T U1799 ( .A1(n1559), .A2(n1306), .ZN(n844) );
  AOI22D1BWP12T U1800 ( .A1(n1742), .A2(DEC_RF_operand_a[3]), .B1(n1308), .B2(
        n1307), .ZN(n1309) );
  CKND2D1BWP12T U1801 ( .A1(n1310), .A2(n1309), .ZN(n812) );
  CKND0BWP12T U1802 ( .I(DEC_RF_operand_b[1]), .ZN(n1317) );
  OAI211D0BWP12T U1803 ( .A1(n1719), .A2(n1313), .B(n1312), .C(n1311), .ZN(
        n1315) );
  NR2XD0BWP12T U1804 ( .A1(n1315), .A2(n1314), .ZN(n1316) );
  OAI222D0BWP12T U1805 ( .A1(n1317), .A2(n1600), .B1(n1602), .B2(n1561), .C1(
        n1743), .C2(n1316), .ZN(n843) );
  HICIND1BWP12T U1806 ( .A(RF_pc_out[23]), .CIN(n1318), .CO(n1287), .S(n1319)
         );
  AN2XD0BWP12T U1807 ( .A1(n1319), .A2(n1016), .Z(n1749) );
  CKND0BWP12T U1808 ( .I(n1583), .ZN(n1537) );
  NR4D0BWP12T U1809 ( .A1(n1322), .A2(n1321), .A3(n1320), .A4(n1537), .ZN(
        n1676) );
  AN4D0BWP12T U1810 ( .A1(n1676), .A2(n1640), .A3(n1323), .A4(n1677), .Z(n1324) );
  CKND0BWP12T U1811 ( .I(DEC_IF_stall_to_instructionfetch), .ZN(n1360) );
  OAI22D0BWP12T U1812 ( .A1(n1324), .A2(n1743), .B1(n1360), .B2(n1600), .ZN(
        n845) );
  NR2D1BWP12T U1813 ( .A1(n1326), .A2(n1632), .ZN(n1518) );
  OAI22D0BWP12T U1814 ( .A1(n1518), .A2(n1325), .B1(n1694), .B2(n1633), .ZN(
        n853) );
  AO222D0BWP12T U1815 ( .A1(IF_DEC_instruction[2]), .A2(n1327), .B1(n1632), 
        .B2(irdecode_inst1_itstate_2_), .C1(irdecode_inst1_itstate_1_), .C2(
        n1326), .Z(n858) );
  AO222D0BWP12T U1816 ( .A1(IF_DEC_instruction[3]), .A2(n1327), .B1(n1632), 
        .B2(irdecode_inst1_itstate_3_), .C1(irdecode_inst1_itstate_2_), .C2(
        n1326), .Z(n857) );
  AO222D0BWP12T U1817 ( .A1(IF_DEC_instruction[4]), .A2(n1327), .B1(n1326), 
        .B2(irdecode_inst1_itstate_3_), .C1(irdecode_inst1_itstate_4_), .C2(
        n1632), .Z(n856) );
  AO22XD1BWP12T U1818 ( .A1(n1328), .A2(n1711), .B1(n1742), .B2(
        DEC_RF_memory_store_address_reg[1]), .Z(n834) );
  AO21D0BWP12T U1819 ( .A1(n1742), .A2(DEC_RF_offset_b[29]), .B(n1584), .Z(
        n780) );
  AO21D0BWP12T U1820 ( .A1(n1742), .A2(DEC_RF_offset_b[30]), .B(n1584), .Z(
        n779) );
  AO21D0BWP12T U1821 ( .A1(n1742), .A2(DEC_RF_offset_b[28]), .B(n1584), .Z(
        n781) );
  AO21D0BWP12T U1822 ( .A1(n1742), .A2(DEC_RF_offset_b[27]), .B(n1584), .Z(
        n782) );
  AO21D0BWP12T U1823 ( .A1(n1742), .A2(DEC_RF_offset_b[26]), .B(n1584), .Z(
        n783) );
  AO21D0BWP12T U1824 ( .A1(n1742), .A2(DEC_RF_offset_b[25]), .B(n1584), .Z(
        n784) );
  AO21D0BWP12T U1825 ( .A1(n1742), .A2(DEC_RF_offset_b[23]), .B(n1584), .Z(
        n786) );
  AO21D0BWP12T U1826 ( .A1(n1742), .A2(DEC_RF_offset_b[24]), .B(n1584), .Z(
        n785) );
  TPND2D0BWP12T U1827 ( .A1(n1742), .A2(
        DEC_MEMCTRL_memorycontroller_sign_extend), .ZN(n1331) );
  OAI31D0BWP12T U1828 ( .A1(n1696), .A2(n1743), .A3(n1737), .B(n1331), .ZN(
        n839) );
  AO21D0BWP12T U1829 ( .A1(n1742), .A2(DEC_RF_offset_b[31]), .B(n1584), .Z(
        n777) );
  HICIND2BWP12T U1830 ( .A(RF_pc_out[17]), .CIN(n1332), .CO(n1329), .S(n1333)
         );
  AN2XD0BWP12T U1831 ( .A1(n1333), .A2(n1016), .Z(IF_RF_incremented_pc_out[17]) );
  CKND0BWP12T U1832 ( .I(RF_pc_out[1]), .ZN(n1340) );
  MAOI22D0BWP12T U1833 ( .A1(RF_pc_out[2]), .A2(n1340), .B1(RF_pc_out[2]), 
        .B2(n1340), .ZN(n1500) );
  OR4D0BWP12T U1834 ( .A1(RF_pc_out[15]), .A2(RF_pc_out[18]), .A3(
        RF_pc_out[20]), .A4(RF_pc_out[19]), .Z(n1334) );
  NR4D0BWP12T U1835 ( .A1(n1500), .A2(RF_pc_out[17]), .A3(RF_pc_out[16]), .A4(
        n1334), .ZN(n1354) );
  NR4D0BWP12T U1836 ( .A1(RF_pc_out[14]), .A2(RF_pc_out[13]), .A3(
        RF_pc_out[27]), .A4(RF_pc_out[26]), .ZN(n1353) );
  NR4D0BWP12T U1837 ( .A1(RF_pc_out[25]), .A2(RF_pc_out[24]), .A3(
        RF_pc_out[23]), .A4(RF_pc_out[22]), .ZN(n1352) );
  NR2D1BWP12T U1838 ( .A1(RF_pc_out[6]), .A2(n1335), .ZN(n1343) );
  IND2D1BWP12T U1839 ( .A1(RF_pc_out[7]), .B1(n1343), .ZN(n1345) );
  NR2D1BWP12T U1840 ( .A1(RF_pc_out[8]), .A2(n1345), .ZN(n1344) );
  IND2D1BWP12T U1841 ( .A1(RF_pc_out[9]), .B1(n1344), .ZN(n1338) );
  NR2XD0BWP12T U1842 ( .A1(RF_pc_out[10]), .A2(n1338), .ZN(n1337) );
  IND2D1BWP12T U1843 ( .A1(RF_pc_out[11]), .B1(n1337), .ZN(n1336) );
  MOAI22D0BWP12T U1844 ( .A1(RF_pc_out[12]), .A2(n1336), .B1(RF_pc_out[12]), 
        .B2(n1336), .ZN(n1448) );
  MAOI22D0BWP12T U1845 ( .A1(RF_pc_out[11]), .A2(n1337), .B1(RF_pc_out[11]), 
        .B2(n1337), .ZN(n1456) );
  MOAI22D0BWP12T U1846 ( .A1(RF_pc_out[10]), .A2(n1338), .B1(RF_pc_out[10]), 
        .B2(n1338), .ZN(n1458) );
  NR4D0BWP12T U1847 ( .A1(n1448), .A2(n1456), .A3(n1458), .A4(RF_pc_out[28]), 
        .ZN(n1350) );
  NR4D0BWP12T U1848 ( .A1(RF_pc_out[31]), .A2(RF_pc_out[30]), .A3(
        RF_pc_out[21]), .A4(RF_pc_out[29]), .ZN(n1349) );
  MAOI22D0BWP12T U1849 ( .A1(RF_pc_out[5]), .A2(n1339), .B1(RF_pc_out[5]), 
        .B2(n1339), .ZN(n1488) );
  NR4D0BWP12T U1850 ( .A1(n1342), .A2(n1488), .A3(n1341), .A4(n1340), .ZN(
        n1348) );
  MAOI22D0BWP12T U1851 ( .A1(RF_pc_out[7]), .A2(n1343), .B1(RF_pc_out[7]), 
        .B2(n1343), .ZN(n1477) );
  MAOI22D0BWP12T U1852 ( .A1(RF_pc_out[9]), .A2(n1344), .B1(RF_pc_out[9]), 
        .B2(n1344), .ZN(n1461) );
  MOAI22D0BWP12T U1853 ( .A1(RF_pc_out[8]), .A2(n1345), .B1(RF_pc_out[8]), 
        .B2(n1345), .ZN(n1472) );
  NR4D0BWP12T U1854 ( .A1(n1477), .A2(n1461), .A3(n1346), .A4(n1472), .ZN(
        n1347) );
  AN4XD1BWP12T U1855 ( .A1(n1350), .A2(n1349), .A3(n1348), .A4(n1347), .Z(
        n1351) );
  AN4XD1BWP12T U1856 ( .A1(n1354), .A2(n1353), .A3(n1352), .A4(n1351), .Z(
        n1513) );
  ND3XD0BWP12T U1857 ( .A1(n1513), .A2(n1016), .A3(
        Instruction_Fetch_inst1_first_instruction_fetched), .ZN(n1364) );
  OAI21D0BWP12T U1858 ( .A1(Instruction_Fetch_inst1_currentState_1_), .A2(
        DEC_IF_stall_to_instructionfetch), .B(
        Instruction_Fetch_inst1_currentState_0_), .ZN(n1355) );
  TPND2D0BWP12T U1859 ( .A1(n1364), .A2(n1355), .ZN(n1357) );
  AO21D0BWP12T U1860 ( .A1(n1357), .A2(n1375), .B(n1356), .Z(
        Instruction_Fetch_inst1_N79) );
  HICOND1BWP12T U1861 ( .A(RF_pc_out[16]), .CI(n1358), .CON(n1332), .S(n1359)
         );
  CKND2D0BWP12T U1862 ( .A1(n1361), .A2(n1360), .ZN(n1362) );
  AOI31D0BWP12T U1863 ( .A1(n1364), .A2(n1363), .A3(n1362), .B(reset), .ZN(
        Instruction_Fetch_inst1_N80) );
  HICIND1BWP12T U1864 ( .A(RF_pc_out[15]), .CIN(n1365), .CO(n1358), .S(n1366)
         );
  MUX2ND0BWP12T U1865 ( .I0(MEMCTRL_RF_IF_data_in[8]), .I1(
        Instruction_Fetch_inst1_fetched_instruction_reg_8_), .S(n754), .ZN(
        n1367) );
  CKND2D1BWP12T U1866 ( .A1(n1367), .A2(n1375), .ZN(
        Instruction_Fetch_inst1_N91) );
  MUX2ND0BWP12T U1867 ( .I0(MEMCTRL_RF_IF_data_in[9]), .I1(
        Instruction_Fetch_inst1_fetched_instruction_reg_9_), .S(n754), .ZN(
        n1368) );
  CKND2D1BWP12T U1868 ( .A1(n1368), .A2(n1375), .ZN(
        Instruction_Fetch_inst1_N92) );
  MUX2ND0BWP12T U1869 ( .I0(MEMCTRL_RF_IF_data_in[11]), .I1(
        Instruction_Fetch_inst1_fetched_instruction_reg_11_), .S(n754), .ZN(
        n1369) );
  CKND2D1BWP12T U1870 ( .A1(n1369), .A2(n1375), .ZN(
        Instruction_Fetch_inst1_N94) );
  MUX2ND0BWP12T U1871 ( .I0(MEMCTRL_RF_IF_data_in[10]), .I1(
        Instruction_Fetch_inst1_fetched_instruction_reg_10_), .S(n754), .ZN(
        n1370) );
  CKND2D1BWP12T U1872 ( .A1(n1370), .A2(n1375), .ZN(
        Instruction_Fetch_inst1_N93) );
  MUX2ND0BWP12T U1873 ( .I0(MEMCTRL_RF_IF_data_in[13]), .I1(
        Instruction_Fetch_inst1_fetched_instruction_reg_13_), .S(n754), .ZN(
        n1371) );
  CKND2D1BWP12T U1874 ( .A1(n1371), .A2(n1375), .ZN(
        Instruction_Fetch_inst1_N96) );
  MUX2ND0BWP12T U1875 ( .I0(MEMCTRL_RF_IF_data_in[12]), .I1(
        Instruction_Fetch_inst1_fetched_instruction_reg_12_), .S(n754), .ZN(
        n1372) );
  CKND2D1BWP12T U1876 ( .A1(n1372), .A2(n1375), .ZN(
        Instruction_Fetch_inst1_N95) );
  HICOND1BWP12T U1877 ( .A(RF_pc_out[14]), .CI(n1373), .CON(n1365), .S(n1374)
         );
  MUX2ND0BWP12T U1878 ( .I0(MEMCTRL_RF_IF_data_in[15]), .I1(
        Instruction_Fetch_inst1_fetched_instruction_reg_15_), .S(n754), .ZN(
        n1376) );
  CKND2D1BWP12T U1879 ( .A1(n1376), .A2(n1375), .ZN(
        Instruction_Fetch_inst1_N98) );
  CKND0BWP12T U1880 ( .I(RF_pc_out[10]), .ZN(n1382) );
  XNR2XD0BWP12T U1881 ( .A1(n1383), .A2(n1382), .ZN(n1384) );
  AN2XD0BWP12T U1882 ( .A1(n1384), .A2(n1016), .Z(IF_RF_incremented_pc_out[10]) );
  BUFFD12BWP12T U1883 ( .I(RF_ALU_operand_b[0]), .Z(n1761) );
  OAI22D0BWP12T U1884 ( .A1(n1388), .A2(n1387), .B1(n1386), .B2(n1385), .ZN(
        Instruction_Fetch_inst1_N90) );
  CKND0BWP12T U1885 ( .I(n1391), .ZN(n1393) );
  OAI31D0BWP12T U1886 ( .A1(n1629), .A2(n1628), .A3(n1393), .B(n1392), .ZN(
        memory_interface_inst1_fsm_N32) );
  CKND2D0BWP12T U1887 ( .A1(n1400), .A2(RF_pc_out[4]), .ZN(n1395) );
  CKXOR2D0BWP12T U1888 ( .A1(n1398), .A2(n1397), .Z(n1399) );
  AN2XD0BWP12T U1889 ( .A1(n1399), .A2(n1016), .Z(IF_RF_incremented_pc_out[7])
         );
  BUFFXD4BWP12T U1890 ( .I(RF_ALU_operand_a[21]), .Z(n1765) );
  CKND2D0BWP12T U1891 ( .A1(n1742), .A2(DEC_RF_offset_b[21]), .ZN(n1403) );
  OAI211D0BWP12T U1892 ( .A1(n1687), .A2(n1404), .B(n1403), .C(n1587), .ZN(
        n788) );
  BUFFD6BWP12T U1893 ( .I(RF_ALU_operand_a[19]), .Z(n1764) );
  HICOND1BWP12T U1894 ( .A(RF_pc_out[30]), .CI(n1408), .CON(n1409), .S(n1200)
         );
  INVD1BWP12T U1895 ( .I(MEM_MEMCTRL_from_mem_data[2]), .ZN(n1434) );
  OAI21D1BWP12T U1896 ( .A1(n1434), .A2(n1728), .B(n1730), .ZN(
        MEMCTRL_RF_IF_data_in[26]) );
  IOA21D1BWP12T U1897 ( .A1(n1731), .A2(MEM_MEMCTRL_from_mem_data[14]), .B(
        n1730), .ZN(MEMCTRL_RF_IF_data_in[22]) );
  IOA21D1BWP12T U1898 ( .A1(n1731), .A2(MEM_MEMCTRL_from_mem_data[11]), .B(
        n1730), .ZN(MEMCTRL_RF_IF_data_in[19]) );
  IOA21D1BWP12T U1899 ( .A1(n1731), .A2(MEM_MEMCTRL_from_mem_data[8]), .B(
        n1730), .ZN(MEMCTRL_RF_IF_data_in[16]) );
  IOA21D1BWP12T U1900 ( .A1(n1731), .A2(MEM_MEMCTRL_from_mem_data[10]), .B(
        n1730), .ZN(MEMCTRL_RF_IF_data_in[18]) );
  INVD1BWP12T U1901 ( .I(MEM_MEMCTRL_from_mem_data[1]), .ZN(n1438) );
  OAI21D1BWP12T U1902 ( .A1(n1438), .A2(n1728), .B(n1730), .ZN(
        MEMCTRL_RF_IF_data_in[25]) );
  CKND2D0BWP12T U1903 ( .A1(n1411), .A2(n1410), .ZN(n1415) );
  OAI31D1BWP12T U1904 ( .A1(n1629), .A2(n1511), .A3(n1415), .B(n1412), .ZN(
        MEMCTRL_MEM_to_mem_write_enable) );
  NR2D0BWP12T U1905 ( .A1(n1731), .A2(n1413), .ZN(n1631) );
  INVD1BWP12T U1906 ( .I(n1415), .ZN(n1630) );
  ND2D1BWP12T U1907 ( .A1(n1417), .A2(n1630), .ZN(n1509) );
  INVD1BWP12T U1908 ( .I(n1414), .ZN(n1512) );
  ND2D1BWP12T U1909 ( .A1(n1512), .A2(n1418), .ZN(n1506) );
  NR2D1BWP12T U1910 ( .A1(n1417), .A2(n1415), .ZN(n1508) );
  INVD1BWP12T U1911 ( .I(RF_MEMCTRL_data_reg[15]), .ZN(n1421) );
  INVD1BWP12T U1912 ( .I(n1508), .ZN(n1446) );
  INVD1BWP12T U1913 ( .I(MEM_MEMCTRL_from_mem_data[7]), .ZN(n1619) );
  ND2D1BWP12T U1914 ( .A1(n1417), .A2(n1416), .ZN(n1486) );
  MAOI22D0BWP12T U1915 ( .A1(n1507), .A2(
        memory_interface_inst1_delay_data_in32[31]), .B1(n1619), .B2(n1486), 
        .ZN(n1420) );
  INVD1BWP12T U1916 ( .I(n1418), .ZN(n1443) );
  ND2D1BWP12T U1917 ( .A1(n1443), .A2(
        memory_interface_inst1_delay_data_in32[15]), .ZN(n1419) );
  OAI211D1BWP12T U1918 ( .A1(n1421), .A2(n1446), .B(n1420), .C(n1419), .ZN(
        MEMCTRL_MEM_to_mem_data[7]) );
  INVD1BWP12T U1919 ( .I(RF_MEMCTRL_data_reg[14]), .ZN(n1424) );
  INVD1BWP12T U1920 ( .I(MEM_MEMCTRL_from_mem_data[6]), .ZN(n1623) );
  MAOI22D0BWP12T U1921 ( .A1(n1507), .A2(
        memory_interface_inst1_delay_data_in32[30]), .B1(n1623), .B2(n1486), 
        .ZN(n1423) );
  ND2D1BWP12T U1922 ( .A1(n1443), .A2(
        memory_interface_inst1_delay_data_in32[14]), .ZN(n1422) );
  OAI211D1BWP12T U1923 ( .A1(n1424), .A2(n1446), .B(n1423), .C(n1422), .ZN(
        MEMCTRL_MEM_to_mem_data[6]) );
  INVD1BWP12T U1924 ( .I(RF_MEMCTRL_data_reg[13]), .ZN(n1427) );
  INVD1BWP12T U1925 ( .I(MEM_MEMCTRL_from_mem_data[5]), .ZN(n1620) );
  MAOI22D0BWP12T U1926 ( .A1(n1507), .A2(
        memory_interface_inst1_delay_data_in32[29]), .B1(n1620), .B2(n1486), 
        .ZN(n1426) );
  ND2D1BWP12T U1927 ( .A1(n1443), .A2(
        memory_interface_inst1_delay_data_in32[13]), .ZN(n1425) );
  OAI211D1BWP12T U1928 ( .A1(n1427), .A2(n1446), .B(n1426), .C(n1425), .ZN(
        MEMCTRL_MEM_to_mem_data[5]) );
  INVD1BWP12T U1929 ( .I(RF_MEMCTRL_data_reg[12]), .ZN(n1430) );
  INVD1BWP12T U1930 ( .I(MEM_MEMCTRL_from_mem_data[4]), .ZN(n1622) );
  MAOI22D0BWP12T U1931 ( .A1(n1507), .A2(
        memory_interface_inst1_delay_data_in32[28]), .B1(n1622), .B2(n1486), 
        .ZN(n1429) );
  ND2D1BWP12T U1932 ( .A1(n1443), .A2(
        memory_interface_inst1_delay_data_in32[12]), .ZN(n1428) );
  OAI211D1BWP12T U1933 ( .A1(n1430), .A2(n1446), .B(n1429), .C(n1428), .ZN(
        MEMCTRL_MEM_to_mem_data[4]) );
  INVD1BWP12T U1934 ( .I(RF_MEMCTRL_data_reg[11]), .ZN(n1433) );
  INVD1BWP12T U1935 ( .I(MEM_MEMCTRL_from_mem_data[3]), .ZN(n1729) );
  MAOI22D0BWP12T U1936 ( .A1(n1507), .A2(
        memory_interface_inst1_delay_data_in32[27]), .B1(n1729), .B2(n1486), 
        .ZN(n1432) );
  ND2D1BWP12T U1937 ( .A1(n1443), .A2(
        memory_interface_inst1_delay_data_in32[11]), .ZN(n1431) );
  OAI211D1BWP12T U1938 ( .A1(n1433), .A2(n1446), .B(n1432), .C(n1431), .ZN(
        MEMCTRL_MEM_to_mem_data[3]) );
  INVD1BWP12T U1939 ( .I(RF_MEMCTRL_data_reg[10]), .ZN(n1437) );
  MAOI22D0BWP12T U1940 ( .A1(n1507), .A2(
        memory_interface_inst1_delay_data_in32[26]), .B1(n1434), .B2(n1486), 
        .ZN(n1436) );
  ND2D1BWP12T U1941 ( .A1(n1443), .A2(
        memory_interface_inst1_delay_data_in32[10]), .ZN(n1435) );
  OAI211D1BWP12T U1942 ( .A1(n1437), .A2(n1446), .B(n1436), .C(n1435), .ZN(
        MEMCTRL_MEM_to_mem_data[2]) );
  INVD1BWP12T U1943 ( .I(RF_MEMCTRL_data_reg[9]), .ZN(n1441) );
  MAOI22D0BWP12T U1944 ( .A1(n1507), .A2(
        memory_interface_inst1_delay_data_in32[25]), .B1(n1438), .B2(n1486), 
        .ZN(n1440) );
  ND2D1BWP12T U1945 ( .A1(n1443), .A2(
        memory_interface_inst1_delay_data_in32[9]), .ZN(n1439) );
  OAI211D1BWP12T U1946 ( .A1(n1441), .A2(n1446), .B(n1440), .C(n1439), .ZN(
        MEMCTRL_MEM_to_mem_data[1]) );
  INVD1BWP12T U1947 ( .I(RF_MEMCTRL_data_reg[8]), .ZN(n1447) );
  MAOI22D0BWP12T U1948 ( .A1(n1507), .A2(
        memory_interface_inst1_delay_data_in32[24]), .B1(n1442), .B2(n1486), 
        .ZN(n1445) );
  ND2D1BWP12T U1949 ( .A1(n1443), .A2(
        memory_interface_inst1_delay_data_in32[8]), .ZN(n1444) );
  OAI211D1BWP12T U1950 ( .A1(n1447), .A2(n1446), .B(n1445), .C(n1444), .ZN(
        MEMCTRL_MEM_to_mem_data[0]) );
  AO222D1BWP12T U1951 ( .A1(n1016), .A2(n1448), .B1(n1498), .B2(
        ALU_MISC_OUT_result[12]), .C1(n1499), .C2(RF_MEMCTRL_address_reg[12]), 
        .Z(MEMCTRL_IN_address[11]) );
  INVD1BWP12T U1952 ( .I(MEMCTRL_IN_address[11]), .ZN(n1454) );
  ND2D1BWP12T U1953 ( .A1(n1486), .A2(n1479), .ZN(n1496) );
  ND3D1BWP12T U1954 ( .A1(memory_interface_inst1_delay_addr_for_adder[0]), 
        .A2(memory_interface_inst1_delay_addr_for_adder[1]), .A3(
        memory_interface_inst1_delay_addr_for_adder[2]), .ZN(n1495) );
  INVD1BWP12T U1955 ( .I(n1495), .ZN(n1487) );
  ND2D1BWP12T U1956 ( .A1(n1487), .A2(
        memory_interface_inst1_delay_addr_for_adder[3]), .ZN(n1491) );
  IND2D1BWP12T U1957 ( .A1(n1491), .B1(
        memory_interface_inst1_delay_addr_for_adder[4]), .ZN(n1485) );
  ND3D1BWP12T U1958 ( .A1(n1462), .A2(
        memory_interface_inst1_delay_addr_for_adder[7]), .A3(
        memory_interface_inst1_delay_addr_for_adder[8]), .ZN(n1450) );
  NR2D1BWP12T U1959 ( .A1(n1496), .A2(n1450), .ZN(n1459) );
  IND4D1BWP12T U1960 ( .A1(memory_interface_inst1_delay_addr_for_adder[11]), 
        .B1(memory_interface_inst1_delay_addr_for_adder[10]), .B2(n1459), .B3(
        memory_interface_inst1_delay_addr_for_adder[9]), .ZN(n1453) );
  NR2D1BWP12T U1961 ( .A1(memory_interface_inst1_delay_addr_for_adder[10]), 
        .A2(n1496), .ZN(n1451) );
  INVD1BWP12T U1962 ( .I(n1496), .ZN(n1497) );
  INVD1BWP12T U1963 ( .I(n1486), .ZN(n1467) );
  AOI21D1BWP12T U1964 ( .A1(n1497), .A2(n1450), .B(n1467), .ZN(n1460) );
  OAI21D1BWP12T U1965 ( .A1(memory_interface_inst1_delay_addr_for_adder[9]), 
        .A2(n1496), .B(n1460), .ZN(n1457) );
  OAI21D1BWP12T U1966 ( .A1(n1451), .A2(n1457), .B(
        memory_interface_inst1_delay_addr_for_adder[11]), .ZN(n1452) );
  OAI211D1BWP12T U1967 ( .A1(n1454), .A2(n1479), .B(n1453), .C(n1452), .ZN(
        MEMCTRL_MEM_to_mem_address[11]) );
  INVD1BWP12T U1968 ( .I(n1479), .ZN(n1501) );
  AOI22D1BWP12T U1969 ( .A1(memory_interface_inst1_delay_addr_for_adder[0]), 
        .A2(n1467), .B1(MEMCTRL_IN_address[0]), .B2(n1501), .ZN(n1455) );
  OAI21D1BWP12T U1970 ( .A1(memory_interface_inst1_delay_addr_for_adder[0]), 
        .A2(n1496), .B(n1455), .ZN(MEMCTRL_MEM_to_mem_address[0]) );
  AO222D1BWP12T U1971 ( .A1(n1016), .A2(n1456), .B1(n1499), .B2(
        RF_MEMCTRL_address_reg[11]), .C1(n1498), .C2(ALU_MISC_OUT_result[11]), 
        .Z(MEMCTRL_IN_address[10]) );
  AO222D1BWP12T U1972 ( .A1(n1016), .A2(n1458), .B1(n1499), .B2(
        RF_MEMCTRL_address_reg[10]), .C1(n1498), .C2(ALU_MISC_OUT_result[10]), 
        .Z(MEMCTRL_IN_address[9]) );
  AO222D1BWP12T U1973 ( .A1(n1016), .A2(n1461), .B1(n1499), .B2(
        RF_MEMCTRL_address_reg[9]), .C1(n1498), .C2(ALU_MISC_OUT_result[9]), 
        .Z(MEMCTRL_IN_address[8]) );
  INVD1BWP12T U1974 ( .I(MEMCTRL_IN_address[8]), .ZN(n1466) );
  IND4D1BWP12T U1975 ( .A1(memory_interface_inst1_delay_addr_for_adder[8]), 
        .B1(n1462), .B2(n1497), .B3(
        memory_interface_inst1_delay_addr_for_adder[7]), .ZN(n1465) );
  NR2D1BWP12T U1976 ( .A1(memory_interface_inst1_delay_addr_for_adder[7]), 
        .A2(n1501), .ZN(n1463) );
  INVD1BWP12T U1977 ( .I(n1462), .ZN(n1475) );
  OAI21D1BWP12T U1978 ( .A1(n1463), .A2(n1473), .B(
        memory_interface_inst1_delay_addr_for_adder[8]), .ZN(n1464) );
  OAI211D1BWP12T U1979 ( .A1(n1479), .A2(n1466), .B(n1465), .C(n1464), .ZN(
        MEMCTRL_MEM_to_mem_address[8]) );
  ND2D1BWP12T U1980 ( .A1(memory_interface_inst1_delay_addr_for_adder[0]), 
        .A2(memory_interface_inst1_delay_addr_for_adder[1]), .ZN(n1471) );
  INVD1BWP12T U1981 ( .I(memory_interface_inst1_delay_addr_for_adder[0]), .ZN(
        n1468) );
  AOI21D1BWP12T U1982 ( .A1(n1479), .A2(n1468), .B(n1467), .ZN(n1505) );
  OAI21D1BWP12T U1983 ( .A1(memory_interface_inst1_delay_addr_for_adder[1]), 
        .A2(n1501), .B(n1505), .ZN(n1469) );
  AOI22D1BWP12T U1984 ( .A1(memory_interface_inst1_delay_addr_for_adder[2]), 
        .A2(n1469), .B1(n1501), .B2(MEMCTRL_IN_address[2]), .ZN(n1470) );
  OAI31D1BWP12T U1985 ( .A1(memory_interface_inst1_delay_addr_for_adder[2]), 
        .A2(n1496), .A3(n1471), .B(n1470), .ZN(MEMCTRL_MEM_to_mem_address[2])
         );
  AO222D1BWP12T U1986 ( .A1(n1016), .A2(n1472), .B1(n1499), .B2(
        RF_MEMCTRL_address_reg[8]), .C1(n1498), .C2(ALU_MISC_OUT_result[8]), 
        .Z(MEMCTRL_IN_address[7]) );
  ND2D1BWP12T U1987 ( .A1(memory_interface_inst1_delay_addr_for_adder[7]), 
        .A2(n1473), .ZN(n1474) );
  OAI31D1BWP12T U1988 ( .A1(memory_interface_inst1_delay_addr_for_adder[7]), 
        .A2(n1475), .A3(n1496), .B(n1474), .ZN(n1476) );
  AO21D1BWP12T U1989 ( .A1(n1501), .A2(MEMCTRL_IN_address[7]), .B(n1476), .Z(
        MEMCTRL_MEM_to_mem_address[7]) );
  NR3D1BWP12T U1990 ( .A1(n1496), .A2(n1478), .A3(
        memory_interface_inst1_delay_addr_for_adder[6]), .ZN(n1482) );
  NR2D1BWP12T U1991 ( .A1(n1501), .A2(
        memory_interface_inst1_delay_addr_for_adder[5]), .ZN(n1480) );
  OA21D1BWP12T U1992 ( .A1(n1483), .A2(n1480), .B(
        memory_interface_inst1_delay_addr_for_adder[6]), .Z(n1481) );
  AO211D1BWP12T U1993 ( .A1(MEMCTRL_IN_address[6]), .A2(n1501), .B(n1482), .C(
        n1481), .Z(MEMCTRL_MEM_to_mem_address[6]) );
  AOI22D1BWP12T U1994 ( .A1(memory_interface_inst1_delay_addr_for_adder[5]), 
        .A2(n1483), .B1(n1501), .B2(MEMCTRL_IN_address[5]), .ZN(n1484) );
  OAI31D1BWP12T U1995 ( .A1(memory_interface_inst1_delay_addr_for_adder[5]), 
        .A2(n1496), .A3(n1485), .B(n1484), .ZN(MEMCTRL_MEM_to_mem_address[5])
         );
  OA21D1BWP12T U1996 ( .A1(n1487), .A2(n1501), .B(n1486), .Z(n1492) );
  OAI21D1BWP12T U1997 ( .A1(memory_interface_inst1_delay_addr_for_adder[3]), 
        .A2(n1501), .B(n1492), .ZN(n1489) );
  AO222D1BWP12T U1998 ( .A1(n1016), .A2(n1488), .B1(n1499), .B2(
        RF_MEMCTRL_address_reg[5]), .C1(n1498), .C2(ALU_MISC_OUT_result[5]), 
        .Z(MEMCTRL_IN_address[4]) );
  AOI22D1BWP12T U1999 ( .A1(memory_interface_inst1_delay_addr_for_adder[4]), 
        .A2(n1489), .B1(n1501), .B2(MEMCTRL_IN_address[4]), .ZN(n1490) );
  OAI31D1BWP12T U2000 ( .A1(memory_interface_inst1_delay_addr_for_adder[4]), 
        .A2(n1496), .A3(n1491), .B(n1490), .ZN(MEMCTRL_MEM_to_mem_address[4])
         );
  INVD1BWP12T U2001 ( .I(n1492), .ZN(n1493) );
  AOI22D1BWP12T U2002 ( .A1(memory_interface_inst1_delay_addr_for_adder[3]), 
        .A2(n1493), .B1(n1501), .B2(MEMCTRL_IN_address[3]), .ZN(n1494) );
  OAI31D1BWP12T U2003 ( .A1(memory_interface_inst1_delay_addr_for_adder[3]), 
        .A2(n1496), .A3(n1495), .B(n1494), .ZN(MEMCTRL_MEM_to_mem_address[3])
         );
  INVD1BWP12T U2004 ( .I(memory_interface_inst1_delay_addr_for_adder[1]), .ZN(
        n1504) );
  ND3D1BWP12T U2005 ( .A1(n1497), .A2(
        memory_interface_inst1_delay_addr_for_adder[0]), .A3(n1504), .ZN(n1503) );
  AO222D1BWP12T U2006 ( .A1(n1016), .A2(n1500), .B1(n1499), .B2(
        RF_MEMCTRL_address_reg[2]), .C1(n1498), .C2(ALU_MISC_OUT_result[2]), 
        .Z(MEMCTRL_IN_address[1]) );
  ND2D1BWP12T U2007 ( .A1(n1501), .A2(MEMCTRL_IN_address[1]), .ZN(n1502) );
  OAI211D1BWP12T U2008 ( .A1(n1505), .A2(n1504), .B(n1503), .C(n1502), .ZN(
        MEMCTRL_MEM_to_mem_address[1]) );
  AOI21D0BWP12T U2009 ( .A1(n1514), .A2(n1513), .B(
        Instruction_Fetch_inst1_first_instruction_fetched), .ZN(n1515) );
  NR2D1BWP12T U2010 ( .A1(n1515), .A2(reset), .ZN(n862) );
  OAI22D1BWP12T U2011 ( .A1(n1518), .A2(n1516), .B1(n1555), .B2(n1633), .ZN(
        n855) );
  OAI22D1BWP12T U2012 ( .A1(n1518), .A2(n1517), .B1(n1722), .B2(n1633), .ZN(
        n854) );
  AO21D1BWP12T U2013 ( .A1(n1742), .A2(DEC_RF_operand_a[4]), .B(n1519), .Z(
        n810) );
  NR3D0BWP12T U2014 ( .A1(n1721), .A2(n1523), .A3(n1738), .ZN(n1673) );
  NR2D0BWP12T U2015 ( .A1(n1546), .A2(n1567), .ZN(n1572) );
  NR2D0BWP12T U2016 ( .A1(n1668), .A2(n1634), .ZN(n1577) );
  NR2D0BWP12T U2017 ( .A1(n1603), .A2(n1668), .ZN(n1576) );
  OR2XD1BWP12T U2018 ( .A1(n1548), .A2(n1547), .Z(n1656) );
  ND2D1BWP12T U2019 ( .A1(n1563), .A2(n1552), .ZN(n1569) );
  CKND0BWP12T U2020 ( .I(n1576), .ZN(n1560) );
  NR2D0BWP12T U2021 ( .A1(n1668), .A2(n1555), .ZN(n1556) );
  AOI22D0BWP12T U2022 ( .A1(n1557), .A2(n1556), .B1(n1742), .B2(
        DEC_RF_operand_b[2]), .ZN(n1558) );
  OAI211D1BWP12T U2023 ( .A1(n1561), .A2(n1560), .B(n1559), .C(n1558), .ZN(
        n842) );
  IOA21D0BWP12T U2024 ( .A1(n1742), .A2(irdecode_inst1_step[7]), .B(n1567), 
        .ZN(n1565) );
  AO211D1BWP12T U2025 ( .A1(n1570), .A2(n1566), .B(n1665), .C(n1565), .Z(
        irdecode_inst1_next_step_7_) );
  OA21XD1BWP12T U2026 ( .A1(n1568), .A2(n1567), .B(n1656), .Z(n1573) );
  AOI22D0BWP12T U2027 ( .A1(n1742), .A2(irdecode_inst1_step[3]), .B1(n1570), 
        .B2(n1569), .ZN(n1571) );
  ND2D1BWP12T U2028 ( .A1(n1573), .A2(n1571), .ZN(irdecode_inst1_next_step_3_)
         );
  AOI22D0BWP12T U2029 ( .A1(n1644), .A2(n1576), .B1(n1742), .B2(
        DEC_RF_memory_store_data_reg[0]), .ZN(n1579) );
  TPND2D0BWP12T U2030 ( .A1(n1650), .A2(n1577), .ZN(n1578) );
  ND4D1BWP12T U2031 ( .A1(n1581), .A2(n1580), .A3(n1579), .A4(n1578), .ZN(n830) );
  AOI21D0BWP12T U2032 ( .A1(n1583), .A2(n1582), .B(n1602), .ZN(n1585) );
  AOI211D0BWP12T U2033 ( .A1(n1742), .A2(DEC_RF_offset_b[9]), .B(n1585), .C(
        n1584), .ZN(n1586) );
  OAI21D1BWP12T U2034 ( .A1(n1589), .A2(n1603), .B(n1586), .ZN(n800) );
  CKND2D1BWP12T U2035 ( .A1(n1742), .A2(DEC_RF_offset_b[11]), .ZN(n1588) );
  OAI211D1BWP12T U2036 ( .A1(n1739), .A2(n1589), .B(n1588), .C(n1587), .ZN(
        n798) );
  INVD1BWP12T U2037 ( .I(n1726), .ZN(n1615) );
  TPNR2D0BWP12T U2038 ( .A1(n1743), .A2(n1722), .ZN(n1590) );
  TPAOI22D0BWP12T U2039 ( .A1(n1606), .A2(n1590), .B1(n1742), .B2(
        DEC_RF_offset_b[8]), .ZN(n1591) );
  OAI21D1BWP12T U2040 ( .A1(n1615), .A2(n1602), .B(n1591), .ZN(n801) );
  AOI21D0BWP12T U2041 ( .A1(n1740), .A2(IF_DEC_instruction[6]), .B(n1735), 
        .ZN(n1592) );
  OAI211D0BWP12T U2042 ( .A1(n1608), .A2(n1721), .B(n1640), .C(n1592), .ZN(
        n1593) );
  AOI211D1BWP12T U2043 ( .A1(n1726), .A2(IF_DEC_instruction[0]), .B(n1733), 
        .C(n1593), .ZN(n1595) );
  CKND0BWP12T U2044 ( .I(DEC_RF_offset_b[1]), .ZN(n1594) );
  OAI222D1BWP12T U2045 ( .A1(n1635), .A2(n1602), .B1(n1743), .B2(n1595), .C1(
        n1600), .C2(n1594), .ZN(n808) );
  INVD1BWP12T U2046 ( .I(n1708), .ZN(n1723) );
  INVD1BWP12T U2047 ( .I(n1606), .ZN(n1720) );
  NR2D1BWP12T U2048 ( .A1(n1720), .A2(n1608), .ZN(n1598) );
  AOI22D0BWP12T U2049 ( .A1(n1709), .A2(IF_DEC_instruction[3]), .B1(n1740), 
        .B2(n1707), .ZN(n1596) );
  OAI31D0BWP12T U2050 ( .A1(n1687), .A2(n1710), .A3(n1688), .B(n1596), .ZN(
        n1597) );
  AOI211D1BWP12T U2051 ( .A1(n1726), .A2(IF_DEC_instruction[2]), .B(n1598), 
        .C(n1597), .ZN(n1601) );
  CKND0BWP12T U2052 ( .I(DEC_RF_offset_b[3]), .ZN(n1599) );
  OAI222D1BWP12T U2053 ( .A1(n1602), .A2(n1723), .B1(n1743), .B2(n1601), .C1(
        n1600), .C2(n1599), .ZN(n806) );
  NR2D0BWP12T U2054 ( .A1(n1635), .A2(n1603), .ZN(n1605) );
  OAI22D0BWP12T U2055 ( .A1(n1723), .A2(n1722), .B1(n1716), .B2(n1721), .ZN(
        n1604) );
  AOI211D0BWP12T U2056 ( .A1(n1606), .A2(IF_DEC_instruction[0]), .B(n1605), 
        .C(n1604), .ZN(n1607) );
  OAI21D1BWP12T U2057 ( .A1(n1615), .A2(n1608), .B(n1607), .ZN(n1610) );
  AO222D1BWP12T U2058 ( .A1(n1610), .A2(n1682), .B1(n1740), .B2(n1609), .C1(
        n1742), .C2(DEC_RF_offset_b[2]), .Z(n807) );
  MUX2D1BWP12T U2059 ( .I0(RF_OUT_n), .I1(ALU_OUT_n), .S(
        DEC_CPSR_update_flag_n), .Z(new_n) );
  MUX2D1BWP12T U2060 ( .I0(RF_OUT_c), .I1(ALU_OUT_c), .S(
        DEC_CPSR_update_flag_c), .Z(new_c) );
  TPOAI21D0BWP12T U2061 ( .A1(n1707), .A2(n1677), .B(n1611), .ZN(n1667) );
  INVD1BWP12T U2062 ( .I(n1612), .ZN(n1666) );
  AOI22D0BWP12T U2063 ( .A1(n1667), .A2(IF_DEC_instruction[0]), .B1(n1707), 
        .B2(n1666), .ZN(n1613) );
  TPAOI31D0BWP12T U2064 ( .A1(n1615), .A2(n1614), .A3(n1613), .B(n1668), .ZN(
        n1617) );
  AO211D1BWP12T U2065 ( .A1(n1742), .A2(DEC_RF_alu_write_to_reg[0]), .B(n1617), 
        .C(n1616), .Z(n816) );
  INVD1BWP12T U2066 ( .I(n1768), .ZN(irdecode_inst1_next_step_0_) );
  MUX2D1BWP12T U2067 ( .I0(RF_OUT_z), .I1(ALU_OUT_z), .S(
        DEC_CPSR_update_flag_z), .Z(new_z) );
  INR2D1BWP12T U2068 ( .A1(RF_OUT_v), .B1(DEC_CPSR_update_flag_v), .ZN(n1618)
         );
  AO21D1BWP12T U2069 ( .A1(ALU_OUT_v), .A2(DEC_CPSR_update_flag_v), .B(n1618), 
        .Z(new_v) );
  OAI21D1BWP12T U2070 ( .A1(n1619), .A2(n1728), .B(n1730), .ZN(
        MEMCTRL_RF_IF_data_in[31]) );
  OAI21D1BWP12T U2071 ( .A1(n1620), .A2(n1728), .B(n1730), .ZN(
        MEMCTRL_RF_IF_data_in[29]) );
  INVD1BWP12T U2072 ( .I(MEM_MEMCTRL_from_mem_data[15]), .ZN(n1621) );
  OAI21D1BWP12T U2073 ( .A1(n1728), .A2(n1621), .B(n1730), .ZN(
        MEMCTRL_RF_IF_data_in[23]) );
  OAI21D1BWP12T U2074 ( .A1(n1622), .A2(n1728), .B(n1730), .ZN(
        MEMCTRL_RF_IF_data_in[28]) );
  OAI21D1BWP12T U2075 ( .A1(n1623), .A2(n1728), .B(n1730), .ZN(
        MEMCTRL_RF_IF_data_in[30]) );
  IND3D0BWP12T U2076 ( .A1(DEC_ALU_alu_opcode[3]), .B1(DEC_ALU_alu_opcode[1]), 
        .B2(DEC_ALU_alu_opcode[4]), .ZN(n1627) );
  CKND0BWP12T U2077 ( .I(DEC_ALU_alu_opcode[0]), .ZN(n1624) );
  CKND2D0BWP12T U2078 ( .A1(n1624), .A2(DEC_ALU_alu_opcode[2]), .ZN(n1626) );
  OAI22D1BWP12T U2079 ( .A1(n1627), .A2(n1626), .B1(DEC_ALU_alu_opcode[4]), 
        .B2(n1625), .ZN(ALU_IN_c) );
  MOAI22D0BWP12T U2080 ( .A1(n1634), .A2(n1633), .B1(n1632), .B2(
        irdecode_inst1_itstate_0_), .ZN(n860) );
  OAI22D0BWP12T U2081 ( .A1(n1635), .A2(n1722), .B1(n1634), .B2(n1721), .ZN(
        n1636) );
  TPNR2D0BWP12T U2082 ( .A1(n1637), .A2(n1636), .ZN(n1638) );
  MOAI22D0BWP12T U2083 ( .A1(n1638), .A2(n1743), .B1(n1742), .B2(
        DEC_RF_offset_b[0]), .ZN(n809) );
  CKND0BWP12T U2084 ( .I(n1639), .ZN(n1642) );
  AO31D0BWP12T U2085 ( .A1(n1643), .A2(n1642), .A3(n1641), .B(n1640), .Z(n1647) );
  AOI22D0BWP12T U2086 ( .A1(n1645), .A2(IF_DEC_instruction[1]), .B1(n1644), 
        .B2(n1711), .ZN(n1646) );
  OAI211D1BWP12T U2087 ( .A1(n1649), .A2(n1648), .B(n1647), .C(n1646), .ZN(
        n1654) );
  AOI22D0BWP12T U2088 ( .A1(n1654), .A2(n1696), .B1(n1650), .B2(
        IF_DEC_instruction[1]), .ZN(n1651) );
  MOAI22D0BWP12T U2089 ( .A1(n1651), .A2(n1743), .B1(n1742), .B2(
        DEC_RF_memory_store_data_reg[1]), .ZN(n829) );
  AOI222D0BWP12T U2090 ( .A1(n1654), .A2(n1738), .B1(n1711), .B2(n1653), .C1(
        IF_DEC_instruction[1]), .C2(n1652), .ZN(n1655) );
  MOAI22D0BWP12T U2091 ( .A1(n1655), .A2(n1743), .B1(n1742), .B2(
        DEC_RF_memory_write_to_reg[1]), .ZN(n823) );
  IOA21D1BWP12T U2092 ( .A1(n1742), .A2(DEC_RF_memory_store_address_reg[4]), 
        .B(n1656), .ZN(n831) );
  IOA21D1BWP12T U2093 ( .A1(n1742), .A2(DEC_RF_memory_store_address_reg[3]), 
        .B(n1657), .ZN(n832) );
  AO211D0BWP12T U2094 ( .A1(n1711), .A2(n1666), .B(n1659), .C(n1658), .Z(n1660) );
  AOI21D0BWP12T U2095 ( .A1(IF_DEC_instruction[1]), .A2(n1667), .B(n1660), 
        .ZN(n1661) );
  MOAI22D0BWP12T U2096 ( .A1(n1661), .A2(n1743), .B1(n1742), .B2(
        DEC_RF_alu_write_to_reg[1]), .ZN(n819) );
  AOI22D0BWP12T U2097 ( .A1(n1667), .A2(IF_DEC_instruction[2]), .B1(n1701), 
        .B2(n1666), .ZN(n1669) );
  AOI21D0BWP12T U2098 ( .A1(n1670), .A2(n1669), .B(n1668), .ZN(n1672) );
  AO211D0BWP12T U2099 ( .A1(n1742), .A2(DEC_RF_alu_write_to_reg[2]), .B(n1672), 
        .C(n1671), .Z(n818) );
  TPNR2D0BWP12T U2100 ( .A1(n1674), .A2(n1673), .ZN(n1675) );
  OAI211D1BWP12T U2101 ( .A1(n1678), .A2(n1677), .B(n1676), .C(n1675), .ZN(
        n1692) );
  TPND3D0BWP12T U2102 ( .A1(n1681), .A2(n1680), .A3(n1679), .ZN(n1684) );
  TPOAI31D0BWP12T U2103 ( .A1(n1692), .A2(n1684), .A3(n1683), .B(n1682), .ZN(
        n1685) );
  IOA21D1BWP12T U2104 ( .A1(DEC_ALU_alu_opcode[4]), .A2(n1742), .B(n1685), 
        .ZN(n848) );
  AOI21D0BWP12T U2105 ( .A1(n1687), .A2(n1738), .B(n1686), .ZN(n1689) );
  OAI22D0BWP12T U2106 ( .A1(n1690), .A2(n1722), .B1(n1689), .B2(n1688), .ZN(
        n1691) );
  RCAOI211D0BWP12T U2107 ( .A1(n1694), .A2(n1693), .B(n1692), .C(n1691), .ZN(
        n1695) );
  TPOAI21D0BWP12T U2108 ( .A1(n1697), .A2(n1696), .B(n1695), .ZN(n1698) );
  TPAOI31D0BWP12T U2109 ( .A1(irdecode_inst1_next_step_1_), .A2(n1699), .A3(
        n1768), .B(n1698), .ZN(n1700) );
  MOAI22D0BWP12T U2110 ( .A1(n1700), .A2(n1743), .B1(n1742), .B2(
        DEC_ALU_alu_opcode[0]), .ZN(n851) );
  AOI22D0BWP12T U2111 ( .A1(n1740), .A2(n1701), .B1(n1708), .B2(n1711), .ZN(
        n1703) );
  ND2XD0BWP12T U2112 ( .A1(n1709), .A2(IF_DEC_instruction[5]), .ZN(n1702) );
  OAI211D1BWP12T U2113 ( .A1(n1704), .A2(n1720), .B(n1703), .C(n1702), .ZN(
        n1705) );
  TPAOI21D0BWP12T U2114 ( .A1(IF_DEC_instruction[4]), .A2(n1726), .B(n1705), 
        .ZN(n1706) );
  MOAI22D0BWP12T U2115 ( .A1(n1706), .A2(n1743), .B1(n1742), .B2(
        DEC_RF_offset_b[5]), .ZN(n804) );
  AOI22D0BWP12T U2116 ( .A1(n1709), .A2(IF_DEC_instruction[4]), .B1(n1708), 
        .B2(n1707), .ZN(n1715) );
  NR2D0BWP12T U2117 ( .A1(n1710), .A2(n1739), .ZN(n1712) );
  AOI22D0BWP12T U2118 ( .A1(n1713), .A2(n1712), .B1(n1740), .B2(n1711), .ZN(
        n1714) );
  OAI211D1BWP12T U2119 ( .A1(n1716), .A2(n1720), .B(n1715), .C(n1714), .ZN(
        n1717) );
  TPAOI21D0BWP12T U2120 ( .A1(IF_DEC_instruction[3]), .A2(n1726), .B(n1717), 
        .ZN(n1718) );
  MOAI22D0BWP12T U2121 ( .A1(n1718), .A2(n1743), .B1(n1742), .B2(
        DEC_RF_offset_b[4]), .ZN(n805) );
  NR2D1BWP12T U2122 ( .A1(n1720), .A2(n1719), .ZN(n1725) );
  OAI22D0BWP12T U2123 ( .A1(n1723), .A2(n1739), .B1(n1722), .B2(n1721), .ZN(
        n1724) );
  AOI211D1BWP12T U2124 ( .A1(n1726), .A2(IF_DEC_instruction[5]), .B(n1725), 
        .C(n1724), .ZN(n1727) );
  MOAI22D0BWP12T U2125 ( .A1(n1727), .A2(n1743), .B1(n1742), .B2(
        DEC_RF_offset_b[6]), .ZN(n803) );
  OAI21D1BWP12T U2126 ( .A1(n1729), .A2(n1728), .B(n1730), .ZN(
        MEMCTRL_RF_IF_data_in[27]) );
  IOA21D1BWP12T U2127 ( .A1(n1731), .A2(MEM_MEMCTRL_from_mem_data[13]), .B(
        n1730), .ZN(MEMCTRL_RF_IF_data_in[21]) );
  IOA21D1BWP12T U2128 ( .A1(n1731), .A2(MEM_MEMCTRL_from_mem_data[12]), .B(
        n1730), .ZN(MEMCTRL_RF_IF_data_in[20]) );
  IOA21D1BWP12T U2129 ( .A1(n1731), .A2(MEM_MEMCTRL_from_mem_data[9]), .B(
        n1730), .ZN(MEMCTRL_RF_IF_data_in[17]) );
  AOI211D0BWP12T U2130 ( .A1(n1735), .A2(n1734), .B(n1733), .C(n1732), .ZN(
        n1736) );
  MOAI22D0BWP12T U2131 ( .A1(n1736), .A2(n1743), .B1(
        irdecode_inst1_split_instruction), .B2(n1742), .ZN(n847) );
  AOI21D0BWP12T U2132 ( .A1(n1739), .A2(n1738), .B(n1737), .ZN(n1741) );
  NR2D0BWP12T U2133 ( .A1(n1741), .A2(n1740), .ZN(n1744) );
  MOAI22D0BWP12T U2134 ( .A1(n1744), .A2(n1743), .B1(n1742), .B2(
        DEC_MEMCTRL_load_store_width[0]), .ZN(n838) );
endmodule

