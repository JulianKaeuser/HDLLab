
module memory_interface ( address, data_in, load, store, clk, reset, is_signed, 
        word_type, from_mem_data, to_mem_read_enable, to_mem_write_enable, 
        to_mem_mem_enable, to_mem_address, to_mem_data, data_out, write_ready, 
        output_valid, busy );
  input [11:0] address;
  input [31:0] data_in;
  input [1:0] word_type;
  input [15:0] from_mem_data;
  output [11:0] to_mem_address;
  output [15:0] to_mem_data;
  output [31:0] data_out;
  input load, store, clk, reset, is_signed;
  output to_mem_read_enable, to_mem_write_enable, to_mem_mem_enable,
         write_ready, output_valid, busy;
  wire   delayed_is_signed, fsm_N35, fsm_N34, fsm_N33, fsm_N32, fsm_state_0_,
         fsm_state_1_, fsm_state_2_, fsm_state_3_, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254;
  wire   [11:0] delay_addr_single;
  wire   [31:0] delay_data_in32;
  wire   [15:0] delay_first_two_bytes_out;

  DFQD1BWP12T delay_first_two_bytes_out_reg_15_ ( .D(from_mem_data[15]), .CP(
        clk), .Q(delay_first_two_bytes_out[15]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_14_ ( .D(from_mem_data[14]), .CP(
        clk), .Q(delay_first_two_bytes_out[14]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_13_ ( .D(from_mem_data[13]), .CP(
        clk), .Q(delay_first_two_bytes_out[13]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_12_ ( .D(from_mem_data[12]), .CP(
        clk), .Q(delay_first_two_bytes_out[12]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_11_ ( .D(from_mem_data[11]), .CP(
        clk), .Q(delay_first_two_bytes_out[11]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_10_ ( .D(from_mem_data[10]), .CP(
        clk), .Q(delay_first_two_bytes_out[10]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_9_ ( .D(from_mem_data[9]), .CP(clk), .Q(delay_first_two_bytes_out[9]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_8_ ( .D(from_mem_data[8]), .CP(clk), .Q(delay_first_two_bytes_out[8]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_7_ ( .D(from_mem_data[7]), .CP(clk), .Q(delay_first_two_bytes_out[7]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_6_ ( .D(from_mem_data[6]), .CP(clk), .Q(delay_first_two_bytes_out[6]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_5_ ( .D(from_mem_data[5]), .CP(clk), .Q(delay_first_two_bytes_out[5]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_4_ ( .D(from_mem_data[4]), .CP(clk), .Q(delay_first_two_bytes_out[4]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_3_ ( .D(from_mem_data[3]), .CP(clk), .Q(delay_first_two_bytes_out[3]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_2_ ( .D(from_mem_data[2]), .CP(clk), .Q(delay_first_two_bytes_out[2]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_1_ ( .D(from_mem_data[1]), .CP(clk), .Q(delay_first_two_bytes_out[1]) );
  DFQD1BWP12T delay_first_two_bytes_out_reg_0_ ( .D(from_mem_data[0]), .CP(clk), .Q(delay_first_two_bytes_out[0]) );
  DFQD1BWP12T delay_data_in32_reg_31_ ( .D(data_in[31]), .CP(clk), .Q(
        delay_data_in32[31]) );
  DFQD1BWP12T delay_data_in32_reg_30_ ( .D(data_in[30]), .CP(clk), .Q(
        delay_data_in32[30]) );
  DFQD1BWP12T delay_data_in32_reg_29_ ( .D(data_in[29]), .CP(clk), .Q(
        delay_data_in32[29]) );
  DFQD1BWP12T delay_data_in32_reg_28_ ( .D(data_in[28]), .CP(clk), .Q(
        delay_data_in32[28]) );
  DFQD1BWP12T delay_data_in32_reg_27_ ( .D(data_in[27]), .CP(clk), .Q(
        delay_data_in32[27]) );
  DFQD1BWP12T delay_data_in32_reg_26_ ( .D(data_in[26]), .CP(clk), .Q(
        delay_data_in32[26]) );
  DFQD1BWP12T delay_data_in32_reg_25_ ( .D(data_in[25]), .CP(clk), .Q(
        delay_data_in32[25]) );
  DFQD1BWP12T delay_data_in32_reg_24_ ( .D(data_in[24]), .CP(clk), .Q(
        delay_data_in32[24]) );
  DFQD1BWP12T delay_data_in32_reg_23_ ( .D(data_in[23]), .CP(clk), .Q(
        delay_data_in32[23]) );
  DFQD1BWP12T delay_data_in32_reg_22_ ( .D(data_in[22]), .CP(clk), .Q(
        delay_data_in32[22]) );
  DFQD1BWP12T delay_data_in32_reg_21_ ( .D(data_in[21]), .CP(clk), .Q(
        delay_data_in32[21]) );
  DFQD1BWP12T delay_data_in32_reg_20_ ( .D(data_in[20]), .CP(clk), .Q(
        delay_data_in32[20]) );
  DFQD1BWP12T delay_data_in32_reg_19_ ( .D(data_in[19]), .CP(clk), .Q(
        delay_data_in32[19]) );
  DFQD1BWP12T delay_data_in32_reg_18_ ( .D(data_in[18]), .CP(clk), .Q(
        delay_data_in32[18]) );
  DFQD1BWP12T delay_data_in32_reg_17_ ( .D(data_in[17]), .CP(clk), .Q(
        delay_data_in32[17]) );
  DFQD1BWP12T delay_data_in32_reg_16_ ( .D(data_in[16]), .CP(clk), .Q(
        delay_data_in32[16]) );
  DFQD1BWP12T delay_data_in32_reg_15_ ( .D(data_in[15]), .CP(clk), .Q(
        delay_data_in32[15]) );
  DFQD1BWP12T delay_data_in32_reg_14_ ( .D(data_in[14]), .CP(clk), .Q(
        delay_data_in32[14]) );
  DFQD1BWP12T delay_data_in32_reg_13_ ( .D(data_in[13]), .CP(clk), .Q(
        delay_data_in32[13]) );
  DFQD1BWP12T delay_data_in32_reg_12_ ( .D(data_in[12]), .CP(clk), .Q(
        delay_data_in32[12]) );
  DFQD1BWP12T delay_data_in32_reg_11_ ( .D(data_in[11]), .CP(clk), .Q(
        delay_data_in32[11]) );
  DFQD1BWP12T delay_data_in32_reg_10_ ( .D(data_in[10]), .CP(clk), .Q(
        delay_data_in32[10]) );
  DFQD1BWP12T delay_data_in32_reg_9_ ( .D(data_in[9]), .CP(clk), .Q(
        delay_data_in32[9]) );
  DFQD1BWP12T delay_data_in32_reg_8_ ( .D(data_in[8]), .CP(clk), .Q(
        delay_data_in32[8]) );
  DFQD1BWP12T delay_data_in32_reg_7_ ( .D(data_in[7]), .CP(clk), .Q(
        delay_data_in32[7]) );
  DFQD1BWP12T delay_data_in32_reg_6_ ( .D(data_in[6]), .CP(clk), .Q(
        delay_data_in32[6]) );
  DFQD1BWP12T delay_data_in32_reg_5_ ( .D(data_in[5]), .CP(clk), .Q(
        delay_data_in32[5]) );
  DFQD1BWP12T delay_data_in32_reg_4_ ( .D(data_in[4]), .CP(clk), .Q(
        delay_data_in32[4]) );
  DFQD1BWP12T delay_data_in32_reg_3_ ( .D(data_in[3]), .CP(clk), .Q(
        delay_data_in32[3]) );
  DFQD1BWP12T delay_data_in32_reg_2_ ( .D(data_in[2]), .CP(clk), .Q(
        delay_data_in32[2]) );
  DFQD1BWP12T delay_data_in32_reg_1_ ( .D(data_in[1]), .CP(clk), .Q(
        delay_data_in32[1]) );
  DFQD1BWP12T delay_data_in32_reg_0_ ( .D(data_in[0]), .CP(clk), .Q(
        delay_data_in32[0]) );
  DFQD1BWP12T delay_addr_single_reg_11_ ( .D(address[11]), .CP(clk), .Q(
        delay_addr_single[11]) );
  DFQD1BWP12T delay_addr_single_reg_10_ ( .D(address[10]), .CP(clk), .Q(
        delay_addr_single[10]) );
  DFQD1BWP12T delay_addr_single_reg_9_ ( .D(address[9]), .CP(clk), .Q(
        delay_addr_single[9]) );
  DFQD1BWP12T delay_addr_single_reg_8_ ( .D(address[8]), .CP(clk), .Q(
        delay_addr_single[8]) );
  DFQD1BWP12T delay_addr_single_reg_7_ ( .D(address[7]), .CP(clk), .Q(
        delay_addr_single[7]) );
  DFQD1BWP12T delay_addr_single_reg_6_ ( .D(address[6]), .CP(clk), .Q(
        delay_addr_single[6]) );
  DFQD1BWP12T delay_addr_single_reg_5_ ( .D(address[5]), .CP(clk), .Q(
        delay_addr_single[5]) );
  DFQD1BWP12T delay_addr_single_reg_4_ ( .D(address[4]), .CP(clk), .Q(
        delay_addr_single[4]) );
  DFQD1BWP12T delay_addr_single_reg_3_ ( .D(address[3]), .CP(clk), .Q(
        delay_addr_single[3]) );
  DFQD1BWP12T delay_addr_single_reg_2_ ( .D(address[2]), .CP(clk), .Q(
        delay_addr_single[2]) );
  DFQD1BWP12T delay_addr_single_reg_1_ ( .D(address[1]), .CP(clk), .Q(
        delay_addr_single[1]) );
  DFQD1BWP12T delay_addr_single_reg_0_ ( .D(address[0]), .CP(clk), .Q(
        delay_addr_single[0]) );
  DFQD1BWP12T delayed_is_signed_reg ( .D(is_signed), .CP(clk), .Q(
        delayed_is_signed) );
  DFXD1BWP12T fsm_state_reg_1_ ( .D(fsm_N33), .CP(clk), .Q(fsm_state_1_), .QN(
        n252) );
  DFXD1BWP12T fsm_state_reg_2_ ( .D(fsm_N34), .CP(clk), .Q(fsm_state_2_), .QN(
        n254) );
  DFXD1BWP12T fsm_state_reg_3_ ( .D(fsm_N35), .CP(clk), .Q(fsm_state_3_), .QN(
        n253) );
  DFXD1BWP12T fsm_state_reg_0_ ( .D(fsm_N32), .CP(clk), .Q(fsm_state_0_), .QN(
        n251) );
  TIELBWP12T U191 ( .ZN(n120) );
  INVD1BWP12T U192 ( .I(n120), .ZN(to_mem_mem_enable) );
  NR3D1BWP12T U193 ( .A1(fsm_state_1_), .A2(fsm_state_2_), .A3(fsm_state_3_), 
        .ZN(n134) );
  INVD1BWP12T U194 ( .I(n134), .ZN(n216) );
  INVD1BWP12T U195 ( .I(n206), .ZN(n215) );
  NR2D1BWP12T U196 ( .A1(fsm_state_0_), .A2(n216), .ZN(n206) );
  INVD1BWP12T U197 ( .I(store), .ZN(n132) );
  NR2D1BWP12T U198 ( .A1(fsm_state_2_), .A2(n252), .ZN(n131) );
  MAOI22D0BWP12T U199 ( .A1(word_type[0]), .A2(n133), .B1(word_type[0]), .B2(
        n133), .ZN(n234) );
  NR3D1BWP12T U200 ( .A1(load), .A2(n132), .A3(n215), .ZN(n230) );
  INVD1BWP12T U201 ( .I(word_type[1]), .ZN(n133) );
  OA211D0BWP12T U202 ( .A1(n219), .A2(delayed_is_signed), .B(n249), .C(n218), 
        .Z(n121) );
  CKND2D0BWP12T U203 ( .A1(n217), .A2(n121), .ZN(n228) );
  CKND0BWP12T U204 ( .I(delayed_is_signed), .ZN(n122) );
  OAI211D0BWP12T U205 ( .A1(n219), .A2(n122), .B(n217), .C(n215), .ZN(n123) );
  CKND2D0BWP12T U206 ( .A1(from_mem_data[15]), .A2(delayed_is_signed), .ZN(
        n124) );
  NR2D0BWP12T U207 ( .A1(n214), .A2(n124), .ZN(n125) );
  MOAI22D0BWP12T U208 ( .A1(n123), .A2(n125), .B1(n123), .B2(n249), .ZN(n240)
         );
  IND3D0BWP12T U209 ( .A1(write_ready), .B1(n219), .B2(n218), .ZN(n236) );
  IOA21D0BWP12T U210 ( .A1(word_type[1]), .A2(word_type[0]), .B(n230), .ZN(
        n233) );
  INR2D0BWP12T U211 ( .A1(n230), .B1(n234), .ZN(n126) );
  AOI31D0BWP12T U212 ( .A1(fsm_state_0_), .A2(n253), .A3(n131), .B(n126), .ZN(
        n127) );
  AOI21D0BWP12T U213 ( .A1(n127), .A2(n232), .B(reset), .ZN(fsm_N34) );
  AO222D0BWP12T U214 ( .A1(delay_addr_single[9]), .A2(n239), .B1(n236), .B2(
        address[9]), .C1(n238), .C2(n237), .Z(to_mem_address[9]) );
  MAOI22D0BWP12T U215 ( .A1(n230), .A2(n133), .B1(word_type[0]), .B2(n235), 
        .ZN(n128) );
  AOI21D0BWP12T U216 ( .A1(n231), .A2(n128), .B(reset), .ZN(fsm_N33) );
  CKND2D0BWP12T U217 ( .A1(n131), .A2(n251), .ZN(n129) );
  OR2XD0BWP12T U218 ( .A1(n129), .A2(fsm_state_3_), .Z(n219) );
  NR4D0BWP12T U219 ( .A1(fsm_state_1_), .A2(fsm_state_0_), .A3(fsm_state_3_), 
        .A4(n254), .ZN(n241) );
  INVD1BWP12T U220 ( .I(n241), .ZN(n250) );
  CKND2D0BWP12T U221 ( .A1(fsm_state_0_), .A2(n134), .ZN(n214) );
  ND3D1BWP12T U222 ( .A1(n219), .A2(n250), .A3(n214), .ZN(output_valid) );
  ND4D1BWP12T U223 ( .A1(fsm_state_2_), .A2(fsm_state_0_), .A3(fsm_state_3_), 
        .A4(n252), .ZN(n232) );
  CKND1BWP12T U224 ( .I(n232), .ZN(n208) );
  OAI221D0BWP12T U225 ( .A1(fsm_state_1_), .A2(n251), .B1(n252), .B2(
        fsm_state_0_), .C(fsm_state_2_), .ZN(n130) );
  AOI21D0BWP12T U226 ( .A1(n130), .A2(n129), .B(n253), .ZN(write_ready) );
  RCAOI211D0BWP12T U227 ( .A1(fsm_state_0_), .A2(n131), .B(n208), .C(
        write_ready), .ZN(n217) );
  IND2D1BWP12T U228 ( .A1(output_valid), .B1(n217), .ZN(busy) );
  INVD1BWP12T U229 ( .I(busy), .ZN(n213) );
  OAI21D1BWP12T U230 ( .A1(word_type[0]), .A2(word_type[1]), .B(n213), .ZN(
        n211) );
  ND3D1BWP12T U231 ( .A1(fsm_state_0_), .A2(fsm_state_3_), .A3(n131), .ZN(n231) );
  OAI211D0BWP12T U232 ( .A1(n211), .A2(n132), .B(n232), .C(n231), .ZN(
        to_mem_write_enable) );
  CKND2D1BWP12T U233 ( .A1(n206), .A2(load), .ZN(n235) );
  INVD1BWP12T U234 ( .I(delay_addr_single[10]), .ZN(n141) );
  ND3D1BWP12T U235 ( .A1(delay_addr_single[0]), .A2(delay_addr_single[1]), 
        .A3(delay_addr_single[2]), .ZN(n163) );
  INVD1BWP12T U236 ( .I(n163), .ZN(n160) );
  ND2D1BWP12T U237 ( .A1(n160), .A2(delay_addr_single[3]), .ZN(n159) );
  IND2D1BWP12T U238 ( .A1(n159), .B1(delay_addr_single[4]), .ZN(n156) );
  INVD1BWP12T U239 ( .I(n156), .ZN(n153) );
  ND2D1BWP12T U240 ( .A1(n153), .A2(delay_addr_single[5]), .ZN(n152) );
  IND2D1BWP12T U241 ( .A1(n152), .B1(delay_addr_single[6]), .ZN(n149) );
  INVD1BWP12T U242 ( .I(n149), .ZN(n146) );
  ND2D1BWP12T U243 ( .A1(n146), .A2(delay_addr_single[7]), .ZN(n145) );
  INR2D1BWP12T U244 ( .A1(delay_addr_single[8]), .B1(n145), .ZN(n135) );
  NR2D0BWP12T U245 ( .A1(n134), .A2(n241), .ZN(n218) );
  OAI32D0BWP12T U246 ( .A1(fsm_state_3_), .A2(fsm_state_1_), .A3(fsm_state_0_), 
        .B1(fsm_state_2_), .B2(fsm_state_3_), .ZN(n212) );
  NR2D1BWP12T U247 ( .A1(write_ready), .A2(n212), .ZN(n190) );
  CKND2D1BWP12T U248 ( .A1(n190), .A2(n232), .ZN(n167) );
  INVD1BWP12T U249 ( .I(n167), .ZN(n187) );
  NR2D1BWP12T U250 ( .A1(n236), .A2(n187), .ZN(n136) );
  INVD1BWP12T U251 ( .I(n136), .ZN(n171) );
  INR2D1BWP12T U252 ( .A1(n135), .B1(n171), .ZN(n238) );
  ND2D1BWP12T U253 ( .A1(delay_addr_single[9]), .A2(n238), .ZN(n142) );
  INVD1BWP12T U254 ( .I(delay_addr_single[9]), .ZN(n237) );
  OAI21D1BWP12T U255 ( .A1(n135), .A2(n171), .B(n167), .ZN(n239) );
  AOI21D1BWP12T U256 ( .A1(n136), .A2(n237), .B(n239), .ZN(n140) );
  OAI21D1BWP12T U257 ( .A1(delay_addr_single[10]), .A2(n171), .B(n140), .ZN(
        n137) );
  AOI22D1BWP12T U258 ( .A1(delay_addr_single[11]), .A2(n137), .B1(address[11]), 
        .B2(n236), .ZN(n138) );
  OAI31D1BWP12T U259 ( .A1(delay_addr_single[11]), .A2(n141), .A3(n142), .B(
        n138), .ZN(to_mem_address[11]) );
  ND2D1BWP12T U260 ( .A1(address[10]), .A2(n236), .ZN(n139) );
  OAI221D1BWP12T U261 ( .A1(delay_addr_single[10]), .A2(n142), .B1(n141), .B2(
        n140), .C(n139), .ZN(to_mem_address[10]) );
  AOI31D1BWP12T U262 ( .A1(n146), .A2(delay_addr_single[7]), .A3(n167), .B(
        n236), .ZN(n143) );
  AOI22D1BWP12T U263 ( .A1(delay_addr_single[8]), .A2(n143), .B1(address[8]), 
        .B2(n236), .ZN(n144) );
  OAI31D1BWP12T U264 ( .A1(delay_addr_single[8]), .A2(n171), .A3(n145), .B(
        n144), .ZN(to_mem_address[8]) );
  OAI21D1BWP12T U265 ( .A1(n236), .A2(n146), .B(n167), .ZN(n147) );
  AOI22D1BWP12T U266 ( .A1(delay_addr_single[7]), .A2(n147), .B1(address[7]), 
        .B2(n236), .ZN(n148) );
  OAI31D1BWP12T U267 ( .A1(delay_addr_single[7]), .A2(n171), .A3(n149), .B(
        n148), .ZN(to_mem_address[7]) );
  AOI31D1BWP12T U268 ( .A1(n153), .A2(delay_addr_single[5]), .A3(n167), .B(
        n236), .ZN(n150) );
  AOI22D1BWP12T U269 ( .A1(delay_addr_single[6]), .A2(n150), .B1(address[6]), 
        .B2(n236), .ZN(n151) );
  OAI31D1BWP12T U270 ( .A1(delay_addr_single[6]), .A2(n171), .A3(n152), .B(
        n151), .ZN(to_mem_address[6]) );
  OAI21D1BWP12T U271 ( .A1(n236), .A2(n153), .B(n167), .ZN(n154) );
  AOI22D1BWP12T U272 ( .A1(delay_addr_single[5]), .A2(n154), .B1(address[5]), 
        .B2(n236), .ZN(n155) );
  OAI31D1BWP12T U273 ( .A1(delay_addr_single[5]), .A2(n171), .A3(n156), .B(
        n155), .ZN(to_mem_address[5]) );
  AOI31D1BWP12T U274 ( .A1(n160), .A2(delay_addr_single[3]), .A3(n167), .B(
        n236), .ZN(n157) );
  AOI22D1BWP12T U275 ( .A1(delay_addr_single[4]), .A2(n157), .B1(address[4]), 
        .B2(n236), .ZN(n158) );
  OAI31D1BWP12T U276 ( .A1(delay_addr_single[4]), .A2(n171), .A3(n159), .B(
        n158), .ZN(to_mem_address[4]) );
  OAI21D1BWP12T U277 ( .A1(n236), .A2(n160), .B(n167), .ZN(n161) );
  AOI22D1BWP12T U278 ( .A1(delay_addr_single[3]), .A2(n161), .B1(address[3]), 
        .B2(n236), .ZN(n162) );
  OAI31D1BWP12T U279 ( .A1(delay_addr_single[3]), .A2(n171), .A3(n163), .B(
        n162), .ZN(to_mem_address[3]) );
  ND2D1BWP12T U280 ( .A1(delay_addr_single[0]), .A2(delay_addr_single[1]), 
        .ZN(n166) );
  AOI31D1BWP12T U281 ( .A1(delay_addr_single[0]), .A2(delay_addr_single[1]), 
        .A3(n167), .B(n236), .ZN(n164) );
  AOI22D1BWP12T U282 ( .A1(delay_addr_single[2]), .A2(n164), .B1(address[2]), 
        .B2(n236), .ZN(n165) );
  OAI31D1BWP12T U283 ( .A1(delay_addr_single[2]), .A2(n171), .A3(n166), .B(
        n165), .ZN(to_mem_address[2]) );
  OAI21D1BWP12T U284 ( .A1(delay_addr_single[0]), .A2(n236), .B(n167), .ZN(
        n169) );
  NR2D1BWP12T U285 ( .A1(delay_addr_single[1]), .A2(n171), .ZN(n168) );
  AO222D1BWP12T U286 ( .A1(n169), .A2(delay_addr_single[1]), .B1(n236), .B2(
        address[1]), .C1(delay_addr_single[0]), .C2(n168), .Z(
        to_mem_address[1]) );
  AOI22D1BWP12T U287 ( .A1(n187), .A2(delay_addr_single[0]), .B1(address[0]), 
        .B2(n236), .ZN(n170) );
  OAI21D1BWP12T U288 ( .A1(delay_addr_single[0]), .A2(n171), .B(n170), .ZN(
        to_mem_address[0]) );
  RCAOI21D0BWP12T U289 ( .A1(n190), .A2(n231), .B(n213), .ZN(n205) );
  INR2D1BWP12T U290 ( .A1(n205), .B1(n187), .ZN(n186) );
  AOI22D1BWP12T U291 ( .A1(n187), .A2(from_mem_data[15]), .B1(n186), .B2(
        delay_data_in32[15]), .ZN(n173) );
  AOI22D0BWP12T U292 ( .A1(n208), .A2(delay_data_in32[31]), .B1(n206), .B2(
        data_in[15]), .ZN(n172) );
  ND2D1BWP12T U293 ( .A1(n173), .A2(n172), .ZN(to_mem_data[15]) );
  AOI22D1BWP12T U294 ( .A1(n187), .A2(from_mem_data[14]), .B1(n186), .B2(
        delay_data_in32[14]), .ZN(n175) );
  AOI22D0BWP12T U295 ( .A1(n208), .A2(delay_data_in32[30]), .B1(n206), .B2(
        data_in[14]), .ZN(n174) );
  ND2D1BWP12T U296 ( .A1(n175), .A2(n174), .ZN(to_mem_data[14]) );
  AOI22D1BWP12T U297 ( .A1(n187), .A2(from_mem_data[13]), .B1(n186), .B2(
        delay_data_in32[13]), .ZN(n177) );
  AOI22D0BWP12T U298 ( .A1(n208), .A2(delay_data_in32[29]), .B1(n206), .B2(
        data_in[13]), .ZN(n176) );
  ND2D1BWP12T U299 ( .A1(n177), .A2(n176), .ZN(to_mem_data[13]) );
  AOI22D1BWP12T U300 ( .A1(n187), .A2(from_mem_data[12]), .B1(n186), .B2(
        delay_data_in32[12]), .ZN(n179) );
  AOI22D0BWP12T U301 ( .A1(n208), .A2(delay_data_in32[28]), .B1(n206), .B2(
        data_in[12]), .ZN(n178) );
  ND2D1BWP12T U302 ( .A1(n179), .A2(n178), .ZN(to_mem_data[12]) );
  AOI22D1BWP12T U303 ( .A1(n187), .A2(from_mem_data[11]), .B1(n186), .B2(
        delay_data_in32[11]), .ZN(n181) );
  AOI22D0BWP12T U304 ( .A1(n208), .A2(delay_data_in32[27]), .B1(n206), .B2(
        data_in[11]), .ZN(n180) );
  ND2D1BWP12T U305 ( .A1(n181), .A2(n180), .ZN(to_mem_data[11]) );
  AOI22D1BWP12T U306 ( .A1(n187), .A2(from_mem_data[10]), .B1(n186), .B2(
        delay_data_in32[10]), .ZN(n183) );
  AOI22D0BWP12T U307 ( .A1(n208), .A2(delay_data_in32[26]), .B1(n206), .B2(
        data_in[10]), .ZN(n182) );
  ND2D1BWP12T U308 ( .A1(n183), .A2(n182), .ZN(to_mem_data[10]) );
  AOI22D1BWP12T U309 ( .A1(n187), .A2(from_mem_data[9]), .B1(n186), .B2(
        delay_data_in32[9]), .ZN(n185) );
  AOI22D0BWP12T U310 ( .A1(n208), .A2(delay_data_in32[25]), .B1(n206), .B2(
        data_in[9]), .ZN(n184) );
  ND2D1BWP12T U311 ( .A1(n185), .A2(n184), .ZN(to_mem_data[9]) );
  AOI22D1BWP12T U312 ( .A1(n187), .A2(from_mem_data[8]), .B1(n186), .B2(
        delay_data_in32[8]), .ZN(n189) );
  AOI22D0BWP12T U313 ( .A1(n208), .A2(delay_data_in32[24]), .B1(n206), .B2(
        data_in[8]), .ZN(n188) );
  ND2D1BWP12T U314 ( .A1(n189), .A2(n188), .ZN(to_mem_data[8]) );
  AOI22D0BWP12T U315 ( .A1(n206), .A2(data_in[7]), .B1(n205), .B2(
        delay_data_in32[7]), .ZN(n192) );
  AN2D1BWP12T U316 ( .A1(n190), .A2(n213), .Z(n207) );
  AOI22D1BWP12T U317 ( .A1(n208), .A2(delay_data_in32[23]), .B1(n207), .B2(
        data_in[23]), .ZN(n191) );
  ND2D1BWP12T U318 ( .A1(n192), .A2(n191), .ZN(to_mem_data[7]) );
  AOI22D0BWP12T U319 ( .A1(n206), .A2(data_in[6]), .B1(n205), .B2(
        delay_data_in32[6]), .ZN(n194) );
  AOI22D1BWP12T U320 ( .A1(n208), .A2(delay_data_in32[22]), .B1(n207), .B2(
        data_in[22]), .ZN(n193) );
  ND2D1BWP12T U321 ( .A1(n194), .A2(n193), .ZN(to_mem_data[6]) );
  AOI22D0BWP12T U322 ( .A1(n206), .A2(data_in[5]), .B1(n205), .B2(
        delay_data_in32[5]), .ZN(n196) );
  AOI22D1BWP12T U323 ( .A1(n208), .A2(delay_data_in32[21]), .B1(n207), .B2(
        data_in[21]), .ZN(n195) );
  ND2D1BWP12T U324 ( .A1(n196), .A2(n195), .ZN(to_mem_data[5]) );
  AOI22D0BWP12T U325 ( .A1(n206), .A2(data_in[4]), .B1(n205), .B2(
        delay_data_in32[4]), .ZN(n198) );
  AOI22D1BWP12T U326 ( .A1(n208), .A2(delay_data_in32[20]), .B1(n207), .B2(
        data_in[20]), .ZN(n197) );
  ND2D1BWP12T U327 ( .A1(n198), .A2(n197), .ZN(to_mem_data[4]) );
  AOI22D0BWP12T U328 ( .A1(n206), .A2(data_in[3]), .B1(n205), .B2(
        delay_data_in32[3]), .ZN(n200) );
  AOI22D1BWP12T U329 ( .A1(n208), .A2(delay_data_in32[19]), .B1(n207), .B2(
        data_in[19]), .ZN(n199) );
  ND2D1BWP12T U330 ( .A1(n200), .A2(n199), .ZN(to_mem_data[3]) );
  AOI22D0BWP12T U331 ( .A1(n206), .A2(data_in[2]), .B1(n205), .B2(
        delay_data_in32[2]), .ZN(n202) );
  AOI22D1BWP12T U332 ( .A1(n208), .A2(delay_data_in32[18]), .B1(n207), .B2(
        data_in[18]), .ZN(n201) );
  ND2D1BWP12T U333 ( .A1(n202), .A2(n201), .ZN(to_mem_data[2]) );
  AOI22D0BWP12T U334 ( .A1(n206), .A2(data_in[1]), .B1(n205), .B2(
        delay_data_in32[1]), .ZN(n204) );
  AOI22D1BWP12T U335 ( .A1(n208), .A2(delay_data_in32[17]), .B1(n207), .B2(
        data_in[17]), .ZN(n203) );
  ND2D1BWP12T U336 ( .A1(n204), .A2(n203), .ZN(to_mem_data[1]) );
  AOI22D0BWP12T U337 ( .A1(n206), .A2(data_in[0]), .B1(n205), .B2(
        delay_data_in32[0]), .ZN(n210) );
  AOI22D1BWP12T U338 ( .A1(n208), .A2(delay_data_in32[16]), .B1(n207), .B2(
        data_in[16]), .ZN(n209) );
  ND2D1BWP12T U339 ( .A1(n210), .A2(n209), .ZN(to_mem_data[0]) );
  OA22D1BWP12T U340 ( .A1(n213), .A2(n212), .B1(load), .B2(n211), .Z(
        to_mem_read_enable) );
  INVD1BWP12T U341 ( .I(from_mem_data[7]), .ZN(n249) );
  OAI21D1BWP12T U342 ( .A1(n249), .A2(n250), .B(n240), .ZN(data_out[23]) );
  INVD1BWP12T U343 ( .I(from_mem_data[6]), .ZN(n248) );
  OAI21D1BWP12T U344 ( .A1(n250), .A2(n248), .B(n240), .ZN(data_out[22]) );
  INVD1BWP12T U345 ( .I(from_mem_data[5]), .ZN(n247) );
  OAI21D1BWP12T U346 ( .A1(n250), .A2(n247), .B(n240), .ZN(data_out[21]) );
  INVD1BWP12T U347 ( .I(from_mem_data[4]), .ZN(n246) );
  OAI21D1BWP12T U348 ( .A1(n250), .A2(n246), .B(n240), .ZN(data_out[20]) );
  INVD1BWP12T U349 ( .I(from_mem_data[3]), .ZN(n245) );
  OAI21D1BWP12T U350 ( .A1(n250), .A2(n245), .B(n240), .ZN(data_out[19]) );
  INVD1BWP12T U351 ( .I(from_mem_data[2]), .ZN(n244) );
  OAI21D1BWP12T U352 ( .A1(n250), .A2(n244), .B(n240), .ZN(data_out[18]) );
  INVD1BWP12T U353 ( .I(from_mem_data[1]), .ZN(n243) );
  OAI21D1BWP12T U354 ( .A1(n250), .A2(n243), .B(n240), .ZN(data_out[17]) );
  INVD1BWP12T U355 ( .I(from_mem_data[0]), .ZN(n242) );
  OAI21D1BWP12T U356 ( .A1(n250), .A2(n242), .B(n240), .ZN(data_out[16]) );
  CKND2D1BWP12T U357 ( .A1(n216), .A2(n217), .ZN(n227) );
  AOI22D1BWP12T U358 ( .A1(n241), .A2(delay_first_two_bytes_out[15]), .B1(
        from_mem_data[15]), .B2(n227), .ZN(n220) );
  ND2D1BWP12T U359 ( .A1(n220), .A2(n228), .ZN(data_out[15]) );
  AOI22D1BWP12T U360 ( .A1(n241), .A2(delay_first_two_bytes_out[14]), .B1(
        from_mem_data[14]), .B2(n227), .ZN(n221) );
  ND2D1BWP12T U361 ( .A1(n221), .A2(n228), .ZN(data_out[14]) );
  AOI22D1BWP12T U362 ( .A1(n241), .A2(delay_first_two_bytes_out[13]), .B1(
        from_mem_data[13]), .B2(n227), .ZN(n222) );
  ND2D1BWP12T U363 ( .A1(n222), .A2(n228), .ZN(data_out[13]) );
  AOI22D1BWP12T U364 ( .A1(n241), .A2(delay_first_two_bytes_out[12]), .B1(
        from_mem_data[12]), .B2(n227), .ZN(n223) );
  ND2D1BWP12T U365 ( .A1(n223), .A2(n228), .ZN(data_out[12]) );
  AOI22D1BWP12T U366 ( .A1(n241), .A2(delay_first_two_bytes_out[11]), .B1(
        from_mem_data[11]), .B2(n227), .ZN(n224) );
  ND2D1BWP12T U367 ( .A1(n224), .A2(n228), .ZN(data_out[11]) );
  AOI22D1BWP12T U368 ( .A1(n241), .A2(delay_first_two_bytes_out[10]), .B1(
        from_mem_data[10]), .B2(n227), .ZN(n225) );
  ND2D1BWP12T U369 ( .A1(n225), .A2(n228), .ZN(data_out[10]) );
  AOI22D1BWP12T U370 ( .A1(n241), .A2(delay_first_two_bytes_out[9]), .B1(
        from_mem_data[9]), .B2(n227), .ZN(n226) );
  ND2D1BWP12T U371 ( .A1(n226), .A2(n228), .ZN(data_out[9]) );
  AOI22D1BWP12T U372 ( .A1(n241), .A2(delay_first_two_bytes_out[8]), .B1(
        from_mem_data[8]), .B2(n227), .ZN(n229) );
  ND2D1BWP12T U373 ( .A1(n229), .A2(n228), .ZN(data_out[8]) );
  AOI31D1BWP12T U374 ( .A1(n232), .A2(n231), .A3(n233), .B(reset), .ZN(fsm_N35) );
  OAI32D1BWP12T U375 ( .A1(reset), .A2(n235), .A3(n234), .B1(n233), .B2(reset), 
        .ZN(fsm_N32) );
  IOA21D1BWP12T U376 ( .A1(from_mem_data[15]), .A2(n241), .B(n240), .ZN(
        data_out[31]) );
  IOA21D1BWP12T U377 ( .A1(from_mem_data[14]), .A2(n241), .B(n240), .ZN(
        data_out[30]) );
  IOA21D1BWP12T U378 ( .A1(from_mem_data[13]), .A2(n241), .B(n240), .ZN(
        data_out[29]) );
  IOA21D1BWP12T U379 ( .A1(from_mem_data[12]), .A2(n241), .B(n240), .ZN(
        data_out[28]) );
  IOA21D1BWP12T U380 ( .A1(from_mem_data[11]), .A2(n241), .B(n240), .ZN(
        data_out[27]) );
  IOA21D1BWP12T U381 ( .A1(from_mem_data[10]), .A2(n241), .B(n240), .ZN(
        data_out[26]) );
  IOA21D1BWP12T U382 ( .A1(from_mem_data[9]), .A2(n241), .B(n240), .ZN(
        data_out[25]) );
  IOA21D1BWP12T U383 ( .A1(from_mem_data[8]), .A2(n241), .B(n240), .ZN(
        data_out[24]) );
  MAOI22D0BWP12T U384 ( .A1(n250), .A2(n242), .B1(n250), .B2(
        delay_first_two_bytes_out[0]), .ZN(data_out[0]) );
  MAOI22D0BWP12T U385 ( .A1(n250), .A2(n243), .B1(n250), .B2(
        delay_first_two_bytes_out[1]), .ZN(data_out[1]) );
  MAOI22D0BWP12T U386 ( .A1(n250), .A2(n244), .B1(n250), .B2(
        delay_first_two_bytes_out[2]), .ZN(data_out[2]) );
  MAOI22D0BWP12T U387 ( .A1(n250), .A2(n245), .B1(n250), .B2(
        delay_first_two_bytes_out[3]), .ZN(data_out[3]) );
  MAOI22D0BWP12T U388 ( .A1(n250), .A2(n246), .B1(n250), .B2(
        delay_first_two_bytes_out[4]), .ZN(data_out[4]) );
  MAOI22D0BWP12T U389 ( .A1(n250), .A2(n247), .B1(n250), .B2(
        delay_first_two_bytes_out[5]), .ZN(data_out[5]) );
  MAOI22D0BWP12T U390 ( .A1(n250), .A2(n248), .B1(n250), .B2(
        delay_first_two_bytes_out[6]), .ZN(data_out[6]) );
  MAOI22D0BWP12T U391 ( .A1(n250), .A2(n249), .B1(n250), .B2(
        delay_first_two_bytes_out[7]), .ZN(data_out[7]) );
endmodule

