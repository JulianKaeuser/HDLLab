module register_file_tb ();


// some test cases
endmodule
