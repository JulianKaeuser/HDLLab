`define BIT_SIZE 16
`timescale 1ns/100ps

module ALU_VARIABLE_tb();
	reg signed [`BIT_SIZE-1:0] a, b;
	reg c_in;
	reg [3:0] op;
	wire c_out, z, n, v;
	wire [`BIT_SIZE-1:0] result;

ALU_VARIABLE alu_inst(
	.a(a), .b(b), .c_in(c_in), .op(op), .c_out(c_out), .z(z), .n(n), .v(v), .result(result)
);

initial begin
	$monitor("%g\t a: %b b: %b c_in: %b op: %b | c_out: %b z: %b n: %b v: %b result: %b", $time, a, b, c_in, op, c_out, z, n, v, result);
	
	a = 16'b0101110010110001;

	b = 16'b1000111010011011;

	/*op = 4'b1100; // ORR
	#1;
	op = 4'b0000; // AND
	#1;
	op = 4'b1110; //BIC
	#1;
	op = 4'b0001; //EOR
	#1;
	$display("=================================================================================================");
	
	b = 16'b0000000000001011;
	op = 4'b0010; //LSL
	#1;
	op = 4'b0011; //LSR
	#1;
	op = 4'b0100; //ASR
	#1;
	op = 4'b0111; //ROR
	#1;
	$display("=================================================================================================");
	op = 4'b1111; // MVN
	#1;
	op = 4'b1001; //NEG
	#1;
	$display("=================================================================================================");
	c_in = 0;
	op = 4'b0101; // ADC
	#1;
	c_in = 1;
	#1;
	//b = 16'b1100111010011011;
	#1;
	c_in = 0;
	op = 4'b0110; // SBC
	#1;
	c_in = 1;
	//a =  16'b0000000000000001;
	//b = 16'b0111111111111111;
	#1;
	op = 4'b1000; //TST
	#1;
	op = 4'b1010; //CMP
	#1;
	op = 4'b1011; //CMN
	#1;*/
	$display("=================================================================================================");
	//a = 16'b1111111111111111;
	//sb = 16'b0111111111111111;
	a = a[`BIT_SIZE / 2 - 1:0];

	b = b[`BIT_SIZE / 2 - 1:0];
	op = 4'b1101; // MUL
	#1;
	$display("=================================================================================================");

end

endmodule